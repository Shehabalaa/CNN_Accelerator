LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY DFFZ IS
	PORT(
		D: in std_logic;
		clk, rst, en: in std_logic;
		Q: out std_logic
		);
END DFFZ;

Architecture DFFZArch OF DFFZ IS 
BEGIN

END ARCHITECTURE;
