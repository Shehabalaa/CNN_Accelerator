library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity IODFF is
   port (
      D : IN std_logic ;
      clk : IN std_logic ;
      rst : IN std_logic ;
      en : IN std_logic ;
      Q : OUT std_logic) ;
end IODFF ;

architecture IODFFArch of IODFF is
begin
end IODFFArch ;
