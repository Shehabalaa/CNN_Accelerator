//
// Verilog description for cell CNNMuls, 
// Thu Apr 11 12:57:10 2019
//
// LeonardoSpectrum Level 3, 2018a.2 
//


module CNNMuls ( filter_24__7, filter_24__6, filter_24__5, filter_24__4, 
                 filter_24__3, filter_24__2, filter_24__1, filter_24__0, 
                 filter_23__7, filter_23__6, filter_23__5, filter_23__4, 
                 filter_23__3, filter_23__2, filter_23__1, filter_23__0, 
                 filter_22__7, filter_22__6, filter_22__5, filter_22__4, 
                 filter_22__3, filter_22__2, filter_22__1, filter_22__0, 
                 filter_21__7, filter_21__6, filter_21__5, filter_21__4, 
                 filter_21__3, filter_21__2, filter_21__1, filter_21__0, 
                 filter_20__7, filter_20__6, filter_20__5, filter_20__4, 
                 filter_20__3, filter_20__2, filter_20__1, filter_20__0, 
                 filter_19__7, filter_19__6, filter_19__5, filter_19__4, 
                 filter_19__3, filter_19__2, filter_19__1, filter_19__0, 
                 filter_18__7, filter_18__6, filter_18__5, filter_18__4, 
                 filter_18__3, filter_18__2, filter_18__1, filter_18__0, 
                 filter_17__7, filter_17__6, filter_17__5, filter_17__4, 
                 filter_17__3, filter_17__2, filter_17__1, filter_17__0, 
                 filter_16__7, filter_16__6, filter_16__5, filter_16__4, 
                 filter_16__3, filter_16__2, filter_16__1, filter_16__0, 
                 filter_15__7, filter_15__6, filter_15__5, filter_15__4, 
                 filter_15__3, filter_15__2, filter_15__1, filter_15__0, 
                 filter_14__7, filter_14__6, filter_14__5, filter_14__4, 
                 filter_14__3, filter_14__2, filter_14__1, filter_14__0, 
                 filter_13__7, filter_13__6, filter_13__5, filter_13__4, 
                 filter_13__3, filter_13__2, filter_13__1, filter_13__0, 
                 filter_12__7, filter_12__6, filter_12__5, filter_12__4, 
                 filter_12__3, filter_12__2, filter_12__1, filter_12__0, 
                 filter_11__7, filter_11__6, filter_11__5, filter_11__4, 
                 filter_11__3, filter_11__2, filter_11__1, filter_11__0, 
                 filter_10__7, filter_10__6, filter_10__5, filter_10__4, 
                 filter_10__3, filter_10__2, filter_10__1, filter_10__0, 
                 filter_9__7, filter_9__6, filter_9__5, filter_9__4, filter_9__3, 
                 filter_9__2, filter_9__1, filter_9__0, filter_8__7, filter_8__6, 
                 filter_8__5, filter_8__4, filter_8__3, filter_8__2, filter_8__1, 
                 filter_8__0, filter_7__7, filter_7__6, filter_7__5, filter_7__4, 
                 filter_7__3, filter_7__2, filter_7__1, filter_7__0, filter_6__7, 
                 filter_6__6, filter_6__5, filter_6__4, filter_6__3, filter_6__2, 
                 filter_6__1, filter_6__0, filter_5__7, filter_5__6, filter_5__5, 
                 filter_5__4, filter_5__3, filter_5__2, filter_5__1, filter_5__0, 
                 filter_4__7, filter_4__6, filter_4__5, filter_4__4, filter_4__3, 
                 filter_4__2, filter_4__1, filter_4__0, filter_3__7, filter_3__6, 
                 filter_3__5, filter_3__4, filter_3__3, filter_3__2, filter_3__1, 
                 filter_3__0, filter_2__7, filter_2__6, filter_2__5, filter_2__4, 
                 filter_2__3, filter_2__2, filter_2__1, filter_2__0, filter_1__7, 
                 filter_1__6, filter_1__5, filter_1__4, filter_1__3, filter_1__2, 
                 filter_1__1, filter_1__0, filter_0__7, filter_0__6, filter_0__5, 
                 filter_0__4, filter_0__3, filter_0__2, filter_0__1, filter_0__0, 
                 window_24__15, window_24__14, window_24__13, window_24__12, 
                 window_24__11, window_24__10, window_24__9, window_24__8, 
                 window_24__7, window_24__6, window_24__5, window_24__4, 
                 window_24__3, window_24__2, window_24__1, window_24__0, 
                 window_23__15, window_23__14, window_23__13, window_23__12, 
                 window_23__11, window_23__10, window_23__9, window_23__8, 
                 window_23__7, window_23__6, window_23__5, window_23__4, 
                 window_23__3, window_23__2, window_23__1, window_23__0, 
                 window_22__15, window_22__14, window_22__13, window_22__12, 
                 window_22__11, window_22__10, window_22__9, window_22__8, 
                 window_22__7, window_22__6, window_22__5, window_22__4, 
                 window_22__3, window_22__2, window_22__1, window_22__0, 
                 window_21__15, window_21__14, window_21__13, window_21__12, 
                 window_21__11, window_21__10, window_21__9, window_21__8, 
                 window_21__7, window_21__6, window_21__5, window_21__4, 
                 window_21__3, window_21__2, window_21__1, window_21__0, 
                 window_20__15, window_20__14, window_20__13, window_20__12, 
                 window_20__11, window_20__10, window_20__9, window_20__8, 
                 window_20__7, window_20__6, window_20__5, window_20__4, 
                 window_20__3, window_20__2, window_20__1, window_20__0, 
                 window_19__15, window_19__14, window_19__13, window_19__12, 
                 window_19__11, window_19__10, window_19__9, window_19__8, 
                 window_19__7, window_19__6, window_19__5, window_19__4, 
                 window_19__3, window_19__2, window_19__1, window_19__0, 
                 window_18__15, window_18__14, window_18__13, window_18__12, 
                 window_18__11, window_18__10, window_18__9, window_18__8, 
                 window_18__7, window_18__6, window_18__5, window_18__4, 
                 window_18__3, window_18__2, window_18__1, window_18__0, 
                 window_17__15, window_17__14, window_17__13, window_17__12, 
                 window_17__11, window_17__10, window_17__9, window_17__8, 
                 window_17__7, window_17__6, window_17__5, window_17__4, 
                 window_17__3, window_17__2, window_17__1, window_17__0, 
                 window_16__15, window_16__14, window_16__13, window_16__12, 
                 window_16__11, window_16__10, window_16__9, window_16__8, 
                 window_16__7, window_16__6, window_16__5, window_16__4, 
                 window_16__3, window_16__2, window_16__1, window_16__0, 
                 window_15__15, window_15__14, window_15__13, window_15__12, 
                 window_15__11, window_15__10, window_15__9, window_15__8, 
                 window_15__7, window_15__6, window_15__5, window_15__4, 
                 window_15__3, window_15__2, window_15__1, window_15__0, 
                 window_14__15, window_14__14, window_14__13, window_14__12, 
                 window_14__11, window_14__10, window_14__9, window_14__8, 
                 window_14__7, window_14__6, window_14__5, window_14__4, 
                 window_14__3, window_14__2, window_14__1, window_14__0, 
                 window_13__15, window_13__14, window_13__13, window_13__12, 
                 window_13__11, window_13__10, window_13__9, window_13__8, 
                 window_13__7, window_13__6, window_13__5, window_13__4, 
                 window_13__3, window_13__2, window_13__1, window_13__0, 
                 window_12__15, window_12__14, window_12__13, window_12__12, 
                 window_12__11, window_12__10, window_12__9, window_12__8, 
                 window_12__7, window_12__6, window_12__5, window_12__4, 
                 window_12__3, window_12__2, window_12__1, window_12__0, 
                 window_11__15, window_11__14, window_11__13, window_11__12, 
                 window_11__11, window_11__10, window_11__9, window_11__8, 
                 window_11__7, window_11__6, window_11__5, window_11__4, 
                 window_11__3, window_11__2, window_11__1, window_11__0, 
                 window_10__15, window_10__14, window_10__13, window_10__12, 
                 window_10__11, window_10__10, window_10__9, window_10__8, 
                 window_10__7, window_10__6, window_10__5, window_10__4, 
                 window_10__3, window_10__2, window_10__1, window_10__0, 
                 window_9__15, window_9__14, window_9__13, window_9__12, 
                 window_9__11, window_9__10, window_9__9, window_9__8, 
                 window_9__7, window_9__6, window_9__5, window_9__4, window_9__3, 
                 window_9__2, window_9__1, window_9__0, window_8__15, 
                 window_8__14, window_8__13, window_8__12, window_8__11, 
                 window_8__10, window_8__9, window_8__8, window_8__7, 
                 window_8__6, window_8__5, window_8__4, window_8__3, window_8__2, 
                 window_8__1, window_8__0, window_7__15, window_7__14, 
                 window_7__13, window_7__12, window_7__11, window_7__10, 
                 window_7__9, window_7__8, window_7__7, window_7__6, window_7__5, 
                 window_7__4, window_7__3, window_7__2, window_7__1, window_7__0, 
                 window_6__15, window_6__14, window_6__13, window_6__12, 
                 window_6__11, window_6__10, window_6__9, window_6__8, 
                 window_6__7, window_6__6, window_6__5, window_6__4, window_6__3, 
                 window_6__2, window_6__1, window_6__0, window_5__15, 
                 window_5__14, window_5__13, window_5__12, window_5__11, 
                 window_5__10, window_5__9, window_5__8, window_5__7, 
                 window_5__6, window_5__5, window_5__4, window_5__3, window_5__2, 
                 window_5__1, window_5__0, window_4__15, window_4__14, 
                 window_4__13, window_4__12, window_4__11, window_4__10, 
                 window_4__9, window_4__8, window_4__7, window_4__6, window_4__5, 
                 window_4__4, window_4__3, window_4__2, window_4__1, window_4__0, 
                 window_3__15, window_3__14, window_3__13, window_3__12, 
                 window_3__11, window_3__10, window_3__9, window_3__8, 
                 window_3__7, window_3__6, window_3__5, window_3__4, window_3__3, 
                 window_3__2, window_3__1, window_3__0, window_2__15, 
                 window_2__14, window_2__13, window_2__12, window_2__11, 
                 window_2__10, window_2__9, window_2__8, window_2__7, 
                 window_2__6, window_2__5, window_2__4, window_2__3, window_2__2, 
                 window_2__1, window_2__0, window_1__15, window_1__14, 
                 window_1__13, window_1__12, window_1__11, window_1__10, 
                 window_1__9, window_1__8, window_1__7, window_1__6, window_1__5, 
                 window_1__4, window_1__3, window_1__2, window_1__1, window_1__0, 
                 window_0__15, window_0__14, window_0__13, window_0__12, 
                 window_0__11, window_0__10, window_0__9, window_0__8, 
                 window_0__7, window_0__6, window_0__5, window_0__4, window_0__3, 
                 window_0__2, window_0__1, window_0__0, outputs_24__15, 
                 outputs_24__14, outputs_24__13, outputs_24__12, outputs_24__11, 
                 outputs_24__10, outputs_24__9, outputs_24__8, outputs_24__7, 
                 outputs_24__6, outputs_24__5, outputs_24__4, outputs_24__3, 
                 outputs_24__2, outputs_24__1, outputs_24__0, outputs_23__15, 
                 outputs_23__14, outputs_23__13, outputs_23__12, outputs_23__11, 
                 outputs_23__10, outputs_23__9, outputs_23__8, outputs_23__7, 
                 outputs_23__6, outputs_23__5, outputs_23__4, outputs_23__3, 
                 outputs_23__2, outputs_23__1, outputs_23__0, outputs_22__15, 
                 outputs_22__14, outputs_22__13, outputs_22__12, outputs_22__11, 
                 outputs_22__10, outputs_22__9, outputs_22__8, outputs_22__7, 
                 outputs_22__6, outputs_22__5, outputs_22__4, outputs_22__3, 
                 outputs_22__2, outputs_22__1, outputs_22__0, outputs_21__15, 
                 outputs_21__14, outputs_21__13, outputs_21__12, outputs_21__11, 
                 outputs_21__10, outputs_21__9, outputs_21__8, outputs_21__7, 
                 outputs_21__6, outputs_21__5, outputs_21__4, outputs_21__3, 
                 outputs_21__2, outputs_21__1, outputs_21__0, outputs_20__15, 
                 outputs_20__14, outputs_20__13, outputs_20__12, outputs_20__11, 
                 outputs_20__10, outputs_20__9, outputs_20__8, outputs_20__7, 
                 outputs_20__6, outputs_20__5, outputs_20__4, outputs_20__3, 
                 outputs_20__2, outputs_20__1, outputs_20__0, outputs_19__15, 
                 outputs_19__14, outputs_19__13, outputs_19__12, outputs_19__11, 
                 outputs_19__10, outputs_19__9, outputs_19__8, outputs_19__7, 
                 outputs_19__6, outputs_19__5, outputs_19__4, outputs_19__3, 
                 outputs_19__2, outputs_19__1, outputs_19__0, outputs_18__15, 
                 outputs_18__14, outputs_18__13, outputs_18__12, outputs_18__11, 
                 outputs_18__10, outputs_18__9, outputs_18__8, outputs_18__7, 
                 outputs_18__6, outputs_18__5, outputs_18__4, outputs_18__3, 
                 outputs_18__2, outputs_18__1, outputs_18__0, outputs_17__15, 
                 outputs_17__14, outputs_17__13, outputs_17__12, outputs_17__11, 
                 outputs_17__10, outputs_17__9, outputs_17__8, outputs_17__7, 
                 outputs_17__6, outputs_17__5, outputs_17__4, outputs_17__3, 
                 outputs_17__2, outputs_17__1, outputs_17__0, outputs_16__15, 
                 outputs_16__14, outputs_16__13, outputs_16__12, outputs_16__11, 
                 outputs_16__10, outputs_16__9, outputs_16__8, outputs_16__7, 
                 outputs_16__6, outputs_16__5, outputs_16__4, outputs_16__3, 
                 outputs_16__2, outputs_16__1, outputs_16__0, outputs_15__15, 
                 outputs_15__14, outputs_15__13, outputs_15__12, outputs_15__11, 
                 outputs_15__10, outputs_15__9, outputs_15__8, outputs_15__7, 
                 outputs_15__6, outputs_15__5, outputs_15__4, outputs_15__3, 
                 outputs_15__2, outputs_15__1, outputs_15__0, outputs_14__15, 
                 outputs_14__14, outputs_14__13, outputs_14__12, outputs_14__11, 
                 outputs_14__10, outputs_14__9, outputs_14__8, outputs_14__7, 
                 outputs_14__6, outputs_14__5, outputs_14__4, outputs_14__3, 
                 outputs_14__2, outputs_14__1, outputs_14__0, outputs_13__15, 
                 outputs_13__14, outputs_13__13, outputs_13__12, outputs_13__11, 
                 outputs_13__10, outputs_13__9, outputs_13__8, outputs_13__7, 
                 outputs_13__6, outputs_13__5, outputs_13__4, outputs_13__3, 
                 outputs_13__2, outputs_13__1, outputs_13__0, outputs_12__15, 
                 outputs_12__14, outputs_12__13, outputs_12__12, outputs_12__11, 
                 outputs_12__10, outputs_12__9, outputs_12__8, outputs_12__7, 
                 outputs_12__6, outputs_12__5, outputs_12__4, outputs_12__3, 
                 outputs_12__2, outputs_12__1, outputs_12__0, outputs_11__15, 
                 outputs_11__14, outputs_11__13, outputs_11__12, outputs_11__11, 
                 outputs_11__10, outputs_11__9, outputs_11__8, outputs_11__7, 
                 outputs_11__6, outputs_11__5, outputs_11__4, outputs_11__3, 
                 outputs_11__2, outputs_11__1, outputs_11__0, outputs_10__15, 
                 outputs_10__14, outputs_10__13, outputs_10__12, outputs_10__11, 
                 outputs_10__10, outputs_10__9, outputs_10__8, outputs_10__7, 
                 outputs_10__6, outputs_10__5, outputs_10__4, outputs_10__3, 
                 outputs_10__2, outputs_10__1, outputs_10__0, outputs_9__15, 
                 outputs_9__14, outputs_9__13, outputs_9__12, outputs_9__11, 
                 outputs_9__10, outputs_9__9, outputs_9__8, outputs_9__7, 
                 outputs_9__6, outputs_9__5, outputs_9__4, outputs_9__3, 
                 outputs_9__2, outputs_9__1, outputs_9__0, outputs_8__15, 
                 outputs_8__14, outputs_8__13, outputs_8__12, outputs_8__11, 
                 outputs_8__10, outputs_8__9, outputs_8__8, outputs_8__7, 
                 outputs_8__6, outputs_8__5, outputs_8__4, outputs_8__3, 
                 outputs_8__2, outputs_8__1, outputs_8__0, outputs_7__15, 
                 outputs_7__14, outputs_7__13, outputs_7__12, outputs_7__11, 
                 outputs_7__10, outputs_7__9, outputs_7__8, outputs_7__7, 
                 outputs_7__6, outputs_7__5, outputs_7__4, outputs_7__3, 
                 outputs_7__2, outputs_7__1, outputs_7__0, outputs_6__15, 
                 outputs_6__14, outputs_6__13, outputs_6__12, outputs_6__11, 
                 outputs_6__10, outputs_6__9, outputs_6__8, outputs_6__7, 
                 outputs_6__6, outputs_6__5, outputs_6__4, outputs_6__3, 
                 outputs_6__2, outputs_6__1, outputs_6__0, outputs_5__15, 
                 outputs_5__14, outputs_5__13, outputs_5__12, outputs_5__11, 
                 outputs_5__10, outputs_5__9, outputs_5__8, outputs_5__7, 
                 outputs_5__6, outputs_5__5, outputs_5__4, outputs_5__3, 
                 outputs_5__2, outputs_5__1, outputs_5__0, outputs_4__15, 
                 outputs_4__14, outputs_4__13, outputs_4__12, outputs_4__11, 
                 outputs_4__10, outputs_4__9, outputs_4__8, outputs_4__7, 
                 outputs_4__6, outputs_4__5, outputs_4__4, outputs_4__3, 
                 outputs_4__2, outputs_4__1, outputs_4__0, outputs_3__15, 
                 outputs_3__14, outputs_3__13, outputs_3__12, outputs_3__11, 
                 outputs_3__10, outputs_3__9, outputs_3__8, outputs_3__7, 
                 outputs_3__6, outputs_3__5, outputs_3__4, outputs_3__3, 
                 outputs_3__2, outputs_3__1, outputs_3__0, outputs_2__15, 
                 outputs_2__14, outputs_2__13, outputs_2__12, outputs_2__11, 
                 outputs_2__10, outputs_2__9, outputs_2__8, outputs_2__7, 
                 outputs_2__6, outputs_2__5, outputs_2__4, outputs_2__3, 
                 outputs_2__2, outputs_2__1, outputs_2__0, outputs_1__15, 
                 outputs_1__14, outputs_1__13, outputs_1__12, outputs_1__11, 
                 outputs_1__10, outputs_1__9, outputs_1__8, outputs_1__7, 
                 outputs_1__6, outputs_1__5, outputs_1__4, outputs_1__3, 
                 outputs_1__2, outputs_1__1, outputs_1__0, outputs_0__15, 
                 outputs_0__14, outputs_0__13, outputs_0__12, outputs_0__11, 
                 outputs_0__10, outputs_0__9, outputs_0__8, outputs_0__7, 
                 outputs_0__6, outputs_0__5, outputs_0__4, outputs_0__3, 
                 outputs_0__2, outputs_0__1, outputs_0__0, clk, start, rst, done, 
                 working ) ;

    input filter_24__7 ;
    input filter_24__6 ;
    input filter_24__5 ;
    input filter_24__4 ;
    input filter_24__3 ;
    input filter_24__2 ;
    input filter_24__1 ;
    input filter_24__0 ;
    input filter_23__7 ;
    input filter_23__6 ;
    input filter_23__5 ;
    input filter_23__4 ;
    input filter_23__3 ;
    input filter_23__2 ;
    input filter_23__1 ;
    input filter_23__0 ;
    input filter_22__7 ;
    input filter_22__6 ;
    input filter_22__5 ;
    input filter_22__4 ;
    input filter_22__3 ;
    input filter_22__2 ;
    input filter_22__1 ;
    input filter_22__0 ;
    input filter_21__7 ;
    input filter_21__6 ;
    input filter_21__5 ;
    input filter_21__4 ;
    input filter_21__3 ;
    input filter_21__2 ;
    input filter_21__1 ;
    input filter_21__0 ;
    input filter_20__7 ;
    input filter_20__6 ;
    input filter_20__5 ;
    input filter_20__4 ;
    input filter_20__3 ;
    input filter_20__2 ;
    input filter_20__1 ;
    input filter_20__0 ;
    input filter_19__7 ;
    input filter_19__6 ;
    input filter_19__5 ;
    input filter_19__4 ;
    input filter_19__3 ;
    input filter_19__2 ;
    input filter_19__1 ;
    input filter_19__0 ;
    input filter_18__7 ;
    input filter_18__6 ;
    input filter_18__5 ;
    input filter_18__4 ;
    input filter_18__3 ;
    input filter_18__2 ;
    input filter_18__1 ;
    input filter_18__0 ;
    input filter_17__7 ;
    input filter_17__6 ;
    input filter_17__5 ;
    input filter_17__4 ;
    input filter_17__3 ;
    input filter_17__2 ;
    input filter_17__1 ;
    input filter_17__0 ;
    input filter_16__7 ;
    input filter_16__6 ;
    input filter_16__5 ;
    input filter_16__4 ;
    input filter_16__3 ;
    input filter_16__2 ;
    input filter_16__1 ;
    input filter_16__0 ;
    input filter_15__7 ;
    input filter_15__6 ;
    input filter_15__5 ;
    input filter_15__4 ;
    input filter_15__3 ;
    input filter_15__2 ;
    input filter_15__1 ;
    input filter_15__0 ;
    input filter_14__7 ;
    input filter_14__6 ;
    input filter_14__5 ;
    input filter_14__4 ;
    input filter_14__3 ;
    input filter_14__2 ;
    input filter_14__1 ;
    input filter_14__0 ;
    input filter_13__7 ;
    input filter_13__6 ;
    input filter_13__5 ;
    input filter_13__4 ;
    input filter_13__3 ;
    input filter_13__2 ;
    input filter_13__1 ;
    input filter_13__0 ;
    input filter_12__7 ;
    input filter_12__6 ;
    input filter_12__5 ;
    input filter_12__4 ;
    input filter_12__3 ;
    input filter_12__2 ;
    input filter_12__1 ;
    input filter_12__0 ;
    input filter_11__7 ;
    input filter_11__6 ;
    input filter_11__5 ;
    input filter_11__4 ;
    input filter_11__3 ;
    input filter_11__2 ;
    input filter_11__1 ;
    input filter_11__0 ;
    input filter_10__7 ;
    input filter_10__6 ;
    input filter_10__5 ;
    input filter_10__4 ;
    input filter_10__3 ;
    input filter_10__2 ;
    input filter_10__1 ;
    input filter_10__0 ;
    input filter_9__7 ;
    input filter_9__6 ;
    input filter_9__5 ;
    input filter_9__4 ;
    input filter_9__3 ;
    input filter_9__2 ;
    input filter_9__1 ;
    input filter_9__0 ;
    input filter_8__7 ;
    input filter_8__6 ;
    input filter_8__5 ;
    input filter_8__4 ;
    input filter_8__3 ;
    input filter_8__2 ;
    input filter_8__1 ;
    input filter_8__0 ;
    input filter_7__7 ;
    input filter_7__6 ;
    input filter_7__5 ;
    input filter_7__4 ;
    input filter_7__3 ;
    input filter_7__2 ;
    input filter_7__1 ;
    input filter_7__0 ;
    input filter_6__7 ;
    input filter_6__6 ;
    input filter_6__5 ;
    input filter_6__4 ;
    input filter_6__3 ;
    input filter_6__2 ;
    input filter_6__1 ;
    input filter_6__0 ;
    input filter_5__7 ;
    input filter_5__6 ;
    input filter_5__5 ;
    input filter_5__4 ;
    input filter_5__3 ;
    input filter_5__2 ;
    input filter_5__1 ;
    input filter_5__0 ;
    input filter_4__7 ;
    input filter_4__6 ;
    input filter_4__5 ;
    input filter_4__4 ;
    input filter_4__3 ;
    input filter_4__2 ;
    input filter_4__1 ;
    input filter_4__0 ;
    input filter_3__7 ;
    input filter_3__6 ;
    input filter_3__5 ;
    input filter_3__4 ;
    input filter_3__3 ;
    input filter_3__2 ;
    input filter_3__1 ;
    input filter_3__0 ;
    input filter_2__7 ;
    input filter_2__6 ;
    input filter_2__5 ;
    input filter_2__4 ;
    input filter_2__3 ;
    input filter_2__2 ;
    input filter_2__1 ;
    input filter_2__0 ;
    input filter_1__7 ;
    input filter_1__6 ;
    input filter_1__5 ;
    input filter_1__4 ;
    input filter_1__3 ;
    input filter_1__2 ;
    input filter_1__1 ;
    input filter_1__0 ;
    input filter_0__7 ;
    input filter_0__6 ;
    input filter_0__5 ;
    input filter_0__4 ;
    input filter_0__3 ;
    input filter_0__2 ;
    input filter_0__1 ;
    input filter_0__0 ;
    input window_24__15 ;
    input window_24__14 ;
    input window_24__13 ;
    input window_24__12 ;
    input window_24__11 ;
    input window_24__10 ;
    input window_24__9 ;
    input window_24__8 ;
    input window_24__7 ;
    input window_24__6 ;
    input window_24__5 ;
    input window_24__4 ;
    input window_24__3 ;
    input window_24__2 ;
    input window_24__1 ;
    input window_24__0 ;
    input window_23__15 ;
    input window_23__14 ;
    input window_23__13 ;
    input window_23__12 ;
    input window_23__11 ;
    input window_23__10 ;
    input window_23__9 ;
    input window_23__8 ;
    input window_23__7 ;
    input window_23__6 ;
    input window_23__5 ;
    input window_23__4 ;
    input window_23__3 ;
    input window_23__2 ;
    input window_23__1 ;
    input window_23__0 ;
    input window_22__15 ;
    input window_22__14 ;
    input window_22__13 ;
    input window_22__12 ;
    input window_22__11 ;
    input window_22__10 ;
    input window_22__9 ;
    input window_22__8 ;
    input window_22__7 ;
    input window_22__6 ;
    input window_22__5 ;
    input window_22__4 ;
    input window_22__3 ;
    input window_22__2 ;
    input window_22__1 ;
    input window_22__0 ;
    input window_21__15 ;
    input window_21__14 ;
    input window_21__13 ;
    input window_21__12 ;
    input window_21__11 ;
    input window_21__10 ;
    input window_21__9 ;
    input window_21__8 ;
    input window_21__7 ;
    input window_21__6 ;
    input window_21__5 ;
    input window_21__4 ;
    input window_21__3 ;
    input window_21__2 ;
    input window_21__1 ;
    input window_21__0 ;
    input window_20__15 ;
    input window_20__14 ;
    input window_20__13 ;
    input window_20__12 ;
    input window_20__11 ;
    input window_20__10 ;
    input window_20__9 ;
    input window_20__8 ;
    input window_20__7 ;
    input window_20__6 ;
    input window_20__5 ;
    input window_20__4 ;
    input window_20__3 ;
    input window_20__2 ;
    input window_20__1 ;
    input window_20__0 ;
    input window_19__15 ;
    input window_19__14 ;
    input window_19__13 ;
    input window_19__12 ;
    input window_19__11 ;
    input window_19__10 ;
    input window_19__9 ;
    input window_19__8 ;
    input window_19__7 ;
    input window_19__6 ;
    input window_19__5 ;
    input window_19__4 ;
    input window_19__3 ;
    input window_19__2 ;
    input window_19__1 ;
    input window_19__0 ;
    input window_18__15 ;
    input window_18__14 ;
    input window_18__13 ;
    input window_18__12 ;
    input window_18__11 ;
    input window_18__10 ;
    input window_18__9 ;
    input window_18__8 ;
    input window_18__7 ;
    input window_18__6 ;
    input window_18__5 ;
    input window_18__4 ;
    input window_18__3 ;
    input window_18__2 ;
    input window_18__1 ;
    input window_18__0 ;
    input window_17__15 ;
    input window_17__14 ;
    input window_17__13 ;
    input window_17__12 ;
    input window_17__11 ;
    input window_17__10 ;
    input window_17__9 ;
    input window_17__8 ;
    input window_17__7 ;
    input window_17__6 ;
    input window_17__5 ;
    input window_17__4 ;
    input window_17__3 ;
    input window_17__2 ;
    input window_17__1 ;
    input window_17__0 ;
    input window_16__15 ;
    input window_16__14 ;
    input window_16__13 ;
    input window_16__12 ;
    input window_16__11 ;
    input window_16__10 ;
    input window_16__9 ;
    input window_16__8 ;
    input window_16__7 ;
    input window_16__6 ;
    input window_16__5 ;
    input window_16__4 ;
    input window_16__3 ;
    input window_16__2 ;
    input window_16__1 ;
    input window_16__0 ;
    input window_15__15 ;
    input window_15__14 ;
    input window_15__13 ;
    input window_15__12 ;
    input window_15__11 ;
    input window_15__10 ;
    input window_15__9 ;
    input window_15__8 ;
    input window_15__7 ;
    input window_15__6 ;
    input window_15__5 ;
    input window_15__4 ;
    input window_15__3 ;
    input window_15__2 ;
    input window_15__1 ;
    input window_15__0 ;
    input window_14__15 ;
    input window_14__14 ;
    input window_14__13 ;
    input window_14__12 ;
    input window_14__11 ;
    input window_14__10 ;
    input window_14__9 ;
    input window_14__8 ;
    input window_14__7 ;
    input window_14__6 ;
    input window_14__5 ;
    input window_14__4 ;
    input window_14__3 ;
    input window_14__2 ;
    input window_14__1 ;
    input window_14__0 ;
    input window_13__15 ;
    input window_13__14 ;
    input window_13__13 ;
    input window_13__12 ;
    input window_13__11 ;
    input window_13__10 ;
    input window_13__9 ;
    input window_13__8 ;
    input window_13__7 ;
    input window_13__6 ;
    input window_13__5 ;
    input window_13__4 ;
    input window_13__3 ;
    input window_13__2 ;
    input window_13__1 ;
    input window_13__0 ;
    input window_12__15 ;
    input window_12__14 ;
    input window_12__13 ;
    input window_12__12 ;
    input window_12__11 ;
    input window_12__10 ;
    input window_12__9 ;
    input window_12__8 ;
    input window_12__7 ;
    input window_12__6 ;
    input window_12__5 ;
    input window_12__4 ;
    input window_12__3 ;
    input window_12__2 ;
    input window_12__1 ;
    input window_12__0 ;
    input window_11__15 ;
    input window_11__14 ;
    input window_11__13 ;
    input window_11__12 ;
    input window_11__11 ;
    input window_11__10 ;
    input window_11__9 ;
    input window_11__8 ;
    input window_11__7 ;
    input window_11__6 ;
    input window_11__5 ;
    input window_11__4 ;
    input window_11__3 ;
    input window_11__2 ;
    input window_11__1 ;
    input window_11__0 ;
    input window_10__15 ;
    input window_10__14 ;
    input window_10__13 ;
    input window_10__12 ;
    input window_10__11 ;
    input window_10__10 ;
    input window_10__9 ;
    input window_10__8 ;
    input window_10__7 ;
    input window_10__6 ;
    input window_10__5 ;
    input window_10__4 ;
    input window_10__3 ;
    input window_10__2 ;
    input window_10__1 ;
    input window_10__0 ;
    input window_9__15 ;
    input window_9__14 ;
    input window_9__13 ;
    input window_9__12 ;
    input window_9__11 ;
    input window_9__10 ;
    input window_9__9 ;
    input window_9__8 ;
    input window_9__7 ;
    input window_9__6 ;
    input window_9__5 ;
    input window_9__4 ;
    input window_9__3 ;
    input window_9__2 ;
    input window_9__1 ;
    input window_9__0 ;
    input window_8__15 ;
    input window_8__14 ;
    input window_8__13 ;
    input window_8__12 ;
    input window_8__11 ;
    input window_8__10 ;
    input window_8__9 ;
    input window_8__8 ;
    input window_8__7 ;
    input window_8__6 ;
    input window_8__5 ;
    input window_8__4 ;
    input window_8__3 ;
    input window_8__2 ;
    input window_8__1 ;
    input window_8__0 ;
    input window_7__15 ;
    input window_7__14 ;
    input window_7__13 ;
    input window_7__12 ;
    input window_7__11 ;
    input window_7__10 ;
    input window_7__9 ;
    input window_7__8 ;
    input window_7__7 ;
    input window_7__6 ;
    input window_7__5 ;
    input window_7__4 ;
    input window_7__3 ;
    input window_7__2 ;
    input window_7__1 ;
    input window_7__0 ;
    input window_6__15 ;
    input window_6__14 ;
    input window_6__13 ;
    input window_6__12 ;
    input window_6__11 ;
    input window_6__10 ;
    input window_6__9 ;
    input window_6__8 ;
    input window_6__7 ;
    input window_6__6 ;
    input window_6__5 ;
    input window_6__4 ;
    input window_6__3 ;
    input window_6__2 ;
    input window_6__1 ;
    input window_6__0 ;
    input window_5__15 ;
    input window_5__14 ;
    input window_5__13 ;
    input window_5__12 ;
    input window_5__11 ;
    input window_5__10 ;
    input window_5__9 ;
    input window_5__8 ;
    input window_5__7 ;
    input window_5__6 ;
    input window_5__5 ;
    input window_5__4 ;
    input window_5__3 ;
    input window_5__2 ;
    input window_5__1 ;
    input window_5__0 ;
    input window_4__15 ;
    input window_4__14 ;
    input window_4__13 ;
    input window_4__12 ;
    input window_4__11 ;
    input window_4__10 ;
    input window_4__9 ;
    input window_4__8 ;
    input window_4__7 ;
    input window_4__6 ;
    input window_4__5 ;
    input window_4__4 ;
    input window_4__3 ;
    input window_4__2 ;
    input window_4__1 ;
    input window_4__0 ;
    input window_3__15 ;
    input window_3__14 ;
    input window_3__13 ;
    input window_3__12 ;
    input window_3__11 ;
    input window_3__10 ;
    input window_3__9 ;
    input window_3__8 ;
    input window_3__7 ;
    input window_3__6 ;
    input window_3__5 ;
    input window_3__4 ;
    input window_3__3 ;
    input window_3__2 ;
    input window_3__1 ;
    input window_3__0 ;
    input window_2__15 ;
    input window_2__14 ;
    input window_2__13 ;
    input window_2__12 ;
    input window_2__11 ;
    input window_2__10 ;
    input window_2__9 ;
    input window_2__8 ;
    input window_2__7 ;
    input window_2__6 ;
    input window_2__5 ;
    input window_2__4 ;
    input window_2__3 ;
    input window_2__2 ;
    input window_2__1 ;
    input window_2__0 ;
    input window_1__15 ;
    input window_1__14 ;
    input window_1__13 ;
    input window_1__12 ;
    input window_1__11 ;
    input window_1__10 ;
    input window_1__9 ;
    input window_1__8 ;
    input window_1__7 ;
    input window_1__6 ;
    input window_1__5 ;
    input window_1__4 ;
    input window_1__3 ;
    input window_1__2 ;
    input window_1__1 ;
    input window_1__0 ;
    input window_0__15 ;
    input window_0__14 ;
    input window_0__13 ;
    input window_0__12 ;
    input window_0__11 ;
    input window_0__10 ;
    input window_0__9 ;
    input window_0__8 ;
    input window_0__7 ;
    input window_0__6 ;
    input window_0__5 ;
    input window_0__4 ;
    input window_0__3 ;
    input window_0__2 ;
    input window_0__1 ;
    input window_0__0 ;
    inout outputs_24__15 ;
    inout outputs_24__14 ;
    inout outputs_24__13 ;
    inout outputs_24__12 ;
    inout outputs_24__11 ;
    inout outputs_24__10 ;
    inout outputs_24__9 ;
    inout outputs_24__8 ;
    inout outputs_24__7 ;
    inout outputs_24__6 ;
    inout outputs_24__5 ;
    inout outputs_24__4 ;
    inout outputs_24__3 ;
    inout outputs_24__2 ;
    inout outputs_24__1 ;
    inout outputs_24__0 ;
    inout outputs_23__15 ;
    inout outputs_23__14 ;
    inout outputs_23__13 ;
    inout outputs_23__12 ;
    inout outputs_23__11 ;
    inout outputs_23__10 ;
    inout outputs_23__9 ;
    inout outputs_23__8 ;
    inout outputs_23__7 ;
    inout outputs_23__6 ;
    inout outputs_23__5 ;
    inout outputs_23__4 ;
    inout outputs_23__3 ;
    inout outputs_23__2 ;
    inout outputs_23__1 ;
    inout outputs_23__0 ;
    inout outputs_22__15 ;
    inout outputs_22__14 ;
    inout outputs_22__13 ;
    inout outputs_22__12 ;
    inout outputs_22__11 ;
    inout outputs_22__10 ;
    inout outputs_22__9 ;
    inout outputs_22__8 ;
    inout outputs_22__7 ;
    inout outputs_22__6 ;
    inout outputs_22__5 ;
    inout outputs_22__4 ;
    inout outputs_22__3 ;
    inout outputs_22__2 ;
    inout outputs_22__1 ;
    inout outputs_22__0 ;
    inout outputs_21__15 ;
    inout outputs_21__14 ;
    inout outputs_21__13 ;
    inout outputs_21__12 ;
    inout outputs_21__11 ;
    inout outputs_21__10 ;
    inout outputs_21__9 ;
    inout outputs_21__8 ;
    inout outputs_21__7 ;
    inout outputs_21__6 ;
    inout outputs_21__5 ;
    inout outputs_21__4 ;
    inout outputs_21__3 ;
    inout outputs_21__2 ;
    inout outputs_21__1 ;
    inout outputs_21__0 ;
    inout outputs_20__15 ;
    inout outputs_20__14 ;
    inout outputs_20__13 ;
    inout outputs_20__12 ;
    inout outputs_20__11 ;
    inout outputs_20__10 ;
    inout outputs_20__9 ;
    inout outputs_20__8 ;
    inout outputs_20__7 ;
    inout outputs_20__6 ;
    inout outputs_20__5 ;
    inout outputs_20__4 ;
    inout outputs_20__3 ;
    inout outputs_20__2 ;
    inout outputs_20__1 ;
    inout outputs_20__0 ;
    inout outputs_19__15 ;
    inout outputs_19__14 ;
    inout outputs_19__13 ;
    inout outputs_19__12 ;
    inout outputs_19__11 ;
    inout outputs_19__10 ;
    inout outputs_19__9 ;
    inout outputs_19__8 ;
    inout outputs_19__7 ;
    inout outputs_19__6 ;
    inout outputs_19__5 ;
    inout outputs_19__4 ;
    inout outputs_19__3 ;
    inout outputs_19__2 ;
    inout outputs_19__1 ;
    inout outputs_19__0 ;
    inout outputs_18__15 ;
    inout outputs_18__14 ;
    inout outputs_18__13 ;
    inout outputs_18__12 ;
    inout outputs_18__11 ;
    inout outputs_18__10 ;
    inout outputs_18__9 ;
    inout outputs_18__8 ;
    inout outputs_18__7 ;
    inout outputs_18__6 ;
    inout outputs_18__5 ;
    inout outputs_18__4 ;
    inout outputs_18__3 ;
    inout outputs_18__2 ;
    inout outputs_18__1 ;
    inout outputs_18__0 ;
    inout outputs_17__15 ;
    inout outputs_17__14 ;
    inout outputs_17__13 ;
    inout outputs_17__12 ;
    inout outputs_17__11 ;
    inout outputs_17__10 ;
    inout outputs_17__9 ;
    inout outputs_17__8 ;
    inout outputs_17__7 ;
    inout outputs_17__6 ;
    inout outputs_17__5 ;
    inout outputs_17__4 ;
    inout outputs_17__3 ;
    inout outputs_17__2 ;
    inout outputs_17__1 ;
    inout outputs_17__0 ;
    inout outputs_16__15 ;
    inout outputs_16__14 ;
    inout outputs_16__13 ;
    inout outputs_16__12 ;
    inout outputs_16__11 ;
    inout outputs_16__10 ;
    inout outputs_16__9 ;
    inout outputs_16__8 ;
    inout outputs_16__7 ;
    inout outputs_16__6 ;
    inout outputs_16__5 ;
    inout outputs_16__4 ;
    inout outputs_16__3 ;
    inout outputs_16__2 ;
    inout outputs_16__1 ;
    inout outputs_16__0 ;
    inout outputs_15__15 ;
    inout outputs_15__14 ;
    inout outputs_15__13 ;
    inout outputs_15__12 ;
    inout outputs_15__11 ;
    inout outputs_15__10 ;
    inout outputs_15__9 ;
    inout outputs_15__8 ;
    inout outputs_15__7 ;
    inout outputs_15__6 ;
    inout outputs_15__5 ;
    inout outputs_15__4 ;
    inout outputs_15__3 ;
    inout outputs_15__2 ;
    inout outputs_15__1 ;
    inout outputs_15__0 ;
    inout outputs_14__15 ;
    inout outputs_14__14 ;
    inout outputs_14__13 ;
    inout outputs_14__12 ;
    inout outputs_14__11 ;
    inout outputs_14__10 ;
    inout outputs_14__9 ;
    inout outputs_14__8 ;
    inout outputs_14__7 ;
    inout outputs_14__6 ;
    inout outputs_14__5 ;
    inout outputs_14__4 ;
    inout outputs_14__3 ;
    inout outputs_14__2 ;
    inout outputs_14__1 ;
    inout outputs_14__0 ;
    inout outputs_13__15 ;
    inout outputs_13__14 ;
    inout outputs_13__13 ;
    inout outputs_13__12 ;
    inout outputs_13__11 ;
    inout outputs_13__10 ;
    inout outputs_13__9 ;
    inout outputs_13__8 ;
    inout outputs_13__7 ;
    inout outputs_13__6 ;
    inout outputs_13__5 ;
    inout outputs_13__4 ;
    inout outputs_13__3 ;
    inout outputs_13__2 ;
    inout outputs_13__1 ;
    inout outputs_13__0 ;
    inout outputs_12__15 ;
    inout outputs_12__14 ;
    inout outputs_12__13 ;
    inout outputs_12__12 ;
    inout outputs_12__11 ;
    inout outputs_12__10 ;
    inout outputs_12__9 ;
    inout outputs_12__8 ;
    inout outputs_12__7 ;
    inout outputs_12__6 ;
    inout outputs_12__5 ;
    inout outputs_12__4 ;
    inout outputs_12__3 ;
    inout outputs_12__2 ;
    inout outputs_12__1 ;
    inout outputs_12__0 ;
    inout outputs_11__15 ;
    inout outputs_11__14 ;
    inout outputs_11__13 ;
    inout outputs_11__12 ;
    inout outputs_11__11 ;
    inout outputs_11__10 ;
    inout outputs_11__9 ;
    inout outputs_11__8 ;
    inout outputs_11__7 ;
    inout outputs_11__6 ;
    inout outputs_11__5 ;
    inout outputs_11__4 ;
    inout outputs_11__3 ;
    inout outputs_11__2 ;
    inout outputs_11__1 ;
    inout outputs_11__0 ;
    inout outputs_10__15 ;
    inout outputs_10__14 ;
    inout outputs_10__13 ;
    inout outputs_10__12 ;
    inout outputs_10__11 ;
    inout outputs_10__10 ;
    inout outputs_10__9 ;
    inout outputs_10__8 ;
    inout outputs_10__7 ;
    inout outputs_10__6 ;
    inout outputs_10__5 ;
    inout outputs_10__4 ;
    inout outputs_10__3 ;
    inout outputs_10__2 ;
    inout outputs_10__1 ;
    inout outputs_10__0 ;
    inout outputs_9__15 ;
    inout outputs_9__14 ;
    inout outputs_9__13 ;
    inout outputs_9__12 ;
    inout outputs_9__11 ;
    inout outputs_9__10 ;
    inout outputs_9__9 ;
    inout outputs_9__8 ;
    inout outputs_9__7 ;
    inout outputs_9__6 ;
    inout outputs_9__5 ;
    inout outputs_9__4 ;
    inout outputs_9__3 ;
    inout outputs_9__2 ;
    inout outputs_9__1 ;
    inout outputs_9__0 ;
    inout outputs_8__15 ;
    inout outputs_8__14 ;
    inout outputs_8__13 ;
    inout outputs_8__12 ;
    inout outputs_8__11 ;
    inout outputs_8__10 ;
    inout outputs_8__9 ;
    inout outputs_8__8 ;
    inout outputs_8__7 ;
    inout outputs_8__6 ;
    inout outputs_8__5 ;
    inout outputs_8__4 ;
    inout outputs_8__3 ;
    inout outputs_8__2 ;
    inout outputs_8__1 ;
    inout outputs_8__0 ;
    inout outputs_7__15 ;
    inout outputs_7__14 ;
    inout outputs_7__13 ;
    inout outputs_7__12 ;
    inout outputs_7__11 ;
    inout outputs_7__10 ;
    inout outputs_7__9 ;
    inout outputs_7__8 ;
    inout outputs_7__7 ;
    inout outputs_7__6 ;
    inout outputs_7__5 ;
    inout outputs_7__4 ;
    inout outputs_7__3 ;
    inout outputs_7__2 ;
    inout outputs_7__1 ;
    inout outputs_7__0 ;
    inout outputs_6__15 ;
    inout outputs_6__14 ;
    inout outputs_6__13 ;
    inout outputs_6__12 ;
    inout outputs_6__11 ;
    inout outputs_6__10 ;
    inout outputs_6__9 ;
    inout outputs_6__8 ;
    inout outputs_6__7 ;
    inout outputs_6__6 ;
    inout outputs_6__5 ;
    inout outputs_6__4 ;
    inout outputs_6__3 ;
    inout outputs_6__2 ;
    inout outputs_6__1 ;
    inout outputs_6__0 ;
    inout outputs_5__15 ;
    inout outputs_5__14 ;
    inout outputs_5__13 ;
    inout outputs_5__12 ;
    inout outputs_5__11 ;
    inout outputs_5__10 ;
    inout outputs_5__9 ;
    inout outputs_5__8 ;
    inout outputs_5__7 ;
    inout outputs_5__6 ;
    inout outputs_5__5 ;
    inout outputs_5__4 ;
    inout outputs_5__3 ;
    inout outputs_5__2 ;
    inout outputs_5__1 ;
    inout outputs_5__0 ;
    inout outputs_4__15 ;
    inout outputs_4__14 ;
    inout outputs_4__13 ;
    inout outputs_4__12 ;
    inout outputs_4__11 ;
    inout outputs_4__10 ;
    inout outputs_4__9 ;
    inout outputs_4__8 ;
    inout outputs_4__7 ;
    inout outputs_4__6 ;
    inout outputs_4__5 ;
    inout outputs_4__4 ;
    inout outputs_4__3 ;
    inout outputs_4__2 ;
    inout outputs_4__1 ;
    inout outputs_4__0 ;
    inout outputs_3__15 ;
    inout outputs_3__14 ;
    inout outputs_3__13 ;
    inout outputs_3__12 ;
    inout outputs_3__11 ;
    inout outputs_3__10 ;
    inout outputs_3__9 ;
    inout outputs_3__8 ;
    inout outputs_3__7 ;
    inout outputs_3__6 ;
    inout outputs_3__5 ;
    inout outputs_3__4 ;
    inout outputs_3__3 ;
    inout outputs_3__2 ;
    inout outputs_3__1 ;
    inout outputs_3__0 ;
    inout outputs_2__15 ;
    inout outputs_2__14 ;
    inout outputs_2__13 ;
    inout outputs_2__12 ;
    inout outputs_2__11 ;
    inout outputs_2__10 ;
    inout outputs_2__9 ;
    inout outputs_2__8 ;
    inout outputs_2__7 ;
    inout outputs_2__6 ;
    inout outputs_2__5 ;
    inout outputs_2__4 ;
    inout outputs_2__3 ;
    inout outputs_2__2 ;
    inout outputs_2__1 ;
    inout outputs_2__0 ;
    inout outputs_1__15 ;
    inout outputs_1__14 ;
    inout outputs_1__13 ;
    inout outputs_1__12 ;
    inout outputs_1__11 ;
    inout outputs_1__10 ;
    inout outputs_1__9 ;
    inout outputs_1__8 ;
    inout outputs_1__7 ;
    inout outputs_1__6 ;
    inout outputs_1__5 ;
    inout outputs_1__4 ;
    inout outputs_1__3 ;
    inout outputs_1__2 ;
    inout outputs_1__1 ;
    inout outputs_1__0 ;
    inout outputs_0__15 ;
    inout outputs_0__14 ;
    inout outputs_0__13 ;
    inout outputs_0__12 ;
    inout outputs_0__11 ;
    inout outputs_0__10 ;
    inout outputs_0__9 ;
    inout outputs_0__8 ;
    inout outputs_0__7 ;
    inout outputs_0__6 ;
    inout outputs_0__5 ;
    inout outputs_0__4 ;
    inout outputs_0__3 ;
    inout outputs_0__2 ;
    inout outputs_0__1 ;
    inout outputs_0__0 ;
    input clk ;
    input start ;
    input rst ;
    inout done ;
    inout working ;

    wire gen_24_cmp_pBs_30, gen_24_cmp_pBs_29, gen_24_cmp_pBs_28, 
         gen_24_cmp_pBs_27, gen_24_cmp_pBs_26, gen_24_cmp_pBs_25, 
         gen_24_cmp_pBs_24, gen_24_cmp_pBs_23, gen_24_cmp_pMux_30, 
         gen_24_cmp_pMux_29, gen_24_cmp_pMux_28, gen_24_cmp_pMux_27, 
         gen_24_cmp_pMux_26, gen_24_cmp_pMux_25, gen_24_cmp_pMux_24, 
         gen_24_cmp_pMux_23, gen_24_cmp_pMux_22, gen_24_cmp_pMux_21, 
         gen_24_cmp_pMux_20, gen_24_cmp_pMux_19, gen_24_cmp_pMux_18, 
         gen_24_cmp_pMux_17, gen_24_cmp_pMux_16, gen_24_cmp_pMux_15, 
         gen_24_cmp_pMux_14, gen_24_cmp_pMux_13, gen_24_cmp_pMux_12, 
         gen_24_cmp_pMux_11, gen_24_cmp_pMux_10, gen_24_cmp_pMux_9, 
         gen_24_cmp_pMux_8, gen_24_cmp_pMux_7, gen_24_cmp_pMux_6, 
         gen_24_cmp_pMux_5, gen_24_cmp_pMux_4, gen_24_cmp_pMux_3, 
         gen_24_cmp_pMux_2, gen_24_cmp_pMux_1, gen_24_cmp_pMux_0, 
         gen_24_cmp_pReg_30, gen_24_cmp_pReg_29, gen_24_cmp_pReg_28, 
         gen_24_cmp_pReg_27, gen_24_cmp_pReg_26, gen_24_cmp_pReg_25, 
         gen_24_cmp_pReg_24, gen_24_cmp_pReg_23, gen_24_cmp_pReg_22, 
         gen_24_cmp_pReg_21, gen_24_cmp_pReg_20, gen_24_cmp_pReg_19, 
         gen_24_cmp_pReg_18, gen_24_cmp_pReg_17, gen_24_cmp_pReg_16, 
         gen_24_cmp_pReg_15, gen_24_cmp_pReg_14, gen_24_cmp_pReg_13, 
         gen_24_cmp_pReg_12, gen_24_cmp_pReg_11, gen_24_cmp_pReg_10, 
         gen_24_cmp_pReg_9, gen_24_cmp_pReg_8, gen_24_cmp_pReg_7, 
         gen_24_cmp_pReg_6, gen_24_cmp_pReg_5, gen_24_cmp_pReg_4, 
         gen_24_cmp_pReg_3, gen_24_cmp_pReg_2, gen_24_cmp_pReg_1, 
         gen_24_cmp_pReg_0, gen_24_cmp_BSCmp_op2_0, gen_24_cmp_BSCmp_carryIn, 
         gen_23_cmp_pBs_30, gen_23_cmp_pBs_29, gen_23_cmp_pBs_28, 
         gen_23_cmp_pBs_27, gen_23_cmp_pBs_26, gen_23_cmp_pBs_25, 
         gen_23_cmp_pBs_24, gen_23_cmp_pBs_23, gen_23_cmp_pMux_30, 
         gen_23_cmp_pMux_29, gen_23_cmp_pMux_28, gen_23_cmp_pMux_27, 
         gen_23_cmp_pMux_26, gen_23_cmp_pMux_25, gen_23_cmp_pMux_24, 
         gen_23_cmp_pMux_23, gen_23_cmp_pMux_22, gen_23_cmp_pMux_21, 
         gen_23_cmp_pMux_20, gen_23_cmp_pMux_19, gen_23_cmp_pMux_18, 
         gen_23_cmp_pMux_17, gen_23_cmp_pMux_16, gen_23_cmp_pMux_15, 
         gen_23_cmp_pMux_14, gen_23_cmp_pMux_13, gen_23_cmp_pMux_12, 
         gen_23_cmp_pMux_11, gen_23_cmp_pMux_10, gen_23_cmp_pMux_9, 
         gen_23_cmp_pMux_8, gen_23_cmp_pMux_7, gen_23_cmp_pMux_6, 
         gen_23_cmp_pMux_5, gen_23_cmp_pMux_4, gen_23_cmp_pMux_3, 
         gen_23_cmp_pMux_2, gen_23_cmp_pMux_1, gen_23_cmp_pMux_0, 
         gen_23_cmp_pReg_30, gen_23_cmp_pReg_29, gen_23_cmp_pReg_28, 
         gen_23_cmp_pReg_27, gen_23_cmp_pReg_26, gen_23_cmp_pReg_25, 
         gen_23_cmp_pReg_24, gen_23_cmp_pReg_23, gen_23_cmp_pReg_22, 
         gen_23_cmp_pReg_21, gen_23_cmp_pReg_20, gen_23_cmp_pReg_19, 
         gen_23_cmp_pReg_18, gen_23_cmp_pReg_17, gen_23_cmp_pReg_16, 
         gen_23_cmp_pReg_15, gen_23_cmp_pReg_14, gen_23_cmp_pReg_13, 
         gen_23_cmp_pReg_12, gen_23_cmp_pReg_11, gen_23_cmp_pReg_10, 
         gen_23_cmp_pReg_9, gen_23_cmp_pReg_8, gen_23_cmp_pReg_7, 
         gen_23_cmp_pReg_6, gen_23_cmp_pReg_5, gen_23_cmp_pReg_4, 
         gen_23_cmp_pReg_3, gen_23_cmp_pReg_2, gen_23_cmp_pReg_1, 
         gen_23_cmp_pReg_0, gen_23_cmp_BSCmp_op2_0, gen_23_cmp_BSCmp_carryIn, 
         gen_22_cmp_pBs_30, gen_22_cmp_pBs_29, gen_22_cmp_pBs_28, 
         gen_22_cmp_pBs_27, gen_22_cmp_pBs_26, gen_22_cmp_pBs_25, 
         gen_22_cmp_pBs_24, gen_22_cmp_pBs_23, gen_22_cmp_pMux_30, 
         gen_22_cmp_pMux_29, gen_22_cmp_pMux_28, gen_22_cmp_pMux_27, 
         gen_22_cmp_pMux_26, gen_22_cmp_pMux_25, gen_22_cmp_pMux_24, 
         gen_22_cmp_pMux_23, gen_22_cmp_pMux_22, gen_22_cmp_pMux_21, 
         gen_22_cmp_pMux_20, gen_22_cmp_pMux_19, gen_22_cmp_pMux_18, 
         gen_22_cmp_pMux_17, gen_22_cmp_pMux_16, gen_22_cmp_pMux_15, 
         gen_22_cmp_pMux_14, gen_22_cmp_pMux_13, gen_22_cmp_pMux_12, 
         gen_22_cmp_pMux_11, gen_22_cmp_pMux_10, gen_22_cmp_pMux_9, 
         gen_22_cmp_pMux_8, gen_22_cmp_pMux_7, gen_22_cmp_pMux_6, 
         gen_22_cmp_pMux_5, gen_22_cmp_pMux_4, gen_22_cmp_pMux_3, 
         gen_22_cmp_pMux_2, gen_22_cmp_pMux_1, gen_22_cmp_pMux_0, 
         gen_22_cmp_pReg_30, gen_22_cmp_pReg_29, gen_22_cmp_pReg_28, 
         gen_22_cmp_pReg_27, gen_22_cmp_pReg_26, gen_22_cmp_pReg_25, 
         gen_22_cmp_pReg_24, gen_22_cmp_pReg_23, gen_22_cmp_pReg_22, 
         gen_22_cmp_pReg_21, gen_22_cmp_pReg_20, gen_22_cmp_pReg_19, 
         gen_22_cmp_pReg_18, gen_22_cmp_pReg_17, gen_22_cmp_pReg_16, 
         gen_22_cmp_pReg_15, gen_22_cmp_pReg_14, gen_22_cmp_pReg_13, 
         gen_22_cmp_pReg_12, gen_22_cmp_pReg_11, gen_22_cmp_pReg_10, 
         gen_22_cmp_pReg_9, gen_22_cmp_pReg_8, gen_22_cmp_pReg_7, 
         gen_22_cmp_pReg_6, gen_22_cmp_pReg_5, gen_22_cmp_pReg_4, 
         gen_22_cmp_pReg_3, gen_22_cmp_pReg_2, gen_22_cmp_pReg_1, 
         gen_22_cmp_pReg_0, gen_22_cmp_BSCmp_op2_0, gen_22_cmp_BSCmp_carryIn, 
         gen_21_cmp_pBs_30, gen_21_cmp_pBs_29, gen_21_cmp_pBs_28, 
         gen_21_cmp_pBs_27, gen_21_cmp_pBs_26, gen_21_cmp_pBs_25, 
         gen_21_cmp_pBs_24, gen_21_cmp_pBs_23, gen_21_cmp_pMux_30, 
         gen_21_cmp_pMux_29, gen_21_cmp_pMux_28, gen_21_cmp_pMux_27, 
         gen_21_cmp_pMux_26, gen_21_cmp_pMux_25, gen_21_cmp_pMux_24, 
         gen_21_cmp_pMux_23, gen_21_cmp_pMux_22, gen_21_cmp_pMux_21, 
         gen_21_cmp_pMux_20, gen_21_cmp_pMux_19, gen_21_cmp_pMux_18, 
         gen_21_cmp_pMux_17, gen_21_cmp_pMux_16, gen_21_cmp_pMux_15, 
         gen_21_cmp_pMux_14, gen_21_cmp_pMux_13, gen_21_cmp_pMux_12, 
         gen_21_cmp_pMux_11, gen_21_cmp_pMux_10, gen_21_cmp_pMux_9, 
         gen_21_cmp_pMux_8, gen_21_cmp_pMux_7, gen_21_cmp_pMux_6, 
         gen_21_cmp_pMux_5, gen_21_cmp_pMux_4, gen_21_cmp_pMux_3, 
         gen_21_cmp_pMux_2, gen_21_cmp_pMux_1, gen_21_cmp_pMux_0, 
         gen_21_cmp_pReg_30, gen_21_cmp_pReg_29, gen_21_cmp_pReg_28, 
         gen_21_cmp_pReg_27, gen_21_cmp_pReg_26, gen_21_cmp_pReg_25, 
         gen_21_cmp_pReg_24, gen_21_cmp_pReg_23, gen_21_cmp_pReg_22, 
         gen_21_cmp_pReg_21, gen_21_cmp_pReg_20, gen_21_cmp_pReg_19, 
         gen_21_cmp_pReg_18, gen_21_cmp_pReg_17, gen_21_cmp_pReg_16, 
         gen_21_cmp_pReg_15, gen_21_cmp_pReg_14, gen_21_cmp_pReg_13, 
         gen_21_cmp_pReg_12, gen_21_cmp_pReg_11, gen_21_cmp_pReg_10, 
         gen_21_cmp_pReg_9, gen_21_cmp_pReg_8, gen_21_cmp_pReg_7, 
         gen_21_cmp_pReg_6, gen_21_cmp_pReg_5, gen_21_cmp_pReg_4, 
         gen_21_cmp_pReg_3, gen_21_cmp_pReg_2, gen_21_cmp_pReg_1, 
         gen_21_cmp_pReg_0, gen_21_cmp_BSCmp_op2_0, gen_21_cmp_BSCmp_carryIn, 
         gen_20_cmp_pBs_30, gen_20_cmp_pBs_29, gen_20_cmp_pBs_28, 
         gen_20_cmp_pBs_27, gen_20_cmp_pBs_26, gen_20_cmp_pBs_25, 
         gen_20_cmp_pBs_24, gen_20_cmp_pBs_23, gen_20_cmp_pMux_30, 
         gen_20_cmp_pMux_29, gen_20_cmp_pMux_28, gen_20_cmp_pMux_27, 
         gen_20_cmp_pMux_26, gen_20_cmp_pMux_25, gen_20_cmp_pMux_24, 
         gen_20_cmp_pMux_23, gen_20_cmp_pMux_22, gen_20_cmp_pMux_21, 
         gen_20_cmp_pMux_20, gen_20_cmp_pMux_19, gen_20_cmp_pMux_18, 
         gen_20_cmp_pMux_17, gen_20_cmp_pMux_16, gen_20_cmp_pMux_15, 
         gen_20_cmp_pMux_14, gen_20_cmp_pMux_13, gen_20_cmp_pMux_12, 
         gen_20_cmp_pMux_11, gen_20_cmp_pMux_10, gen_20_cmp_pMux_9, 
         gen_20_cmp_pMux_8, gen_20_cmp_pMux_7, gen_20_cmp_pMux_6, 
         gen_20_cmp_pMux_5, gen_20_cmp_pMux_4, gen_20_cmp_pMux_3, 
         gen_20_cmp_pMux_2, gen_20_cmp_pMux_1, gen_20_cmp_pMux_0, 
         gen_20_cmp_pReg_30, gen_20_cmp_pReg_29, gen_20_cmp_pReg_28, 
         gen_20_cmp_pReg_27, gen_20_cmp_pReg_26, gen_20_cmp_pReg_25, 
         gen_20_cmp_pReg_24, gen_20_cmp_pReg_23, gen_20_cmp_pReg_22, 
         gen_20_cmp_pReg_21, gen_20_cmp_pReg_20, gen_20_cmp_pReg_19, 
         gen_20_cmp_pReg_18, gen_20_cmp_pReg_17, gen_20_cmp_pReg_16, 
         gen_20_cmp_pReg_15, gen_20_cmp_pReg_14, gen_20_cmp_pReg_13, 
         gen_20_cmp_pReg_12, gen_20_cmp_pReg_11, gen_20_cmp_pReg_10, 
         gen_20_cmp_pReg_9, gen_20_cmp_pReg_8, gen_20_cmp_pReg_7, 
         gen_20_cmp_pReg_6, gen_20_cmp_pReg_5, gen_20_cmp_pReg_4, 
         gen_20_cmp_pReg_3, gen_20_cmp_pReg_2, gen_20_cmp_pReg_1, 
         gen_20_cmp_pReg_0, gen_20_cmp_BSCmp_op2_0, gen_20_cmp_BSCmp_carryIn, 
         gen_19_cmp_pBs_30, gen_19_cmp_pBs_29, gen_19_cmp_pBs_28, 
         gen_19_cmp_pBs_27, gen_19_cmp_pBs_26, gen_19_cmp_pBs_25, 
         gen_19_cmp_pBs_24, gen_19_cmp_pBs_23, gen_19_cmp_pMux_30, 
         gen_19_cmp_pMux_29, gen_19_cmp_pMux_28, gen_19_cmp_pMux_27, 
         gen_19_cmp_pMux_26, gen_19_cmp_pMux_25, gen_19_cmp_pMux_24, 
         gen_19_cmp_pMux_23, gen_19_cmp_pMux_22, gen_19_cmp_pMux_21, 
         gen_19_cmp_pMux_20, gen_19_cmp_pMux_19, gen_19_cmp_pMux_18, 
         gen_19_cmp_pMux_17, gen_19_cmp_pMux_16, gen_19_cmp_pMux_15, 
         gen_19_cmp_pMux_14, gen_19_cmp_pMux_13, gen_19_cmp_pMux_12, 
         gen_19_cmp_pMux_11, gen_19_cmp_pMux_10, gen_19_cmp_pMux_9, 
         gen_19_cmp_pMux_8, gen_19_cmp_pMux_7, gen_19_cmp_pMux_6, 
         gen_19_cmp_pMux_5, gen_19_cmp_pMux_4, gen_19_cmp_pMux_3, 
         gen_19_cmp_pMux_2, gen_19_cmp_pMux_1, gen_19_cmp_pMux_0, 
         gen_19_cmp_pReg_30, gen_19_cmp_pReg_29, gen_19_cmp_pReg_28, 
         gen_19_cmp_pReg_27, gen_19_cmp_pReg_26, gen_19_cmp_pReg_25, 
         gen_19_cmp_pReg_24, gen_19_cmp_pReg_23, gen_19_cmp_pReg_22, 
         gen_19_cmp_pReg_21, gen_19_cmp_pReg_20, gen_19_cmp_pReg_19, 
         gen_19_cmp_pReg_18, gen_19_cmp_pReg_17, gen_19_cmp_pReg_16, 
         gen_19_cmp_pReg_15, gen_19_cmp_pReg_14, gen_19_cmp_pReg_13, 
         gen_19_cmp_pReg_12, gen_19_cmp_pReg_11, gen_19_cmp_pReg_10, 
         gen_19_cmp_pReg_9, gen_19_cmp_pReg_8, gen_19_cmp_pReg_7, 
         gen_19_cmp_pReg_6, gen_19_cmp_pReg_5, gen_19_cmp_pReg_4, 
         gen_19_cmp_pReg_3, gen_19_cmp_pReg_2, gen_19_cmp_pReg_1, 
         gen_19_cmp_pReg_0, gen_19_cmp_BSCmp_op2_0, gen_19_cmp_BSCmp_carryIn, 
         gen_18_cmp_pBs_30, gen_18_cmp_pBs_29, gen_18_cmp_pBs_28, 
         gen_18_cmp_pBs_27, gen_18_cmp_pBs_26, gen_18_cmp_pBs_25, 
         gen_18_cmp_pBs_24, gen_18_cmp_pBs_23, gen_18_cmp_pMux_30, 
         gen_18_cmp_pMux_29, gen_18_cmp_pMux_28, gen_18_cmp_pMux_27, 
         gen_18_cmp_pMux_26, gen_18_cmp_pMux_25, gen_18_cmp_pMux_24, 
         gen_18_cmp_pMux_23, gen_18_cmp_pMux_22, gen_18_cmp_pMux_21, 
         gen_18_cmp_pMux_20, gen_18_cmp_pMux_19, gen_18_cmp_pMux_18, 
         gen_18_cmp_pMux_17, gen_18_cmp_pMux_16, gen_18_cmp_pMux_15, 
         gen_18_cmp_pMux_14, gen_18_cmp_pMux_13, gen_18_cmp_pMux_12, 
         gen_18_cmp_pMux_11, gen_18_cmp_pMux_10, gen_18_cmp_pMux_9, 
         gen_18_cmp_pMux_8, gen_18_cmp_pMux_7, gen_18_cmp_pMux_6, 
         gen_18_cmp_pMux_5, gen_18_cmp_pMux_4, gen_18_cmp_pMux_3, 
         gen_18_cmp_pMux_2, gen_18_cmp_pMux_1, gen_18_cmp_pMux_0, 
         gen_18_cmp_pReg_30, gen_18_cmp_pReg_29, gen_18_cmp_pReg_28, 
         gen_18_cmp_pReg_27, gen_18_cmp_pReg_26, gen_18_cmp_pReg_25, 
         gen_18_cmp_pReg_24, gen_18_cmp_pReg_23, gen_18_cmp_pReg_22, 
         gen_18_cmp_pReg_21, gen_18_cmp_pReg_20, gen_18_cmp_pReg_19, 
         gen_18_cmp_pReg_18, gen_18_cmp_pReg_17, gen_18_cmp_pReg_16, 
         gen_18_cmp_pReg_15, gen_18_cmp_pReg_14, gen_18_cmp_pReg_13, 
         gen_18_cmp_pReg_12, gen_18_cmp_pReg_11, gen_18_cmp_pReg_10, 
         gen_18_cmp_pReg_9, gen_18_cmp_pReg_8, gen_18_cmp_pReg_7, 
         gen_18_cmp_pReg_6, gen_18_cmp_pReg_5, gen_18_cmp_pReg_4, 
         gen_18_cmp_pReg_3, gen_18_cmp_pReg_2, gen_18_cmp_pReg_1, 
         gen_18_cmp_pReg_0, gen_18_cmp_BSCmp_op2_0, gen_18_cmp_BSCmp_carryIn, 
         gen_17_cmp_pBs_30, gen_17_cmp_pBs_29, gen_17_cmp_pBs_28, 
         gen_17_cmp_pBs_27, gen_17_cmp_pBs_26, gen_17_cmp_pBs_25, 
         gen_17_cmp_pBs_24, gen_17_cmp_pBs_23, gen_17_cmp_pMux_30, 
         gen_17_cmp_pMux_29, gen_17_cmp_pMux_28, gen_17_cmp_pMux_27, 
         gen_17_cmp_pMux_26, gen_17_cmp_pMux_25, gen_17_cmp_pMux_24, 
         gen_17_cmp_pMux_23, gen_17_cmp_pMux_22, gen_17_cmp_pMux_21, 
         gen_17_cmp_pMux_20, gen_17_cmp_pMux_19, gen_17_cmp_pMux_18, 
         gen_17_cmp_pMux_17, gen_17_cmp_pMux_16, gen_17_cmp_pMux_15, 
         gen_17_cmp_pMux_14, gen_17_cmp_pMux_13, gen_17_cmp_pMux_12, 
         gen_17_cmp_pMux_11, gen_17_cmp_pMux_10, gen_17_cmp_pMux_9, 
         gen_17_cmp_pMux_8, gen_17_cmp_pMux_7, gen_17_cmp_pMux_6, 
         gen_17_cmp_pMux_5, gen_17_cmp_pMux_4, gen_17_cmp_pMux_3, 
         gen_17_cmp_pMux_2, gen_17_cmp_pMux_1, gen_17_cmp_pMux_0, 
         gen_17_cmp_pReg_30, gen_17_cmp_pReg_29, gen_17_cmp_pReg_28, 
         gen_17_cmp_pReg_27, gen_17_cmp_pReg_26, gen_17_cmp_pReg_25, 
         gen_17_cmp_pReg_24, gen_17_cmp_pReg_23, gen_17_cmp_pReg_22, 
         gen_17_cmp_pReg_21, gen_17_cmp_pReg_20, gen_17_cmp_pReg_19, 
         gen_17_cmp_pReg_18, gen_17_cmp_pReg_17, gen_17_cmp_pReg_16, 
         gen_17_cmp_pReg_15, gen_17_cmp_pReg_14, gen_17_cmp_pReg_13, 
         gen_17_cmp_pReg_12, gen_17_cmp_pReg_11, gen_17_cmp_pReg_10, 
         gen_17_cmp_pReg_9, gen_17_cmp_pReg_8, gen_17_cmp_pReg_7, 
         gen_17_cmp_pReg_6, gen_17_cmp_pReg_5, gen_17_cmp_pReg_4, 
         gen_17_cmp_pReg_3, gen_17_cmp_pReg_2, gen_17_cmp_pReg_1, 
         gen_17_cmp_pReg_0, gen_17_cmp_BSCmp_op2_0, gen_17_cmp_BSCmp_carryIn, 
         gen_16_cmp_pBs_30, gen_16_cmp_pBs_29, gen_16_cmp_pBs_28, 
         gen_16_cmp_pBs_27, gen_16_cmp_pBs_26, gen_16_cmp_pBs_25, 
         gen_16_cmp_pBs_24, gen_16_cmp_pBs_23, gen_16_cmp_pMux_30, 
         gen_16_cmp_pMux_29, gen_16_cmp_pMux_28, gen_16_cmp_pMux_27, 
         gen_16_cmp_pMux_26, gen_16_cmp_pMux_25, gen_16_cmp_pMux_24, 
         gen_16_cmp_pMux_23, gen_16_cmp_pMux_22, gen_16_cmp_pMux_21, 
         gen_16_cmp_pMux_20, gen_16_cmp_pMux_19, gen_16_cmp_pMux_18, 
         gen_16_cmp_pMux_17, gen_16_cmp_pMux_16, gen_16_cmp_pMux_15, 
         gen_16_cmp_pMux_14, gen_16_cmp_pMux_13, gen_16_cmp_pMux_12, 
         gen_16_cmp_pMux_11, gen_16_cmp_pMux_10, gen_16_cmp_pMux_9, 
         gen_16_cmp_pMux_8, gen_16_cmp_pMux_7, gen_16_cmp_pMux_6, 
         gen_16_cmp_pMux_5, gen_16_cmp_pMux_4, gen_16_cmp_pMux_3, 
         gen_16_cmp_pMux_2, gen_16_cmp_pMux_1, gen_16_cmp_pMux_0, 
         gen_16_cmp_pReg_30, gen_16_cmp_pReg_29, gen_16_cmp_pReg_28, 
         gen_16_cmp_pReg_27, gen_16_cmp_pReg_26, gen_16_cmp_pReg_25, 
         gen_16_cmp_pReg_24, gen_16_cmp_pReg_23, gen_16_cmp_pReg_22, 
         gen_16_cmp_pReg_21, gen_16_cmp_pReg_20, gen_16_cmp_pReg_19, 
         gen_16_cmp_pReg_18, gen_16_cmp_pReg_17, gen_16_cmp_pReg_16, 
         gen_16_cmp_pReg_15, gen_16_cmp_pReg_14, gen_16_cmp_pReg_13, 
         gen_16_cmp_pReg_12, gen_16_cmp_pReg_11, gen_16_cmp_pReg_10, 
         gen_16_cmp_pReg_9, gen_16_cmp_pReg_8, gen_16_cmp_pReg_7, 
         gen_16_cmp_pReg_6, gen_16_cmp_pReg_5, gen_16_cmp_pReg_4, 
         gen_16_cmp_pReg_3, gen_16_cmp_pReg_2, gen_16_cmp_pReg_1, 
         gen_16_cmp_pReg_0, gen_16_cmp_BSCmp_op2_0, gen_16_cmp_BSCmp_carryIn, 
         gen_15_cmp_pBs_30, gen_15_cmp_pBs_29, gen_15_cmp_pBs_28, 
         gen_15_cmp_pBs_27, gen_15_cmp_pBs_26, gen_15_cmp_pBs_25, 
         gen_15_cmp_pBs_24, gen_15_cmp_pBs_23, gen_15_cmp_pMux_30, 
         gen_15_cmp_pMux_29, gen_15_cmp_pMux_28, gen_15_cmp_pMux_27, 
         gen_15_cmp_pMux_26, gen_15_cmp_pMux_25, gen_15_cmp_pMux_24, 
         gen_15_cmp_pMux_23, gen_15_cmp_pMux_22, gen_15_cmp_pMux_21, 
         gen_15_cmp_pMux_20, gen_15_cmp_pMux_19, gen_15_cmp_pMux_18, 
         gen_15_cmp_pMux_17, gen_15_cmp_pMux_16, gen_15_cmp_pMux_15, 
         gen_15_cmp_pMux_14, gen_15_cmp_pMux_13, gen_15_cmp_pMux_12, 
         gen_15_cmp_pMux_11, gen_15_cmp_pMux_10, gen_15_cmp_pMux_9, 
         gen_15_cmp_pMux_8, gen_15_cmp_pMux_7, gen_15_cmp_pMux_6, 
         gen_15_cmp_pMux_5, gen_15_cmp_pMux_4, gen_15_cmp_pMux_3, 
         gen_15_cmp_pMux_2, gen_15_cmp_pMux_1, gen_15_cmp_pMux_0, 
         gen_15_cmp_pReg_30, gen_15_cmp_pReg_29, gen_15_cmp_pReg_28, 
         gen_15_cmp_pReg_27, gen_15_cmp_pReg_26, gen_15_cmp_pReg_25, 
         gen_15_cmp_pReg_24, gen_15_cmp_pReg_23, gen_15_cmp_pReg_22, 
         gen_15_cmp_pReg_21, gen_15_cmp_pReg_20, gen_15_cmp_pReg_19, 
         gen_15_cmp_pReg_18, gen_15_cmp_pReg_17, gen_15_cmp_pReg_16, 
         gen_15_cmp_pReg_15, gen_15_cmp_pReg_14, gen_15_cmp_pReg_13, 
         gen_15_cmp_pReg_12, gen_15_cmp_pReg_11, gen_15_cmp_pReg_10, 
         gen_15_cmp_pReg_9, gen_15_cmp_pReg_8, gen_15_cmp_pReg_7, 
         gen_15_cmp_pReg_6, gen_15_cmp_pReg_5, gen_15_cmp_pReg_4, 
         gen_15_cmp_pReg_3, gen_15_cmp_pReg_2, gen_15_cmp_pReg_1, 
         gen_15_cmp_pReg_0, gen_15_cmp_BSCmp_op2_0, gen_15_cmp_BSCmp_carryIn, 
         gen_14_cmp_pBs_30, gen_14_cmp_pBs_29, gen_14_cmp_pBs_28, 
         gen_14_cmp_pBs_27, gen_14_cmp_pBs_26, gen_14_cmp_pBs_25, 
         gen_14_cmp_pBs_24, gen_14_cmp_pBs_23, gen_14_cmp_pMux_30, 
         gen_14_cmp_pMux_29, gen_14_cmp_pMux_28, gen_14_cmp_pMux_27, 
         gen_14_cmp_pMux_26, gen_14_cmp_pMux_25, gen_14_cmp_pMux_24, 
         gen_14_cmp_pMux_23, gen_14_cmp_pMux_22, gen_14_cmp_pMux_21, 
         gen_14_cmp_pMux_20, gen_14_cmp_pMux_19, gen_14_cmp_pMux_18, 
         gen_14_cmp_pMux_17, gen_14_cmp_pMux_16, gen_14_cmp_pMux_15, 
         gen_14_cmp_pMux_14, gen_14_cmp_pMux_13, gen_14_cmp_pMux_12, 
         gen_14_cmp_pMux_11, gen_14_cmp_pMux_10, gen_14_cmp_pMux_9, 
         gen_14_cmp_pMux_8, gen_14_cmp_pMux_7, gen_14_cmp_pMux_6, 
         gen_14_cmp_pMux_5, gen_14_cmp_pMux_4, gen_14_cmp_pMux_3, 
         gen_14_cmp_pMux_2, gen_14_cmp_pMux_1, gen_14_cmp_pMux_0, 
         gen_14_cmp_pReg_30, gen_14_cmp_pReg_29, gen_14_cmp_pReg_28, 
         gen_14_cmp_pReg_27, gen_14_cmp_pReg_26, gen_14_cmp_pReg_25, 
         gen_14_cmp_pReg_24, gen_14_cmp_pReg_23, gen_14_cmp_pReg_22, 
         gen_14_cmp_pReg_21, gen_14_cmp_pReg_20, gen_14_cmp_pReg_19, 
         gen_14_cmp_pReg_18, gen_14_cmp_pReg_17, gen_14_cmp_pReg_16, 
         gen_14_cmp_pReg_15, gen_14_cmp_pReg_14, gen_14_cmp_pReg_13, 
         gen_14_cmp_pReg_12, gen_14_cmp_pReg_11, gen_14_cmp_pReg_10, 
         gen_14_cmp_pReg_9, gen_14_cmp_pReg_8, gen_14_cmp_pReg_7, 
         gen_14_cmp_pReg_6, gen_14_cmp_pReg_5, gen_14_cmp_pReg_4, 
         gen_14_cmp_pReg_3, gen_14_cmp_pReg_2, gen_14_cmp_pReg_1, 
         gen_14_cmp_pReg_0, gen_14_cmp_BSCmp_op2_0, gen_14_cmp_BSCmp_carryIn, 
         gen_13_cmp_pBs_30, gen_13_cmp_pBs_29, gen_13_cmp_pBs_28, 
         gen_13_cmp_pBs_27, gen_13_cmp_pBs_26, gen_13_cmp_pBs_25, 
         gen_13_cmp_pBs_24, gen_13_cmp_pBs_23, gen_13_cmp_pMux_30, 
         gen_13_cmp_pMux_29, gen_13_cmp_pMux_28, gen_13_cmp_pMux_27, 
         gen_13_cmp_pMux_26, gen_13_cmp_pMux_25, gen_13_cmp_pMux_24, 
         gen_13_cmp_pMux_23, gen_13_cmp_pMux_22, gen_13_cmp_pMux_21, 
         gen_13_cmp_pMux_20, gen_13_cmp_pMux_19, gen_13_cmp_pMux_18, 
         gen_13_cmp_pMux_17, gen_13_cmp_pMux_16, gen_13_cmp_pMux_15, 
         gen_13_cmp_pMux_14, gen_13_cmp_pMux_13, gen_13_cmp_pMux_12, 
         gen_13_cmp_pMux_11, gen_13_cmp_pMux_10, gen_13_cmp_pMux_9, 
         gen_13_cmp_pMux_8, gen_13_cmp_pMux_7, gen_13_cmp_pMux_6, 
         gen_13_cmp_pMux_5, gen_13_cmp_pMux_4, gen_13_cmp_pMux_3, 
         gen_13_cmp_pMux_2, gen_13_cmp_pMux_1, gen_13_cmp_pMux_0, 
         gen_13_cmp_pReg_30, gen_13_cmp_pReg_29, gen_13_cmp_pReg_28, 
         gen_13_cmp_pReg_27, gen_13_cmp_pReg_26, gen_13_cmp_pReg_25, 
         gen_13_cmp_pReg_24, gen_13_cmp_pReg_23, gen_13_cmp_pReg_22, 
         gen_13_cmp_pReg_21, gen_13_cmp_pReg_20, gen_13_cmp_pReg_19, 
         gen_13_cmp_pReg_18, gen_13_cmp_pReg_17, gen_13_cmp_pReg_16, 
         gen_13_cmp_pReg_15, gen_13_cmp_pReg_14, gen_13_cmp_pReg_13, 
         gen_13_cmp_pReg_12, gen_13_cmp_pReg_11, gen_13_cmp_pReg_10, 
         gen_13_cmp_pReg_9, gen_13_cmp_pReg_8, gen_13_cmp_pReg_7, 
         gen_13_cmp_pReg_6, gen_13_cmp_pReg_5, gen_13_cmp_pReg_4, 
         gen_13_cmp_pReg_3, gen_13_cmp_pReg_2, gen_13_cmp_pReg_1, 
         gen_13_cmp_pReg_0, gen_13_cmp_BSCmp_op2_0, gen_13_cmp_BSCmp_carryIn, 
         gen_12_cmp_pBs_30, gen_12_cmp_pBs_29, gen_12_cmp_pBs_28, 
         gen_12_cmp_pBs_27, gen_12_cmp_pBs_26, gen_12_cmp_pBs_25, 
         gen_12_cmp_pBs_24, gen_12_cmp_pBs_23, gen_12_cmp_pMux_30, 
         gen_12_cmp_pMux_29, gen_12_cmp_pMux_28, gen_12_cmp_pMux_27, 
         gen_12_cmp_pMux_26, gen_12_cmp_pMux_25, gen_12_cmp_pMux_24, 
         gen_12_cmp_pMux_23, gen_12_cmp_pMux_22, gen_12_cmp_pMux_21, 
         gen_12_cmp_pMux_20, gen_12_cmp_pMux_19, gen_12_cmp_pMux_18, 
         gen_12_cmp_pMux_17, gen_12_cmp_pMux_16, gen_12_cmp_pMux_15, 
         gen_12_cmp_pMux_14, gen_12_cmp_pMux_13, gen_12_cmp_pMux_12, 
         gen_12_cmp_pMux_11, gen_12_cmp_pMux_10, gen_12_cmp_pMux_9, 
         gen_12_cmp_pMux_8, gen_12_cmp_pMux_7, gen_12_cmp_pMux_6, 
         gen_12_cmp_pMux_5, gen_12_cmp_pMux_4, gen_12_cmp_pMux_3, 
         gen_12_cmp_pMux_2, gen_12_cmp_pMux_1, gen_12_cmp_pMux_0, 
         gen_12_cmp_pReg_30, gen_12_cmp_pReg_29, gen_12_cmp_pReg_28, 
         gen_12_cmp_pReg_27, gen_12_cmp_pReg_26, gen_12_cmp_pReg_25, 
         gen_12_cmp_pReg_24, gen_12_cmp_pReg_23, gen_12_cmp_pReg_22, 
         gen_12_cmp_pReg_21, gen_12_cmp_pReg_20, gen_12_cmp_pReg_19, 
         gen_12_cmp_pReg_18, gen_12_cmp_pReg_17, gen_12_cmp_pReg_16, 
         gen_12_cmp_pReg_15, gen_12_cmp_pReg_14, gen_12_cmp_pReg_13, 
         gen_12_cmp_pReg_12, gen_12_cmp_pReg_11, gen_12_cmp_pReg_10, 
         gen_12_cmp_pReg_9, gen_12_cmp_pReg_8, gen_12_cmp_pReg_7, 
         gen_12_cmp_pReg_6, gen_12_cmp_pReg_5, gen_12_cmp_pReg_4, 
         gen_12_cmp_pReg_3, gen_12_cmp_pReg_2, gen_12_cmp_pReg_1, 
         gen_12_cmp_pReg_0, gen_12_cmp_BSCmp_op2_0, gen_12_cmp_BSCmp_carryIn, 
         gen_11_cmp_pBs_30, gen_11_cmp_pBs_29, gen_11_cmp_pBs_28, 
         gen_11_cmp_pBs_27, gen_11_cmp_pBs_26, gen_11_cmp_pBs_25, 
         gen_11_cmp_pBs_24, gen_11_cmp_pBs_23, gen_11_cmp_pMux_30, 
         gen_11_cmp_pMux_29, gen_11_cmp_pMux_28, gen_11_cmp_pMux_27, 
         gen_11_cmp_pMux_26, gen_11_cmp_pMux_25, gen_11_cmp_pMux_24, 
         gen_11_cmp_pMux_23, gen_11_cmp_pMux_22, gen_11_cmp_pMux_21, 
         gen_11_cmp_pMux_20, gen_11_cmp_pMux_19, gen_11_cmp_pMux_18, 
         gen_11_cmp_pMux_17, gen_11_cmp_pMux_16, gen_11_cmp_pMux_15, 
         gen_11_cmp_pMux_14, gen_11_cmp_pMux_13, gen_11_cmp_pMux_12, 
         gen_11_cmp_pMux_11, gen_11_cmp_pMux_10, gen_11_cmp_pMux_9, 
         gen_11_cmp_pMux_8, gen_11_cmp_pMux_7, gen_11_cmp_pMux_6, 
         gen_11_cmp_pMux_5, gen_11_cmp_pMux_4, gen_11_cmp_pMux_3, 
         gen_11_cmp_pMux_2, gen_11_cmp_pMux_1, gen_11_cmp_pMux_0, 
         gen_11_cmp_pReg_30, gen_11_cmp_pReg_29, gen_11_cmp_pReg_28, 
         gen_11_cmp_pReg_27, gen_11_cmp_pReg_26, gen_11_cmp_pReg_25, 
         gen_11_cmp_pReg_24, gen_11_cmp_pReg_23, gen_11_cmp_pReg_22, 
         gen_11_cmp_pReg_21, gen_11_cmp_pReg_20, gen_11_cmp_pReg_19, 
         gen_11_cmp_pReg_18, gen_11_cmp_pReg_17, gen_11_cmp_pReg_16, 
         gen_11_cmp_pReg_15, gen_11_cmp_pReg_14, gen_11_cmp_pReg_13, 
         gen_11_cmp_pReg_12, gen_11_cmp_pReg_11, gen_11_cmp_pReg_10, 
         gen_11_cmp_pReg_9, gen_11_cmp_pReg_8, gen_11_cmp_pReg_7, 
         gen_11_cmp_pReg_6, gen_11_cmp_pReg_5, gen_11_cmp_pReg_4, 
         gen_11_cmp_pReg_3, gen_11_cmp_pReg_2, gen_11_cmp_pReg_1, 
         gen_11_cmp_pReg_0, gen_11_cmp_BSCmp_op2_0, gen_11_cmp_BSCmp_carryIn, 
         gen_10_cmp_pBs_30, gen_10_cmp_pBs_29, gen_10_cmp_pBs_28, 
         gen_10_cmp_pBs_27, gen_10_cmp_pBs_26, gen_10_cmp_pBs_25, 
         gen_10_cmp_pBs_24, gen_10_cmp_pBs_23, gen_10_cmp_pMux_30, 
         gen_10_cmp_pMux_29, gen_10_cmp_pMux_28, gen_10_cmp_pMux_27, 
         gen_10_cmp_pMux_26, gen_10_cmp_pMux_25, gen_10_cmp_pMux_24, 
         gen_10_cmp_pMux_23, gen_10_cmp_pMux_22, gen_10_cmp_pMux_21, 
         gen_10_cmp_pMux_20, gen_10_cmp_pMux_19, gen_10_cmp_pMux_18, 
         gen_10_cmp_pMux_17, gen_10_cmp_pMux_16, gen_10_cmp_pMux_15, 
         gen_10_cmp_pMux_14, gen_10_cmp_pMux_13, gen_10_cmp_pMux_12, 
         gen_10_cmp_pMux_11, gen_10_cmp_pMux_10, gen_10_cmp_pMux_9, 
         gen_10_cmp_pMux_8, gen_10_cmp_pMux_7, gen_10_cmp_pMux_6, 
         gen_10_cmp_pMux_5, gen_10_cmp_pMux_4, gen_10_cmp_pMux_3, 
         gen_10_cmp_pMux_2, gen_10_cmp_pMux_1, gen_10_cmp_pMux_0, 
         gen_10_cmp_pReg_30, gen_10_cmp_pReg_29, gen_10_cmp_pReg_28, 
         gen_10_cmp_pReg_27, gen_10_cmp_pReg_26, gen_10_cmp_pReg_25, 
         gen_10_cmp_pReg_24, gen_10_cmp_pReg_23, gen_10_cmp_pReg_22, 
         gen_10_cmp_pReg_21, gen_10_cmp_pReg_20, gen_10_cmp_pReg_19, 
         gen_10_cmp_pReg_18, gen_10_cmp_pReg_17, gen_10_cmp_pReg_16, 
         gen_10_cmp_pReg_15, gen_10_cmp_pReg_14, gen_10_cmp_pReg_13, 
         gen_10_cmp_pReg_12, gen_10_cmp_pReg_11, gen_10_cmp_pReg_10, 
         gen_10_cmp_pReg_9, gen_10_cmp_pReg_8, gen_10_cmp_pReg_7, 
         gen_10_cmp_pReg_6, gen_10_cmp_pReg_5, gen_10_cmp_pReg_4, 
         gen_10_cmp_pReg_3, gen_10_cmp_pReg_2, gen_10_cmp_pReg_1, 
         gen_10_cmp_pReg_0, gen_10_cmp_BSCmp_op2_0, gen_10_cmp_BSCmp_carryIn, 
         gen_9_cmp_pBs_30, gen_9_cmp_pBs_29, gen_9_cmp_pBs_28, gen_9_cmp_pBs_27, 
         gen_9_cmp_pBs_26, gen_9_cmp_pBs_25, gen_9_cmp_pBs_24, gen_9_cmp_pBs_23, 
         gen_9_cmp_pMux_30, gen_9_cmp_pMux_29, gen_9_cmp_pMux_28, 
         gen_9_cmp_pMux_27, gen_9_cmp_pMux_26, gen_9_cmp_pMux_25, 
         gen_9_cmp_pMux_24, gen_9_cmp_pMux_23, gen_9_cmp_pMux_22, 
         gen_9_cmp_pMux_21, gen_9_cmp_pMux_20, gen_9_cmp_pMux_19, 
         gen_9_cmp_pMux_18, gen_9_cmp_pMux_17, gen_9_cmp_pMux_16, 
         gen_9_cmp_pMux_15, gen_9_cmp_pMux_14, gen_9_cmp_pMux_13, 
         gen_9_cmp_pMux_12, gen_9_cmp_pMux_11, gen_9_cmp_pMux_10, 
         gen_9_cmp_pMux_9, gen_9_cmp_pMux_8, gen_9_cmp_pMux_7, gen_9_cmp_pMux_6, 
         gen_9_cmp_pMux_5, gen_9_cmp_pMux_4, gen_9_cmp_pMux_3, gen_9_cmp_pMux_2, 
         gen_9_cmp_pMux_1, gen_9_cmp_pMux_0, gen_9_cmp_pReg_30, 
         gen_9_cmp_pReg_29, gen_9_cmp_pReg_28, gen_9_cmp_pReg_27, 
         gen_9_cmp_pReg_26, gen_9_cmp_pReg_25, gen_9_cmp_pReg_24, 
         gen_9_cmp_pReg_23, gen_9_cmp_pReg_22, gen_9_cmp_pReg_21, 
         gen_9_cmp_pReg_20, gen_9_cmp_pReg_19, gen_9_cmp_pReg_18, 
         gen_9_cmp_pReg_17, gen_9_cmp_pReg_16, gen_9_cmp_pReg_15, 
         gen_9_cmp_pReg_14, gen_9_cmp_pReg_13, gen_9_cmp_pReg_12, 
         gen_9_cmp_pReg_11, gen_9_cmp_pReg_10, gen_9_cmp_pReg_9, 
         gen_9_cmp_pReg_8, gen_9_cmp_pReg_7, gen_9_cmp_pReg_6, gen_9_cmp_pReg_5, 
         gen_9_cmp_pReg_4, gen_9_cmp_pReg_3, gen_9_cmp_pReg_2, gen_9_cmp_pReg_1, 
         gen_9_cmp_pReg_0, gen_9_cmp_BSCmp_op2_0, gen_9_cmp_BSCmp_carryIn, 
         gen_8_cmp_pBs_30, gen_8_cmp_pBs_29, gen_8_cmp_pBs_28, gen_8_cmp_pBs_27, 
         gen_8_cmp_pBs_26, gen_8_cmp_pBs_25, gen_8_cmp_pBs_24, gen_8_cmp_pBs_23, 
         gen_8_cmp_pMux_30, gen_8_cmp_pMux_29, gen_8_cmp_pMux_28, 
         gen_8_cmp_pMux_27, gen_8_cmp_pMux_26, gen_8_cmp_pMux_25, 
         gen_8_cmp_pMux_24, gen_8_cmp_pMux_23, gen_8_cmp_pMux_22, 
         gen_8_cmp_pMux_21, gen_8_cmp_pMux_20, gen_8_cmp_pMux_19, 
         gen_8_cmp_pMux_18, gen_8_cmp_pMux_17, gen_8_cmp_pMux_16, 
         gen_8_cmp_pMux_15, gen_8_cmp_pMux_14, gen_8_cmp_pMux_13, 
         gen_8_cmp_pMux_12, gen_8_cmp_pMux_11, gen_8_cmp_pMux_10, 
         gen_8_cmp_pMux_9, gen_8_cmp_pMux_8, gen_8_cmp_pMux_7, gen_8_cmp_pMux_6, 
         gen_8_cmp_pMux_5, gen_8_cmp_pMux_4, gen_8_cmp_pMux_3, gen_8_cmp_pMux_2, 
         gen_8_cmp_pMux_1, gen_8_cmp_pMux_0, gen_8_cmp_pReg_30, 
         gen_8_cmp_pReg_29, gen_8_cmp_pReg_28, gen_8_cmp_pReg_27, 
         gen_8_cmp_pReg_26, gen_8_cmp_pReg_25, gen_8_cmp_pReg_24, 
         gen_8_cmp_pReg_23, gen_8_cmp_pReg_22, gen_8_cmp_pReg_21, 
         gen_8_cmp_pReg_20, gen_8_cmp_pReg_19, gen_8_cmp_pReg_18, 
         gen_8_cmp_pReg_17, gen_8_cmp_pReg_16, gen_8_cmp_pReg_15, 
         gen_8_cmp_pReg_14, gen_8_cmp_pReg_13, gen_8_cmp_pReg_12, 
         gen_8_cmp_pReg_11, gen_8_cmp_pReg_10, gen_8_cmp_pReg_9, 
         gen_8_cmp_pReg_8, gen_8_cmp_pReg_7, gen_8_cmp_pReg_6, gen_8_cmp_pReg_5, 
         gen_8_cmp_pReg_4, gen_8_cmp_pReg_3, gen_8_cmp_pReg_2, gen_8_cmp_pReg_1, 
         gen_8_cmp_pReg_0, gen_8_cmp_BSCmp_op2_0, gen_8_cmp_BSCmp_carryIn, 
         gen_7_cmp_pBs_30, gen_7_cmp_pBs_29, gen_7_cmp_pBs_28, gen_7_cmp_pBs_27, 
         gen_7_cmp_pBs_26, gen_7_cmp_pBs_25, gen_7_cmp_pBs_24, gen_7_cmp_pBs_23, 
         gen_7_cmp_pMux_30, gen_7_cmp_pMux_29, gen_7_cmp_pMux_28, 
         gen_7_cmp_pMux_27, gen_7_cmp_pMux_26, gen_7_cmp_pMux_25, 
         gen_7_cmp_pMux_24, gen_7_cmp_pMux_23, gen_7_cmp_pMux_22, 
         gen_7_cmp_pMux_21, gen_7_cmp_pMux_20, gen_7_cmp_pMux_19, 
         gen_7_cmp_pMux_18, gen_7_cmp_pMux_17, gen_7_cmp_pMux_16, 
         gen_7_cmp_pMux_15, gen_7_cmp_pMux_14, gen_7_cmp_pMux_13, 
         gen_7_cmp_pMux_12, gen_7_cmp_pMux_11, gen_7_cmp_pMux_10, 
         gen_7_cmp_pMux_9, gen_7_cmp_pMux_8, gen_7_cmp_pMux_7, gen_7_cmp_pMux_6, 
         gen_7_cmp_pMux_5, gen_7_cmp_pMux_4, gen_7_cmp_pMux_3, gen_7_cmp_pMux_2, 
         gen_7_cmp_pMux_1, gen_7_cmp_pMux_0, gen_7_cmp_pReg_30, 
         gen_7_cmp_pReg_29, gen_7_cmp_pReg_28, gen_7_cmp_pReg_27, 
         gen_7_cmp_pReg_26, gen_7_cmp_pReg_25, gen_7_cmp_pReg_24, 
         gen_7_cmp_pReg_23, gen_7_cmp_pReg_22, gen_7_cmp_pReg_21, 
         gen_7_cmp_pReg_20, gen_7_cmp_pReg_19, gen_7_cmp_pReg_18, 
         gen_7_cmp_pReg_17, gen_7_cmp_pReg_16, gen_7_cmp_pReg_15, 
         gen_7_cmp_pReg_14, gen_7_cmp_pReg_13, gen_7_cmp_pReg_12, 
         gen_7_cmp_pReg_11, gen_7_cmp_pReg_10, gen_7_cmp_pReg_9, 
         gen_7_cmp_pReg_8, gen_7_cmp_pReg_7, gen_7_cmp_pReg_6, gen_7_cmp_pReg_5, 
         gen_7_cmp_pReg_4, gen_7_cmp_pReg_3, gen_7_cmp_pReg_2, gen_7_cmp_pReg_1, 
         gen_7_cmp_pReg_0, gen_7_cmp_BSCmp_op2_0, gen_7_cmp_BSCmp_carryIn, 
         gen_6_cmp_pBs_30, gen_6_cmp_pBs_29, gen_6_cmp_pBs_28, gen_6_cmp_pBs_27, 
         gen_6_cmp_pBs_26, gen_6_cmp_pBs_25, gen_6_cmp_pBs_24, gen_6_cmp_pBs_23, 
         gen_6_cmp_pMux_30, gen_6_cmp_pMux_29, gen_6_cmp_pMux_28, 
         gen_6_cmp_pMux_27, gen_6_cmp_pMux_26, gen_6_cmp_pMux_25, 
         gen_6_cmp_pMux_24, gen_6_cmp_pMux_23, gen_6_cmp_pMux_22, 
         gen_6_cmp_pMux_21, gen_6_cmp_pMux_20, gen_6_cmp_pMux_19, 
         gen_6_cmp_pMux_18, gen_6_cmp_pMux_17, gen_6_cmp_pMux_16, 
         gen_6_cmp_pMux_15, gen_6_cmp_pMux_14, gen_6_cmp_pMux_13, 
         gen_6_cmp_pMux_12, gen_6_cmp_pMux_11, gen_6_cmp_pMux_10, 
         gen_6_cmp_pMux_9, gen_6_cmp_pMux_8, gen_6_cmp_pMux_7, gen_6_cmp_pMux_6, 
         gen_6_cmp_pMux_5, gen_6_cmp_pMux_4, gen_6_cmp_pMux_3, gen_6_cmp_pMux_2, 
         gen_6_cmp_pMux_1, gen_6_cmp_pMux_0, gen_6_cmp_pReg_30, 
         gen_6_cmp_pReg_29, gen_6_cmp_pReg_28, gen_6_cmp_pReg_27, 
         gen_6_cmp_pReg_26, gen_6_cmp_pReg_25, gen_6_cmp_pReg_24, 
         gen_6_cmp_pReg_23, gen_6_cmp_pReg_22, gen_6_cmp_pReg_21, 
         gen_6_cmp_pReg_20, gen_6_cmp_pReg_19, gen_6_cmp_pReg_18, 
         gen_6_cmp_pReg_17, gen_6_cmp_pReg_16, gen_6_cmp_pReg_15, 
         gen_6_cmp_pReg_14, gen_6_cmp_pReg_13, gen_6_cmp_pReg_12, 
         gen_6_cmp_pReg_11, gen_6_cmp_pReg_10, gen_6_cmp_pReg_9, 
         gen_6_cmp_pReg_8, gen_6_cmp_pReg_7, gen_6_cmp_pReg_6, gen_6_cmp_pReg_5, 
         gen_6_cmp_pReg_4, gen_6_cmp_pReg_3, gen_6_cmp_pReg_2, gen_6_cmp_pReg_1, 
         gen_6_cmp_pReg_0, gen_6_cmp_BSCmp_op2_0, gen_6_cmp_BSCmp_carryIn, 
         gen_5_cmp_pBs_30, gen_5_cmp_pBs_29, gen_5_cmp_pBs_28, gen_5_cmp_pBs_27, 
         gen_5_cmp_pBs_26, gen_5_cmp_pBs_25, gen_5_cmp_pBs_24, gen_5_cmp_pBs_23, 
         gen_5_cmp_pMux_30, gen_5_cmp_pMux_29, gen_5_cmp_pMux_28, 
         gen_5_cmp_pMux_27, gen_5_cmp_pMux_26, gen_5_cmp_pMux_25, 
         gen_5_cmp_pMux_24, gen_5_cmp_pMux_23, gen_5_cmp_pMux_22, 
         gen_5_cmp_pMux_21, gen_5_cmp_pMux_20, gen_5_cmp_pMux_19, 
         gen_5_cmp_pMux_18, gen_5_cmp_pMux_17, gen_5_cmp_pMux_16, 
         gen_5_cmp_pMux_15, gen_5_cmp_pMux_14, gen_5_cmp_pMux_13, 
         gen_5_cmp_pMux_12, gen_5_cmp_pMux_11, gen_5_cmp_pMux_10, 
         gen_5_cmp_pMux_9, gen_5_cmp_pMux_8, gen_5_cmp_pMux_7, gen_5_cmp_pMux_6, 
         gen_5_cmp_pMux_5, gen_5_cmp_pMux_4, gen_5_cmp_pMux_3, gen_5_cmp_pMux_2, 
         gen_5_cmp_pMux_1, gen_5_cmp_pMux_0, gen_5_cmp_pReg_30, 
         gen_5_cmp_pReg_29, gen_5_cmp_pReg_28, gen_5_cmp_pReg_27, 
         gen_5_cmp_pReg_26, gen_5_cmp_pReg_25, gen_5_cmp_pReg_24, 
         gen_5_cmp_pReg_23, gen_5_cmp_pReg_22, gen_5_cmp_pReg_21, 
         gen_5_cmp_pReg_20, gen_5_cmp_pReg_19, gen_5_cmp_pReg_18, 
         gen_5_cmp_pReg_17, gen_5_cmp_pReg_16, gen_5_cmp_pReg_15, 
         gen_5_cmp_pReg_14, gen_5_cmp_pReg_13, gen_5_cmp_pReg_12, 
         gen_5_cmp_pReg_11, gen_5_cmp_pReg_10, gen_5_cmp_pReg_9, 
         gen_5_cmp_pReg_8, gen_5_cmp_pReg_7, gen_5_cmp_pReg_6, gen_5_cmp_pReg_5, 
         gen_5_cmp_pReg_4, gen_5_cmp_pReg_3, gen_5_cmp_pReg_2, gen_5_cmp_pReg_1, 
         gen_5_cmp_pReg_0, gen_5_cmp_BSCmp_op2_0, gen_5_cmp_BSCmp_carryIn, 
         gen_4_cmp_pBs_30, gen_4_cmp_pBs_29, gen_4_cmp_pBs_28, gen_4_cmp_pBs_27, 
         gen_4_cmp_pBs_26, gen_4_cmp_pBs_25, gen_4_cmp_pBs_24, gen_4_cmp_pBs_23, 
         gen_4_cmp_pMux_30, gen_4_cmp_pMux_29, gen_4_cmp_pMux_28, 
         gen_4_cmp_pMux_27, gen_4_cmp_pMux_26, gen_4_cmp_pMux_25, 
         gen_4_cmp_pMux_24, gen_4_cmp_pMux_23, gen_4_cmp_pMux_22, 
         gen_4_cmp_pMux_21, gen_4_cmp_pMux_20, gen_4_cmp_pMux_19, 
         gen_4_cmp_pMux_18, gen_4_cmp_pMux_17, gen_4_cmp_pMux_16, 
         gen_4_cmp_pMux_15, gen_4_cmp_pMux_14, gen_4_cmp_pMux_13, 
         gen_4_cmp_pMux_12, gen_4_cmp_pMux_11, gen_4_cmp_pMux_10, 
         gen_4_cmp_pMux_9, gen_4_cmp_pMux_8, gen_4_cmp_pMux_7, gen_4_cmp_pMux_6, 
         gen_4_cmp_pMux_5, gen_4_cmp_pMux_4, gen_4_cmp_pMux_3, gen_4_cmp_pMux_2, 
         gen_4_cmp_pMux_1, gen_4_cmp_pMux_0, gen_4_cmp_pReg_30, 
         gen_4_cmp_pReg_29, gen_4_cmp_pReg_28, gen_4_cmp_pReg_27, 
         gen_4_cmp_pReg_26, gen_4_cmp_pReg_25, gen_4_cmp_pReg_24, 
         gen_4_cmp_pReg_23, gen_4_cmp_pReg_22, gen_4_cmp_pReg_21, 
         gen_4_cmp_pReg_20, gen_4_cmp_pReg_19, gen_4_cmp_pReg_18, 
         gen_4_cmp_pReg_17, gen_4_cmp_pReg_16, gen_4_cmp_pReg_15, 
         gen_4_cmp_pReg_14, gen_4_cmp_pReg_13, gen_4_cmp_pReg_12, 
         gen_4_cmp_pReg_11, gen_4_cmp_pReg_10, gen_4_cmp_pReg_9, 
         gen_4_cmp_pReg_8, gen_4_cmp_pReg_7, gen_4_cmp_pReg_6, gen_4_cmp_pReg_5, 
         gen_4_cmp_pReg_4, gen_4_cmp_pReg_3, gen_4_cmp_pReg_2, gen_4_cmp_pReg_1, 
         gen_4_cmp_pReg_0, gen_4_cmp_BSCmp_op2_0, gen_4_cmp_BSCmp_carryIn, 
         gen_3_cmp_pBs_30, gen_3_cmp_pBs_29, gen_3_cmp_pBs_28, gen_3_cmp_pBs_27, 
         gen_3_cmp_pBs_26, gen_3_cmp_pBs_25, gen_3_cmp_pBs_24, gen_3_cmp_pBs_23, 
         gen_3_cmp_pMux_30, gen_3_cmp_pMux_29, gen_3_cmp_pMux_28, 
         gen_3_cmp_pMux_27, gen_3_cmp_pMux_26, gen_3_cmp_pMux_25, 
         gen_3_cmp_pMux_24, gen_3_cmp_pMux_23, gen_3_cmp_pMux_22, 
         gen_3_cmp_pMux_21, gen_3_cmp_pMux_20, gen_3_cmp_pMux_19, 
         gen_3_cmp_pMux_18, gen_3_cmp_pMux_17, gen_3_cmp_pMux_16, 
         gen_3_cmp_pMux_15, gen_3_cmp_pMux_14, gen_3_cmp_pMux_13, 
         gen_3_cmp_pMux_12, gen_3_cmp_pMux_11, gen_3_cmp_pMux_10, 
         gen_3_cmp_pMux_9, gen_3_cmp_pMux_8, gen_3_cmp_pMux_7, gen_3_cmp_pMux_6, 
         gen_3_cmp_pMux_5, gen_3_cmp_pMux_4, gen_3_cmp_pMux_3, gen_3_cmp_pMux_2, 
         gen_3_cmp_pMux_1, gen_3_cmp_pMux_0, gen_3_cmp_pReg_30, 
         gen_3_cmp_pReg_29, gen_3_cmp_pReg_28, gen_3_cmp_pReg_27, 
         gen_3_cmp_pReg_26, gen_3_cmp_pReg_25, gen_3_cmp_pReg_24, 
         gen_3_cmp_pReg_23, gen_3_cmp_pReg_22, gen_3_cmp_pReg_21, 
         gen_3_cmp_pReg_20, gen_3_cmp_pReg_19, gen_3_cmp_pReg_18, 
         gen_3_cmp_pReg_17, gen_3_cmp_pReg_16, gen_3_cmp_pReg_15, 
         gen_3_cmp_pReg_14, gen_3_cmp_pReg_13, gen_3_cmp_pReg_12, 
         gen_3_cmp_pReg_11, gen_3_cmp_pReg_10, gen_3_cmp_pReg_9, 
         gen_3_cmp_pReg_8, gen_3_cmp_pReg_7, gen_3_cmp_pReg_6, gen_3_cmp_pReg_5, 
         gen_3_cmp_pReg_4, gen_3_cmp_pReg_3, gen_3_cmp_pReg_2, gen_3_cmp_pReg_1, 
         gen_3_cmp_pReg_0, gen_3_cmp_BSCmp_op2_0, gen_3_cmp_BSCmp_carryIn, 
         gen_2_cmp_pBs_30, gen_2_cmp_pBs_29, gen_2_cmp_pBs_28, gen_2_cmp_pBs_27, 
         gen_2_cmp_pBs_26, gen_2_cmp_pBs_25, gen_2_cmp_pBs_24, gen_2_cmp_pBs_23, 
         gen_2_cmp_pMux_30, gen_2_cmp_pMux_29, gen_2_cmp_pMux_28, 
         gen_2_cmp_pMux_27, gen_2_cmp_pMux_26, gen_2_cmp_pMux_25, 
         gen_2_cmp_pMux_24, gen_2_cmp_pMux_23, gen_2_cmp_pMux_22, 
         gen_2_cmp_pMux_21, gen_2_cmp_pMux_20, gen_2_cmp_pMux_19, 
         gen_2_cmp_pMux_18, gen_2_cmp_pMux_17, gen_2_cmp_pMux_16, 
         gen_2_cmp_pMux_15, gen_2_cmp_pMux_14, gen_2_cmp_pMux_13, 
         gen_2_cmp_pMux_12, gen_2_cmp_pMux_11, gen_2_cmp_pMux_10, 
         gen_2_cmp_pMux_9, gen_2_cmp_pMux_8, gen_2_cmp_pMux_7, gen_2_cmp_pMux_6, 
         gen_2_cmp_pMux_5, gen_2_cmp_pMux_4, gen_2_cmp_pMux_3, gen_2_cmp_pMux_2, 
         gen_2_cmp_pMux_1, gen_2_cmp_pMux_0, gen_2_cmp_pReg_30, 
         gen_2_cmp_pReg_29, gen_2_cmp_pReg_28, gen_2_cmp_pReg_27, 
         gen_2_cmp_pReg_26, gen_2_cmp_pReg_25, gen_2_cmp_pReg_24, 
         gen_2_cmp_pReg_23, gen_2_cmp_pReg_22, gen_2_cmp_pReg_21, 
         gen_2_cmp_pReg_20, gen_2_cmp_pReg_19, gen_2_cmp_pReg_18, 
         gen_2_cmp_pReg_17, gen_2_cmp_pReg_16, gen_2_cmp_pReg_15, 
         gen_2_cmp_pReg_14, gen_2_cmp_pReg_13, gen_2_cmp_pReg_12, 
         gen_2_cmp_pReg_11, gen_2_cmp_pReg_10, gen_2_cmp_pReg_9, 
         gen_2_cmp_pReg_8, gen_2_cmp_pReg_7, gen_2_cmp_pReg_6, gen_2_cmp_pReg_5, 
         gen_2_cmp_pReg_4, gen_2_cmp_pReg_3, gen_2_cmp_pReg_2, gen_2_cmp_pReg_1, 
         gen_2_cmp_pReg_0, gen_2_cmp_BSCmp_op2_0, gen_2_cmp_BSCmp_carryIn, 
         gen_1_cmp_pBs_30, gen_1_cmp_pBs_29, gen_1_cmp_pBs_28, gen_1_cmp_pBs_27, 
         gen_1_cmp_pBs_26, gen_1_cmp_pBs_25, gen_1_cmp_pBs_24, gen_1_cmp_pBs_23, 
         gen_1_cmp_pMux_30, gen_1_cmp_pMux_29, gen_1_cmp_pMux_28, 
         gen_1_cmp_pMux_27, gen_1_cmp_pMux_26, gen_1_cmp_pMux_25, 
         gen_1_cmp_pMux_24, gen_1_cmp_pMux_23, gen_1_cmp_pMux_22, 
         gen_1_cmp_pMux_21, gen_1_cmp_pMux_20, gen_1_cmp_pMux_19, 
         gen_1_cmp_pMux_18, gen_1_cmp_pMux_17, gen_1_cmp_pMux_16, 
         gen_1_cmp_pMux_15, gen_1_cmp_pMux_14, gen_1_cmp_pMux_13, 
         gen_1_cmp_pMux_12, gen_1_cmp_pMux_11, gen_1_cmp_pMux_10, 
         gen_1_cmp_pMux_9, gen_1_cmp_pMux_8, gen_1_cmp_pMux_7, gen_1_cmp_pMux_6, 
         gen_1_cmp_pMux_5, gen_1_cmp_pMux_4, gen_1_cmp_pMux_3, gen_1_cmp_pMux_2, 
         gen_1_cmp_pMux_1, gen_1_cmp_pMux_0, gen_1_cmp_pReg_30, 
         gen_1_cmp_pReg_29, gen_1_cmp_pReg_28, gen_1_cmp_pReg_27, 
         gen_1_cmp_pReg_26, gen_1_cmp_pReg_25, gen_1_cmp_pReg_24, 
         gen_1_cmp_pReg_23, gen_1_cmp_pReg_22, gen_1_cmp_pReg_21, 
         gen_1_cmp_pReg_20, gen_1_cmp_pReg_19, gen_1_cmp_pReg_18, 
         gen_1_cmp_pReg_17, gen_1_cmp_pReg_16, gen_1_cmp_pReg_15, 
         gen_1_cmp_pReg_14, gen_1_cmp_pReg_13, gen_1_cmp_pReg_12, 
         gen_1_cmp_pReg_11, gen_1_cmp_pReg_10, gen_1_cmp_pReg_9, 
         gen_1_cmp_pReg_8, gen_1_cmp_pReg_7, gen_1_cmp_pReg_6, gen_1_cmp_pReg_5, 
         gen_1_cmp_pReg_4, gen_1_cmp_pReg_3, gen_1_cmp_pReg_2, gen_1_cmp_pReg_1, 
         gen_1_cmp_pReg_0, gen_1_cmp_BSCmp_op2_0, gen_1_cmp_BSCmp_carryIn, 
         gen_0_cmp_pBs_30, gen_0_cmp_pBs_29, gen_0_cmp_pBs_28, gen_0_cmp_pBs_27, 
         gen_0_cmp_pBs_26, gen_0_cmp_pBs_25, gen_0_cmp_pBs_24, gen_0_cmp_pBs_23, 
         gen_0_cmp_pMux_30, gen_0_cmp_pMux_29, gen_0_cmp_pMux_28, 
         gen_0_cmp_pMux_27, gen_0_cmp_pMux_26, gen_0_cmp_pMux_25, 
         gen_0_cmp_pMux_24, gen_0_cmp_pMux_23, gen_0_cmp_pMux_22, 
         gen_0_cmp_pMux_21, gen_0_cmp_pMux_20, gen_0_cmp_pMux_19, 
         gen_0_cmp_pMux_18, gen_0_cmp_pMux_17, gen_0_cmp_pMux_16, 
         gen_0_cmp_pMux_15, gen_0_cmp_pMux_14, gen_0_cmp_pMux_13, 
         gen_0_cmp_pMux_12, gen_0_cmp_pMux_11, gen_0_cmp_pMux_10, 
         gen_0_cmp_pMux_9, gen_0_cmp_pMux_8, gen_0_cmp_pMux_7, gen_0_cmp_pMux_6, 
         gen_0_cmp_pMux_5, gen_0_cmp_pMux_4, gen_0_cmp_pMux_3, gen_0_cmp_pMux_2, 
         gen_0_cmp_pMux_1, gen_0_cmp_pMux_0, gen_0_cmp_pReg_30, 
         gen_0_cmp_pReg_29, gen_0_cmp_pReg_28, gen_0_cmp_pReg_27, 
         gen_0_cmp_pReg_26, gen_0_cmp_pReg_25, gen_0_cmp_pReg_24, 
         gen_0_cmp_pReg_23, gen_0_cmp_pReg_22, gen_0_cmp_pReg_21, 
         gen_0_cmp_pReg_20, gen_0_cmp_pReg_19, gen_0_cmp_pReg_18, 
         gen_0_cmp_pReg_17, gen_0_cmp_pReg_16, gen_0_cmp_pReg_15, 
         gen_0_cmp_pReg_14, gen_0_cmp_pReg_13, gen_0_cmp_pReg_12, 
         gen_0_cmp_pReg_11, gen_0_cmp_pReg_10, gen_0_cmp_pReg_9, 
         gen_0_cmp_pReg_8, gen_0_cmp_pReg_7, gen_0_cmp_pReg_6, gen_0_cmp_pReg_5, 
         gen_0_cmp_pReg_4, gen_0_cmp_pReg_3, gen_0_cmp_pReg_2, gen_0_cmp_pReg_1, 
         gen_0_cmp_pReg_0, gen_0_cmp_BSCmp_op2_0, gen_0_cmp_BSCmp_carryIn, 
         gen_24_cmp_BSCmp_op2_16, gen_24_cmp_BSCmp_op2_15, 
         gen_24_cmp_BSCmp_op2_14, gen_24_cmp_BSCmp_op2_13, 
         gen_24_cmp_BSCmp_op2_12, gen_24_cmp_BSCmp_op2_11, 
         gen_24_cmp_BSCmp_op2_10, gen_24_cmp_BSCmp_op2_9, gen_24_cmp_BSCmp_op2_8, 
         gen_24_cmp_BSCmp_op2_7, gen_24_cmp_BSCmp_op2_6, gen_24_cmp_BSCmp_op2_5, 
         gen_24_cmp_BSCmp_op2_4, gen_24_cmp_BSCmp_op2_3, gen_24_cmp_BSCmp_op2_2, 
         gen_24_cmp_BSCmp_op2_1, gen_23_cmp_BSCmp_op2_16, 
         gen_23_cmp_BSCmp_op2_15, gen_23_cmp_BSCmp_op2_14, 
         gen_23_cmp_BSCmp_op2_13, gen_23_cmp_BSCmp_op2_12, 
         gen_23_cmp_BSCmp_op2_11, gen_23_cmp_BSCmp_op2_10, 
         gen_23_cmp_BSCmp_op2_9, gen_23_cmp_BSCmp_op2_8, gen_23_cmp_BSCmp_op2_7, 
         gen_23_cmp_BSCmp_op2_6, gen_23_cmp_BSCmp_op2_5, gen_23_cmp_BSCmp_op2_4, 
         gen_23_cmp_BSCmp_op2_3, gen_23_cmp_BSCmp_op2_2, gen_23_cmp_BSCmp_op2_1, 
         gen_22_cmp_BSCmp_op2_16, gen_22_cmp_BSCmp_op2_15, 
         gen_22_cmp_BSCmp_op2_14, gen_22_cmp_BSCmp_op2_13, 
         gen_22_cmp_BSCmp_op2_12, gen_22_cmp_BSCmp_op2_11, 
         gen_22_cmp_BSCmp_op2_10, gen_22_cmp_BSCmp_op2_9, gen_22_cmp_BSCmp_op2_8, 
         gen_22_cmp_BSCmp_op2_7, gen_22_cmp_BSCmp_op2_6, gen_22_cmp_BSCmp_op2_5, 
         gen_22_cmp_BSCmp_op2_4, gen_22_cmp_BSCmp_op2_3, gen_22_cmp_BSCmp_op2_2, 
         gen_22_cmp_BSCmp_op2_1, gen_21_cmp_BSCmp_op2_16, 
         gen_21_cmp_BSCmp_op2_15, gen_21_cmp_BSCmp_op2_14, 
         gen_21_cmp_BSCmp_op2_13, gen_21_cmp_BSCmp_op2_12, 
         gen_21_cmp_BSCmp_op2_11, gen_21_cmp_BSCmp_op2_10, 
         gen_21_cmp_BSCmp_op2_9, gen_21_cmp_BSCmp_op2_8, gen_21_cmp_BSCmp_op2_7, 
         gen_21_cmp_BSCmp_op2_6, gen_21_cmp_BSCmp_op2_5, gen_21_cmp_BSCmp_op2_4, 
         gen_21_cmp_BSCmp_op2_3, gen_21_cmp_BSCmp_op2_2, gen_21_cmp_BSCmp_op2_1, 
         gen_20_cmp_BSCmp_op2_16, gen_20_cmp_BSCmp_op2_15, 
         gen_20_cmp_BSCmp_op2_14, gen_20_cmp_BSCmp_op2_13, 
         gen_20_cmp_BSCmp_op2_12, gen_20_cmp_BSCmp_op2_11, 
         gen_20_cmp_BSCmp_op2_10, gen_20_cmp_BSCmp_op2_9, gen_20_cmp_BSCmp_op2_8, 
         gen_20_cmp_BSCmp_op2_7, gen_20_cmp_BSCmp_op2_6, gen_20_cmp_BSCmp_op2_5, 
         gen_20_cmp_BSCmp_op2_4, gen_20_cmp_BSCmp_op2_3, gen_20_cmp_BSCmp_op2_2, 
         gen_20_cmp_BSCmp_op2_1, gen_19_cmp_BSCmp_op2_16, 
         gen_19_cmp_BSCmp_op2_15, gen_19_cmp_BSCmp_op2_14, 
         gen_19_cmp_BSCmp_op2_13, gen_19_cmp_BSCmp_op2_12, 
         gen_19_cmp_BSCmp_op2_11, gen_19_cmp_BSCmp_op2_10, 
         gen_19_cmp_BSCmp_op2_9, gen_19_cmp_BSCmp_op2_8, gen_19_cmp_BSCmp_op2_7, 
         gen_19_cmp_BSCmp_op2_6, gen_19_cmp_BSCmp_op2_5, gen_19_cmp_BSCmp_op2_4, 
         gen_19_cmp_BSCmp_op2_3, gen_19_cmp_BSCmp_op2_2, gen_19_cmp_BSCmp_op2_1, 
         gen_18_cmp_BSCmp_op2_16, gen_18_cmp_BSCmp_op2_15, 
         gen_18_cmp_BSCmp_op2_14, gen_18_cmp_BSCmp_op2_13, 
         gen_18_cmp_BSCmp_op2_12, gen_18_cmp_BSCmp_op2_11, 
         gen_18_cmp_BSCmp_op2_10, gen_18_cmp_BSCmp_op2_9, gen_18_cmp_BSCmp_op2_8, 
         gen_18_cmp_BSCmp_op2_7, gen_18_cmp_BSCmp_op2_6, gen_18_cmp_BSCmp_op2_5, 
         gen_18_cmp_BSCmp_op2_4, gen_18_cmp_BSCmp_op2_3, gen_18_cmp_BSCmp_op2_2, 
         gen_18_cmp_BSCmp_op2_1, gen_17_cmp_BSCmp_op2_16, 
         gen_17_cmp_BSCmp_op2_15, gen_17_cmp_BSCmp_op2_14, 
         gen_17_cmp_BSCmp_op2_13, gen_17_cmp_BSCmp_op2_12, 
         gen_17_cmp_BSCmp_op2_11, gen_17_cmp_BSCmp_op2_10, 
         gen_17_cmp_BSCmp_op2_9, gen_17_cmp_BSCmp_op2_8, gen_17_cmp_BSCmp_op2_7, 
         gen_17_cmp_BSCmp_op2_6, gen_17_cmp_BSCmp_op2_5, gen_17_cmp_BSCmp_op2_4, 
         gen_17_cmp_BSCmp_op2_3, gen_17_cmp_BSCmp_op2_2, gen_17_cmp_BSCmp_op2_1, 
         gen_16_cmp_BSCmp_op2_16, gen_16_cmp_BSCmp_op2_15, 
         gen_16_cmp_BSCmp_op2_14, gen_16_cmp_BSCmp_op2_13, 
         gen_16_cmp_BSCmp_op2_12, gen_16_cmp_BSCmp_op2_11, 
         gen_16_cmp_BSCmp_op2_10, gen_16_cmp_BSCmp_op2_9, gen_16_cmp_BSCmp_op2_8, 
         gen_16_cmp_BSCmp_op2_7, gen_16_cmp_BSCmp_op2_6, gen_16_cmp_BSCmp_op2_5, 
         gen_16_cmp_BSCmp_op2_4, gen_16_cmp_BSCmp_op2_3, gen_16_cmp_BSCmp_op2_2, 
         gen_16_cmp_BSCmp_op2_1, gen_15_cmp_BSCmp_op2_16, 
         gen_15_cmp_BSCmp_op2_15, gen_15_cmp_BSCmp_op2_14, 
         gen_15_cmp_BSCmp_op2_13, gen_15_cmp_BSCmp_op2_12, 
         gen_15_cmp_BSCmp_op2_11, gen_15_cmp_BSCmp_op2_10, 
         gen_15_cmp_BSCmp_op2_9, gen_15_cmp_BSCmp_op2_8, gen_15_cmp_BSCmp_op2_7, 
         gen_15_cmp_BSCmp_op2_6, gen_15_cmp_BSCmp_op2_5, gen_15_cmp_BSCmp_op2_4, 
         gen_15_cmp_BSCmp_op2_3, gen_15_cmp_BSCmp_op2_2, gen_15_cmp_BSCmp_op2_1, 
         gen_14_cmp_BSCmp_op2_16, gen_14_cmp_BSCmp_op2_15, 
         gen_14_cmp_BSCmp_op2_14, gen_14_cmp_BSCmp_op2_13, 
         gen_14_cmp_BSCmp_op2_12, gen_14_cmp_BSCmp_op2_11, 
         gen_14_cmp_BSCmp_op2_10, gen_14_cmp_BSCmp_op2_9, gen_14_cmp_BSCmp_op2_8, 
         gen_14_cmp_BSCmp_op2_7, gen_14_cmp_BSCmp_op2_6, gen_14_cmp_BSCmp_op2_5, 
         gen_14_cmp_BSCmp_op2_4, gen_14_cmp_BSCmp_op2_3, gen_14_cmp_BSCmp_op2_2, 
         gen_14_cmp_BSCmp_op2_1, gen_13_cmp_BSCmp_op2_16, 
         gen_13_cmp_BSCmp_op2_15, gen_13_cmp_BSCmp_op2_14, 
         gen_13_cmp_BSCmp_op2_13, gen_13_cmp_BSCmp_op2_12, 
         gen_13_cmp_BSCmp_op2_11, gen_13_cmp_BSCmp_op2_10, 
         gen_13_cmp_BSCmp_op2_9, gen_13_cmp_BSCmp_op2_8, gen_13_cmp_BSCmp_op2_7, 
         gen_13_cmp_BSCmp_op2_6, gen_13_cmp_BSCmp_op2_5, gen_13_cmp_BSCmp_op2_4, 
         gen_13_cmp_BSCmp_op2_3, gen_13_cmp_BSCmp_op2_2, gen_13_cmp_BSCmp_op2_1, 
         gen_12_cmp_BSCmp_op2_16, gen_12_cmp_BSCmp_op2_15, 
         gen_12_cmp_BSCmp_op2_14, gen_12_cmp_BSCmp_op2_13, 
         gen_12_cmp_BSCmp_op2_12, gen_12_cmp_BSCmp_op2_11, 
         gen_12_cmp_BSCmp_op2_10, gen_12_cmp_BSCmp_op2_9, gen_12_cmp_BSCmp_op2_8, 
         gen_12_cmp_BSCmp_op2_7, gen_12_cmp_BSCmp_op2_6, gen_12_cmp_BSCmp_op2_5, 
         gen_12_cmp_BSCmp_op2_4, gen_12_cmp_BSCmp_op2_3, gen_12_cmp_BSCmp_op2_2, 
         gen_12_cmp_BSCmp_op2_1, gen_11_cmp_BSCmp_op2_16, 
         gen_11_cmp_BSCmp_op2_15, gen_11_cmp_BSCmp_op2_14, 
         gen_11_cmp_BSCmp_op2_13, gen_11_cmp_BSCmp_op2_12, 
         gen_11_cmp_BSCmp_op2_11, gen_11_cmp_BSCmp_op2_10, 
         gen_11_cmp_BSCmp_op2_9, gen_11_cmp_BSCmp_op2_8, gen_11_cmp_BSCmp_op2_7, 
         gen_11_cmp_BSCmp_op2_6, gen_11_cmp_BSCmp_op2_5, gen_11_cmp_BSCmp_op2_4, 
         gen_11_cmp_BSCmp_op2_3, gen_11_cmp_BSCmp_op2_2, gen_11_cmp_BSCmp_op2_1, 
         gen_10_cmp_BSCmp_op2_16, gen_10_cmp_BSCmp_op2_15, 
         gen_10_cmp_BSCmp_op2_14, gen_10_cmp_BSCmp_op2_13, 
         gen_10_cmp_BSCmp_op2_12, gen_10_cmp_BSCmp_op2_11, 
         gen_10_cmp_BSCmp_op2_10, gen_10_cmp_BSCmp_op2_9, gen_10_cmp_BSCmp_op2_8, 
         gen_10_cmp_BSCmp_op2_7, gen_10_cmp_BSCmp_op2_6, gen_10_cmp_BSCmp_op2_5, 
         gen_10_cmp_BSCmp_op2_4, gen_10_cmp_BSCmp_op2_3, gen_10_cmp_BSCmp_op2_2, 
         gen_10_cmp_BSCmp_op2_1, gen_9_cmp_BSCmp_op2_16, gen_9_cmp_BSCmp_op2_15, 
         gen_9_cmp_BSCmp_op2_14, gen_9_cmp_BSCmp_op2_13, gen_9_cmp_BSCmp_op2_12, 
         gen_9_cmp_BSCmp_op2_11, gen_9_cmp_BSCmp_op2_10, gen_9_cmp_BSCmp_op2_9, 
         gen_9_cmp_BSCmp_op2_8, gen_9_cmp_BSCmp_op2_7, gen_9_cmp_BSCmp_op2_6, 
         gen_9_cmp_BSCmp_op2_5, gen_9_cmp_BSCmp_op2_4, gen_9_cmp_BSCmp_op2_3, 
         gen_9_cmp_BSCmp_op2_2, gen_9_cmp_BSCmp_op2_1, gen_8_cmp_BSCmp_op2_16, 
         gen_8_cmp_BSCmp_op2_15, gen_8_cmp_BSCmp_op2_14, gen_8_cmp_BSCmp_op2_13, 
         gen_8_cmp_BSCmp_op2_12, gen_8_cmp_BSCmp_op2_11, gen_8_cmp_BSCmp_op2_10, 
         gen_8_cmp_BSCmp_op2_9, gen_8_cmp_BSCmp_op2_8, gen_8_cmp_BSCmp_op2_7, 
         gen_8_cmp_BSCmp_op2_6, gen_8_cmp_BSCmp_op2_5, gen_8_cmp_BSCmp_op2_4, 
         gen_8_cmp_BSCmp_op2_3, gen_8_cmp_BSCmp_op2_2, gen_8_cmp_BSCmp_op2_1, 
         gen_7_cmp_BSCmp_op2_16, gen_7_cmp_BSCmp_op2_15, gen_7_cmp_BSCmp_op2_14, 
         gen_7_cmp_BSCmp_op2_13, gen_7_cmp_BSCmp_op2_12, gen_7_cmp_BSCmp_op2_11, 
         gen_7_cmp_BSCmp_op2_10, gen_7_cmp_BSCmp_op2_9, gen_7_cmp_BSCmp_op2_8, 
         gen_7_cmp_BSCmp_op2_7, gen_7_cmp_BSCmp_op2_6, gen_7_cmp_BSCmp_op2_5, 
         gen_7_cmp_BSCmp_op2_4, gen_7_cmp_BSCmp_op2_3, gen_7_cmp_BSCmp_op2_2, 
         gen_7_cmp_BSCmp_op2_1, gen_6_cmp_BSCmp_op2_16, gen_6_cmp_BSCmp_op2_15, 
         gen_6_cmp_BSCmp_op2_14, gen_6_cmp_BSCmp_op2_13, gen_6_cmp_BSCmp_op2_12, 
         gen_6_cmp_BSCmp_op2_11, gen_6_cmp_BSCmp_op2_10, gen_6_cmp_BSCmp_op2_9, 
         gen_6_cmp_BSCmp_op2_8, gen_6_cmp_BSCmp_op2_7, gen_6_cmp_BSCmp_op2_6, 
         gen_6_cmp_BSCmp_op2_5, gen_6_cmp_BSCmp_op2_4, gen_6_cmp_BSCmp_op2_3, 
         gen_6_cmp_BSCmp_op2_2, gen_6_cmp_BSCmp_op2_1, gen_5_cmp_BSCmp_op2_16, 
         gen_5_cmp_BSCmp_op2_15, gen_5_cmp_BSCmp_op2_14, gen_5_cmp_BSCmp_op2_13, 
         gen_5_cmp_BSCmp_op2_12, gen_5_cmp_BSCmp_op2_11, gen_5_cmp_BSCmp_op2_10, 
         gen_5_cmp_BSCmp_op2_9, gen_5_cmp_BSCmp_op2_8, gen_5_cmp_BSCmp_op2_7, 
         gen_5_cmp_BSCmp_op2_6, gen_5_cmp_BSCmp_op2_5, gen_5_cmp_BSCmp_op2_4, 
         gen_5_cmp_BSCmp_op2_3, gen_5_cmp_BSCmp_op2_2, gen_5_cmp_BSCmp_op2_1, 
         gen_4_cmp_BSCmp_op2_16, gen_4_cmp_BSCmp_op2_15, gen_4_cmp_BSCmp_op2_14, 
         gen_4_cmp_BSCmp_op2_13, gen_4_cmp_BSCmp_op2_12, gen_4_cmp_BSCmp_op2_11, 
         gen_4_cmp_BSCmp_op2_10, gen_4_cmp_BSCmp_op2_9, gen_4_cmp_BSCmp_op2_8, 
         gen_4_cmp_BSCmp_op2_7, gen_4_cmp_BSCmp_op2_6, gen_4_cmp_BSCmp_op2_5, 
         gen_4_cmp_BSCmp_op2_4, gen_4_cmp_BSCmp_op2_3, gen_4_cmp_BSCmp_op2_2, 
         gen_4_cmp_BSCmp_op2_1, gen_3_cmp_BSCmp_op2_16, gen_3_cmp_BSCmp_op2_15, 
         gen_3_cmp_BSCmp_op2_14, gen_3_cmp_BSCmp_op2_13, gen_3_cmp_BSCmp_op2_12, 
         gen_3_cmp_BSCmp_op2_11, gen_3_cmp_BSCmp_op2_10, gen_3_cmp_BSCmp_op2_9, 
         gen_3_cmp_BSCmp_op2_8, gen_3_cmp_BSCmp_op2_7, gen_3_cmp_BSCmp_op2_6, 
         gen_3_cmp_BSCmp_op2_5, gen_3_cmp_BSCmp_op2_4, gen_3_cmp_BSCmp_op2_3, 
         gen_3_cmp_BSCmp_op2_2, gen_3_cmp_BSCmp_op2_1, gen_2_cmp_BSCmp_op2_16, 
         gen_2_cmp_BSCmp_op2_15, gen_2_cmp_BSCmp_op2_14, gen_2_cmp_BSCmp_op2_13, 
         gen_2_cmp_BSCmp_op2_12, gen_2_cmp_BSCmp_op2_11, gen_2_cmp_BSCmp_op2_10, 
         gen_2_cmp_BSCmp_op2_9, gen_2_cmp_BSCmp_op2_8, gen_2_cmp_BSCmp_op2_7, 
         gen_2_cmp_BSCmp_op2_6, gen_2_cmp_BSCmp_op2_5, gen_2_cmp_BSCmp_op2_4, 
         gen_2_cmp_BSCmp_op2_3, gen_2_cmp_BSCmp_op2_2, gen_2_cmp_BSCmp_op2_1, 
         gen_1_cmp_BSCmp_op2_16, gen_1_cmp_BSCmp_op2_15, gen_1_cmp_BSCmp_op2_14, 
         gen_1_cmp_BSCmp_op2_13, gen_1_cmp_BSCmp_op2_12, gen_1_cmp_BSCmp_op2_11, 
         gen_1_cmp_BSCmp_op2_10, gen_1_cmp_BSCmp_op2_9, gen_1_cmp_BSCmp_op2_8, 
         gen_1_cmp_BSCmp_op2_7, gen_1_cmp_BSCmp_op2_6, gen_1_cmp_BSCmp_op2_5, 
         gen_1_cmp_BSCmp_op2_4, gen_1_cmp_BSCmp_op2_3, gen_1_cmp_BSCmp_op2_2, 
         gen_1_cmp_BSCmp_op2_1, gen_0_cmp_BSCmp_op2_16, gen_0_cmp_BSCmp_op2_15, 
         gen_0_cmp_BSCmp_op2_14, gen_0_cmp_BSCmp_op2_13, gen_0_cmp_BSCmp_op2_12, 
         gen_0_cmp_BSCmp_op2_11, gen_0_cmp_BSCmp_op2_10, gen_0_cmp_BSCmp_op2_9, 
         gen_0_cmp_BSCmp_op2_8, gen_0_cmp_BSCmp_op2_7, gen_0_cmp_BSCmp_op2_6, 
         gen_0_cmp_BSCmp_op2_5, gen_0_cmp_BSCmp_op2_4, gen_0_cmp_BSCmp_op2_3, 
         gen_0_cmp_BSCmp_op2_2, gen_0_cmp_BSCmp_op2_1, gen_24_cmp_pInit_32, nx6, 
         gen_0_cmp_mReg_0, nx26, nx34, gen_0_cmp_mReg_1, nx46, nx48, nx58, nx62, 
         gen_0_cmp_mReg_2, nx74, nx76, nx80, nx84, gen_0_cmp_mReg_3, nx96, nx98, 
         nx102, nx106, gen_0_cmp_mReg_4, nx118, nx120, nx124, nx128, 
         gen_0_cmp_mReg_5, nx140, nx142, nx146, nx150, gen_0_cmp_mReg_6, nx162, 
         nx164, nx168, nx172, gen_0_cmp_mReg_7, nx184, nx186, nx190, nx194, 
         gen_0_cmp_mReg_8, nx206, nx208, nx212, nx216, gen_0_cmp_mReg_9, nx228, 
         nx230, nx234, nx238, gen_0_cmp_mReg_10, nx250, nx252, nx256, nx260, 
         gen_0_cmp_mReg_11, nx272, nx274, nx278, nx282, gen_0_cmp_mReg_12, nx294, 
         nx296, nx300, nx304, gen_0_cmp_mReg_13, nx316, nx318, nx322, nx326, 
         gen_0_cmp_mReg_14, nx338, nx340, nx344, nx348, gen_0_cmp_mReg_15, nx360, 
         nx362, nx366, nx370, nx376, nx380, nx392, gen_1_cmp_mReg_0, nx412, 
         nx420, gen_1_cmp_mReg_1, nx432, nx434, nx444, nx448, gen_1_cmp_mReg_2, 
         nx460, nx462, nx466, nx470, gen_1_cmp_mReg_3, nx482, nx484, nx488, 
         nx492, gen_1_cmp_mReg_4, nx504, nx506, nx510, nx514, gen_1_cmp_mReg_5, 
         nx526, nx528, nx532, nx536, gen_1_cmp_mReg_6, nx548, nx550, nx554, 
         nx558, gen_1_cmp_mReg_7, nx570, nx572, nx576, nx580, gen_1_cmp_mReg_8, 
         nx592, nx594, nx598, nx602, gen_1_cmp_mReg_9, nx614, nx616, nx620, 
         nx624, gen_1_cmp_mReg_10, nx636, nx638, nx642, nx646, gen_1_cmp_mReg_11, 
         nx658, nx660, nx664, nx668, gen_1_cmp_mReg_12, nx680, nx682, nx686, 
         nx690, gen_1_cmp_mReg_13, nx702, nx704, nx708, nx712, gen_1_cmp_mReg_14, 
         nx724, nx726, nx730, nx734, gen_1_cmp_mReg_15, nx746, nx748, nx752, 
         nx756, nx762, nx766, nx778, gen_2_cmp_mReg_0, nx798, nx806, 
         gen_2_cmp_mReg_1, nx818, nx820, nx830, nx834, gen_2_cmp_mReg_2, nx846, 
         nx848, nx852, nx856, gen_2_cmp_mReg_3, nx868, nx870, nx874, nx878, 
         gen_2_cmp_mReg_4, nx890, nx892, nx896, nx900, gen_2_cmp_mReg_5, nx912, 
         nx914, nx918, nx922, gen_2_cmp_mReg_6, nx934, nx936, nx940, nx944, 
         gen_2_cmp_mReg_7, nx956, nx958, nx962, nx966, gen_2_cmp_mReg_8, nx978, 
         nx980, nx984, nx988, gen_2_cmp_mReg_9, nx1000, nx1002, nx1006, nx1010, 
         gen_2_cmp_mReg_10, nx1022, nx1024, nx1028, nx1032, gen_2_cmp_mReg_11, 
         nx1044, nx1046, nx1050, nx1054, gen_2_cmp_mReg_12, nx1066, nx1068, 
         nx1072, nx1076, gen_2_cmp_mReg_13, nx1088, nx1090, nx1094, nx1098, 
         gen_2_cmp_mReg_14, nx1110, nx1112, nx1116, nx1120, gen_2_cmp_mReg_15, 
         nx1132, nx1134, nx1138, nx1142, nx1148, nx1152, nx1164, 
         gen_3_cmp_mReg_0, nx1184, nx1192, gen_3_cmp_mReg_1, nx1204, nx1206, 
         nx1216, nx1220, gen_3_cmp_mReg_2, nx1232, nx1234, nx1238, nx1242, 
         gen_3_cmp_mReg_3, nx1254, nx1256, nx1260, nx1264, gen_3_cmp_mReg_4, 
         nx1276, nx1278, nx1282, nx1286, gen_3_cmp_mReg_5, nx1298, nx1300, 
         nx1304, nx1308, gen_3_cmp_mReg_6, nx1320, nx1322, nx1326, nx1330, 
         gen_3_cmp_mReg_7, nx1342, nx1344, nx1348, nx1352, gen_3_cmp_mReg_8, 
         nx1364, nx1366, nx1370, nx1374, gen_3_cmp_mReg_9, nx1386, nx1388, 
         nx1392, nx1396, gen_3_cmp_mReg_10, nx1408, nx1410, nx1414, nx1418, 
         gen_3_cmp_mReg_11, nx1430, nx1432, nx1436, nx1440, gen_3_cmp_mReg_12, 
         nx1452, nx1454, nx1458, nx1462, gen_3_cmp_mReg_13, nx1474, nx1476, 
         nx1480, nx1484, gen_3_cmp_mReg_14, nx1496, nx1498, nx1502, nx1506, 
         gen_3_cmp_mReg_15, nx1518, nx1520, nx1524, nx1528, nx1534, nx1538, 
         nx1550, gen_4_cmp_mReg_0, nx1570, nx1578, gen_4_cmp_mReg_1, nx1590, 
         nx1592, nx1602, nx1606, gen_4_cmp_mReg_2, nx1618, nx1620, nx1624, 
         nx1628, gen_4_cmp_mReg_3, nx1640, nx1642, nx1646, nx1650, 
         gen_4_cmp_mReg_4, nx1662, nx1664, nx1668, nx1672, gen_4_cmp_mReg_5, 
         nx1684, nx1686, nx1690, nx1694, gen_4_cmp_mReg_6, nx1706, nx1708, 
         nx1712, nx1716, gen_4_cmp_mReg_7, nx1728, nx1730, nx1734, nx1738, 
         gen_4_cmp_mReg_8, nx1750, nx1752, nx1756, nx1760, gen_4_cmp_mReg_9, 
         nx1772, nx1774, nx1778, nx1782, gen_4_cmp_mReg_10, nx1794, nx1796, 
         nx1800, nx1804, gen_4_cmp_mReg_11, nx1816, nx1818, nx1822, nx1826, 
         gen_4_cmp_mReg_12, nx1838, nx1840, nx1844, nx1848, gen_4_cmp_mReg_13, 
         nx1860, nx1862, nx1866, nx1870, gen_4_cmp_mReg_14, nx1882, nx1884, 
         nx1888, nx1892, gen_4_cmp_mReg_15, nx1904, nx1906, nx1910, nx1914, 
         nx1920, nx1924, nx1936, gen_5_cmp_mReg_0, nx1956, nx1964, 
         gen_5_cmp_mReg_1, nx1976, nx1978, nx1988, nx1992, gen_5_cmp_mReg_2, 
         nx2004, nx2006, nx2010, nx2014, gen_5_cmp_mReg_3, nx2026, nx2028, 
         nx2032, nx2036, gen_5_cmp_mReg_4, nx2048, nx2050, nx2054, nx2058, 
         gen_5_cmp_mReg_5, nx2070, nx2072, nx2076, nx2080, gen_5_cmp_mReg_6, 
         nx2092, nx2094, nx2098, nx2102, gen_5_cmp_mReg_7, nx2114, nx2116, 
         nx2120, nx2124, gen_5_cmp_mReg_8, nx2136, nx2138, nx2142, nx2146, 
         gen_5_cmp_mReg_9, nx2158, nx2160, nx2164, nx2168, gen_5_cmp_mReg_10, 
         nx2180, nx2182, nx2186, nx2190, gen_5_cmp_mReg_11, nx2202, nx2204, 
         nx2208, nx2212, gen_5_cmp_mReg_12, nx2224, nx2226, nx2230, nx2234, 
         gen_5_cmp_mReg_13, nx2246, nx2248, nx2252, nx2256, gen_5_cmp_mReg_14, 
         nx2268, nx2270, nx2274, nx2278, gen_5_cmp_mReg_15, nx2290, nx2292, 
         nx2296, nx2300, nx2306, nx2310, nx2322, gen_6_cmp_mReg_0, nx2342, 
         nx2350, gen_6_cmp_mReg_1, nx2362, nx2364, nx2374, nx2378, 
         gen_6_cmp_mReg_2, nx2390, nx2392, nx2396, nx2400, gen_6_cmp_mReg_3, 
         nx2412, nx2414, nx2418, nx2422, gen_6_cmp_mReg_4, nx2434, nx2436, 
         nx2440, nx2444, gen_6_cmp_mReg_5, nx2456, nx2458, nx2462, nx2466, 
         gen_6_cmp_mReg_6, nx2478, nx2480, nx2484, nx2488, gen_6_cmp_mReg_7, 
         nx2500, nx2502, nx2506, nx2510, gen_6_cmp_mReg_8, nx2522, nx2524, 
         nx2528, nx2532, gen_6_cmp_mReg_9, nx2544, nx2546, nx2550, nx2554, 
         gen_6_cmp_mReg_10, nx2566, nx2568, nx2572, nx2576, gen_6_cmp_mReg_11, 
         nx2588, nx2590, nx2594, nx2598, gen_6_cmp_mReg_12, nx2610, nx2612, 
         nx2616, nx2620, gen_6_cmp_mReg_13, nx2632, nx2634, nx2638, nx2642, 
         gen_6_cmp_mReg_14, nx2654, nx2656, nx2660, nx2664, gen_6_cmp_mReg_15, 
         nx2676, nx2678, nx2682, nx2686, nx2692, nx2696, nx2708, 
         gen_7_cmp_mReg_0, nx2728, nx2736, gen_7_cmp_mReg_1, nx2748, nx2750, 
         nx2760, nx2764, gen_7_cmp_mReg_2, nx2776, nx2778, nx2782, nx2786, 
         gen_7_cmp_mReg_3, nx2798, nx2800, nx2804, nx2808, gen_7_cmp_mReg_4, 
         nx2820, nx2822, nx2826, nx2830, gen_7_cmp_mReg_5, nx2842, nx2844, 
         nx2848, nx2852, gen_7_cmp_mReg_6, nx2864, nx2866, nx2870, nx2874, 
         gen_7_cmp_mReg_7, nx2886, nx2888, nx2892, nx2896, gen_7_cmp_mReg_8, 
         nx2908, nx2910, nx2914, nx2918, gen_7_cmp_mReg_9, nx2930, nx2932, 
         nx2936, nx2940, gen_7_cmp_mReg_10, nx2952, nx2954, nx2958, nx2962, 
         gen_7_cmp_mReg_11, nx2974, nx2976, nx2980, nx2984, gen_7_cmp_mReg_12, 
         nx2996, nx2998, nx3002, nx3006, gen_7_cmp_mReg_13, nx3018, nx3020, 
         nx3024, nx3028, gen_7_cmp_mReg_14, nx3040, nx3042, nx3046, nx3050, 
         gen_7_cmp_mReg_15, nx3062, nx3064, nx3068, nx3072, nx3078, nx3082, 
         nx3094, gen_8_cmp_mReg_0, nx3114, nx3122, gen_8_cmp_mReg_1, nx3134, 
         nx3136, nx3146, nx3150, gen_8_cmp_mReg_2, nx3162, nx3164, nx3168, 
         nx3172, gen_8_cmp_mReg_3, nx3184, nx3186, nx3190, nx3194, 
         gen_8_cmp_mReg_4, nx3206, nx3208, nx3212, nx3216, gen_8_cmp_mReg_5, 
         nx3228, nx3230, nx3234, nx3238, gen_8_cmp_mReg_6, nx3250, nx3252, 
         nx3256, nx3260, gen_8_cmp_mReg_7, nx3272, nx3274, nx3278, nx3282, 
         gen_8_cmp_mReg_8, nx3294, nx3296, nx3300, nx3304, gen_8_cmp_mReg_9, 
         nx3316, nx3318, nx3322, nx3326, gen_8_cmp_mReg_10, nx3338, nx3340, 
         nx3344, nx3348, gen_8_cmp_mReg_11, nx3360, nx3362, nx3366, nx3370, 
         gen_8_cmp_mReg_12, nx3382, nx3384, nx3388, nx3392, gen_8_cmp_mReg_13, 
         nx3404, nx3406, nx3410, nx3414, gen_8_cmp_mReg_14, nx3426, nx3428, 
         nx3432, nx3436, gen_8_cmp_mReg_15, nx3448, nx3450, nx3454, nx3458, 
         nx3464, nx3468, nx3480, gen_9_cmp_mReg_0, nx3500, nx3508, 
         gen_9_cmp_mReg_1, nx3520, nx3522, nx3532, nx3536, gen_9_cmp_mReg_2, 
         nx3548, nx3550, nx3554, nx3558, gen_9_cmp_mReg_3, nx3570, nx3572, 
         nx3576, nx3580, gen_9_cmp_mReg_4, nx3592, nx3594, nx3598, nx3602, 
         gen_9_cmp_mReg_5, nx3614, nx3616, nx3620, nx3624, gen_9_cmp_mReg_6, 
         nx3636, nx3638, nx3642, nx3646, gen_9_cmp_mReg_7, nx3658, nx3660, 
         nx3664, nx3668, gen_9_cmp_mReg_8, nx3680, nx3682, nx3686, nx3690, 
         gen_9_cmp_mReg_9, nx3702, nx3704, nx3708, nx3712, gen_9_cmp_mReg_10, 
         nx3724, nx3726, nx3730, nx3734, gen_9_cmp_mReg_11, nx3746, nx3748, 
         nx3752, nx3756, gen_9_cmp_mReg_12, nx3768, nx3770, nx3774, nx3778, 
         gen_9_cmp_mReg_13, nx3790, nx3792, nx3796, nx3800, gen_9_cmp_mReg_14, 
         nx3812, nx3814, nx3818, nx3822, gen_9_cmp_mReg_15, nx3834, nx3836, 
         nx3840, nx3844, nx3850, nx3854, nx3866, gen_10_cmp_mReg_0, nx3886, 
         nx3894, gen_10_cmp_mReg_1, nx3906, nx3908, nx3918, nx3922, 
         gen_10_cmp_mReg_2, nx3934, nx3936, nx3940, nx3944, gen_10_cmp_mReg_3, 
         nx3956, nx3958, nx3962, nx3966, gen_10_cmp_mReg_4, nx3978, nx3980, 
         nx3984, nx3988, gen_10_cmp_mReg_5, nx4000, nx4002, nx4006, nx4010, 
         gen_10_cmp_mReg_6, nx4022, nx4024, nx4028, nx4032, gen_10_cmp_mReg_7, 
         nx4044, nx4046, nx4050, nx4054, gen_10_cmp_mReg_8, nx4066, nx4068, 
         nx4072, nx4076, gen_10_cmp_mReg_9, nx4088, nx4090, nx4094, nx4098, 
         gen_10_cmp_mReg_10, nx4110, nx4112, nx4116, nx4120, gen_10_cmp_mReg_11, 
         nx4132, nx4134, nx4138, nx4142, gen_10_cmp_mReg_12, nx4154, nx4156, 
         nx4160, nx4164, gen_10_cmp_mReg_13, nx4176, nx4178, nx4182, nx4186, 
         gen_10_cmp_mReg_14, nx4198, nx4200, nx4204, nx4208, gen_10_cmp_mReg_15, 
         nx4220, nx4222, nx4226, nx4230, nx4236, nx4240, nx4252, 
         gen_11_cmp_mReg_0, nx4272, nx4280, gen_11_cmp_mReg_1, nx4292, nx4294, 
         nx4304, nx4308, gen_11_cmp_mReg_2, nx4320, nx4322, nx4326, nx4330, 
         gen_11_cmp_mReg_3, nx4342, nx4344, nx4348, nx4352, gen_11_cmp_mReg_4, 
         nx4364, nx4366, nx4370, nx4374, gen_11_cmp_mReg_5, nx4386, nx4388, 
         nx4392, nx4396, gen_11_cmp_mReg_6, nx4408, nx4410, nx4414, nx4418, 
         gen_11_cmp_mReg_7, nx4430, nx4432, nx4436, nx4440, gen_11_cmp_mReg_8, 
         nx4452, nx4454, nx4458, nx4462, gen_11_cmp_mReg_9, nx4474, nx4476, 
         nx4480, nx4484, gen_11_cmp_mReg_10, nx4496, nx4498, nx4502, nx4506, 
         gen_11_cmp_mReg_11, nx4518, nx4520, nx4524, nx4528, gen_11_cmp_mReg_12, 
         nx4540, nx4542, nx4546, nx4550, gen_11_cmp_mReg_13, nx4562, nx4564, 
         nx4568, nx4572, gen_11_cmp_mReg_14, nx4584, nx4586, nx4590, nx4594, 
         gen_11_cmp_mReg_15, nx4606, nx4608, nx4612, nx4616, nx4622, nx4626, 
         nx4638, gen_12_cmp_mReg_0, nx4658, nx4666, gen_12_cmp_mReg_1, nx4678, 
         nx4680, nx4690, nx4694, gen_12_cmp_mReg_2, nx4706, nx4708, nx4712, 
         nx4716, gen_12_cmp_mReg_3, nx4728, nx4730, nx4734, nx4738, 
         gen_12_cmp_mReg_4, nx4750, nx4752, nx4756, nx4760, gen_12_cmp_mReg_5, 
         nx4772, nx4774, nx4778, nx4782, gen_12_cmp_mReg_6, nx4794, nx4796, 
         nx4800, nx4804, gen_12_cmp_mReg_7, nx4816, nx4818, nx4822, nx4826, 
         gen_12_cmp_mReg_8, nx4838, nx4840, nx4844, nx4848, gen_12_cmp_mReg_9, 
         nx4860, nx4862, nx4866, nx4870, gen_12_cmp_mReg_10, nx4882, nx4884, 
         nx4888, nx4892, gen_12_cmp_mReg_11, nx4904, nx4906, nx4910, nx4914, 
         gen_12_cmp_mReg_12, nx4926, nx4928, nx4932, nx4936, gen_12_cmp_mReg_13, 
         nx4948, nx4950, nx4954, nx4958, gen_12_cmp_mReg_14, nx4970, nx4972, 
         nx4976, nx4980, gen_12_cmp_mReg_15, nx4992, nx4994, nx4998, nx5002, 
         nx5008, nx5012, nx5024, gen_13_cmp_mReg_0, nx5044, nx5052, 
         gen_13_cmp_mReg_1, nx5064, nx5066, nx5076, nx5080, gen_13_cmp_mReg_2, 
         nx5092, nx5094, nx5098, nx5102, gen_13_cmp_mReg_3, nx5114, nx5116, 
         nx5120, nx5124, gen_13_cmp_mReg_4, nx5136, nx5138, nx5142, nx5146, 
         gen_13_cmp_mReg_5, nx5158, nx5160, nx5164, nx5168, gen_13_cmp_mReg_6, 
         nx5180, nx5182, nx5186, nx5190, gen_13_cmp_mReg_7, nx5202, nx5204, 
         nx5208, nx5212, gen_13_cmp_mReg_8, nx5224, nx5226, nx5230, nx5234, 
         gen_13_cmp_mReg_9, nx5246, nx5248, nx5252, nx5256, gen_13_cmp_mReg_10, 
         nx5268, nx5270, nx5274, nx5278, gen_13_cmp_mReg_11, nx5290, nx5292, 
         nx5296, nx5300, gen_13_cmp_mReg_12, nx5312, nx5314, nx5318, nx5322, 
         gen_13_cmp_mReg_13, nx5334, nx5336, nx5340, nx5344, gen_13_cmp_mReg_14, 
         nx5356, nx5358, nx5362, nx5366, gen_13_cmp_mReg_15, nx5378, nx5380, 
         nx5384, nx5388, nx5394, nx5398, nx5410, gen_14_cmp_mReg_0, nx5430, 
         nx5438, gen_14_cmp_mReg_1, nx5450, nx5452, nx5462, nx5466, 
         gen_14_cmp_mReg_2, nx5478, nx5480, nx5484, nx5488, gen_14_cmp_mReg_3, 
         nx5500, nx5502, nx5506, nx5510, gen_14_cmp_mReg_4, nx5522, nx5524, 
         nx5528, nx5532, gen_14_cmp_mReg_5, nx5544, nx5546, nx5550, nx5554, 
         gen_14_cmp_mReg_6, nx5566, nx5568, nx5572, nx5576, gen_14_cmp_mReg_7, 
         nx5588, nx5590, nx5594, nx5598, gen_14_cmp_mReg_8, nx5610, nx5612, 
         nx5616, nx5620, gen_14_cmp_mReg_9, nx5632, nx5634, nx5638, nx5642, 
         gen_14_cmp_mReg_10, nx5654, nx5656, nx5660, nx5664, gen_14_cmp_mReg_11, 
         nx5676, nx5678, nx5682, nx5686, gen_14_cmp_mReg_12, nx5698, nx5700, 
         nx5704, nx5708, gen_14_cmp_mReg_13, nx5720, nx5722, nx5726, nx5730, 
         gen_14_cmp_mReg_14, nx5742, nx5744, nx5748, nx5752, gen_14_cmp_mReg_15, 
         nx5764, nx5766, nx5770, nx5774, nx5780, nx5784, nx5796, 
         gen_15_cmp_mReg_0, nx5816, nx5824, gen_15_cmp_mReg_1, nx5836, nx5838, 
         nx5848, nx5852, gen_15_cmp_mReg_2, nx5864, nx5866, nx5870, nx5874, 
         gen_15_cmp_mReg_3, nx5886, nx5888, nx5892, nx5896, gen_15_cmp_mReg_4, 
         nx5908, nx5910, nx5914, nx5918, gen_15_cmp_mReg_5, nx5930, nx5932, 
         nx5936, nx5940, gen_15_cmp_mReg_6, nx5952, nx5954, nx5958, nx5962, 
         gen_15_cmp_mReg_7, nx5974, nx5976, nx5980, nx5984, gen_15_cmp_mReg_8, 
         nx5996, nx5998, nx6002, nx6006, gen_15_cmp_mReg_9, nx6018, nx6020, 
         nx6024, nx6028, gen_15_cmp_mReg_10, nx6040, nx6042, nx6046, nx6050, 
         gen_15_cmp_mReg_11, nx6062, nx6064, nx6068, nx6072, gen_15_cmp_mReg_12, 
         nx6084, nx6086, nx6090, nx6094, gen_15_cmp_mReg_13, nx6106, nx6108, 
         nx6112, nx6116, gen_15_cmp_mReg_14, nx6128, nx6130, nx6134, nx6138, 
         gen_15_cmp_mReg_15, nx6150, nx6152, nx6156, nx6160, nx6166, nx6170, 
         nx6182, gen_16_cmp_mReg_0, nx6202, nx6210, gen_16_cmp_mReg_1, nx6222, 
         nx6224, nx6234, nx6238, gen_16_cmp_mReg_2, nx6250, nx6252, nx6256, 
         nx6260, gen_16_cmp_mReg_3, nx6272, nx6274, nx6278, nx6282, 
         gen_16_cmp_mReg_4, nx6294, nx6296, nx6300, nx6304, gen_16_cmp_mReg_5, 
         nx6316, nx6318, nx6322, nx6326, gen_16_cmp_mReg_6, nx6338, nx6340, 
         nx6344, nx6348, gen_16_cmp_mReg_7, nx6360, nx6362, nx6366, nx6370, 
         gen_16_cmp_mReg_8, nx6382, nx6384, nx6388, nx6392, gen_16_cmp_mReg_9, 
         nx6404, nx6406, nx6410, nx6414, gen_16_cmp_mReg_10, nx6426, nx6428, 
         nx6432, nx6436, gen_16_cmp_mReg_11, nx6448, nx6450, nx6454, nx6458, 
         gen_16_cmp_mReg_12, nx6470, nx6472, nx6476, nx6480, gen_16_cmp_mReg_13, 
         nx6492, nx6494, nx6498, nx6502, gen_16_cmp_mReg_14, nx6514, nx6516, 
         nx6520, nx6524, gen_16_cmp_mReg_15, nx6536, nx6538, nx6542, nx6546, 
         nx6552, nx6556, nx6568, gen_17_cmp_mReg_0, nx6588, nx6596, 
         gen_17_cmp_mReg_1, nx6608, nx6610, nx6620, nx6624, gen_17_cmp_mReg_2, 
         nx6636, nx6638, nx6642, nx6646, gen_17_cmp_mReg_3, nx6658, nx6660, 
         nx6664, nx6668, gen_17_cmp_mReg_4, nx6680, nx6682, nx6686, nx6690, 
         gen_17_cmp_mReg_5, nx6702, nx6704, nx6708, nx6712, gen_17_cmp_mReg_6, 
         nx6724, nx6726, nx6730, nx6734, gen_17_cmp_mReg_7, nx6746, nx6748, 
         nx6752, nx6756, gen_17_cmp_mReg_8, nx6768, nx6770, nx6774, nx6778, 
         gen_17_cmp_mReg_9, nx6790, nx6792, nx6796, nx6800, gen_17_cmp_mReg_10, 
         nx6812, nx6814, nx6818, nx6822, gen_17_cmp_mReg_11, nx6834, nx6836, 
         nx6840, nx6844, gen_17_cmp_mReg_12, nx6856, nx6858, nx6862, nx6866, 
         gen_17_cmp_mReg_13, nx6878, nx6880, nx6884, nx6888, gen_17_cmp_mReg_14, 
         nx6900, nx6902, nx6906, nx6910, gen_17_cmp_mReg_15, nx6922, nx6924, 
         nx6928, nx6932, nx6938, nx6942, nx6954, gen_18_cmp_mReg_0, nx6974, 
         nx6982, gen_18_cmp_mReg_1, nx6994, nx6996, nx7006, nx7010, 
         gen_18_cmp_mReg_2, nx7022, nx7024, nx7028, nx7032, gen_18_cmp_mReg_3, 
         nx7044, nx7046, nx7050, nx7054, gen_18_cmp_mReg_4, nx7066, nx7068, 
         nx7072, nx7076, gen_18_cmp_mReg_5, nx7088, nx7090, nx7094, nx7098, 
         gen_18_cmp_mReg_6, nx7110, nx7112, nx7116, nx7120, gen_18_cmp_mReg_7, 
         nx7132, nx7134, nx7138, nx7142, gen_18_cmp_mReg_8, nx7154, nx7156, 
         nx7160, nx7164, gen_18_cmp_mReg_9, nx7176, nx7178, nx7182, nx7186, 
         gen_18_cmp_mReg_10, nx7198, nx7200, nx7204, nx7208, gen_18_cmp_mReg_11, 
         nx7220, nx7222, nx7226, nx7230, gen_18_cmp_mReg_12, nx7242, nx7244, 
         nx7248, nx7252, gen_18_cmp_mReg_13, nx7264, nx7266, nx7270, nx7274, 
         gen_18_cmp_mReg_14, nx7286, nx7288, nx7292, nx7296, gen_18_cmp_mReg_15, 
         nx7308, nx7310, nx7314, nx7318, nx7324, nx7328, nx7340, 
         gen_19_cmp_mReg_0, nx7360, nx7368, gen_19_cmp_mReg_1, nx7380, nx7382, 
         nx7392, nx7396, gen_19_cmp_mReg_2, nx7408, nx7410, nx7414, nx7418, 
         gen_19_cmp_mReg_3, nx7430, nx7432, nx7436, nx7440, gen_19_cmp_mReg_4, 
         nx7452, nx7454, nx7458, nx7462, gen_19_cmp_mReg_5, nx7474, nx7476, 
         nx7480, nx7484, gen_19_cmp_mReg_6, nx7496, nx7498, nx7502, nx7506, 
         gen_19_cmp_mReg_7, nx7518, nx7520, nx7524, nx7528, gen_19_cmp_mReg_8, 
         nx7540, nx7542, nx7546, nx7550, gen_19_cmp_mReg_9, nx7562, nx7564, 
         nx7568, nx7572, gen_19_cmp_mReg_10, nx7584, nx7586, nx7590, nx7594, 
         gen_19_cmp_mReg_11, nx7606, nx7608, nx7612, nx7616, gen_19_cmp_mReg_12, 
         nx7628, nx7630, nx7634, nx7638, gen_19_cmp_mReg_13, nx7650, nx7652, 
         nx7656, nx7660, gen_19_cmp_mReg_14, nx7672, nx7674, nx7678, nx7682, 
         gen_19_cmp_mReg_15, nx7694, nx7696, nx7700, nx7704, nx7710, nx7714, 
         nx7726, gen_20_cmp_mReg_0, nx7746, nx7754, gen_20_cmp_mReg_1, nx7766, 
         nx7768, nx7778, nx7782, gen_20_cmp_mReg_2, nx7794, nx7796, nx7800, 
         nx7804, gen_20_cmp_mReg_3, nx7816, nx7818, nx7822, nx7826, 
         gen_20_cmp_mReg_4, nx7838, nx7840, nx7844, nx7848, gen_20_cmp_mReg_5, 
         nx7860, nx7862, nx7866, nx7870, gen_20_cmp_mReg_6, nx7882, nx7884, 
         nx7888, nx7892, gen_20_cmp_mReg_7, nx7904, nx7906, nx7910, nx7914, 
         gen_20_cmp_mReg_8, nx7926, nx7928, nx7932, nx7936, gen_20_cmp_mReg_9, 
         nx7948, nx7950, nx7954, nx7958, gen_20_cmp_mReg_10, nx7970, nx7972, 
         nx7976, nx7980, gen_20_cmp_mReg_11, nx7992, nx7994, nx7998, nx8002, 
         gen_20_cmp_mReg_12, nx8014, nx8016, nx8020, nx8024, gen_20_cmp_mReg_13, 
         nx8036, nx8038, nx8042, nx8046, gen_20_cmp_mReg_14, nx8058, nx8060, 
         nx8064, nx8068, gen_20_cmp_mReg_15, nx8080, nx8082, nx8086, nx8090, 
         nx8096, nx8100, nx8112, gen_21_cmp_mReg_0, nx8132, nx8140, 
         gen_21_cmp_mReg_1, nx8152, nx8154, nx8164, nx8168, gen_21_cmp_mReg_2, 
         nx8180, nx8182, nx8186, nx8190, gen_21_cmp_mReg_3, nx8202, nx8204, 
         nx8208, nx8212, gen_21_cmp_mReg_4, nx8224, nx8226, nx8230, nx8234, 
         gen_21_cmp_mReg_5, nx8246, nx8248, nx8252, nx8256, gen_21_cmp_mReg_6, 
         nx8268, nx8270, nx8274, nx8278, gen_21_cmp_mReg_7, nx8290, nx8292, 
         nx8296, nx8300, gen_21_cmp_mReg_8, nx8312, nx8314, nx8318, nx8322, 
         gen_21_cmp_mReg_9, nx8334, nx8336, nx8340, nx8344, gen_21_cmp_mReg_10, 
         nx8356, nx8358, nx8362, nx8366, gen_21_cmp_mReg_11, nx8378, nx8380, 
         nx8384, nx8388, gen_21_cmp_mReg_12, nx8400, nx8402, nx8406, nx8410, 
         gen_21_cmp_mReg_13, nx8422, nx8424, nx8428, nx8432, gen_21_cmp_mReg_14, 
         nx8444, nx8446, nx8450, nx8454, gen_21_cmp_mReg_15, nx8466, nx8468, 
         nx8472, nx8476, nx8482, nx8486, nx8498, gen_22_cmp_mReg_0, nx8518, 
         nx8526, gen_22_cmp_mReg_1, nx8538, nx8540, nx8550, nx8554, 
         gen_22_cmp_mReg_2, nx8566, nx8568, nx8572, nx8576, gen_22_cmp_mReg_3, 
         nx8588, nx8590, nx8594, nx8598, gen_22_cmp_mReg_4, nx8610, nx8612, 
         nx8616, nx8620, gen_22_cmp_mReg_5, nx8632, nx8634, nx8638, nx8642, 
         gen_22_cmp_mReg_6, nx8654, nx8656, nx8660, nx8664, gen_22_cmp_mReg_7, 
         nx8676, nx8678, nx8682, nx8686, gen_22_cmp_mReg_8, nx8698, nx8700, 
         nx8704, nx8708, gen_22_cmp_mReg_9, nx8720, nx8722, nx8726, nx8730, 
         gen_22_cmp_mReg_10, nx8742, nx8744, nx8748, nx8752, gen_22_cmp_mReg_11, 
         nx8764, nx8766, nx8770, nx8774, gen_22_cmp_mReg_12, nx8786, nx8788, 
         nx8792, nx8796, gen_22_cmp_mReg_13, nx8808, nx8810, nx8814, nx8818, 
         gen_22_cmp_mReg_14, nx8830, nx8832, nx8836, nx8840, gen_22_cmp_mReg_15, 
         nx8852, nx8854, nx8858, nx8862, nx8868, nx8872, nx8884, 
         gen_23_cmp_mReg_0, nx8904, nx8912, gen_23_cmp_mReg_1, nx8924, nx8926, 
         nx8936, nx8940, gen_23_cmp_mReg_2, nx8952, nx8954, nx8958, nx8962, 
         gen_23_cmp_mReg_3, nx8974, nx8976, nx8980, nx8984, gen_23_cmp_mReg_4, 
         nx8996, nx8998, nx9002, nx9006, gen_23_cmp_mReg_5, nx9018, nx9020, 
         nx9024, nx9028, gen_23_cmp_mReg_6, nx9040, nx9042, nx9046, nx9050, 
         gen_23_cmp_mReg_7, nx9062, nx9064, nx9068, nx9072, gen_23_cmp_mReg_8, 
         nx9084, nx9086, nx9090, nx9094, gen_23_cmp_mReg_9, nx9106, nx9108, 
         nx9112, nx9116, gen_23_cmp_mReg_10, nx9128, nx9130, nx9134, nx9138, 
         gen_23_cmp_mReg_11, nx9150, nx9152, nx9156, nx9160, gen_23_cmp_mReg_12, 
         nx9172, nx9174, nx9178, nx9182, gen_23_cmp_mReg_13, nx9194, nx9196, 
         nx9200, nx9204, gen_23_cmp_mReg_14, nx9216, nx9218, nx9222, nx9226, 
         gen_23_cmp_mReg_15, nx9238, nx9240, nx9244, nx9248, nx9254, nx9258, 
         nx9270, gen_24_cmp_mReg_0, nx9290, nx9298, gen_24_cmp_mReg_1, nx9310, 
         nx9312, nx9322, nx9326, gen_24_cmp_mReg_2, nx9338, nx9340, nx9344, 
         nx9348, gen_24_cmp_mReg_3, nx9360, nx9362, nx9366, nx9370, 
         gen_24_cmp_mReg_4, nx9382, nx9384, nx9388, nx9392, gen_24_cmp_mReg_5, 
         nx9404, nx9406, nx9410, nx9414, gen_24_cmp_mReg_6, nx9426, nx9428, 
         nx9432, nx9436, gen_24_cmp_mReg_7, nx9448, nx9450, nx9454, nx9458, 
         gen_24_cmp_mReg_8, nx9470, nx9472, nx9476, nx9480, gen_24_cmp_mReg_9, 
         nx9492, nx9494, nx9498, nx9502, gen_24_cmp_mReg_10, nx9514, nx9516, 
         nx9520, nx9524, gen_24_cmp_mReg_11, nx9536, nx9538, nx9542, nx9546, 
         gen_24_cmp_mReg_12, nx9558, nx9560, nx9564, nx9568, gen_24_cmp_mReg_13, 
         nx9580, nx9582, nx9586, nx9590, gen_24_cmp_mReg_14, nx9602, nx9604, 
         nx9608, nx9612, gen_24_cmp_mReg_15, nx9624, nx9626, nx9630, nx9634, 
         nx9640, nx9644, CounterCmp_outp_1, restartDetection, nx9650, 
         StartCaptuerCmp_d, nx9660, nx9666, nx3671, nx3681, nx3691, nx3697, 
         nx3713, nx3720, nx3729, nx3733, nx3737, nx3741, nx3745, nx3751, nx3757, 
         nx3761, nx3769, nx3771, nx3775, nx3786, nx3791, nx3795, nx3801, nx3807, 
         nx3810, nx3817, nx3823, nx3827, nx3831, nx3837, nx3841, nx3845, nx3851, 
         nx3855, nx3861, nx3867, nx3870, nx3874, nx3879, nx3883, nx3889, nx3895, 
         nx3899, nx3903, nx3909, nx3913, nx3919, nx3923, nx3927, nx3931, nx3937, 
         nx3941, nx3945, nx3951, nx3954, nx3961, nx3967, nx3971, nx3975, nx3981, 
         nx3985, nx3989, nx3996, nx4001, nx4005, nx4013, nx4015, nx4018, nx4031, 
         nx4037, nx4040, nx4045, nx4051, nx4055, nx4061, nx4065, nx4069, nx4075, 
         nx4081, nx4084, nx4089, nx4095, nx4099, nx4105, nx4109, nx4113, nx4119, 
         nx4125, nx4128, nx4133, nx4139, nx4143, nx4149, nx4153, nx4157, nx4163, 
         nx4169, nx4172, nx4177, nx4183, nx4187, nx4193, nx4197, nx4201, nx4207, 
         nx4213, nx4216, nx4221, nx4227, nx4231, nx4237, nx4243, nx4249, nx4253, 
         nx4260, nx4263, nx4267, nx4279, nx4285, nx4288, nx4293, nx4299, nx4303, 
         nx4309, nx4315, nx4318, nx4325, nx4331, nx4335, nx4339, nx4345, nx4349, 
         nx4353, nx4359, nx4362, nx4369, nx4375, nx4379, nx4383, nx4389, nx4393, 
         nx4397, nx4403, nx4406, nx4413, nx4419, nx4423, nx4427, nx4433, nx4437, 
         nx4441, nx4447, nx4450, nx4457, nx4463, nx4467, nx4471, nx4477, nx4481, 
         nx4485, nx4492, nx4497, nx4501, nx4509, nx4511, nx4514, nx4527, nx4533, 
         nx4536, nx4541, nx4547, nx4551, nx4557, nx4561, nx4565, nx4571, nx4577, 
         nx4580, nx4585, nx4591, nx4595, nx4601, nx4605, nx4609, nx4615, nx4621, 
         nx4625, nx4631, nx4637, nx4641, nx4645, nx4649, nx4653, nx4659, nx4665, 
         nx4669, nx4674, nx4679, nx4683, nx4687, nx4693, nx4697, nx4702, nx4707, 
         nx4711, nx4717, nx4723, nx4726, nx4733, nx4739, nx4745, nx4748, nx4757, 
         nx4759, nx4763, nx4773, nx4779, nx4783, nx4789, nx4793, nx4797, nx4803, 
         nx4809, nx4812, nx4817, nx4823, nx4827, nx4833, nx4837, nx4841, nx4847, 
         nx4853, nx4856, nx4861, nx4867, nx4871, nx4877, nx4881, nx4885, nx4891, 
         nx4897, nx4900, nx4905, nx4911, nx4915, nx4921, nx4925, nx4929, nx4935, 
         nx4941, nx4944, nx4949, nx4955, nx4959, nx4965, nx4969, nx4973, nx4979, 
         nx4987, nx4991, nx4995, nx5003, nx5005, nx5009, nx5021, nx5027, nx5030, 
         nx5035, nx5041, nx5045, nx5051, nx5057, nx5060, nx5065, nx5071, nx5075, 
         nx5081, nx5087, nx5090, nx5097, nx5103, nx5107, nx5111, nx5117, nx5121, 
         nx5125, nx5131, nx5134, nx5141, nx5147, nx5151, nx5155, nx5161, nx5165, 
         nx5169, nx5175, nx5178, nx5185, nx5191, nx5195, nx5199, nx5205, nx5209, 
         nx5213, nx5219, nx5222, nx5229, nx5235, nx5241, nx5244, nx5253, nx5255, 
         nx5259, nx5269, nx5275, nx5279, nx5285, nx5289, nx5293, nx5299, nx5305, 
         nx5308, nx5313, nx5319, nx5323, nx5329, nx5333, nx5337, nx5343, nx5349, 
         nx5352, nx5357, nx5363, nx5367, nx5373, nx5377, nx5381, nx5387, nx5393, 
         nx5397, nx5403, nx5409, nx5413, nx5417, nx5421, nx5425, nx5431, nx5437, 
         nx5441, nx5446, nx5451, nx5455, nx5459, nx5465, nx5469, nx5474, nx5481, 
         nx5487, nx5491, nx5499, nx5501, nx5505, nx5515, nx5519, nx5523, nx5529, 
         nx5533, nx5537, nx5541, nx5547, nx5551, nx5555, nx5561, nx5564, nx5571, 
         nx5577, nx5581, nx5585, nx5591, nx5595, nx5599, nx5605, nx5608, nx5615, 
         nx5621, nx5625, nx5629, nx5635, nx5639, nx5643, nx5649, nx5652, nx5659, 
         nx5665, nx5669, nx5673, nx5679, nx5683, nx5687, nx5693, nx5696, nx5703, 
         nx5709, nx5713, nx5717, nx5725, nx5731, nx5735, nx5743, nx5745, nx5749, 
         nx5760, nx5765, nx5769, nx5775, nx5781, nx5785, nx5791, nx5797, nx5800, 
         nx5804, nx5809, nx5813, nx5819, nx5825, nx5829, nx5833, nx5839, nx5843, 
         nx5849, nx5853, nx5857, nx5861, nx5867, nx5871, nx5875, nx5881, nx5884, 
         nx5891, nx5897, nx5901, nx5905, nx5911, nx5915, nx5919, nx5925, nx5928, 
         nx5935, nx5941, nx5945, nx5949, nx5955, nx5959, nx5963, nx5970, nx5975, 
         nx5979, nx5987, nx5989, nx5992, nx6005, nx6011, nx6014, nx6019, nx6025, 
         nx6029, nx6035, nx6039, nx6043, nx6049, nx6055, nx6058, nx6063, nx6069, 
         nx6073, nx6079, nx6083, nx6087, nx6093, nx6099, nx6102, nx6107, nx6113, 
         nx6117, nx6123, nx6127, nx6131, nx6137, nx6143, nx6146, nx6151, nx6157, 
         nx6161, nx6167, nx6171, nx6175, nx6181, nx6186, nx6189, nx6193, nx6199, 
         nx6203, nx6209, nx6217, nx6221, nx6225, nx6233, nx6235, nx6239, nx6249, 
         nx6255, nx6259, nx6265, nx6269, nx6273, nx6279, nx6283, nx6287, nx6291, 
         nx6297, nx6301, nx6305, nx6311, nx6314, nx6321, nx6327, nx6331, nx6335, 
         nx6341, nx6345, nx6349, nx6355, nx6358, nx6365, nx6371, nx6375, nx6379, 
         nx6385, nx6389, nx6393, nx6399, nx6402, nx6409, nx6415, nx6419, nx6423, 
         nx6429, nx6433, nx6437, nx6443, nx6446, nx6453, nx6459, nx6465, nx6468, 
         nx6477, nx6479, nx6483, nx6493, nx6499, nx6503, nx6509, nx6513, nx6517, 
         nx6523, nx6529, nx6532, nx6537, nx6543, nx6547, nx6553, nx6557, nx6561, 
         nx6567, nx6572, nx6575, nx6579, nx6585, nx6589, nx6595, nx6601, nx6604, 
         nx6609, nx6615, nx6619, nx6625, nx6631, nx6634, nx6641, nx6647, nx6651, 
         nx6655, nx6661, nx6665, nx6669, nx6675, nx6678, nx6685, nx6691, nx6695, 
         nx6699, nx6707, nx6713, nx6717, nx6725, nx6727, nx6731, nx6742, nx6747, 
         nx6751, nx6757, nx6763, nx6766, nx6773, nx6779, nx6783, nx6787, nx6793, 
         nx6797, nx6801, nx6807, nx6810, nx6817, nx6823, nx6827, nx6831, nx6837, 
         nx6841, nx6845, nx6851, nx6854, nx6861, nx6867, nx6871, nx6875, nx6881, 
         nx6885, nx6889, nx6895, nx6898, nx6905, nx6911, nx6915, nx6919, nx6925, 
         nx6929, nx6933, nx6939, nx6943, nx6949, nx6957, nx6961, nx6965, nx6973, 
         nx6975, nx6979, nx6990, nx6995, nx6999, nx7003, nx7009, nx7013, nx7018, 
         nx7023, nx7027, nx7033, nx7039, nx7042, nx7049, nx7055, nx7059, nx7063, 
         nx7069, nx7073, nx7077, nx7083, nx7086, nx7093, nx7099, nx7103, nx7107, 
         nx7113, nx7117, nx7121, nx7127, nx7130, nx7137, nx7143, nx7147, nx7151, 
         nx7157, nx7161, nx7165, nx7171, nx7174, nx7181, nx7187, nx7191, nx7195, 
         nx7203, nx7209, nx7213, nx7221, nx7223, nx7227, nx7238, nx7243, nx7247, 
         nx7253, nx7259, nx7262, nx7269, nx7275, nx7279, nx7283, nx7289, nx7293, 
         nx7297, nx7303, nx7306, nx7313, nx7319, nx7323, nx7329, nx7335, nx7339, 
         nx7344, nx7348, nx7351, nx7357, nx7363, nx7367, nx7373, nx7377, nx7381, 
         nx7387, nx7393, nx7397, nx7403, nx7407, nx7411, nx7417, nx7423, nx7426, 
         nx7431, nx7437, nx7441, nx7447, nx7453, nx7459, nx7463, nx7471, nx7473, 
         nx7477, nx7489, nx7493, nx7497, nx7503, nx7507, nx7511, nx7515, nx7521, 
         nx7525, nx7529, nx7535, nx7538, nx7545, nx7551, nx7555, nx7559, nx7565, 
         nx7569, nx7573, nx7579, nx7582, nx7589, nx7595, nx7599, nx7603, nx7609, 
         nx7613, nx7617, nx7623, nx7626, nx7633, nx7639, nx7643, nx7647, nx7653, 
         nx7657, nx7661, nx7667, nx7670, nx7677, nx7683, nx7687, nx7691, nx7699, 
         nx7705, nx7709, nx7717, nx7719, nx7723, nx7733, nx7737, nx7741, nx7747, 
         nx7753, nx7757, nx7762, nx7767, nx7771, nx7775, nx7781, nx7785, nx7790, 
         nx7795, nx7799, nx7805, nx7811, nx7814, nx7821, nx7827, nx7831, nx7835, 
         nx7841, nx7845, nx7849, nx7855, nx7858, nx7865, nx7871, nx7875, nx7879, 
         nx7885, nx7889, nx7893, nx7899, nx7902, nx7909, nx7915, nx7919, nx7923, 
         nx7929, nx7933, nx7937, nx7944, nx7949, nx7953, nx7961, nx7963, nx7966, 
         nx7979, nx7985, nx7988, nx7993, nx7999, nx8003, nx8009, nx8013, nx8017, 
         nx8023, nx8029, nx8032, nx8037, nx8043, nx8047, nx8053, nx8057, nx8061, 
         nx8067, nx8073, nx8076, nx8081, nx8087, nx8091, nx8097, nx8101, nx8105, 
         nx8111, nx8116, nx8119, nx8123, nx8129, nx8133, nx8139, nx8145, nx8148, 
         nx8153, nx8159, nx8163, nx8169, nx8175, nx8178, nx8185, nx8191, nx8197, 
         nx8200, nx8209, nx8211, nx8215, nx8225, nx8231, nx8235, nx8241, nx8245, 
         nx8249, nx8255, nx8261, nx8264, nx8269, nx8275, nx8279, nx8285, nx8289, 
         nx8293, nx8299, nx8305, nx8308, nx8313, nx8319, nx8323, nx8329, nx8333, 
         nx8337, nx8343, nx8349, nx8352, nx8357, nx8363, nx8367, nx8373, nx8377, 
         nx8381, nx8387, nx8393, nx8396, nx8401, nx8407, nx8411, nx8417, nx8421, 
         nx8425, nx8431, nx8439, nx8443, nx8447, nx8455, nx8457, nx8461, nx8473, 
         nx8477, nx8481, nx8487, nx8493, nx8497, nx8502, nx8506, nx8509, nx8515, 
         nx8521, nx8525, nx8531, nx8535, nx8539, nx8545, nx8551, nx8555, nx8561, 
         nx8565, nx8569, nx8575, nx8581, nx8584, nx8589, nx8595, nx8599, nx8605, 
         nx8609, nx8613, nx8619, nx8625, nx8628, nx8633, nx8639, nx8643, nx8649, 
         nx8653, nx8657, nx8663, nx8669, nx8672, nx8677, nx8685, nx8691, nx8694, 
         nx8701, nx8703, nx8707, nx8718, nx8725, nx8729, nx8735, nx8739, nx8743, 
         nx8749, nx8753, nx8757, nx8761, nx8767, nx8771, nx8775, nx8781, nx8784, 
         nx8791, nx8797, nx8801, nx8805, nx8811, nx8815, nx8819, nx8825, nx8828, 
         nx8835, nx8841, nx8845, nx8849, nx8855, nx8859, nx8863, nx8869, nx8873, 
         nx8879, nx8885, nx8888, nx8892, nx8897, nx8901, nx8907, nx8913, nx8917, 
         nx8921, nx8929, nx8933, nx8937, nx8945, nx8947, nx8950, nx8963, nx8969, 
         nx8972, nx8979, nx8985, nx8989, nx8993, nx8999, nx9003, nx9007, nx9013, 
         nx9016, nx9023, nx9029, nx9033, nx9037, nx9043, nx9047, nx9051, nx9057, 
         nx9060, nx9067, nx9073, nx9077, nx9081, nx9087, nx9091, nx9095, nx9101, 
         nx9104, nx9111, nx9117, nx9121, nx9125, nx9131, nx9135, nx9139, nx9145, 
         nx9148, nx9155, nx9161, nx9165, nx9169, nx9177, nx9183, nx9187, nx9195, 
         nx9197, nx9201, nx9212, nx9217, nx9221, nx9227, nx9233, nx9236, nx9243, 
         nx9249, nx9253, nx9259, nx9265, nx9269, nx9274, nx9278, nx9281, nx9287, 
         nx9293, nx9297, nx9303, nx9307, nx9311, nx9317, nx9323, nx9327, nx9333, 
         nx9337, nx9341, nx9347, nx9353, nx9356, nx9361, nx9367, nx9371, nx9377, 
         nx9381, nx9385, nx9391, nx9397, nx9400, nx9405, nx9411, nx9415, nx9421, 
         nx9427, nx9433, nx9437, nx9445, nx9447, nx9451, nx9463, nx9467, nx9471, 
         nx9477, nx9481, nx9485, nx9489, nx9495, nx9499, nx9503, nx9509, nx9512, 
         nx9519, nx9525, nx9529, nx9533, nx9539, nx9543, nx9547, nx9553, nx9556, 
         nx9563, nx9569, nx9573, nx9577, nx9583, nx9587, nx9591, nx9597, nx9600, 
         nx9607, nx9613, nx9617, nx9621, nx9627, nx9631, nx9635, nx9641, nx9645, 
         nx9651, nx9655, nx9658, nx9663, nx9669, nx9673, nx9676, nx9683, nx9685, 
         nx9688, nx9698, nx9702, nx9705, nx9709, nx9713, nx9716, nx9720, nx9724, 
         nx9727, nx9731, nx9735, nx9738, nx9742, nx9746, nx9749, nx9753, nx9757, 
         nx9760, nx9764, nx9768, nx9771, nx9775, nx9779, nx9782, nx9786, nx9790, 
         nx9793, nx9797, nx9801, nx9804, nx9808, nx9812, nx9815, nx9819, nx9823, 
         nx9826, nx9830, nx9834, nx9837, nx9841, nx9845, nx9848, nx9852, nx9857, 
         nx9860, nx9864, nx9867, nx9870, nx9874, nx9877, nx9880, nx9884, nx9887, 
         nx9890, nx9894, nx9897, nx9900, nx9904, nx9907, nx9910, nx9914, nx9917, 
         nx9920, nx9924, nx9927, nx9930, nx9934, nx9937, nx9940, nx9944, nx9947, 
         nx9950, nx9954, nx9957, nx9960, nx9964, nx9967, nx9970, nx9974, nx9977, 
         nx9980, nx9984, nx9987, nx9990, nx9994, nx9997, nx10000, nx10004, 
         nx10007, nx10010, nx10014, nx10017, nx10020, nx10024, nx10027, nx10030, 
         nx10034, nx10037, nx10040, nx10044, nx10047, nx10050, nx10054, nx10057, 
         nx10060, nx10064, nx10067, nx10070, nx10074, nx10077, nx10080, nx10084, 
         nx10087, nx10090, nx10094, nx10097, nx10100, nx10104, nx10107, nx10120, 
         nx10122, nx10124, nx10126, nx10128, nx10130, nx10132, nx10134, nx10136, 
         nx10138, nx10140, nx10142, nx10144, nx10146, nx10148, nx10150, nx10152, 
         nx10154, nx10156, nx10158, nx10160, nx10162, nx10164, nx10166, nx10168, 
         nx10170, nx10172, nx10174, nx10176, nx10178, nx10180, nx10182, nx10184, 
         nx10186, nx10188, nx10190, nx10192, nx10194, nx10196, nx10198, nx10200, 
         nx10202, nx10204, nx10206, nx10208, nx10210, nx10212, nx10214, nx10216, 
         nx10218, nx10220, nx10222, nx10224, nx10226, nx10228, nx10230, nx10232, 
         nx10234, nx10236, nx10238, nx10240, nx10242, nx10244, nx10246, nx10248, 
         nx10250, nx10252, nx10254, nx10256, nx10258, nx10260, nx10262, nx10264, 
         nx10266, nx10268, nx10270, nx10272, nx10274, nx10276, nx10278, nx10280, 
         nx10282, nx10284, nx10286, nx10288, nx10290, nx10292, nx10294, nx10296, 
         nx10298, nx10300, nx10302, nx10304, nx10306, nx10308, nx10310, nx10312, 
         nx10314, nx10316, nx10318, nx10320, nx10322, nx10324, nx10326, nx10328, 
         nx10330, nx10332, nx10334, nx10336, nx10338, nx10340, nx10342, nx10344, 
         nx10346, nx10348, nx10350, nx10352, nx10354, nx10356, nx10358, nx10360, 
         nx10362, nx10364, nx10366, nx10368, nx10370, nx10372, nx10374, nx10376, 
         nx10378, nx10380, nx10382, nx10384, nx10386, nx10388, nx10390, nx10392, 
         nx10394, nx10396, nx10398, nx10400, nx10402, nx10404, nx10406, nx10408, 
         nx10410, nx10412, nx10414, nx10416, nx10418, nx10420, nx10422, nx10424, 
         nx10426, nx10428, nx10430, nx10432, nx10434, nx10436, nx10438, nx10440, 
         nx10442, nx10444, nx10446, nx10448, nx10450, nx10452, nx10454, nx10456, 
         nx10458, nx10460, nx10462, nx10464, nx10466, nx10468, nx10470, nx10472, 
         nx10474, nx10476, nx10478, nx10480, nx10482, nx10484, nx10486, nx10488, 
         nx10490, nx10492, nx10494, nx10496, nx10498, nx10500, nx10502, nx10504, 
         nx10506, nx10508, nx10510, nx10512, nx10514, nx10516, nx10518, nx10520, 
         nx10522, nx10524, nx10526, nx10528, nx10530, nx10532, nx10534, nx10536, 
         nx10538, nx10540, nx10542, nx10544, nx10546, nx10548, nx10550, nx10552, 
         nx10554, nx10556, nx10558, nx10560, nx10562, nx10564, nx10566, nx10568, 
         nx10570, nx10572, nx10574, nx10576, nx10578, nx10580, nx10582, nx10584, 
         nx10586, nx10588, nx10590, nx10592, nx10594, nx10596, nx10598, nx10600, 
         nx10602, nx10604, nx10606, nx10608, nx10610, nx10612, nx10614, nx10616, 
         nx10618, nx10620, nx10622, nx10624, nx10626, nx10628, nx10630, nx10632, 
         nx10634, nx10636, nx10638, nx10640, nx10642, nx10644, nx10646, nx10648, 
         nx10650, nx10652, nx10654, nx10656, nx10658, nx10660, nx10662, nx10664, 
         nx10666, nx10668, nx10670, nx10672, nx10674, nx10676, nx10678, nx10680, 
         nx10682, nx10684, nx10686, nx10688, nx10690, nx10692, nx10694, nx10696, 
         nx10698, nx10700, nx10702, nx10704, nx10706, nx10708, nx10710, nx10712, 
         nx10714, nx10716, nx10718, nx10720, nx10722, nx10724, nx10726, nx10728, 
         nx10730, nx10732, nx10734, nx10736, nx10738, nx10740, nx10742, nx10744, 
         nx10746, nx10748, nx10750, nx10752, nx10754, nx10756, nx10758, nx10760, 
         nx10762, nx10764, nx10766, nx10768, nx10770, nx10772, nx10774, nx10776, 
         nx10778, nx10780, nx10782, nx10784, nx10786, nx10788, nx10790, nx10792, 
         nx10794, nx10796, nx10798, nx10800, nx10802, nx10804, nx10806, nx10808, 
         nx10810, nx10812, nx10814, nx10816, nx10818, nx10820, nx10822, nx10824, 
         nx10826, nx10828, nx10830, nx10832, nx10834, nx10836, nx10838, nx10840, 
         nx10842, nx10844, nx10846, nx10848, nx10850, nx10852, nx10854, nx10856, 
         nx10858, nx10860, nx10862, nx10864, nx10866, nx10868, nx10870, nx10872, 
         nx10874, nx10876, nx10878, nx10880, nx10882, nx10884, nx10886, nx10888, 
         nx10890, nx10892, nx10894, nx10896, nx10898, nx10900, nx10902, nx10904, 
         nx10906, nx10908, nx10910, nx10912, nx10914, nx10916, nx10918, nx10920, 
         nx10922, nx10924, nx10926, nx10928, nx10930, nx10932, nx10934, nx10936, 
         nx10938, nx10940, nx10942, nx10944, nx10946, nx10948, nx10950, nx10952, 
         nx10954, nx10956, nx10958, nx10960, nx10962, nx10964, nx10966, nx10968, 
         nx10970, nx10972, nx10974, nx10976, nx10978, nx10980, nx10982, nx10984, 
         nx10986, nx10988, nx10990, nx10992, nx10994, nx10996, nx10998, nx11000, 
         nx11002, nx11004, nx11006, nx11008, nx11010, nx11012, nx11014, nx11016, 
         nx11018, nx11020, nx11022, nx11024, nx11026, nx11028, nx11030, nx11032, 
         nx11034, nx11036, nx11038, nx11040, nx11042, nx11044, nx11046, nx11048, 
         nx11050, nx11052, nx11054, nx11056, nx11058, nx11060, nx11062, nx11064, 
         nx11066, nx11068, nx11070, nx11072, nx11074, nx11076, nx11078, nx11080, 
         nx11082, nx11084, nx11086, nx11088, nx11090, nx11092, nx11094, nx11096, 
         nx11098, nx11100, nx11102, nx11104, nx11106, nx11108, nx11110, nx11112, 
         nx11114, nx11116, nx11118, nx11120, nx11122, nx11124, nx11126, nx11128, 
         nx11130, nx11132, nx11134, nx11136, nx11138, nx11140, nx11142, nx11144, 
         nx11146, nx11148, nx11150, nx11152, nx11154, nx11156, nx11158, nx11160, 
         nx11162, nx11164, nx11166, nx11168, nx11170, nx11172, nx11174, nx11176, 
         nx11178, nx11180, nx11182, nx11184, nx11186, nx11188, nx11190, nx11192, 
         nx11194, nx11196, nx11198, nx11200, nx11202, nx11204, nx11206, nx11208, 
         nx11210, nx11212, nx11214, nx11216, nx11218, nx11220, nx11222, nx11224, 
         nx11226, nx11228, nx11230, nx11232, nx11234, nx11236, nx11238, nx11240, 
         nx11242, nx11244, nx11246, nx11248, nx11250, nx11252, nx11254, nx11256, 
         nx11258, nx11260, nx11262, nx11264, nx11266, nx11268, nx11270, nx11272, 
         nx11274, nx11276, nx11278, nx11280, nx11282, nx11284, nx11286, nx11288, 
         nx11290, nx11292, nx11294, nx11296, nx11298, nx11300, nx11302, nx11304, 
         nx11306, nx11308, nx11310, nx11312, nx11314, nx11316, nx11318, nx11320, 
         nx11322, nx11324, nx11326, nx11328, nx11330, nx11332, nx11334, nx11336, 
         nx11338, nx11340, nx11342, nx11344, nx11346, nx11348, nx11350, nx11352, 
         nx11354, nx11356, nx11358, nx11360, nx11362, nx11364, nx11366, nx11368, 
         nx11370, nx11372, nx11374, nx11376, nx11378, nx11380, nx11382, nx11384, 
         nx11386, nx11388, nx11390, nx11392, nx11394, nx11396, nx11398, nx11400, 
         nx11402, nx11404, nx11406, nx11408, nx11410, nx11412, nx11414, nx11416, 
         nx11418, nx11420, nx11422, nx11424, nx11426, nx11428, nx11430, nx11432, 
         nx11434, nx11436, nx11438, nx11440, nx11442, nx11444, nx11446, nx11448, 
         nx11450, nx11452, nx11454, nx11456, nx11458, nx11460, nx11462, nx11464, 
         nx11466, nx11468, nx11470, nx11472, nx11474, nx11476, nx11478, nx11480, 
         nx11482, nx11484, nx11486, nx11488, nx11490, nx11492, nx11494, nx11496, 
         nx11498, nx11500, nx11502, nx11504, nx11506, nx11508, nx11510, nx11512, 
         nx11514, nx11516, nx11518, nx11520, nx11522, nx11524, nx11526, nx11528, 
         nx11530, nx11532, nx11534, nx11536, nx11538, nx11540, nx11542, nx11544, 
         nx11546, nx11548, nx11550, nx11552, nx11554, nx11556, nx11558, nx11560, 
         nx11562, nx11564, nx11566, nx11568, nx11570, nx11572, nx11574, nx11576, 
         nx11578, nx11580, nx11582, nx11584, nx11586, nx11588, nx11590, nx11592, 
         nx11594, nx11596, nx11598, nx11600, nx11602, nx11604, nx11606, nx11608, 
         nx11610, nx11612, nx11614, nx11616, nx11618, nx11620, nx11622, nx11624, 
         nx11626, nx11628, nx11630, nx11632, nx11634, nx11636, nx11638, nx11640, 
         nx11642, nx11644, nx11646, nx11648, nx11650, nx11652, nx11654, nx11656, 
         nx11658, nx11660, nx11662, nx11664, nx11666, nx11668, nx11670, nx11672, 
         nx11674, nx11676, nx11678, nx11680, nx11682, nx11684, nx11686, nx11688, 
         nx11690, nx11692, nx11694, nx11696, nx11698, nx11700, nx11702, nx11704, 
         nx11706, nx11708, nx11710, nx11712, nx11714, nx11716, nx11718, nx11720, 
         nx11722, nx11724, nx11726, nx11728, nx11730, nx11732, nx11734, nx11736, 
         nx11738, nx11740, nx11742, nx11744, nx11746, nx11748, nx11750, nx11752, 
         nx11754, nx11756, nx11758, nx11760, nx11762, nx11764, nx11766, nx11768, 
         nx11770, nx11772, nx11774, nx11776, nx11778, nx11780, nx11782, nx11784, 
         nx11786, nx11788, nx11790, nx11792, nx11794, nx11796, nx11798, nx11800, 
         nx11802, nx11804, nx11806, nx11808, nx11810, nx11812, nx11814, nx11816, 
         nx11818, nx11820, nx11822, nx11824, nx11826, nx11828, nx11830, nx11832, 
         nx11834, nx11836, nx11838, nx11840, nx11842, nx11844, nx11846, nx11848, 
         nx11850, nx11852, nx11854, nx11856, nx11858, nx11860, nx11862, nx11864, 
         nx11866, nx11868, nx11870, nx11872, nx11874, nx11876, nx11878, nx11880, 
         nx11882, nx11884, nx11886, nx11896, nx11898, nx11900, nx11902, nx11904, 
         nx11906, nx11908, nx11910, nx11912, nx11914, nx11916, nx11918, nx11920, 
         nx11922, nx11924, nx11926, nx11928, nx11934, nx11936, nx11938, nx11940;
    wire [130:0] \$dummy ;




    Reg_33 gen_24_cmp_pRegCmp (.D ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
           gen_24_cmp_pBs_30,gen_24_cmp_pBs_29,gen_24_cmp_pBs_28,
           gen_24_cmp_pBs_27,gen_24_cmp_pBs_26,gen_24_cmp_pBs_25,
           gen_24_cmp_pBs_24,gen_24_cmp_pBs_23,outputs_24__15,outputs_24__14,
           outputs_24__13,outputs_24__12,outputs_24__11,outputs_24__10,
           outputs_24__9,outputs_24__8,outputs_24__7,outputs_24__6,outputs_24__5
           ,outputs_24__4,outputs_24__3,outputs_24__2,outputs_24__1,
           outputs_24__0,gen_24_cmp_pMux_8,gen_24_cmp_pMux_7,gen_24_cmp_pMux_6,
           gen_24_cmp_pMux_5,gen_24_cmp_pMux_4,gen_24_cmp_pMux_3,nx10130}), .en (
           nx11916), .clk (nx10122), .rst (rst), .Q ({\$dummy [0],\$dummy [1],
           gen_24_cmp_pReg_30,gen_24_cmp_pReg_29,gen_24_cmp_pReg_28,
           gen_24_cmp_pReg_27,gen_24_cmp_pReg_26,gen_24_cmp_pReg_25,
           gen_24_cmp_pReg_24,gen_24_cmp_pReg_23,gen_24_cmp_pReg_22,
           gen_24_cmp_pReg_21,gen_24_cmp_pReg_20,gen_24_cmp_pReg_19,
           gen_24_cmp_pReg_18,gen_24_cmp_pReg_17,gen_24_cmp_pReg_16,
           gen_24_cmp_pReg_15,gen_24_cmp_pReg_14,gen_24_cmp_pReg_13,
           gen_24_cmp_pReg_12,gen_24_cmp_pReg_11,gen_24_cmp_pReg_10,
           gen_24_cmp_pReg_9,gen_24_cmp_pReg_8,gen_24_cmp_pReg_7,
           gen_24_cmp_pReg_6,gen_24_cmp_pReg_5,gen_24_cmp_pReg_4,
           gen_24_cmp_pReg_3,gen_24_cmp_pReg_2,gen_24_cmp_pReg_1,
           gen_24_cmp_pReg_0})) ;
    BinaryMux_33 gen_24_cmp_MuxCmp (.a ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32
                 ,gen_24_cmp_pReg_30,gen_24_cmp_pReg_29,gen_24_cmp_pReg_28,
                 gen_24_cmp_pReg_27,gen_24_cmp_pReg_26,gen_24_cmp_pReg_25,
                 gen_24_cmp_pReg_24,gen_24_cmp_pReg_23,gen_24_cmp_pReg_22,
                 gen_24_cmp_pReg_21,gen_24_cmp_pReg_20,gen_24_cmp_pReg_19,
                 gen_24_cmp_pReg_18,gen_24_cmp_pReg_17,gen_24_cmp_pReg_16,
                 gen_24_cmp_pReg_15,gen_24_cmp_pReg_14,gen_24_cmp_pReg_13,
                 gen_24_cmp_pReg_12,gen_24_cmp_pReg_11,gen_24_cmp_pReg_10,
                 gen_24_cmp_pReg_9,gen_24_cmp_pReg_8,gen_24_cmp_pReg_7,
                 gen_24_cmp_pReg_6,gen_24_cmp_pReg_5,gen_24_cmp_pReg_4,
                 gen_24_cmp_pReg_3,gen_24_cmp_pReg_2,gen_24_cmp_pReg_1,
                 gen_24_cmp_pReg_0}), .b ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,filter_24__7,
                 filter_24__6,filter_24__5,filter_24__4,filter_24__3,
                 filter_24__2,filter_24__1,filter_24__0,gen_24_cmp_pInit_32}), .sel (
                 nx11896), .f ({\$dummy [2],\$dummy [3],gen_24_cmp_pMux_30,
                 gen_24_cmp_pMux_29,gen_24_cmp_pMux_28,gen_24_cmp_pMux_27,
                 gen_24_cmp_pMux_26,gen_24_cmp_pMux_25,gen_24_cmp_pMux_24,
                 gen_24_cmp_pMux_23,gen_24_cmp_pMux_22,gen_24_cmp_pMux_21,
                 gen_24_cmp_pMux_20,gen_24_cmp_pMux_19,gen_24_cmp_pMux_18,
                 gen_24_cmp_pMux_17,gen_24_cmp_pMux_16,gen_24_cmp_pMux_15,
                 gen_24_cmp_pMux_14,gen_24_cmp_pMux_13,gen_24_cmp_pMux_12,
                 gen_24_cmp_pMux_11,gen_24_cmp_pMux_10,gen_24_cmp_pMux_9,
                 gen_24_cmp_pMux_8,gen_24_cmp_pMux_7,gen_24_cmp_pMux_6,
                 gen_24_cmp_pMux_5,gen_24_cmp_pMux_4,gen_24_cmp_pMux_3,
                 gen_24_cmp_pMux_2,gen_24_cmp_pMux_1,gen_24_cmp_pMux_0})) ;
    NBitAdder_24 gen_24_cmp_BSCmp_AdderCmp (.a ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pMux_30,gen_24_cmp_pMux_29,
                 gen_24_cmp_pMux_28,gen_24_cmp_pMux_27,gen_24_cmp_pMux_26,
                 gen_24_cmp_pMux_25,gen_24_cmp_pMux_24,gen_24_cmp_pMux_23,
                 gen_24_cmp_pMux_22,gen_24_cmp_pMux_21,gen_24_cmp_pMux_20,
                 gen_24_cmp_pMux_19,gen_24_cmp_pMux_18,gen_24_cmp_pMux_17,
                 gen_24_cmp_pMux_16,gen_24_cmp_pMux_15,gen_24_cmp_pMux_14,
                 gen_24_cmp_pMux_13,gen_24_cmp_pMux_12,gen_24_cmp_pMux_11,
                 gen_24_cmp_pMux_10,gen_24_cmp_pMux_9}), .b ({nx10434,nx10434,
                 nx10432,nx10440,nx10438,nx10436,nx10434,nx10432,
                 gen_24_cmp_BSCmp_op2_15,gen_24_cmp_BSCmp_op2_14,
                 gen_24_cmp_BSCmp_op2_13,gen_24_cmp_BSCmp_op2_12,
                 gen_24_cmp_BSCmp_op2_11,gen_24_cmp_BSCmp_op2_10,
                 gen_24_cmp_BSCmp_op2_9,gen_24_cmp_BSCmp_op2_8,
                 gen_24_cmp_BSCmp_op2_7,gen_24_cmp_BSCmp_op2_6,
                 gen_24_cmp_BSCmp_op2_5,gen_24_cmp_BSCmp_op2_4,
                 gen_24_cmp_BSCmp_op2_3,gen_24_cmp_BSCmp_op2_2,
                 gen_24_cmp_BSCmp_op2_1,gen_24_cmp_BSCmp_op2_0}), .carryIn (
                 gen_24_cmp_BSCmp_carryIn), .sum ({gen_24_cmp_pBs_30,
                 gen_24_cmp_pBs_29,gen_24_cmp_pBs_28,gen_24_cmp_pBs_27,
                 gen_24_cmp_pBs_26,gen_24_cmp_pBs_25,gen_24_cmp_pBs_24,
                 gen_24_cmp_pBs_23,outputs_24__15,outputs_24__14,outputs_24__13,
                 outputs_24__12,outputs_24__11,outputs_24__10,outputs_24__9,
                 outputs_24__8,outputs_24__7,outputs_24__6,outputs_24__5,
                 outputs_24__4,outputs_24__3,outputs_24__2,outputs_24__1,
                 outputs_24__0}), .carryOut (\$dummy [4])) ;
    Reg_33 gen_23_cmp_pRegCmp (.D ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
           gen_23_cmp_pBs_30,gen_23_cmp_pBs_29,gen_23_cmp_pBs_28,
           gen_23_cmp_pBs_27,gen_23_cmp_pBs_26,gen_23_cmp_pBs_25,
           gen_23_cmp_pBs_24,gen_23_cmp_pBs_23,outputs_23__15,outputs_23__14,
           outputs_23__13,outputs_23__12,outputs_23__11,outputs_23__10,
           outputs_23__9,outputs_23__8,outputs_23__7,outputs_23__6,outputs_23__5
           ,outputs_23__4,outputs_23__3,outputs_23__2,outputs_23__1,
           outputs_23__0,gen_23_cmp_pMux_8,gen_23_cmp_pMux_7,gen_23_cmp_pMux_6,
           gen_23_cmp_pMux_5,gen_23_cmp_pMux_4,gen_23_cmp_pMux_3,nx10142}), .en (
           nx11916), .clk (nx10122), .rst (rst), .Q ({\$dummy [5],\$dummy [6],
           gen_23_cmp_pReg_30,gen_23_cmp_pReg_29,gen_23_cmp_pReg_28,
           gen_23_cmp_pReg_27,gen_23_cmp_pReg_26,gen_23_cmp_pReg_25,
           gen_23_cmp_pReg_24,gen_23_cmp_pReg_23,gen_23_cmp_pReg_22,
           gen_23_cmp_pReg_21,gen_23_cmp_pReg_20,gen_23_cmp_pReg_19,
           gen_23_cmp_pReg_18,gen_23_cmp_pReg_17,gen_23_cmp_pReg_16,
           gen_23_cmp_pReg_15,gen_23_cmp_pReg_14,gen_23_cmp_pReg_13,
           gen_23_cmp_pReg_12,gen_23_cmp_pReg_11,gen_23_cmp_pReg_10,
           gen_23_cmp_pReg_9,gen_23_cmp_pReg_8,gen_23_cmp_pReg_7,
           gen_23_cmp_pReg_6,gen_23_cmp_pReg_5,gen_23_cmp_pReg_4,
           gen_23_cmp_pReg_3,gen_23_cmp_pReg_2,gen_23_cmp_pReg_1,
           gen_23_cmp_pReg_0})) ;
    BinaryMux_33 gen_23_cmp_MuxCmp (.a ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32
                 ,gen_23_cmp_pReg_30,gen_23_cmp_pReg_29,gen_23_cmp_pReg_28,
                 gen_23_cmp_pReg_27,gen_23_cmp_pReg_26,gen_23_cmp_pReg_25,
                 gen_23_cmp_pReg_24,gen_23_cmp_pReg_23,gen_23_cmp_pReg_22,
                 gen_23_cmp_pReg_21,gen_23_cmp_pReg_20,gen_23_cmp_pReg_19,
                 gen_23_cmp_pReg_18,gen_23_cmp_pReg_17,gen_23_cmp_pReg_16,
                 gen_23_cmp_pReg_15,gen_23_cmp_pReg_14,gen_23_cmp_pReg_13,
                 gen_23_cmp_pReg_12,gen_23_cmp_pReg_11,gen_23_cmp_pReg_10,
                 gen_23_cmp_pReg_9,gen_23_cmp_pReg_8,gen_23_cmp_pReg_7,
                 gen_23_cmp_pReg_6,gen_23_cmp_pReg_5,gen_23_cmp_pReg_4,
                 gen_23_cmp_pReg_3,gen_23_cmp_pReg_2,gen_23_cmp_pReg_1,
                 gen_23_cmp_pReg_0}), .b ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,filter_23__7,
                 filter_23__6,filter_23__5,filter_23__4,filter_23__3,
                 filter_23__2,filter_23__1,filter_23__0,gen_24_cmp_pInit_32}), .sel (
                 nx11896), .f ({\$dummy [7],\$dummy [8],gen_23_cmp_pMux_30,
                 gen_23_cmp_pMux_29,gen_23_cmp_pMux_28,gen_23_cmp_pMux_27,
                 gen_23_cmp_pMux_26,gen_23_cmp_pMux_25,gen_23_cmp_pMux_24,
                 gen_23_cmp_pMux_23,gen_23_cmp_pMux_22,gen_23_cmp_pMux_21,
                 gen_23_cmp_pMux_20,gen_23_cmp_pMux_19,gen_23_cmp_pMux_18,
                 gen_23_cmp_pMux_17,gen_23_cmp_pMux_16,gen_23_cmp_pMux_15,
                 gen_23_cmp_pMux_14,gen_23_cmp_pMux_13,gen_23_cmp_pMux_12,
                 gen_23_cmp_pMux_11,gen_23_cmp_pMux_10,gen_23_cmp_pMux_9,
                 gen_23_cmp_pMux_8,gen_23_cmp_pMux_7,gen_23_cmp_pMux_6,
                 gen_23_cmp_pMux_5,gen_23_cmp_pMux_4,gen_23_cmp_pMux_3,
                 gen_23_cmp_pMux_2,gen_23_cmp_pMux_1,gen_23_cmp_pMux_0})) ;
    NBitAdder_24 gen_23_cmp_BSCmp_AdderCmp (.a ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_23_cmp_pMux_30,gen_23_cmp_pMux_29,
                 gen_23_cmp_pMux_28,gen_23_cmp_pMux_27,gen_23_cmp_pMux_26,
                 gen_23_cmp_pMux_25,gen_23_cmp_pMux_24,gen_23_cmp_pMux_23,
                 gen_23_cmp_pMux_22,gen_23_cmp_pMux_21,gen_23_cmp_pMux_20,
                 gen_23_cmp_pMux_19,gen_23_cmp_pMux_18,gen_23_cmp_pMux_17,
                 gen_23_cmp_pMux_16,gen_23_cmp_pMux_15,gen_23_cmp_pMux_14,
                 gen_23_cmp_pMux_13,gen_23_cmp_pMux_12,gen_23_cmp_pMux_11,
                 gen_23_cmp_pMux_10,gen_23_cmp_pMux_9}), .b ({nx10446,nx10446,
                 nx10444,nx10452,nx10450,nx10448,nx10446,nx10444,
                 gen_23_cmp_BSCmp_op2_15,gen_23_cmp_BSCmp_op2_14,
                 gen_23_cmp_BSCmp_op2_13,gen_23_cmp_BSCmp_op2_12,
                 gen_23_cmp_BSCmp_op2_11,gen_23_cmp_BSCmp_op2_10,
                 gen_23_cmp_BSCmp_op2_9,gen_23_cmp_BSCmp_op2_8,
                 gen_23_cmp_BSCmp_op2_7,gen_23_cmp_BSCmp_op2_6,
                 gen_23_cmp_BSCmp_op2_5,gen_23_cmp_BSCmp_op2_4,
                 gen_23_cmp_BSCmp_op2_3,gen_23_cmp_BSCmp_op2_2,
                 gen_23_cmp_BSCmp_op2_1,gen_23_cmp_BSCmp_op2_0}), .carryIn (
                 gen_23_cmp_BSCmp_carryIn), .sum ({gen_23_cmp_pBs_30,
                 gen_23_cmp_pBs_29,gen_23_cmp_pBs_28,gen_23_cmp_pBs_27,
                 gen_23_cmp_pBs_26,gen_23_cmp_pBs_25,gen_23_cmp_pBs_24,
                 gen_23_cmp_pBs_23,outputs_23__15,outputs_23__14,outputs_23__13,
                 outputs_23__12,outputs_23__11,outputs_23__10,outputs_23__9,
                 outputs_23__8,outputs_23__7,outputs_23__6,outputs_23__5,
                 outputs_23__4,outputs_23__3,outputs_23__2,outputs_23__1,
                 outputs_23__0}), .carryOut (\$dummy [9])) ;
    Reg_33 gen_22_cmp_pRegCmp (.D ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
           gen_22_cmp_pBs_30,gen_22_cmp_pBs_29,gen_22_cmp_pBs_28,
           gen_22_cmp_pBs_27,gen_22_cmp_pBs_26,gen_22_cmp_pBs_25,
           gen_22_cmp_pBs_24,gen_22_cmp_pBs_23,outputs_22__15,outputs_22__14,
           outputs_22__13,outputs_22__12,outputs_22__11,outputs_22__10,
           outputs_22__9,outputs_22__8,outputs_22__7,outputs_22__6,outputs_22__5
           ,outputs_22__4,outputs_22__3,outputs_22__2,outputs_22__1,
           outputs_22__0,gen_22_cmp_pMux_8,gen_22_cmp_pMux_7,gen_22_cmp_pMux_6,
           gen_22_cmp_pMux_5,gen_22_cmp_pMux_4,gen_22_cmp_pMux_3,nx10154}), .en (
           nx11916), .clk (nx10122), .rst (rst), .Q ({\$dummy [10],\$dummy [11],
           gen_22_cmp_pReg_30,gen_22_cmp_pReg_29,gen_22_cmp_pReg_28,
           gen_22_cmp_pReg_27,gen_22_cmp_pReg_26,gen_22_cmp_pReg_25,
           gen_22_cmp_pReg_24,gen_22_cmp_pReg_23,gen_22_cmp_pReg_22,
           gen_22_cmp_pReg_21,gen_22_cmp_pReg_20,gen_22_cmp_pReg_19,
           gen_22_cmp_pReg_18,gen_22_cmp_pReg_17,gen_22_cmp_pReg_16,
           gen_22_cmp_pReg_15,gen_22_cmp_pReg_14,gen_22_cmp_pReg_13,
           gen_22_cmp_pReg_12,gen_22_cmp_pReg_11,gen_22_cmp_pReg_10,
           gen_22_cmp_pReg_9,gen_22_cmp_pReg_8,gen_22_cmp_pReg_7,
           gen_22_cmp_pReg_6,gen_22_cmp_pReg_5,gen_22_cmp_pReg_4,
           gen_22_cmp_pReg_3,gen_22_cmp_pReg_2,gen_22_cmp_pReg_1,
           gen_22_cmp_pReg_0})) ;
    BinaryMux_33 gen_22_cmp_MuxCmp (.a ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32
                 ,gen_22_cmp_pReg_30,gen_22_cmp_pReg_29,gen_22_cmp_pReg_28,
                 gen_22_cmp_pReg_27,gen_22_cmp_pReg_26,gen_22_cmp_pReg_25,
                 gen_22_cmp_pReg_24,gen_22_cmp_pReg_23,gen_22_cmp_pReg_22,
                 gen_22_cmp_pReg_21,gen_22_cmp_pReg_20,gen_22_cmp_pReg_19,
                 gen_22_cmp_pReg_18,gen_22_cmp_pReg_17,gen_22_cmp_pReg_16,
                 gen_22_cmp_pReg_15,gen_22_cmp_pReg_14,gen_22_cmp_pReg_13,
                 gen_22_cmp_pReg_12,gen_22_cmp_pReg_11,gen_22_cmp_pReg_10,
                 gen_22_cmp_pReg_9,gen_22_cmp_pReg_8,gen_22_cmp_pReg_7,
                 gen_22_cmp_pReg_6,gen_22_cmp_pReg_5,gen_22_cmp_pReg_4,
                 gen_22_cmp_pReg_3,gen_22_cmp_pReg_2,gen_22_cmp_pReg_1,
                 gen_22_cmp_pReg_0}), .b ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,filter_22__7,
                 filter_22__6,filter_22__5,filter_22__4,filter_22__3,
                 filter_22__2,filter_22__1,filter_22__0,gen_24_cmp_pInit_32}), .sel (
                 nx11896), .f ({\$dummy [12],\$dummy [13],gen_22_cmp_pMux_30,
                 gen_22_cmp_pMux_29,gen_22_cmp_pMux_28,gen_22_cmp_pMux_27,
                 gen_22_cmp_pMux_26,gen_22_cmp_pMux_25,gen_22_cmp_pMux_24,
                 gen_22_cmp_pMux_23,gen_22_cmp_pMux_22,gen_22_cmp_pMux_21,
                 gen_22_cmp_pMux_20,gen_22_cmp_pMux_19,gen_22_cmp_pMux_18,
                 gen_22_cmp_pMux_17,gen_22_cmp_pMux_16,gen_22_cmp_pMux_15,
                 gen_22_cmp_pMux_14,gen_22_cmp_pMux_13,gen_22_cmp_pMux_12,
                 gen_22_cmp_pMux_11,gen_22_cmp_pMux_10,gen_22_cmp_pMux_9,
                 gen_22_cmp_pMux_8,gen_22_cmp_pMux_7,gen_22_cmp_pMux_6,
                 gen_22_cmp_pMux_5,gen_22_cmp_pMux_4,gen_22_cmp_pMux_3,
                 gen_22_cmp_pMux_2,gen_22_cmp_pMux_1,gen_22_cmp_pMux_0})) ;
    NBitAdder_24 gen_22_cmp_BSCmp_AdderCmp (.a ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_22_cmp_pMux_30,gen_22_cmp_pMux_29,
                 gen_22_cmp_pMux_28,gen_22_cmp_pMux_27,gen_22_cmp_pMux_26,
                 gen_22_cmp_pMux_25,gen_22_cmp_pMux_24,gen_22_cmp_pMux_23,
                 gen_22_cmp_pMux_22,gen_22_cmp_pMux_21,gen_22_cmp_pMux_20,
                 gen_22_cmp_pMux_19,gen_22_cmp_pMux_18,gen_22_cmp_pMux_17,
                 gen_22_cmp_pMux_16,gen_22_cmp_pMux_15,gen_22_cmp_pMux_14,
                 gen_22_cmp_pMux_13,gen_22_cmp_pMux_12,gen_22_cmp_pMux_11,
                 gen_22_cmp_pMux_10,gen_22_cmp_pMux_9}), .b ({nx10458,nx10458,
                 nx10456,nx10464,nx10462,nx10460,nx10458,nx10456,
                 gen_22_cmp_BSCmp_op2_15,gen_22_cmp_BSCmp_op2_14,
                 gen_22_cmp_BSCmp_op2_13,gen_22_cmp_BSCmp_op2_12,
                 gen_22_cmp_BSCmp_op2_11,gen_22_cmp_BSCmp_op2_10,
                 gen_22_cmp_BSCmp_op2_9,gen_22_cmp_BSCmp_op2_8,
                 gen_22_cmp_BSCmp_op2_7,gen_22_cmp_BSCmp_op2_6,
                 gen_22_cmp_BSCmp_op2_5,gen_22_cmp_BSCmp_op2_4,
                 gen_22_cmp_BSCmp_op2_3,gen_22_cmp_BSCmp_op2_2,
                 gen_22_cmp_BSCmp_op2_1,gen_22_cmp_BSCmp_op2_0}), .carryIn (
                 gen_22_cmp_BSCmp_carryIn), .sum ({gen_22_cmp_pBs_30,
                 gen_22_cmp_pBs_29,gen_22_cmp_pBs_28,gen_22_cmp_pBs_27,
                 gen_22_cmp_pBs_26,gen_22_cmp_pBs_25,gen_22_cmp_pBs_24,
                 gen_22_cmp_pBs_23,outputs_22__15,outputs_22__14,outputs_22__13,
                 outputs_22__12,outputs_22__11,outputs_22__10,outputs_22__9,
                 outputs_22__8,outputs_22__7,outputs_22__6,outputs_22__5,
                 outputs_22__4,outputs_22__3,outputs_22__2,outputs_22__1,
                 outputs_22__0}), .carryOut (\$dummy [14])) ;
    Reg_33 gen_21_cmp_pRegCmp (.D ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
           gen_21_cmp_pBs_30,gen_21_cmp_pBs_29,gen_21_cmp_pBs_28,
           gen_21_cmp_pBs_27,gen_21_cmp_pBs_26,gen_21_cmp_pBs_25,
           gen_21_cmp_pBs_24,gen_21_cmp_pBs_23,outputs_21__15,outputs_21__14,
           outputs_21__13,outputs_21__12,outputs_21__11,outputs_21__10,
           outputs_21__9,outputs_21__8,outputs_21__7,outputs_21__6,outputs_21__5
           ,outputs_21__4,outputs_21__3,outputs_21__2,outputs_21__1,
           outputs_21__0,gen_21_cmp_pMux_8,gen_21_cmp_pMux_7,gen_21_cmp_pMux_6,
           gen_21_cmp_pMux_5,gen_21_cmp_pMux_4,gen_21_cmp_pMux_3,nx10166}), .en (
           nx11918), .clk (nx10122), .rst (rst), .Q ({\$dummy [15],\$dummy [16],
           gen_21_cmp_pReg_30,gen_21_cmp_pReg_29,gen_21_cmp_pReg_28,
           gen_21_cmp_pReg_27,gen_21_cmp_pReg_26,gen_21_cmp_pReg_25,
           gen_21_cmp_pReg_24,gen_21_cmp_pReg_23,gen_21_cmp_pReg_22,
           gen_21_cmp_pReg_21,gen_21_cmp_pReg_20,gen_21_cmp_pReg_19,
           gen_21_cmp_pReg_18,gen_21_cmp_pReg_17,gen_21_cmp_pReg_16,
           gen_21_cmp_pReg_15,gen_21_cmp_pReg_14,gen_21_cmp_pReg_13,
           gen_21_cmp_pReg_12,gen_21_cmp_pReg_11,gen_21_cmp_pReg_10,
           gen_21_cmp_pReg_9,gen_21_cmp_pReg_8,gen_21_cmp_pReg_7,
           gen_21_cmp_pReg_6,gen_21_cmp_pReg_5,gen_21_cmp_pReg_4,
           gen_21_cmp_pReg_3,gen_21_cmp_pReg_2,gen_21_cmp_pReg_1,
           gen_21_cmp_pReg_0})) ;
    BinaryMux_33 gen_21_cmp_MuxCmp (.a ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32
                 ,gen_21_cmp_pReg_30,gen_21_cmp_pReg_29,gen_21_cmp_pReg_28,
                 gen_21_cmp_pReg_27,gen_21_cmp_pReg_26,gen_21_cmp_pReg_25,
                 gen_21_cmp_pReg_24,gen_21_cmp_pReg_23,gen_21_cmp_pReg_22,
                 gen_21_cmp_pReg_21,gen_21_cmp_pReg_20,gen_21_cmp_pReg_19,
                 gen_21_cmp_pReg_18,gen_21_cmp_pReg_17,gen_21_cmp_pReg_16,
                 gen_21_cmp_pReg_15,gen_21_cmp_pReg_14,gen_21_cmp_pReg_13,
                 gen_21_cmp_pReg_12,gen_21_cmp_pReg_11,gen_21_cmp_pReg_10,
                 gen_21_cmp_pReg_9,gen_21_cmp_pReg_8,gen_21_cmp_pReg_7,
                 gen_21_cmp_pReg_6,gen_21_cmp_pReg_5,gen_21_cmp_pReg_4,
                 gen_21_cmp_pReg_3,gen_21_cmp_pReg_2,gen_21_cmp_pReg_1,
                 gen_21_cmp_pReg_0}), .b ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,filter_21__7,
                 filter_21__6,filter_21__5,filter_21__4,filter_21__3,
                 filter_21__2,filter_21__1,filter_21__0,gen_24_cmp_pInit_32}), .sel (
                 nx11898), .f ({\$dummy [17],\$dummy [18],gen_21_cmp_pMux_30,
                 gen_21_cmp_pMux_29,gen_21_cmp_pMux_28,gen_21_cmp_pMux_27,
                 gen_21_cmp_pMux_26,gen_21_cmp_pMux_25,gen_21_cmp_pMux_24,
                 gen_21_cmp_pMux_23,gen_21_cmp_pMux_22,gen_21_cmp_pMux_21,
                 gen_21_cmp_pMux_20,gen_21_cmp_pMux_19,gen_21_cmp_pMux_18,
                 gen_21_cmp_pMux_17,gen_21_cmp_pMux_16,gen_21_cmp_pMux_15,
                 gen_21_cmp_pMux_14,gen_21_cmp_pMux_13,gen_21_cmp_pMux_12,
                 gen_21_cmp_pMux_11,gen_21_cmp_pMux_10,gen_21_cmp_pMux_9,
                 gen_21_cmp_pMux_8,gen_21_cmp_pMux_7,gen_21_cmp_pMux_6,
                 gen_21_cmp_pMux_5,gen_21_cmp_pMux_4,gen_21_cmp_pMux_3,
                 gen_21_cmp_pMux_2,gen_21_cmp_pMux_1,gen_21_cmp_pMux_0})) ;
    NBitAdder_24 gen_21_cmp_BSCmp_AdderCmp (.a ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_21_cmp_pMux_30,gen_21_cmp_pMux_29,
                 gen_21_cmp_pMux_28,gen_21_cmp_pMux_27,gen_21_cmp_pMux_26,
                 gen_21_cmp_pMux_25,gen_21_cmp_pMux_24,gen_21_cmp_pMux_23,
                 gen_21_cmp_pMux_22,gen_21_cmp_pMux_21,gen_21_cmp_pMux_20,
                 gen_21_cmp_pMux_19,gen_21_cmp_pMux_18,gen_21_cmp_pMux_17,
                 gen_21_cmp_pMux_16,gen_21_cmp_pMux_15,gen_21_cmp_pMux_14,
                 gen_21_cmp_pMux_13,gen_21_cmp_pMux_12,gen_21_cmp_pMux_11,
                 gen_21_cmp_pMux_10,gen_21_cmp_pMux_9}), .b ({nx10470,nx10470,
                 nx10468,nx10476,nx10474,nx10472,nx10470,nx10468,
                 gen_21_cmp_BSCmp_op2_15,gen_21_cmp_BSCmp_op2_14,
                 gen_21_cmp_BSCmp_op2_13,gen_21_cmp_BSCmp_op2_12,
                 gen_21_cmp_BSCmp_op2_11,gen_21_cmp_BSCmp_op2_10,
                 gen_21_cmp_BSCmp_op2_9,gen_21_cmp_BSCmp_op2_8,
                 gen_21_cmp_BSCmp_op2_7,gen_21_cmp_BSCmp_op2_6,
                 gen_21_cmp_BSCmp_op2_5,gen_21_cmp_BSCmp_op2_4,
                 gen_21_cmp_BSCmp_op2_3,gen_21_cmp_BSCmp_op2_2,
                 gen_21_cmp_BSCmp_op2_1,gen_21_cmp_BSCmp_op2_0}), .carryIn (
                 gen_21_cmp_BSCmp_carryIn), .sum ({gen_21_cmp_pBs_30,
                 gen_21_cmp_pBs_29,gen_21_cmp_pBs_28,gen_21_cmp_pBs_27,
                 gen_21_cmp_pBs_26,gen_21_cmp_pBs_25,gen_21_cmp_pBs_24,
                 gen_21_cmp_pBs_23,outputs_21__15,outputs_21__14,outputs_21__13,
                 outputs_21__12,outputs_21__11,outputs_21__10,outputs_21__9,
                 outputs_21__8,outputs_21__7,outputs_21__6,outputs_21__5,
                 outputs_21__4,outputs_21__3,outputs_21__2,outputs_21__1,
                 outputs_21__0}), .carryOut (\$dummy [19])) ;
    Reg_33 gen_20_cmp_pRegCmp (.D ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
           gen_20_cmp_pBs_30,gen_20_cmp_pBs_29,gen_20_cmp_pBs_28,
           gen_20_cmp_pBs_27,gen_20_cmp_pBs_26,gen_20_cmp_pBs_25,
           gen_20_cmp_pBs_24,gen_20_cmp_pBs_23,outputs_20__15,outputs_20__14,
           outputs_20__13,outputs_20__12,outputs_20__11,outputs_20__10,
           outputs_20__9,outputs_20__8,outputs_20__7,outputs_20__6,outputs_20__5
           ,outputs_20__4,outputs_20__3,outputs_20__2,outputs_20__1,
           outputs_20__0,gen_20_cmp_pMux_8,gen_20_cmp_pMux_7,gen_20_cmp_pMux_6,
           gen_20_cmp_pMux_5,gen_20_cmp_pMux_4,gen_20_cmp_pMux_3,nx10178}), .en (
           nx11918), .clk (nx10122), .rst (rst), .Q ({\$dummy [20],\$dummy [21],
           gen_20_cmp_pReg_30,gen_20_cmp_pReg_29,gen_20_cmp_pReg_28,
           gen_20_cmp_pReg_27,gen_20_cmp_pReg_26,gen_20_cmp_pReg_25,
           gen_20_cmp_pReg_24,gen_20_cmp_pReg_23,gen_20_cmp_pReg_22,
           gen_20_cmp_pReg_21,gen_20_cmp_pReg_20,gen_20_cmp_pReg_19,
           gen_20_cmp_pReg_18,gen_20_cmp_pReg_17,gen_20_cmp_pReg_16,
           gen_20_cmp_pReg_15,gen_20_cmp_pReg_14,gen_20_cmp_pReg_13,
           gen_20_cmp_pReg_12,gen_20_cmp_pReg_11,gen_20_cmp_pReg_10,
           gen_20_cmp_pReg_9,gen_20_cmp_pReg_8,gen_20_cmp_pReg_7,
           gen_20_cmp_pReg_6,gen_20_cmp_pReg_5,gen_20_cmp_pReg_4,
           gen_20_cmp_pReg_3,gen_20_cmp_pReg_2,gen_20_cmp_pReg_1,
           gen_20_cmp_pReg_0})) ;
    BinaryMux_33 gen_20_cmp_MuxCmp (.a ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32
                 ,gen_20_cmp_pReg_30,gen_20_cmp_pReg_29,gen_20_cmp_pReg_28,
                 gen_20_cmp_pReg_27,gen_20_cmp_pReg_26,gen_20_cmp_pReg_25,
                 gen_20_cmp_pReg_24,gen_20_cmp_pReg_23,gen_20_cmp_pReg_22,
                 gen_20_cmp_pReg_21,gen_20_cmp_pReg_20,gen_20_cmp_pReg_19,
                 gen_20_cmp_pReg_18,gen_20_cmp_pReg_17,gen_20_cmp_pReg_16,
                 gen_20_cmp_pReg_15,gen_20_cmp_pReg_14,gen_20_cmp_pReg_13,
                 gen_20_cmp_pReg_12,gen_20_cmp_pReg_11,gen_20_cmp_pReg_10,
                 gen_20_cmp_pReg_9,gen_20_cmp_pReg_8,gen_20_cmp_pReg_7,
                 gen_20_cmp_pReg_6,gen_20_cmp_pReg_5,gen_20_cmp_pReg_4,
                 gen_20_cmp_pReg_3,gen_20_cmp_pReg_2,gen_20_cmp_pReg_1,
                 gen_20_cmp_pReg_0}), .b ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,filter_20__7,
                 filter_20__6,filter_20__5,filter_20__4,filter_20__3,
                 filter_20__2,filter_20__1,filter_20__0,gen_24_cmp_pInit_32}), .sel (
                 nx11898), .f ({\$dummy [22],\$dummy [23],gen_20_cmp_pMux_30,
                 gen_20_cmp_pMux_29,gen_20_cmp_pMux_28,gen_20_cmp_pMux_27,
                 gen_20_cmp_pMux_26,gen_20_cmp_pMux_25,gen_20_cmp_pMux_24,
                 gen_20_cmp_pMux_23,gen_20_cmp_pMux_22,gen_20_cmp_pMux_21,
                 gen_20_cmp_pMux_20,gen_20_cmp_pMux_19,gen_20_cmp_pMux_18,
                 gen_20_cmp_pMux_17,gen_20_cmp_pMux_16,gen_20_cmp_pMux_15,
                 gen_20_cmp_pMux_14,gen_20_cmp_pMux_13,gen_20_cmp_pMux_12,
                 gen_20_cmp_pMux_11,gen_20_cmp_pMux_10,gen_20_cmp_pMux_9,
                 gen_20_cmp_pMux_8,gen_20_cmp_pMux_7,gen_20_cmp_pMux_6,
                 gen_20_cmp_pMux_5,gen_20_cmp_pMux_4,gen_20_cmp_pMux_3,
                 gen_20_cmp_pMux_2,gen_20_cmp_pMux_1,gen_20_cmp_pMux_0})) ;
    NBitAdder_24 gen_20_cmp_BSCmp_AdderCmp (.a ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_20_cmp_pMux_30,gen_20_cmp_pMux_29,
                 gen_20_cmp_pMux_28,gen_20_cmp_pMux_27,gen_20_cmp_pMux_26,
                 gen_20_cmp_pMux_25,gen_20_cmp_pMux_24,gen_20_cmp_pMux_23,
                 gen_20_cmp_pMux_22,gen_20_cmp_pMux_21,gen_20_cmp_pMux_20,
                 gen_20_cmp_pMux_19,gen_20_cmp_pMux_18,gen_20_cmp_pMux_17,
                 gen_20_cmp_pMux_16,gen_20_cmp_pMux_15,gen_20_cmp_pMux_14,
                 gen_20_cmp_pMux_13,gen_20_cmp_pMux_12,gen_20_cmp_pMux_11,
                 gen_20_cmp_pMux_10,gen_20_cmp_pMux_9}), .b ({nx10482,nx10482,
                 nx10480,nx10488,nx10486,nx10484,nx10482,nx10480,
                 gen_20_cmp_BSCmp_op2_15,gen_20_cmp_BSCmp_op2_14,
                 gen_20_cmp_BSCmp_op2_13,gen_20_cmp_BSCmp_op2_12,
                 gen_20_cmp_BSCmp_op2_11,gen_20_cmp_BSCmp_op2_10,
                 gen_20_cmp_BSCmp_op2_9,gen_20_cmp_BSCmp_op2_8,
                 gen_20_cmp_BSCmp_op2_7,gen_20_cmp_BSCmp_op2_6,
                 gen_20_cmp_BSCmp_op2_5,gen_20_cmp_BSCmp_op2_4,
                 gen_20_cmp_BSCmp_op2_3,gen_20_cmp_BSCmp_op2_2,
                 gen_20_cmp_BSCmp_op2_1,gen_20_cmp_BSCmp_op2_0}), .carryIn (
                 gen_20_cmp_BSCmp_carryIn), .sum ({gen_20_cmp_pBs_30,
                 gen_20_cmp_pBs_29,gen_20_cmp_pBs_28,gen_20_cmp_pBs_27,
                 gen_20_cmp_pBs_26,gen_20_cmp_pBs_25,gen_20_cmp_pBs_24,
                 gen_20_cmp_pBs_23,outputs_20__15,outputs_20__14,outputs_20__13,
                 outputs_20__12,outputs_20__11,outputs_20__10,outputs_20__9,
                 outputs_20__8,outputs_20__7,outputs_20__6,outputs_20__5,
                 outputs_20__4,outputs_20__3,outputs_20__2,outputs_20__1,
                 outputs_20__0}), .carryOut (\$dummy [24])) ;
    Reg_33 gen_19_cmp_pRegCmp (.D ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
           gen_19_cmp_pBs_30,gen_19_cmp_pBs_29,gen_19_cmp_pBs_28,
           gen_19_cmp_pBs_27,gen_19_cmp_pBs_26,gen_19_cmp_pBs_25,
           gen_19_cmp_pBs_24,gen_19_cmp_pBs_23,outputs_19__15,outputs_19__14,
           outputs_19__13,outputs_19__12,outputs_19__11,outputs_19__10,
           outputs_19__9,outputs_19__8,outputs_19__7,outputs_19__6,outputs_19__5
           ,outputs_19__4,outputs_19__3,outputs_19__2,outputs_19__1,
           outputs_19__0,gen_19_cmp_pMux_8,gen_19_cmp_pMux_7,gen_19_cmp_pMux_6,
           gen_19_cmp_pMux_5,gen_19_cmp_pMux_4,gen_19_cmp_pMux_3,nx10190}), .en (
           nx11918), .clk (nx10122), .rst (rst), .Q ({\$dummy [25],\$dummy [26],
           gen_19_cmp_pReg_30,gen_19_cmp_pReg_29,gen_19_cmp_pReg_28,
           gen_19_cmp_pReg_27,gen_19_cmp_pReg_26,gen_19_cmp_pReg_25,
           gen_19_cmp_pReg_24,gen_19_cmp_pReg_23,gen_19_cmp_pReg_22,
           gen_19_cmp_pReg_21,gen_19_cmp_pReg_20,gen_19_cmp_pReg_19,
           gen_19_cmp_pReg_18,gen_19_cmp_pReg_17,gen_19_cmp_pReg_16,
           gen_19_cmp_pReg_15,gen_19_cmp_pReg_14,gen_19_cmp_pReg_13,
           gen_19_cmp_pReg_12,gen_19_cmp_pReg_11,gen_19_cmp_pReg_10,
           gen_19_cmp_pReg_9,gen_19_cmp_pReg_8,gen_19_cmp_pReg_7,
           gen_19_cmp_pReg_6,gen_19_cmp_pReg_5,gen_19_cmp_pReg_4,
           gen_19_cmp_pReg_3,gen_19_cmp_pReg_2,gen_19_cmp_pReg_1,
           gen_19_cmp_pReg_0})) ;
    BinaryMux_33 gen_19_cmp_MuxCmp (.a ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32
                 ,gen_19_cmp_pReg_30,gen_19_cmp_pReg_29,gen_19_cmp_pReg_28,
                 gen_19_cmp_pReg_27,gen_19_cmp_pReg_26,gen_19_cmp_pReg_25,
                 gen_19_cmp_pReg_24,gen_19_cmp_pReg_23,gen_19_cmp_pReg_22,
                 gen_19_cmp_pReg_21,gen_19_cmp_pReg_20,gen_19_cmp_pReg_19,
                 gen_19_cmp_pReg_18,gen_19_cmp_pReg_17,gen_19_cmp_pReg_16,
                 gen_19_cmp_pReg_15,gen_19_cmp_pReg_14,gen_19_cmp_pReg_13,
                 gen_19_cmp_pReg_12,gen_19_cmp_pReg_11,gen_19_cmp_pReg_10,
                 gen_19_cmp_pReg_9,gen_19_cmp_pReg_8,gen_19_cmp_pReg_7,
                 gen_19_cmp_pReg_6,gen_19_cmp_pReg_5,gen_19_cmp_pReg_4,
                 gen_19_cmp_pReg_3,gen_19_cmp_pReg_2,gen_19_cmp_pReg_1,
                 gen_19_cmp_pReg_0}), .b ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,filter_19__7,
                 filter_19__6,filter_19__5,filter_19__4,filter_19__3,
                 filter_19__2,filter_19__1,filter_19__0,gen_24_cmp_pInit_32}), .sel (
                 nx11898), .f ({\$dummy [27],\$dummy [28],gen_19_cmp_pMux_30,
                 gen_19_cmp_pMux_29,gen_19_cmp_pMux_28,gen_19_cmp_pMux_27,
                 gen_19_cmp_pMux_26,gen_19_cmp_pMux_25,gen_19_cmp_pMux_24,
                 gen_19_cmp_pMux_23,gen_19_cmp_pMux_22,gen_19_cmp_pMux_21,
                 gen_19_cmp_pMux_20,gen_19_cmp_pMux_19,gen_19_cmp_pMux_18,
                 gen_19_cmp_pMux_17,gen_19_cmp_pMux_16,gen_19_cmp_pMux_15,
                 gen_19_cmp_pMux_14,gen_19_cmp_pMux_13,gen_19_cmp_pMux_12,
                 gen_19_cmp_pMux_11,gen_19_cmp_pMux_10,gen_19_cmp_pMux_9,
                 gen_19_cmp_pMux_8,gen_19_cmp_pMux_7,gen_19_cmp_pMux_6,
                 gen_19_cmp_pMux_5,gen_19_cmp_pMux_4,gen_19_cmp_pMux_3,
                 gen_19_cmp_pMux_2,gen_19_cmp_pMux_1,gen_19_cmp_pMux_0})) ;
    NBitAdder_24 gen_19_cmp_BSCmp_AdderCmp (.a ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_19_cmp_pMux_30,gen_19_cmp_pMux_29,
                 gen_19_cmp_pMux_28,gen_19_cmp_pMux_27,gen_19_cmp_pMux_26,
                 gen_19_cmp_pMux_25,gen_19_cmp_pMux_24,gen_19_cmp_pMux_23,
                 gen_19_cmp_pMux_22,gen_19_cmp_pMux_21,gen_19_cmp_pMux_20,
                 gen_19_cmp_pMux_19,gen_19_cmp_pMux_18,gen_19_cmp_pMux_17,
                 gen_19_cmp_pMux_16,gen_19_cmp_pMux_15,gen_19_cmp_pMux_14,
                 gen_19_cmp_pMux_13,gen_19_cmp_pMux_12,gen_19_cmp_pMux_11,
                 gen_19_cmp_pMux_10,gen_19_cmp_pMux_9}), .b ({nx10494,nx10494,
                 nx10492,nx10500,nx10498,nx10496,nx10494,nx10492,
                 gen_19_cmp_BSCmp_op2_15,gen_19_cmp_BSCmp_op2_14,
                 gen_19_cmp_BSCmp_op2_13,gen_19_cmp_BSCmp_op2_12,
                 gen_19_cmp_BSCmp_op2_11,gen_19_cmp_BSCmp_op2_10,
                 gen_19_cmp_BSCmp_op2_9,gen_19_cmp_BSCmp_op2_8,
                 gen_19_cmp_BSCmp_op2_7,gen_19_cmp_BSCmp_op2_6,
                 gen_19_cmp_BSCmp_op2_5,gen_19_cmp_BSCmp_op2_4,
                 gen_19_cmp_BSCmp_op2_3,gen_19_cmp_BSCmp_op2_2,
                 gen_19_cmp_BSCmp_op2_1,gen_19_cmp_BSCmp_op2_0}), .carryIn (
                 gen_19_cmp_BSCmp_carryIn), .sum ({gen_19_cmp_pBs_30,
                 gen_19_cmp_pBs_29,gen_19_cmp_pBs_28,gen_19_cmp_pBs_27,
                 gen_19_cmp_pBs_26,gen_19_cmp_pBs_25,gen_19_cmp_pBs_24,
                 gen_19_cmp_pBs_23,outputs_19__15,outputs_19__14,outputs_19__13,
                 outputs_19__12,outputs_19__11,outputs_19__10,outputs_19__9,
                 outputs_19__8,outputs_19__7,outputs_19__6,outputs_19__5,
                 outputs_19__4,outputs_19__3,outputs_19__2,outputs_19__1,
                 outputs_19__0}), .carryOut (\$dummy [29])) ;
    Reg_33 gen_18_cmp_pRegCmp (.D ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
           gen_18_cmp_pBs_30,gen_18_cmp_pBs_29,gen_18_cmp_pBs_28,
           gen_18_cmp_pBs_27,gen_18_cmp_pBs_26,gen_18_cmp_pBs_25,
           gen_18_cmp_pBs_24,gen_18_cmp_pBs_23,outputs_18__15,outputs_18__14,
           outputs_18__13,outputs_18__12,outputs_18__11,outputs_18__10,
           outputs_18__9,outputs_18__8,outputs_18__7,outputs_18__6,outputs_18__5
           ,outputs_18__4,outputs_18__3,outputs_18__2,outputs_18__1,
           outputs_18__0,gen_18_cmp_pMux_8,gen_18_cmp_pMux_7,gen_18_cmp_pMux_6,
           gen_18_cmp_pMux_5,gen_18_cmp_pMux_4,gen_18_cmp_pMux_3,nx10202}), .en (
           nx10880), .clk (nx10122), .rst (rst), .Q ({\$dummy [30],\$dummy [31],
           gen_18_cmp_pReg_30,gen_18_cmp_pReg_29,gen_18_cmp_pReg_28,
           gen_18_cmp_pReg_27,gen_18_cmp_pReg_26,gen_18_cmp_pReg_25,
           gen_18_cmp_pReg_24,gen_18_cmp_pReg_23,gen_18_cmp_pReg_22,
           gen_18_cmp_pReg_21,gen_18_cmp_pReg_20,gen_18_cmp_pReg_19,
           gen_18_cmp_pReg_18,gen_18_cmp_pReg_17,gen_18_cmp_pReg_16,
           gen_18_cmp_pReg_15,gen_18_cmp_pReg_14,gen_18_cmp_pReg_13,
           gen_18_cmp_pReg_12,gen_18_cmp_pReg_11,gen_18_cmp_pReg_10,
           gen_18_cmp_pReg_9,gen_18_cmp_pReg_8,gen_18_cmp_pReg_7,
           gen_18_cmp_pReg_6,gen_18_cmp_pReg_5,gen_18_cmp_pReg_4,
           gen_18_cmp_pReg_3,gen_18_cmp_pReg_2,gen_18_cmp_pReg_1,
           gen_18_cmp_pReg_0})) ;
    BinaryMux_33 gen_18_cmp_MuxCmp (.a ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32
                 ,gen_18_cmp_pReg_30,gen_18_cmp_pReg_29,gen_18_cmp_pReg_28,
                 gen_18_cmp_pReg_27,gen_18_cmp_pReg_26,gen_18_cmp_pReg_25,
                 gen_18_cmp_pReg_24,gen_18_cmp_pReg_23,gen_18_cmp_pReg_22,
                 gen_18_cmp_pReg_21,gen_18_cmp_pReg_20,gen_18_cmp_pReg_19,
                 gen_18_cmp_pReg_18,gen_18_cmp_pReg_17,gen_18_cmp_pReg_16,
                 gen_18_cmp_pReg_15,gen_18_cmp_pReg_14,gen_18_cmp_pReg_13,
                 gen_18_cmp_pReg_12,gen_18_cmp_pReg_11,gen_18_cmp_pReg_10,
                 gen_18_cmp_pReg_9,gen_18_cmp_pReg_8,gen_18_cmp_pReg_7,
                 gen_18_cmp_pReg_6,gen_18_cmp_pReg_5,gen_18_cmp_pReg_4,
                 gen_18_cmp_pReg_3,gen_18_cmp_pReg_2,gen_18_cmp_pReg_1,
                 gen_18_cmp_pReg_0}), .b ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,filter_18__7,
                 filter_18__6,filter_18__5,filter_18__4,filter_18__3,
                 filter_18__2,filter_18__1,filter_18__0,gen_24_cmp_pInit_32}), .sel (
                 nx11900), .f ({\$dummy [32],\$dummy [33],gen_18_cmp_pMux_30,
                 gen_18_cmp_pMux_29,gen_18_cmp_pMux_28,gen_18_cmp_pMux_27,
                 gen_18_cmp_pMux_26,gen_18_cmp_pMux_25,gen_18_cmp_pMux_24,
                 gen_18_cmp_pMux_23,gen_18_cmp_pMux_22,gen_18_cmp_pMux_21,
                 gen_18_cmp_pMux_20,gen_18_cmp_pMux_19,gen_18_cmp_pMux_18,
                 gen_18_cmp_pMux_17,gen_18_cmp_pMux_16,gen_18_cmp_pMux_15,
                 gen_18_cmp_pMux_14,gen_18_cmp_pMux_13,gen_18_cmp_pMux_12,
                 gen_18_cmp_pMux_11,gen_18_cmp_pMux_10,gen_18_cmp_pMux_9,
                 gen_18_cmp_pMux_8,gen_18_cmp_pMux_7,gen_18_cmp_pMux_6,
                 gen_18_cmp_pMux_5,gen_18_cmp_pMux_4,gen_18_cmp_pMux_3,
                 gen_18_cmp_pMux_2,gen_18_cmp_pMux_1,gen_18_cmp_pMux_0})) ;
    NBitAdder_24 gen_18_cmp_BSCmp_AdderCmp (.a ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_18_cmp_pMux_30,gen_18_cmp_pMux_29,
                 gen_18_cmp_pMux_28,gen_18_cmp_pMux_27,gen_18_cmp_pMux_26,
                 gen_18_cmp_pMux_25,gen_18_cmp_pMux_24,gen_18_cmp_pMux_23,
                 gen_18_cmp_pMux_22,gen_18_cmp_pMux_21,gen_18_cmp_pMux_20,
                 gen_18_cmp_pMux_19,gen_18_cmp_pMux_18,gen_18_cmp_pMux_17,
                 gen_18_cmp_pMux_16,gen_18_cmp_pMux_15,gen_18_cmp_pMux_14,
                 gen_18_cmp_pMux_13,gen_18_cmp_pMux_12,gen_18_cmp_pMux_11,
                 gen_18_cmp_pMux_10,gen_18_cmp_pMux_9}), .b ({nx10506,nx10506,
                 nx10504,nx10512,nx10510,nx10508,nx10506,nx10504,
                 gen_18_cmp_BSCmp_op2_15,gen_18_cmp_BSCmp_op2_14,
                 gen_18_cmp_BSCmp_op2_13,gen_18_cmp_BSCmp_op2_12,
                 gen_18_cmp_BSCmp_op2_11,gen_18_cmp_BSCmp_op2_10,
                 gen_18_cmp_BSCmp_op2_9,gen_18_cmp_BSCmp_op2_8,
                 gen_18_cmp_BSCmp_op2_7,gen_18_cmp_BSCmp_op2_6,
                 gen_18_cmp_BSCmp_op2_5,gen_18_cmp_BSCmp_op2_4,
                 gen_18_cmp_BSCmp_op2_3,gen_18_cmp_BSCmp_op2_2,
                 gen_18_cmp_BSCmp_op2_1,gen_18_cmp_BSCmp_op2_0}), .carryIn (
                 gen_18_cmp_BSCmp_carryIn), .sum ({gen_18_cmp_pBs_30,
                 gen_18_cmp_pBs_29,gen_18_cmp_pBs_28,gen_18_cmp_pBs_27,
                 gen_18_cmp_pBs_26,gen_18_cmp_pBs_25,gen_18_cmp_pBs_24,
                 gen_18_cmp_pBs_23,outputs_18__15,outputs_18__14,outputs_18__13,
                 outputs_18__12,outputs_18__11,outputs_18__10,outputs_18__9,
                 outputs_18__8,outputs_18__7,outputs_18__6,outputs_18__5,
                 outputs_18__4,outputs_18__3,outputs_18__2,outputs_18__1,
                 outputs_18__0}), .carryOut (\$dummy [34])) ;
    Reg_33 gen_17_cmp_pRegCmp (.D ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
           gen_17_cmp_pBs_30,gen_17_cmp_pBs_29,gen_17_cmp_pBs_28,
           gen_17_cmp_pBs_27,gen_17_cmp_pBs_26,gen_17_cmp_pBs_25,
           gen_17_cmp_pBs_24,gen_17_cmp_pBs_23,outputs_17__15,outputs_17__14,
           outputs_17__13,outputs_17__12,outputs_17__11,outputs_17__10,
           outputs_17__9,outputs_17__8,outputs_17__7,outputs_17__6,outputs_17__5
           ,outputs_17__4,outputs_17__3,outputs_17__2,outputs_17__1,
           outputs_17__0,gen_17_cmp_pMux_8,gen_17_cmp_pMux_7,gen_17_cmp_pMux_6,
           gen_17_cmp_pMux_5,gen_17_cmp_pMux_4,gen_17_cmp_pMux_3,nx10214}), .en (
           nx11920), .clk (nx10124), .rst (rst), .Q ({\$dummy [35],\$dummy [36],
           gen_17_cmp_pReg_30,gen_17_cmp_pReg_29,gen_17_cmp_pReg_28,
           gen_17_cmp_pReg_27,gen_17_cmp_pReg_26,gen_17_cmp_pReg_25,
           gen_17_cmp_pReg_24,gen_17_cmp_pReg_23,gen_17_cmp_pReg_22,
           gen_17_cmp_pReg_21,gen_17_cmp_pReg_20,gen_17_cmp_pReg_19,
           gen_17_cmp_pReg_18,gen_17_cmp_pReg_17,gen_17_cmp_pReg_16,
           gen_17_cmp_pReg_15,gen_17_cmp_pReg_14,gen_17_cmp_pReg_13,
           gen_17_cmp_pReg_12,gen_17_cmp_pReg_11,gen_17_cmp_pReg_10,
           gen_17_cmp_pReg_9,gen_17_cmp_pReg_8,gen_17_cmp_pReg_7,
           gen_17_cmp_pReg_6,gen_17_cmp_pReg_5,gen_17_cmp_pReg_4,
           gen_17_cmp_pReg_3,gen_17_cmp_pReg_2,gen_17_cmp_pReg_1,
           gen_17_cmp_pReg_0})) ;
    BinaryMux_33 gen_17_cmp_MuxCmp (.a ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32
                 ,gen_17_cmp_pReg_30,gen_17_cmp_pReg_29,gen_17_cmp_pReg_28,
                 gen_17_cmp_pReg_27,gen_17_cmp_pReg_26,gen_17_cmp_pReg_25,
                 gen_17_cmp_pReg_24,gen_17_cmp_pReg_23,gen_17_cmp_pReg_22,
                 gen_17_cmp_pReg_21,gen_17_cmp_pReg_20,gen_17_cmp_pReg_19,
                 gen_17_cmp_pReg_18,gen_17_cmp_pReg_17,gen_17_cmp_pReg_16,
                 gen_17_cmp_pReg_15,gen_17_cmp_pReg_14,gen_17_cmp_pReg_13,
                 gen_17_cmp_pReg_12,gen_17_cmp_pReg_11,gen_17_cmp_pReg_10,
                 gen_17_cmp_pReg_9,gen_17_cmp_pReg_8,gen_17_cmp_pReg_7,
                 gen_17_cmp_pReg_6,gen_17_cmp_pReg_5,gen_17_cmp_pReg_4,
                 gen_17_cmp_pReg_3,gen_17_cmp_pReg_2,gen_17_cmp_pReg_1,
                 gen_17_cmp_pReg_0}), .b ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,filter_17__7,
                 filter_17__6,filter_17__5,filter_17__4,filter_17__3,
                 filter_17__2,filter_17__1,filter_17__0,gen_24_cmp_pInit_32}), .sel (
                 nx11902), .f ({\$dummy [37],\$dummy [38],gen_17_cmp_pMux_30,
                 gen_17_cmp_pMux_29,gen_17_cmp_pMux_28,gen_17_cmp_pMux_27,
                 gen_17_cmp_pMux_26,gen_17_cmp_pMux_25,gen_17_cmp_pMux_24,
                 gen_17_cmp_pMux_23,gen_17_cmp_pMux_22,gen_17_cmp_pMux_21,
                 gen_17_cmp_pMux_20,gen_17_cmp_pMux_19,gen_17_cmp_pMux_18,
                 gen_17_cmp_pMux_17,gen_17_cmp_pMux_16,gen_17_cmp_pMux_15,
                 gen_17_cmp_pMux_14,gen_17_cmp_pMux_13,gen_17_cmp_pMux_12,
                 gen_17_cmp_pMux_11,gen_17_cmp_pMux_10,gen_17_cmp_pMux_9,
                 gen_17_cmp_pMux_8,gen_17_cmp_pMux_7,gen_17_cmp_pMux_6,
                 gen_17_cmp_pMux_5,gen_17_cmp_pMux_4,gen_17_cmp_pMux_3,
                 gen_17_cmp_pMux_2,gen_17_cmp_pMux_1,gen_17_cmp_pMux_0})) ;
    NBitAdder_24 gen_17_cmp_BSCmp_AdderCmp (.a ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_17_cmp_pMux_30,gen_17_cmp_pMux_29,
                 gen_17_cmp_pMux_28,gen_17_cmp_pMux_27,gen_17_cmp_pMux_26,
                 gen_17_cmp_pMux_25,gen_17_cmp_pMux_24,gen_17_cmp_pMux_23,
                 gen_17_cmp_pMux_22,gen_17_cmp_pMux_21,gen_17_cmp_pMux_20,
                 gen_17_cmp_pMux_19,gen_17_cmp_pMux_18,gen_17_cmp_pMux_17,
                 gen_17_cmp_pMux_16,gen_17_cmp_pMux_15,gen_17_cmp_pMux_14,
                 gen_17_cmp_pMux_13,gen_17_cmp_pMux_12,gen_17_cmp_pMux_11,
                 gen_17_cmp_pMux_10,gen_17_cmp_pMux_9}), .b ({nx10518,nx10518,
                 nx10516,nx10524,nx10522,nx10520,nx10518,nx10516,
                 gen_17_cmp_BSCmp_op2_15,gen_17_cmp_BSCmp_op2_14,
                 gen_17_cmp_BSCmp_op2_13,gen_17_cmp_BSCmp_op2_12,
                 gen_17_cmp_BSCmp_op2_11,gen_17_cmp_BSCmp_op2_10,
                 gen_17_cmp_BSCmp_op2_9,gen_17_cmp_BSCmp_op2_8,
                 gen_17_cmp_BSCmp_op2_7,gen_17_cmp_BSCmp_op2_6,
                 gen_17_cmp_BSCmp_op2_5,gen_17_cmp_BSCmp_op2_4,
                 gen_17_cmp_BSCmp_op2_3,gen_17_cmp_BSCmp_op2_2,
                 gen_17_cmp_BSCmp_op2_1,gen_17_cmp_BSCmp_op2_0}), .carryIn (
                 gen_17_cmp_BSCmp_carryIn), .sum ({gen_17_cmp_pBs_30,
                 gen_17_cmp_pBs_29,gen_17_cmp_pBs_28,gen_17_cmp_pBs_27,
                 gen_17_cmp_pBs_26,gen_17_cmp_pBs_25,gen_17_cmp_pBs_24,
                 gen_17_cmp_pBs_23,outputs_17__15,outputs_17__14,outputs_17__13,
                 outputs_17__12,outputs_17__11,outputs_17__10,outputs_17__9,
                 outputs_17__8,outputs_17__7,outputs_17__6,outputs_17__5,
                 outputs_17__4,outputs_17__3,outputs_17__2,outputs_17__1,
                 outputs_17__0}), .carryOut (\$dummy [39])) ;
    Reg_33 gen_16_cmp_pRegCmp (.D ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
           gen_16_cmp_pBs_30,gen_16_cmp_pBs_29,gen_16_cmp_pBs_28,
           gen_16_cmp_pBs_27,gen_16_cmp_pBs_26,gen_16_cmp_pBs_25,
           gen_16_cmp_pBs_24,gen_16_cmp_pBs_23,outputs_16__15,outputs_16__14,
           outputs_16__13,outputs_16__12,outputs_16__11,outputs_16__10,
           outputs_16__9,outputs_16__8,outputs_16__7,outputs_16__6,outputs_16__5
           ,outputs_16__4,outputs_16__3,outputs_16__2,outputs_16__1,
           outputs_16__0,gen_16_cmp_pMux_8,gen_16_cmp_pMux_7,gen_16_cmp_pMux_6,
           gen_16_cmp_pMux_5,gen_16_cmp_pMux_4,gen_16_cmp_pMux_3,nx10226}), .en (
           nx11920), .clk (nx10124), .rst (rst), .Q ({\$dummy [40],\$dummy [41],
           gen_16_cmp_pReg_30,gen_16_cmp_pReg_29,gen_16_cmp_pReg_28,
           gen_16_cmp_pReg_27,gen_16_cmp_pReg_26,gen_16_cmp_pReg_25,
           gen_16_cmp_pReg_24,gen_16_cmp_pReg_23,gen_16_cmp_pReg_22,
           gen_16_cmp_pReg_21,gen_16_cmp_pReg_20,gen_16_cmp_pReg_19,
           gen_16_cmp_pReg_18,gen_16_cmp_pReg_17,gen_16_cmp_pReg_16,
           gen_16_cmp_pReg_15,gen_16_cmp_pReg_14,gen_16_cmp_pReg_13,
           gen_16_cmp_pReg_12,gen_16_cmp_pReg_11,gen_16_cmp_pReg_10,
           gen_16_cmp_pReg_9,gen_16_cmp_pReg_8,gen_16_cmp_pReg_7,
           gen_16_cmp_pReg_6,gen_16_cmp_pReg_5,gen_16_cmp_pReg_4,
           gen_16_cmp_pReg_3,gen_16_cmp_pReg_2,gen_16_cmp_pReg_1,
           gen_16_cmp_pReg_0})) ;
    BinaryMux_33 gen_16_cmp_MuxCmp (.a ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32
                 ,gen_16_cmp_pReg_30,gen_16_cmp_pReg_29,gen_16_cmp_pReg_28,
                 gen_16_cmp_pReg_27,gen_16_cmp_pReg_26,gen_16_cmp_pReg_25,
                 gen_16_cmp_pReg_24,gen_16_cmp_pReg_23,gen_16_cmp_pReg_22,
                 gen_16_cmp_pReg_21,gen_16_cmp_pReg_20,gen_16_cmp_pReg_19,
                 gen_16_cmp_pReg_18,gen_16_cmp_pReg_17,gen_16_cmp_pReg_16,
                 gen_16_cmp_pReg_15,gen_16_cmp_pReg_14,gen_16_cmp_pReg_13,
                 gen_16_cmp_pReg_12,gen_16_cmp_pReg_11,gen_16_cmp_pReg_10,
                 gen_16_cmp_pReg_9,gen_16_cmp_pReg_8,gen_16_cmp_pReg_7,
                 gen_16_cmp_pReg_6,gen_16_cmp_pReg_5,gen_16_cmp_pReg_4,
                 gen_16_cmp_pReg_3,gen_16_cmp_pReg_2,gen_16_cmp_pReg_1,
                 gen_16_cmp_pReg_0}), .b ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,filter_16__7,
                 filter_16__6,filter_16__5,filter_16__4,filter_16__3,
                 filter_16__2,filter_16__1,filter_16__0,gen_24_cmp_pInit_32}), .sel (
                 nx11902), .f ({\$dummy [42],\$dummy [43],gen_16_cmp_pMux_30,
                 gen_16_cmp_pMux_29,gen_16_cmp_pMux_28,gen_16_cmp_pMux_27,
                 gen_16_cmp_pMux_26,gen_16_cmp_pMux_25,gen_16_cmp_pMux_24,
                 gen_16_cmp_pMux_23,gen_16_cmp_pMux_22,gen_16_cmp_pMux_21,
                 gen_16_cmp_pMux_20,gen_16_cmp_pMux_19,gen_16_cmp_pMux_18,
                 gen_16_cmp_pMux_17,gen_16_cmp_pMux_16,gen_16_cmp_pMux_15,
                 gen_16_cmp_pMux_14,gen_16_cmp_pMux_13,gen_16_cmp_pMux_12,
                 gen_16_cmp_pMux_11,gen_16_cmp_pMux_10,gen_16_cmp_pMux_9,
                 gen_16_cmp_pMux_8,gen_16_cmp_pMux_7,gen_16_cmp_pMux_6,
                 gen_16_cmp_pMux_5,gen_16_cmp_pMux_4,gen_16_cmp_pMux_3,
                 gen_16_cmp_pMux_2,gen_16_cmp_pMux_1,gen_16_cmp_pMux_0})) ;
    NBitAdder_24 gen_16_cmp_BSCmp_AdderCmp (.a ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_16_cmp_pMux_30,gen_16_cmp_pMux_29,
                 gen_16_cmp_pMux_28,gen_16_cmp_pMux_27,gen_16_cmp_pMux_26,
                 gen_16_cmp_pMux_25,gen_16_cmp_pMux_24,gen_16_cmp_pMux_23,
                 gen_16_cmp_pMux_22,gen_16_cmp_pMux_21,gen_16_cmp_pMux_20,
                 gen_16_cmp_pMux_19,gen_16_cmp_pMux_18,gen_16_cmp_pMux_17,
                 gen_16_cmp_pMux_16,gen_16_cmp_pMux_15,gen_16_cmp_pMux_14,
                 gen_16_cmp_pMux_13,gen_16_cmp_pMux_12,gen_16_cmp_pMux_11,
                 gen_16_cmp_pMux_10,gen_16_cmp_pMux_9}), .b ({nx10530,nx10530,
                 nx10528,nx10536,nx10534,nx10532,nx10530,nx10528,
                 gen_16_cmp_BSCmp_op2_15,gen_16_cmp_BSCmp_op2_14,
                 gen_16_cmp_BSCmp_op2_13,gen_16_cmp_BSCmp_op2_12,
                 gen_16_cmp_BSCmp_op2_11,gen_16_cmp_BSCmp_op2_10,
                 gen_16_cmp_BSCmp_op2_9,gen_16_cmp_BSCmp_op2_8,
                 gen_16_cmp_BSCmp_op2_7,gen_16_cmp_BSCmp_op2_6,
                 gen_16_cmp_BSCmp_op2_5,gen_16_cmp_BSCmp_op2_4,
                 gen_16_cmp_BSCmp_op2_3,gen_16_cmp_BSCmp_op2_2,
                 gen_16_cmp_BSCmp_op2_1,gen_16_cmp_BSCmp_op2_0}), .carryIn (
                 gen_16_cmp_BSCmp_carryIn), .sum ({gen_16_cmp_pBs_30,
                 gen_16_cmp_pBs_29,gen_16_cmp_pBs_28,gen_16_cmp_pBs_27,
                 gen_16_cmp_pBs_26,gen_16_cmp_pBs_25,gen_16_cmp_pBs_24,
                 gen_16_cmp_pBs_23,outputs_16__15,outputs_16__14,outputs_16__13,
                 outputs_16__12,outputs_16__11,outputs_16__10,outputs_16__9,
                 outputs_16__8,outputs_16__7,outputs_16__6,outputs_16__5,
                 outputs_16__4,outputs_16__3,outputs_16__2,outputs_16__1,
                 outputs_16__0}), .carryOut (\$dummy [44])) ;
    Reg_33 gen_15_cmp_pRegCmp (.D ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
           gen_15_cmp_pBs_30,gen_15_cmp_pBs_29,gen_15_cmp_pBs_28,
           gen_15_cmp_pBs_27,gen_15_cmp_pBs_26,gen_15_cmp_pBs_25,
           gen_15_cmp_pBs_24,gen_15_cmp_pBs_23,outputs_15__15,outputs_15__14,
           outputs_15__13,outputs_15__12,outputs_15__11,outputs_15__10,
           outputs_15__9,outputs_15__8,outputs_15__7,outputs_15__6,outputs_15__5
           ,outputs_15__4,outputs_15__3,outputs_15__2,outputs_15__1,
           outputs_15__0,gen_15_cmp_pMux_8,gen_15_cmp_pMux_7,gen_15_cmp_pMux_6,
           gen_15_cmp_pMux_5,gen_15_cmp_pMux_4,gen_15_cmp_pMux_3,nx10238}), .en (
           nx11920), .clk (nx10124), .rst (rst), .Q ({\$dummy [45],\$dummy [46],
           gen_15_cmp_pReg_30,gen_15_cmp_pReg_29,gen_15_cmp_pReg_28,
           gen_15_cmp_pReg_27,gen_15_cmp_pReg_26,gen_15_cmp_pReg_25,
           gen_15_cmp_pReg_24,gen_15_cmp_pReg_23,gen_15_cmp_pReg_22,
           gen_15_cmp_pReg_21,gen_15_cmp_pReg_20,gen_15_cmp_pReg_19,
           gen_15_cmp_pReg_18,gen_15_cmp_pReg_17,gen_15_cmp_pReg_16,
           gen_15_cmp_pReg_15,gen_15_cmp_pReg_14,gen_15_cmp_pReg_13,
           gen_15_cmp_pReg_12,gen_15_cmp_pReg_11,gen_15_cmp_pReg_10,
           gen_15_cmp_pReg_9,gen_15_cmp_pReg_8,gen_15_cmp_pReg_7,
           gen_15_cmp_pReg_6,gen_15_cmp_pReg_5,gen_15_cmp_pReg_4,
           gen_15_cmp_pReg_3,gen_15_cmp_pReg_2,gen_15_cmp_pReg_1,
           gen_15_cmp_pReg_0})) ;
    BinaryMux_33 gen_15_cmp_MuxCmp (.a ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32
                 ,gen_15_cmp_pReg_30,gen_15_cmp_pReg_29,gen_15_cmp_pReg_28,
                 gen_15_cmp_pReg_27,gen_15_cmp_pReg_26,gen_15_cmp_pReg_25,
                 gen_15_cmp_pReg_24,gen_15_cmp_pReg_23,gen_15_cmp_pReg_22,
                 gen_15_cmp_pReg_21,gen_15_cmp_pReg_20,gen_15_cmp_pReg_19,
                 gen_15_cmp_pReg_18,gen_15_cmp_pReg_17,gen_15_cmp_pReg_16,
                 gen_15_cmp_pReg_15,gen_15_cmp_pReg_14,gen_15_cmp_pReg_13,
                 gen_15_cmp_pReg_12,gen_15_cmp_pReg_11,gen_15_cmp_pReg_10,
                 gen_15_cmp_pReg_9,gen_15_cmp_pReg_8,gen_15_cmp_pReg_7,
                 gen_15_cmp_pReg_6,gen_15_cmp_pReg_5,gen_15_cmp_pReg_4,
                 gen_15_cmp_pReg_3,gen_15_cmp_pReg_2,gen_15_cmp_pReg_1,
                 gen_15_cmp_pReg_0}), .b ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,filter_15__7,
                 filter_15__6,filter_15__5,filter_15__4,filter_15__3,
                 filter_15__2,filter_15__1,filter_15__0,gen_24_cmp_pInit_32}), .sel (
                 nx11902), .f ({\$dummy [47],\$dummy [48],gen_15_cmp_pMux_30,
                 gen_15_cmp_pMux_29,gen_15_cmp_pMux_28,gen_15_cmp_pMux_27,
                 gen_15_cmp_pMux_26,gen_15_cmp_pMux_25,gen_15_cmp_pMux_24,
                 gen_15_cmp_pMux_23,gen_15_cmp_pMux_22,gen_15_cmp_pMux_21,
                 gen_15_cmp_pMux_20,gen_15_cmp_pMux_19,gen_15_cmp_pMux_18,
                 gen_15_cmp_pMux_17,gen_15_cmp_pMux_16,gen_15_cmp_pMux_15,
                 gen_15_cmp_pMux_14,gen_15_cmp_pMux_13,gen_15_cmp_pMux_12,
                 gen_15_cmp_pMux_11,gen_15_cmp_pMux_10,gen_15_cmp_pMux_9,
                 gen_15_cmp_pMux_8,gen_15_cmp_pMux_7,gen_15_cmp_pMux_6,
                 gen_15_cmp_pMux_5,gen_15_cmp_pMux_4,gen_15_cmp_pMux_3,
                 gen_15_cmp_pMux_2,gen_15_cmp_pMux_1,gen_15_cmp_pMux_0})) ;
    NBitAdder_24 gen_15_cmp_BSCmp_AdderCmp (.a ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_15_cmp_pMux_30,gen_15_cmp_pMux_29,
                 gen_15_cmp_pMux_28,gen_15_cmp_pMux_27,gen_15_cmp_pMux_26,
                 gen_15_cmp_pMux_25,gen_15_cmp_pMux_24,gen_15_cmp_pMux_23,
                 gen_15_cmp_pMux_22,gen_15_cmp_pMux_21,gen_15_cmp_pMux_20,
                 gen_15_cmp_pMux_19,gen_15_cmp_pMux_18,gen_15_cmp_pMux_17,
                 gen_15_cmp_pMux_16,gen_15_cmp_pMux_15,gen_15_cmp_pMux_14,
                 gen_15_cmp_pMux_13,gen_15_cmp_pMux_12,gen_15_cmp_pMux_11,
                 gen_15_cmp_pMux_10,gen_15_cmp_pMux_9}), .b ({nx10542,nx10542,
                 nx10540,nx10548,nx10546,nx10544,nx10542,nx10540,
                 gen_15_cmp_BSCmp_op2_15,gen_15_cmp_BSCmp_op2_14,
                 gen_15_cmp_BSCmp_op2_13,gen_15_cmp_BSCmp_op2_12,
                 gen_15_cmp_BSCmp_op2_11,gen_15_cmp_BSCmp_op2_10,
                 gen_15_cmp_BSCmp_op2_9,gen_15_cmp_BSCmp_op2_8,
                 gen_15_cmp_BSCmp_op2_7,gen_15_cmp_BSCmp_op2_6,
                 gen_15_cmp_BSCmp_op2_5,gen_15_cmp_BSCmp_op2_4,
                 gen_15_cmp_BSCmp_op2_3,gen_15_cmp_BSCmp_op2_2,
                 gen_15_cmp_BSCmp_op2_1,gen_15_cmp_BSCmp_op2_0}), .carryIn (
                 gen_15_cmp_BSCmp_carryIn), .sum ({gen_15_cmp_pBs_30,
                 gen_15_cmp_pBs_29,gen_15_cmp_pBs_28,gen_15_cmp_pBs_27,
                 gen_15_cmp_pBs_26,gen_15_cmp_pBs_25,gen_15_cmp_pBs_24,
                 gen_15_cmp_pBs_23,outputs_15__15,outputs_15__14,outputs_15__13,
                 outputs_15__12,outputs_15__11,outputs_15__10,outputs_15__9,
                 outputs_15__8,outputs_15__7,outputs_15__6,outputs_15__5,
                 outputs_15__4,outputs_15__3,outputs_15__2,outputs_15__1,
                 outputs_15__0}), .carryOut (\$dummy [49])) ;
    Reg_33 gen_14_cmp_pRegCmp (.D ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
           gen_14_cmp_pBs_30,gen_14_cmp_pBs_29,gen_14_cmp_pBs_28,
           gen_14_cmp_pBs_27,gen_14_cmp_pBs_26,gen_14_cmp_pBs_25,
           gen_14_cmp_pBs_24,gen_14_cmp_pBs_23,outputs_14__15,outputs_14__14,
           outputs_14__13,outputs_14__12,outputs_14__11,outputs_14__10,
           outputs_14__9,outputs_14__8,outputs_14__7,outputs_14__6,outputs_14__5
           ,outputs_14__4,outputs_14__3,outputs_14__2,outputs_14__1,
           outputs_14__0,gen_14_cmp_pMux_8,gen_14_cmp_pMux_7,gen_14_cmp_pMux_6,
           gen_14_cmp_pMux_5,gen_14_cmp_pMux_4,gen_14_cmp_pMux_3,nx10250}), .en (
           nx11922), .clk (nx10124), .rst (rst), .Q ({\$dummy [50],\$dummy [51],
           gen_14_cmp_pReg_30,gen_14_cmp_pReg_29,gen_14_cmp_pReg_28,
           gen_14_cmp_pReg_27,gen_14_cmp_pReg_26,gen_14_cmp_pReg_25,
           gen_14_cmp_pReg_24,gen_14_cmp_pReg_23,gen_14_cmp_pReg_22,
           gen_14_cmp_pReg_21,gen_14_cmp_pReg_20,gen_14_cmp_pReg_19,
           gen_14_cmp_pReg_18,gen_14_cmp_pReg_17,gen_14_cmp_pReg_16,
           gen_14_cmp_pReg_15,gen_14_cmp_pReg_14,gen_14_cmp_pReg_13,
           gen_14_cmp_pReg_12,gen_14_cmp_pReg_11,gen_14_cmp_pReg_10,
           gen_14_cmp_pReg_9,gen_14_cmp_pReg_8,gen_14_cmp_pReg_7,
           gen_14_cmp_pReg_6,gen_14_cmp_pReg_5,gen_14_cmp_pReg_4,
           gen_14_cmp_pReg_3,gen_14_cmp_pReg_2,gen_14_cmp_pReg_1,
           gen_14_cmp_pReg_0})) ;
    BinaryMux_33 gen_14_cmp_MuxCmp (.a ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32
                 ,gen_14_cmp_pReg_30,gen_14_cmp_pReg_29,gen_14_cmp_pReg_28,
                 gen_14_cmp_pReg_27,gen_14_cmp_pReg_26,gen_14_cmp_pReg_25,
                 gen_14_cmp_pReg_24,gen_14_cmp_pReg_23,gen_14_cmp_pReg_22,
                 gen_14_cmp_pReg_21,gen_14_cmp_pReg_20,gen_14_cmp_pReg_19,
                 gen_14_cmp_pReg_18,gen_14_cmp_pReg_17,gen_14_cmp_pReg_16,
                 gen_14_cmp_pReg_15,gen_14_cmp_pReg_14,gen_14_cmp_pReg_13,
                 gen_14_cmp_pReg_12,gen_14_cmp_pReg_11,gen_14_cmp_pReg_10,
                 gen_14_cmp_pReg_9,gen_14_cmp_pReg_8,gen_14_cmp_pReg_7,
                 gen_14_cmp_pReg_6,gen_14_cmp_pReg_5,gen_14_cmp_pReg_4,
                 gen_14_cmp_pReg_3,gen_14_cmp_pReg_2,gen_14_cmp_pReg_1,
                 gen_14_cmp_pReg_0}), .b ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,filter_14__7,
                 filter_14__6,filter_14__5,filter_14__4,filter_14__3,
                 filter_14__2,filter_14__1,filter_14__0,gen_24_cmp_pInit_32}), .sel (
                 nx11904), .f ({\$dummy [52],\$dummy [53],gen_14_cmp_pMux_30,
                 gen_14_cmp_pMux_29,gen_14_cmp_pMux_28,gen_14_cmp_pMux_27,
                 gen_14_cmp_pMux_26,gen_14_cmp_pMux_25,gen_14_cmp_pMux_24,
                 gen_14_cmp_pMux_23,gen_14_cmp_pMux_22,gen_14_cmp_pMux_21,
                 gen_14_cmp_pMux_20,gen_14_cmp_pMux_19,gen_14_cmp_pMux_18,
                 gen_14_cmp_pMux_17,gen_14_cmp_pMux_16,gen_14_cmp_pMux_15,
                 gen_14_cmp_pMux_14,gen_14_cmp_pMux_13,gen_14_cmp_pMux_12,
                 gen_14_cmp_pMux_11,gen_14_cmp_pMux_10,gen_14_cmp_pMux_9,
                 gen_14_cmp_pMux_8,gen_14_cmp_pMux_7,gen_14_cmp_pMux_6,
                 gen_14_cmp_pMux_5,gen_14_cmp_pMux_4,gen_14_cmp_pMux_3,
                 gen_14_cmp_pMux_2,gen_14_cmp_pMux_1,gen_14_cmp_pMux_0})) ;
    NBitAdder_24 gen_14_cmp_BSCmp_AdderCmp (.a ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_14_cmp_pMux_30,gen_14_cmp_pMux_29,
                 gen_14_cmp_pMux_28,gen_14_cmp_pMux_27,gen_14_cmp_pMux_26,
                 gen_14_cmp_pMux_25,gen_14_cmp_pMux_24,gen_14_cmp_pMux_23,
                 gen_14_cmp_pMux_22,gen_14_cmp_pMux_21,gen_14_cmp_pMux_20,
                 gen_14_cmp_pMux_19,gen_14_cmp_pMux_18,gen_14_cmp_pMux_17,
                 gen_14_cmp_pMux_16,gen_14_cmp_pMux_15,gen_14_cmp_pMux_14,
                 gen_14_cmp_pMux_13,gen_14_cmp_pMux_12,gen_14_cmp_pMux_11,
                 gen_14_cmp_pMux_10,gen_14_cmp_pMux_9}), .b ({nx10554,nx10554,
                 nx10552,nx10560,nx10558,nx10556,nx10554,nx10552,
                 gen_14_cmp_BSCmp_op2_15,gen_14_cmp_BSCmp_op2_14,
                 gen_14_cmp_BSCmp_op2_13,gen_14_cmp_BSCmp_op2_12,
                 gen_14_cmp_BSCmp_op2_11,gen_14_cmp_BSCmp_op2_10,
                 gen_14_cmp_BSCmp_op2_9,gen_14_cmp_BSCmp_op2_8,
                 gen_14_cmp_BSCmp_op2_7,gen_14_cmp_BSCmp_op2_6,
                 gen_14_cmp_BSCmp_op2_5,gen_14_cmp_BSCmp_op2_4,
                 gen_14_cmp_BSCmp_op2_3,gen_14_cmp_BSCmp_op2_2,
                 gen_14_cmp_BSCmp_op2_1,gen_14_cmp_BSCmp_op2_0}), .carryIn (
                 gen_14_cmp_BSCmp_carryIn), .sum ({gen_14_cmp_pBs_30,
                 gen_14_cmp_pBs_29,gen_14_cmp_pBs_28,gen_14_cmp_pBs_27,
                 gen_14_cmp_pBs_26,gen_14_cmp_pBs_25,gen_14_cmp_pBs_24,
                 gen_14_cmp_pBs_23,outputs_14__15,outputs_14__14,outputs_14__13,
                 outputs_14__12,outputs_14__11,outputs_14__10,outputs_14__9,
                 outputs_14__8,outputs_14__7,outputs_14__6,outputs_14__5,
                 outputs_14__4,outputs_14__3,outputs_14__2,outputs_14__1,
                 outputs_14__0}), .carryOut (\$dummy [54])) ;
    Reg_33 gen_13_cmp_pRegCmp (.D ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
           gen_13_cmp_pBs_30,gen_13_cmp_pBs_29,gen_13_cmp_pBs_28,
           gen_13_cmp_pBs_27,gen_13_cmp_pBs_26,gen_13_cmp_pBs_25,
           gen_13_cmp_pBs_24,gen_13_cmp_pBs_23,outputs_13__15,outputs_13__14,
           outputs_13__13,outputs_13__12,outputs_13__11,outputs_13__10,
           outputs_13__9,outputs_13__8,outputs_13__7,outputs_13__6,outputs_13__5
           ,outputs_13__4,outputs_13__3,outputs_13__2,outputs_13__1,
           outputs_13__0,gen_13_cmp_pMux_8,gen_13_cmp_pMux_7,gen_13_cmp_pMux_6,
           gen_13_cmp_pMux_5,gen_13_cmp_pMux_4,gen_13_cmp_pMux_3,nx10262}), .en (
           nx11922), .clk (nx10124), .rst (rst), .Q ({\$dummy [55],\$dummy [56],
           gen_13_cmp_pReg_30,gen_13_cmp_pReg_29,gen_13_cmp_pReg_28,
           gen_13_cmp_pReg_27,gen_13_cmp_pReg_26,gen_13_cmp_pReg_25,
           gen_13_cmp_pReg_24,gen_13_cmp_pReg_23,gen_13_cmp_pReg_22,
           gen_13_cmp_pReg_21,gen_13_cmp_pReg_20,gen_13_cmp_pReg_19,
           gen_13_cmp_pReg_18,gen_13_cmp_pReg_17,gen_13_cmp_pReg_16,
           gen_13_cmp_pReg_15,gen_13_cmp_pReg_14,gen_13_cmp_pReg_13,
           gen_13_cmp_pReg_12,gen_13_cmp_pReg_11,gen_13_cmp_pReg_10,
           gen_13_cmp_pReg_9,gen_13_cmp_pReg_8,gen_13_cmp_pReg_7,
           gen_13_cmp_pReg_6,gen_13_cmp_pReg_5,gen_13_cmp_pReg_4,
           gen_13_cmp_pReg_3,gen_13_cmp_pReg_2,gen_13_cmp_pReg_1,
           gen_13_cmp_pReg_0})) ;
    BinaryMux_33 gen_13_cmp_MuxCmp (.a ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32
                 ,gen_13_cmp_pReg_30,gen_13_cmp_pReg_29,gen_13_cmp_pReg_28,
                 gen_13_cmp_pReg_27,gen_13_cmp_pReg_26,gen_13_cmp_pReg_25,
                 gen_13_cmp_pReg_24,gen_13_cmp_pReg_23,gen_13_cmp_pReg_22,
                 gen_13_cmp_pReg_21,gen_13_cmp_pReg_20,gen_13_cmp_pReg_19,
                 gen_13_cmp_pReg_18,gen_13_cmp_pReg_17,gen_13_cmp_pReg_16,
                 gen_13_cmp_pReg_15,gen_13_cmp_pReg_14,gen_13_cmp_pReg_13,
                 gen_13_cmp_pReg_12,gen_13_cmp_pReg_11,gen_13_cmp_pReg_10,
                 gen_13_cmp_pReg_9,gen_13_cmp_pReg_8,gen_13_cmp_pReg_7,
                 gen_13_cmp_pReg_6,gen_13_cmp_pReg_5,gen_13_cmp_pReg_4,
                 gen_13_cmp_pReg_3,gen_13_cmp_pReg_2,gen_13_cmp_pReg_1,
                 gen_13_cmp_pReg_0}), .b ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,filter_13__7,
                 filter_13__6,filter_13__5,filter_13__4,filter_13__3,
                 filter_13__2,filter_13__1,filter_13__0,gen_24_cmp_pInit_32}), .sel (
                 nx11904), .f ({\$dummy [57],\$dummy [58],gen_13_cmp_pMux_30,
                 gen_13_cmp_pMux_29,gen_13_cmp_pMux_28,gen_13_cmp_pMux_27,
                 gen_13_cmp_pMux_26,gen_13_cmp_pMux_25,gen_13_cmp_pMux_24,
                 gen_13_cmp_pMux_23,gen_13_cmp_pMux_22,gen_13_cmp_pMux_21,
                 gen_13_cmp_pMux_20,gen_13_cmp_pMux_19,gen_13_cmp_pMux_18,
                 gen_13_cmp_pMux_17,gen_13_cmp_pMux_16,gen_13_cmp_pMux_15,
                 gen_13_cmp_pMux_14,gen_13_cmp_pMux_13,gen_13_cmp_pMux_12,
                 gen_13_cmp_pMux_11,gen_13_cmp_pMux_10,gen_13_cmp_pMux_9,
                 gen_13_cmp_pMux_8,gen_13_cmp_pMux_7,gen_13_cmp_pMux_6,
                 gen_13_cmp_pMux_5,gen_13_cmp_pMux_4,gen_13_cmp_pMux_3,
                 gen_13_cmp_pMux_2,gen_13_cmp_pMux_1,gen_13_cmp_pMux_0})) ;
    NBitAdder_24 gen_13_cmp_BSCmp_AdderCmp (.a ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_13_cmp_pMux_30,gen_13_cmp_pMux_29,
                 gen_13_cmp_pMux_28,gen_13_cmp_pMux_27,gen_13_cmp_pMux_26,
                 gen_13_cmp_pMux_25,gen_13_cmp_pMux_24,gen_13_cmp_pMux_23,
                 gen_13_cmp_pMux_22,gen_13_cmp_pMux_21,gen_13_cmp_pMux_20,
                 gen_13_cmp_pMux_19,gen_13_cmp_pMux_18,gen_13_cmp_pMux_17,
                 gen_13_cmp_pMux_16,gen_13_cmp_pMux_15,gen_13_cmp_pMux_14,
                 gen_13_cmp_pMux_13,gen_13_cmp_pMux_12,gen_13_cmp_pMux_11,
                 gen_13_cmp_pMux_10,gen_13_cmp_pMux_9}), .b ({nx10566,nx10566,
                 nx10564,nx10572,nx10570,nx10568,nx10566,nx10564,
                 gen_13_cmp_BSCmp_op2_15,gen_13_cmp_BSCmp_op2_14,
                 gen_13_cmp_BSCmp_op2_13,gen_13_cmp_BSCmp_op2_12,
                 gen_13_cmp_BSCmp_op2_11,gen_13_cmp_BSCmp_op2_10,
                 gen_13_cmp_BSCmp_op2_9,gen_13_cmp_BSCmp_op2_8,
                 gen_13_cmp_BSCmp_op2_7,gen_13_cmp_BSCmp_op2_6,
                 gen_13_cmp_BSCmp_op2_5,gen_13_cmp_BSCmp_op2_4,
                 gen_13_cmp_BSCmp_op2_3,gen_13_cmp_BSCmp_op2_2,
                 gen_13_cmp_BSCmp_op2_1,gen_13_cmp_BSCmp_op2_0}), .carryIn (
                 gen_13_cmp_BSCmp_carryIn), .sum ({gen_13_cmp_pBs_30,
                 gen_13_cmp_pBs_29,gen_13_cmp_pBs_28,gen_13_cmp_pBs_27,
                 gen_13_cmp_pBs_26,gen_13_cmp_pBs_25,gen_13_cmp_pBs_24,
                 gen_13_cmp_pBs_23,outputs_13__15,outputs_13__14,outputs_13__13,
                 outputs_13__12,outputs_13__11,outputs_13__10,outputs_13__9,
                 outputs_13__8,outputs_13__7,outputs_13__6,outputs_13__5,
                 outputs_13__4,outputs_13__3,outputs_13__2,outputs_13__1,
                 outputs_13__0}), .carryOut (\$dummy [59])) ;
    Reg_33 gen_12_cmp_pRegCmp (.D ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
           gen_12_cmp_pBs_30,gen_12_cmp_pBs_29,gen_12_cmp_pBs_28,
           gen_12_cmp_pBs_27,gen_12_cmp_pBs_26,gen_12_cmp_pBs_25,
           gen_12_cmp_pBs_24,gen_12_cmp_pBs_23,outputs_12__15,outputs_12__14,
           outputs_12__13,outputs_12__12,outputs_12__11,outputs_12__10,
           outputs_12__9,outputs_12__8,outputs_12__7,outputs_12__6,outputs_12__5
           ,outputs_12__4,outputs_12__3,outputs_12__2,outputs_12__1,
           outputs_12__0,gen_12_cmp_pMux_8,gen_12_cmp_pMux_7,gen_12_cmp_pMux_6,
           gen_12_cmp_pMux_5,gen_12_cmp_pMux_4,gen_12_cmp_pMux_3,nx10274}), .en (
           nx11922), .clk (nx10124), .rst (rst), .Q ({\$dummy [60],\$dummy [61],
           gen_12_cmp_pReg_30,gen_12_cmp_pReg_29,gen_12_cmp_pReg_28,
           gen_12_cmp_pReg_27,gen_12_cmp_pReg_26,gen_12_cmp_pReg_25,
           gen_12_cmp_pReg_24,gen_12_cmp_pReg_23,gen_12_cmp_pReg_22,
           gen_12_cmp_pReg_21,gen_12_cmp_pReg_20,gen_12_cmp_pReg_19,
           gen_12_cmp_pReg_18,gen_12_cmp_pReg_17,gen_12_cmp_pReg_16,
           gen_12_cmp_pReg_15,gen_12_cmp_pReg_14,gen_12_cmp_pReg_13,
           gen_12_cmp_pReg_12,gen_12_cmp_pReg_11,gen_12_cmp_pReg_10,
           gen_12_cmp_pReg_9,gen_12_cmp_pReg_8,gen_12_cmp_pReg_7,
           gen_12_cmp_pReg_6,gen_12_cmp_pReg_5,gen_12_cmp_pReg_4,
           gen_12_cmp_pReg_3,gen_12_cmp_pReg_2,gen_12_cmp_pReg_1,
           gen_12_cmp_pReg_0})) ;
    BinaryMux_33 gen_12_cmp_MuxCmp (.a ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32
                 ,gen_12_cmp_pReg_30,gen_12_cmp_pReg_29,gen_12_cmp_pReg_28,
                 gen_12_cmp_pReg_27,gen_12_cmp_pReg_26,gen_12_cmp_pReg_25,
                 gen_12_cmp_pReg_24,gen_12_cmp_pReg_23,gen_12_cmp_pReg_22,
                 gen_12_cmp_pReg_21,gen_12_cmp_pReg_20,gen_12_cmp_pReg_19,
                 gen_12_cmp_pReg_18,gen_12_cmp_pReg_17,gen_12_cmp_pReg_16,
                 gen_12_cmp_pReg_15,gen_12_cmp_pReg_14,gen_12_cmp_pReg_13,
                 gen_12_cmp_pReg_12,gen_12_cmp_pReg_11,gen_12_cmp_pReg_10,
                 gen_12_cmp_pReg_9,gen_12_cmp_pReg_8,gen_12_cmp_pReg_7,
                 gen_12_cmp_pReg_6,gen_12_cmp_pReg_5,gen_12_cmp_pReg_4,
                 gen_12_cmp_pReg_3,gen_12_cmp_pReg_2,gen_12_cmp_pReg_1,
                 gen_12_cmp_pReg_0}), .b ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,filter_12__7,
                 filter_12__6,filter_12__5,filter_12__4,filter_12__3,
                 filter_12__2,filter_12__1,filter_12__0,gen_24_cmp_pInit_32}), .sel (
                 nx11904), .f ({\$dummy [62],\$dummy [63],gen_12_cmp_pMux_30,
                 gen_12_cmp_pMux_29,gen_12_cmp_pMux_28,gen_12_cmp_pMux_27,
                 gen_12_cmp_pMux_26,gen_12_cmp_pMux_25,gen_12_cmp_pMux_24,
                 gen_12_cmp_pMux_23,gen_12_cmp_pMux_22,gen_12_cmp_pMux_21,
                 gen_12_cmp_pMux_20,gen_12_cmp_pMux_19,gen_12_cmp_pMux_18,
                 gen_12_cmp_pMux_17,gen_12_cmp_pMux_16,gen_12_cmp_pMux_15,
                 gen_12_cmp_pMux_14,gen_12_cmp_pMux_13,gen_12_cmp_pMux_12,
                 gen_12_cmp_pMux_11,gen_12_cmp_pMux_10,gen_12_cmp_pMux_9,
                 gen_12_cmp_pMux_8,gen_12_cmp_pMux_7,gen_12_cmp_pMux_6,
                 gen_12_cmp_pMux_5,gen_12_cmp_pMux_4,gen_12_cmp_pMux_3,
                 gen_12_cmp_pMux_2,gen_12_cmp_pMux_1,gen_12_cmp_pMux_0})) ;
    NBitAdder_24 gen_12_cmp_BSCmp_AdderCmp (.a ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_12_cmp_pMux_30,gen_12_cmp_pMux_29,
                 gen_12_cmp_pMux_28,gen_12_cmp_pMux_27,gen_12_cmp_pMux_26,
                 gen_12_cmp_pMux_25,gen_12_cmp_pMux_24,gen_12_cmp_pMux_23,
                 gen_12_cmp_pMux_22,gen_12_cmp_pMux_21,gen_12_cmp_pMux_20,
                 gen_12_cmp_pMux_19,gen_12_cmp_pMux_18,gen_12_cmp_pMux_17,
                 gen_12_cmp_pMux_16,gen_12_cmp_pMux_15,gen_12_cmp_pMux_14,
                 gen_12_cmp_pMux_13,gen_12_cmp_pMux_12,gen_12_cmp_pMux_11,
                 gen_12_cmp_pMux_10,gen_12_cmp_pMux_9}), .b ({nx10578,nx10578,
                 nx10576,nx10584,nx10582,nx10580,nx10578,nx10576,
                 gen_12_cmp_BSCmp_op2_15,gen_12_cmp_BSCmp_op2_14,
                 gen_12_cmp_BSCmp_op2_13,gen_12_cmp_BSCmp_op2_12,
                 gen_12_cmp_BSCmp_op2_11,gen_12_cmp_BSCmp_op2_10,
                 gen_12_cmp_BSCmp_op2_9,gen_12_cmp_BSCmp_op2_8,
                 gen_12_cmp_BSCmp_op2_7,gen_12_cmp_BSCmp_op2_6,
                 gen_12_cmp_BSCmp_op2_5,gen_12_cmp_BSCmp_op2_4,
                 gen_12_cmp_BSCmp_op2_3,gen_12_cmp_BSCmp_op2_2,
                 gen_12_cmp_BSCmp_op2_1,gen_12_cmp_BSCmp_op2_0}), .carryIn (
                 gen_12_cmp_BSCmp_carryIn), .sum ({gen_12_cmp_pBs_30,
                 gen_12_cmp_pBs_29,gen_12_cmp_pBs_28,gen_12_cmp_pBs_27,
                 gen_12_cmp_pBs_26,gen_12_cmp_pBs_25,gen_12_cmp_pBs_24,
                 gen_12_cmp_pBs_23,outputs_12__15,outputs_12__14,outputs_12__13,
                 outputs_12__12,outputs_12__11,outputs_12__10,outputs_12__9,
                 outputs_12__8,outputs_12__7,outputs_12__6,outputs_12__5,
                 outputs_12__4,outputs_12__3,outputs_12__2,outputs_12__1,
                 outputs_12__0}), .carryOut (\$dummy [64])) ;
    Reg_33 gen_11_cmp_pRegCmp (.D ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
           gen_11_cmp_pBs_30,gen_11_cmp_pBs_29,gen_11_cmp_pBs_28,
           gen_11_cmp_pBs_27,gen_11_cmp_pBs_26,gen_11_cmp_pBs_25,
           gen_11_cmp_pBs_24,gen_11_cmp_pBs_23,outputs_11__15,outputs_11__14,
           outputs_11__13,outputs_11__12,outputs_11__11,outputs_11__10,
           outputs_11__9,outputs_11__8,outputs_11__7,outputs_11__6,outputs_11__5
           ,outputs_11__4,outputs_11__3,outputs_11__2,outputs_11__1,
           outputs_11__0,gen_11_cmp_pMux_8,gen_11_cmp_pMux_7,gen_11_cmp_pMux_6,
           gen_11_cmp_pMux_5,gen_11_cmp_pMux_4,gen_11_cmp_pMux_3,nx10286}), .en (
           nx10882), .clk (nx10124), .rst (rst), .Q ({\$dummy [65],\$dummy [66],
           gen_11_cmp_pReg_30,gen_11_cmp_pReg_29,gen_11_cmp_pReg_28,
           gen_11_cmp_pReg_27,gen_11_cmp_pReg_26,gen_11_cmp_pReg_25,
           gen_11_cmp_pReg_24,gen_11_cmp_pReg_23,gen_11_cmp_pReg_22,
           gen_11_cmp_pReg_21,gen_11_cmp_pReg_20,gen_11_cmp_pReg_19,
           gen_11_cmp_pReg_18,gen_11_cmp_pReg_17,gen_11_cmp_pReg_16,
           gen_11_cmp_pReg_15,gen_11_cmp_pReg_14,gen_11_cmp_pReg_13,
           gen_11_cmp_pReg_12,gen_11_cmp_pReg_11,gen_11_cmp_pReg_10,
           gen_11_cmp_pReg_9,gen_11_cmp_pReg_8,gen_11_cmp_pReg_7,
           gen_11_cmp_pReg_6,gen_11_cmp_pReg_5,gen_11_cmp_pReg_4,
           gen_11_cmp_pReg_3,gen_11_cmp_pReg_2,gen_11_cmp_pReg_1,
           gen_11_cmp_pReg_0})) ;
    BinaryMux_33 gen_11_cmp_MuxCmp (.a ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32
                 ,gen_11_cmp_pReg_30,gen_11_cmp_pReg_29,gen_11_cmp_pReg_28,
                 gen_11_cmp_pReg_27,gen_11_cmp_pReg_26,gen_11_cmp_pReg_25,
                 gen_11_cmp_pReg_24,gen_11_cmp_pReg_23,gen_11_cmp_pReg_22,
                 gen_11_cmp_pReg_21,gen_11_cmp_pReg_20,gen_11_cmp_pReg_19,
                 gen_11_cmp_pReg_18,gen_11_cmp_pReg_17,gen_11_cmp_pReg_16,
                 gen_11_cmp_pReg_15,gen_11_cmp_pReg_14,gen_11_cmp_pReg_13,
                 gen_11_cmp_pReg_12,gen_11_cmp_pReg_11,gen_11_cmp_pReg_10,
                 gen_11_cmp_pReg_9,gen_11_cmp_pReg_8,gen_11_cmp_pReg_7,
                 gen_11_cmp_pReg_6,gen_11_cmp_pReg_5,gen_11_cmp_pReg_4,
                 gen_11_cmp_pReg_3,gen_11_cmp_pReg_2,gen_11_cmp_pReg_1,
                 gen_11_cmp_pReg_0}), .b ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,filter_11__7,
                 filter_11__6,filter_11__5,filter_11__4,filter_11__3,
                 filter_11__2,filter_11__1,filter_11__0,gen_24_cmp_pInit_32}), .sel (
                 nx11906), .f ({\$dummy [67],\$dummy [68],gen_11_cmp_pMux_30,
                 gen_11_cmp_pMux_29,gen_11_cmp_pMux_28,gen_11_cmp_pMux_27,
                 gen_11_cmp_pMux_26,gen_11_cmp_pMux_25,gen_11_cmp_pMux_24,
                 gen_11_cmp_pMux_23,gen_11_cmp_pMux_22,gen_11_cmp_pMux_21,
                 gen_11_cmp_pMux_20,gen_11_cmp_pMux_19,gen_11_cmp_pMux_18,
                 gen_11_cmp_pMux_17,gen_11_cmp_pMux_16,gen_11_cmp_pMux_15,
                 gen_11_cmp_pMux_14,gen_11_cmp_pMux_13,gen_11_cmp_pMux_12,
                 gen_11_cmp_pMux_11,gen_11_cmp_pMux_10,gen_11_cmp_pMux_9,
                 gen_11_cmp_pMux_8,gen_11_cmp_pMux_7,gen_11_cmp_pMux_6,
                 gen_11_cmp_pMux_5,gen_11_cmp_pMux_4,gen_11_cmp_pMux_3,
                 gen_11_cmp_pMux_2,gen_11_cmp_pMux_1,gen_11_cmp_pMux_0})) ;
    NBitAdder_24 gen_11_cmp_BSCmp_AdderCmp (.a ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_11_cmp_pMux_30,gen_11_cmp_pMux_29,
                 gen_11_cmp_pMux_28,gen_11_cmp_pMux_27,gen_11_cmp_pMux_26,
                 gen_11_cmp_pMux_25,gen_11_cmp_pMux_24,gen_11_cmp_pMux_23,
                 gen_11_cmp_pMux_22,gen_11_cmp_pMux_21,gen_11_cmp_pMux_20,
                 gen_11_cmp_pMux_19,gen_11_cmp_pMux_18,gen_11_cmp_pMux_17,
                 gen_11_cmp_pMux_16,gen_11_cmp_pMux_15,gen_11_cmp_pMux_14,
                 gen_11_cmp_pMux_13,gen_11_cmp_pMux_12,gen_11_cmp_pMux_11,
                 gen_11_cmp_pMux_10,gen_11_cmp_pMux_9}), .b ({nx10590,nx10590,
                 nx10588,nx10596,nx10594,nx10592,nx10590,nx10588,
                 gen_11_cmp_BSCmp_op2_15,gen_11_cmp_BSCmp_op2_14,
                 gen_11_cmp_BSCmp_op2_13,gen_11_cmp_BSCmp_op2_12,
                 gen_11_cmp_BSCmp_op2_11,gen_11_cmp_BSCmp_op2_10,
                 gen_11_cmp_BSCmp_op2_9,gen_11_cmp_BSCmp_op2_8,
                 gen_11_cmp_BSCmp_op2_7,gen_11_cmp_BSCmp_op2_6,
                 gen_11_cmp_BSCmp_op2_5,gen_11_cmp_BSCmp_op2_4,
                 gen_11_cmp_BSCmp_op2_3,gen_11_cmp_BSCmp_op2_2,
                 gen_11_cmp_BSCmp_op2_1,gen_11_cmp_BSCmp_op2_0}), .carryIn (
                 gen_11_cmp_BSCmp_carryIn), .sum ({gen_11_cmp_pBs_30,
                 gen_11_cmp_pBs_29,gen_11_cmp_pBs_28,gen_11_cmp_pBs_27,
                 gen_11_cmp_pBs_26,gen_11_cmp_pBs_25,gen_11_cmp_pBs_24,
                 gen_11_cmp_pBs_23,outputs_11__15,outputs_11__14,outputs_11__13,
                 outputs_11__12,outputs_11__11,outputs_11__10,outputs_11__9,
                 outputs_11__8,outputs_11__7,outputs_11__6,outputs_11__5,
                 outputs_11__4,outputs_11__3,outputs_11__2,outputs_11__1,
                 outputs_11__0}), .carryOut (\$dummy [69])) ;
    Reg_33 gen_10_cmp_pRegCmp (.D ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
           gen_10_cmp_pBs_30,gen_10_cmp_pBs_29,gen_10_cmp_pBs_28,
           gen_10_cmp_pBs_27,gen_10_cmp_pBs_26,gen_10_cmp_pBs_25,
           gen_10_cmp_pBs_24,gen_10_cmp_pBs_23,outputs_10__15,outputs_10__14,
           outputs_10__13,outputs_10__12,outputs_10__11,outputs_10__10,
           outputs_10__9,outputs_10__8,outputs_10__7,outputs_10__6,outputs_10__5
           ,outputs_10__4,outputs_10__3,outputs_10__2,outputs_10__1,
           outputs_10__0,gen_10_cmp_pMux_8,gen_10_cmp_pMux_7,gen_10_cmp_pMux_6,
           gen_10_cmp_pMux_5,gen_10_cmp_pMux_4,gen_10_cmp_pMux_3,nx10298}), .en (
           nx11924), .clk (nx10126), .rst (rst), .Q ({\$dummy [70],\$dummy [71],
           gen_10_cmp_pReg_30,gen_10_cmp_pReg_29,gen_10_cmp_pReg_28,
           gen_10_cmp_pReg_27,gen_10_cmp_pReg_26,gen_10_cmp_pReg_25,
           gen_10_cmp_pReg_24,gen_10_cmp_pReg_23,gen_10_cmp_pReg_22,
           gen_10_cmp_pReg_21,gen_10_cmp_pReg_20,gen_10_cmp_pReg_19,
           gen_10_cmp_pReg_18,gen_10_cmp_pReg_17,gen_10_cmp_pReg_16,
           gen_10_cmp_pReg_15,gen_10_cmp_pReg_14,gen_10_cmp_pReg_13,
           gen_10_cmp_pReg_12,gen_10_cmp_pReg_11,gen_10_cmp_pReg_10,
           gen_10_cmp_pReg_9,gen_10_cmp_pReg_8,gen_10_cmp_pReg_7,
           gen_10_cmp_pReg_6,gen_10_cmp_pReg_5,gen_10_cmp_pReg_4,
           gen_10_cmp_pReg_3,gen_10_cmp_pReg_2,gen_10_cmp_pReg_1,
           gen_10_cmp_pReg_0})) ;
    BinaryMux_33 gen_10_cmp_MuxCmp (.a ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32
                 ,gen_10_cmp_pReg_30,gen_10_cmp_pReg_29,gen_10_cmp_pReg_28,
                 gen_10_cmp_pReg_27,gen_10_cmp_pReg_26,gen_10_cmp_pReg_25,
                 gen_10_cmp_pReg_24,gen_10_cmp_pReg_23,gen_10_cmp_pReg_22,
                 gen_10_cmp_pReg_21,gen_10_cmp_pReg_20,gen_10_cmp_pReg_19,
                 gen_10_cmp_pReg_18,gen_10_cmp_pReg_17,gen_10_cmp_pReg_16,
                 gen_10_cmp_pReg_15,gen_10_cmp_pReg_14,gen_10_cmp_pReg_13,
                 gen_10_cmp_pReg_12,gen_10_cmp_pReg_11,gen_10_cmp_pReg_10,
                 gen_10_cmp_pReg_9,gen_10_cmp_pReg_8,gen_10_cmp_pReg_7,
                 gen_10_cmp_pReg_6,gen_10_cmp_pReg_5,gen_10_cmp_pReg_4,
                 gen_10_cmp_pReg_3,gen_10_cmp_pReg_2,gen_10_cmp_pReg_1,
                 gen_10_cmp_pReg_0}), .b ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,filter_10__7,
                 filter_10__6,filter_10__5,filter_10__4,filter_10__3,
                 filter_10__2,filter_10__1,filter_10__0,gen_24_cmp_pInit_32}), .sel (
                 nx11908), .f ({\$dummy [72],\$dummy [73],gen_10_cmp_pMux_30,
                 gen_10_cmp_pMux_29,gen_10_cmp_pMux_28,gen_10_cmp_pMux_27,
                 gen_10_cmp_pMux_26,gen_10_cmp_pMux_25,gen_10_cmp_pMux_24,
                 gen_10_cmp_pMux_23,gen_10_cmp_pMux_22,gen_10_cmp_pMux_21,
                 gen_10_cmp_pMux_20,gen_10_cmp_pMux_19,gen_10_cmp_pMux_18,
                 gen_10_cmp_pMux_17,gen_10_cmp_pMux_16,gen_10_cmp_pMux_15,
                 gen_10_cmp_pMux_14,gen_10_cmp_pMux_13,gen_10_cmp_pMux_12,
                 gen_10_cmp_pMux_11,gen_10_cmp_pMux_10,gen_10_cmp_pMux_9,
                 gen_10_cmp_pMux_8,gen_10_cmp_pMux_7,gen_10_cmp_pMux_6,
                 gen_10_cmp_pMux_5,gen_10_cmp_pMux_4,gen_10_cmp_pMux_3,
                 gen_10_cmp_pMux_2,gen_10_cmp_pMux_1,gen_10_cmp_pMux_0})) ;
    NBitAdder_24 gen_10_cmp_BSCmp_AdderCmp (.a ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_10_cmp_pMux_30,gen_10_cmp_pMux_29,
                 gen_10_cmp_pMux_28,gen_10_cmp_pMux_27,gen_10_cmp_pMux_26,
                 gen_10_cmp_pMux_25,gen_10_cmp_pMux_24,gen_10_cmp_pMux_23,
                 gen_10_cmp_pMux_22,gen_10_cmp_pMux_21,gen_10_cmp_pMux_20,
                 gen_10_cmp_pMux_19,gen_10_cmp_pMux_18,gen_10_cmp_pMux_17,
                 gen_10_cmp_pMux_16,gen_10_cmp_pMux_15,gen_10_cmp_pMux_14,
                 gen_10_cmp_pMux_13,gen_10_cmp_pMux_12,gen_10_cmp_pMux_11,
                 gen_10_cmp_pMux_10,gen_10_cmp_pMux_9}), .b ({nx10602,nx10602,
                 nx10600,nx10608,nx10606,nx10604,nx10602,nx10600,
                 gen_10_cmp_BSCmp_op2_15,gen_10_cmp_BSCmp_op2_14,
                 gen_10_cmp_BSCmp_op2_13,gen_10_cmp_BSCmp_op2_12,
                 gen_10_cmp_BSCmp_op2_11,gen_10_cmp_BSCmp_op2_10,
                 gen_10_cmp_BSCmp_op2_9,gen_10_cmp_BSCmp_op2_8,
                 gen_10_cmp_BSCmp_op2_7,gen_10_cmp_BSCmp_op2_6,
                 gen_10_cmp_BSCmp_op2_5,gen_10_cmp_BSCmp_op2_4,
                 gen_10_cmp_BSCmp_op2_3,gen_10_cmp_BSCmp_op2_2,
                 gen_10_cmp_BSCmp_op2_1,gen_10_cmp_BSCmp_op2_0}), .carryIn (
                 gen_10_cmp_BSCmp_carryIn), .sum ({gen_10_cmp_pBs_30,
                 gen_10_cmp_pBs_29,gen_10_cmp_pBs_28,gen_10_cmp_pBs_27,
                 gen_10_cmp_pBs_26,gen_10_cmp_pBs_25,gen_10_cmp_pBs_24,
                 gen_10_cmp_pBs_23,outputs_10__15,outputs_10__14,outputs_10__13,
                 outputs_10__12,outputs_10__11,outputs_10__10,outputs_10__9,
                 outputs_10__8,outputs_10__7,outputs_10__6,outputs_10__5,
                 outputs_10__4,outputs_10__3,outputs_10__2,outputs_10__1,
                 outputs_10__0}), .carryOut (\$dummy [74])) ;
    Reg_33 gen_9_cmp_pRegCmp (.D ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
           gen_9_cmp_pBs_30,gen_9_cmp_pBs_29,gen_9_cmp_pBs_28,gen_9_cmp_pBs_27,
           gen_9_cmp_pBs_26,gen_9_cmp_pBs_25,gen_9_cmp_pBs_24,gen_9_cmp_pBs_23,
           outputs_9__15,outputs_9__14,outputs_9__13,outputs_9__12,outputs_9__11
           ,outputs_9__10,outputs_9__9,outputs_9__8,outputs_9__7,outputs_9__6,
           outputs_9__5,outputs_9__4,outputs_9__3,outputs_9__2,outputs_9__1,
           outputs_9__0,gen_9_cmp_pMux_8,gen_9_cmp_pMux_7,gen_9_cmp_pMux_6,
           gen_9_cmp_pMux_5,gen_9_cmp_pMux_4,gen_9_cmp_pMux_3,nx10310}), .en (
           nx11924), .clk (nx10126), .rst (rst), .Q ({\$dummy [75],\$dummy [76],
           gen_9_cmp_pReg_30,gen_9_cmp_pReg_29,gen_9_cmp_pReg_28,
           gen_9_cmp_pReg_27,gen_9_cmp_pReg_26,gen_9_cmp_pReg_25,
           gen_9_cmp_pReg_24,gen_9_cmp_pReg_23,gen_9_cmp_pReg_22,
           gen_9_cmp_pReg_21,gen_9_cmp_pReg_20,gen_9_cmp_pReg_19,
           gen_9_cmp_pReg_18,gen_9_cmp_pReg_17,gen_9_cmp_pReg_16,
           gen_9_cmp_pReg_15,gen_9_cmp_pReg_14,gen_9_cmp_pReg_13,
           gen_9_cmp_pReg_12,gen_9_cmp_pReg_11,gen_9_cmp_pReg_10,
           gen_9_cmp_pReg_9,gen_9_cmp_pReg_8,gen_9_cmp_pReg_7,gen_9_cmp_pReg_6,
           gen_9_cmp_pReg_5,gen_9_cmp_pReg_4,gen_9_cmp_pReg_3,gen_9_cmp_pReg_2,
           gen_9_cmp_pReg_1,gen_9_cmp_pReg_0})) ;
    BinaryMux_33 gen_9_cmp_MuxCmp (.a ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_9_cmp_pReg_30,gen_9_cmp_pReg_29,gen_9_cmp_pReg_28,
                 gen_9_cmp_pReg_27,gen_9_cmp_pReg_26,gen_9_cmp_pReg_25,
                 gen_9_cmp_pReg_24,gen_9_cmp_pReg_23,gen_9_cmp_pReg_22,
                 gen_9_cmp_pReg_21,gen_9_cmp_pReg_20,gen_9_cmp_pReg_19,
                 gen_9_cmp_pReg_18,gen_9_cmp_pReg_17,gen_9_cmp_pReg_16,
                 gen_9_cmp_pReg_15,gen_9_cmp_pReg_14,gen_9_cmp_pReg_13,
                 gen_9_cmp_pReg_12,gen_9_cmp_pReg_11,gen_9_cmp_pReg_10,
                 gen_9_cmp_pReg_9,gen_9_cmp_pReg_8,gen_9_cmp_pReg_7,
                 gen_9_cmp_pReg_6,gen_9_cmp_pReg_5,gen_9_cmp_pReg_4,
                 gen_9_cmp_pReg_3,gen_9_cmp_pReg_2,gen_9_cmp_pReg_1,
                 gen_9_cmp_pReg_0}), .b ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,filter_9__7,filter_9__6
                 ,filter_9__5,filter_9__4,filter_9__3,filter_9__2,filter_9__1,
                 filter_9__0,gen_24_cmp_pInit_32}), .sel (nx11908), .f ({
                 \$dummy [77],\$dummy [78],gen_9_cmp_pMux_30,gen_9_cmp_pMux_29,
                 gen_9_cmp_pMux_28,gen_9_cmp_pMux_27,gen_9_cmp_pMux_26,
                 gen_9_cmp_pMux_25,gen_9_cmp_pMux_24,gen_9_cmp_pMux_23,
                 gen_9_cmp_pMux_22,gen_9_cmp_pMux_21,gen_9_cmp_pMux_20,
                 gen_9_cmp_pMux_19,gen_9_cmp_pMux_18,gen_9_cmp_pMux_17,
                 gen_9_cmp_pMux_16,gen_9_cmp_pMux_15,gen_9_cmp_pMux_14,
                 gen_9_cmp_pMux_13,gen_9_cmp_pMux_12,gen_9_cmp_pMux_11,
                 gen_9_cmp_pMux_10,gen_9_cmp_pMux_9,gen_9_cmp_pMux_8,
                 gen_9_cmp_pMux_7,gen_9_cmp_pMux_6,gen_9_cmp_pMux_5,
                 gen_9_cmp_pMux_4,gen_9_cmp_pMux_3,gen_9_cmp_pMux_2,
                 gen_9_cmp_pMux_1,gen_9_cmp_pMux_0})) ;
    NBitAdder_24 gen_9_cmp_BSCmp_AdderCmp (.a ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_9_cmp_pMux_30,gen_9_cmp_pMux_29,
                 gen_9_cmp_pMux_28,gen_9_cmp_pMux_27,gen_9_cmp_pMux_26,
                 gen_9_cmp_pMux_25,gen_9_cmp_pMux_24,gen_9_cmp_pMux_23,
                 gen_9_cmp_pMux_22,gen_9_cmp_pMux_21,gen_9_cmp_pMux_20,
                 gen_9_cmp_pMux_19,gen_9_cmp_pMux_18,gen_9_cmp_pMux_17,
                 gen_9_cmp_pMux_16,gen_9_cmp_pMux_15,gen_9_cmp_pMux_14,
                 gen_9_cmp_pMux_13,gen_9_cmp_pMux_12,gen_9_cmp_pMux_11,
                 gen_9_cmp_pMux_10,gen_9_cmp_pMux_9}), .b ({nx10614,nx10614,
                 nx10612,nx10620,nx10618,nx10616,nx10614,nx10612,
                 gen_9_cmp_BSCmp_op2_15,gen_9_cmp_BSCmp_op2_14,
                 gen_9_cmp_BSCmp_op2_13,gen_9_cmp_BSCmp_op2_12,
                 gen_9_cmp_BSCmp_op2_11,gen_9_cmp_BSCmp_op2_10,
                 gen_9_cmp_BSCmp_op2_9,gen_9_cmp_BSCmp_op2_8,
                 gen_9_cmp_BSCmp_op2_7,gen_9_cmp_BSCmp_op2_6,
                 gen_9_cmp_BSCmp_op2_5,gen_9_cmp_BSCmp_op2_4,
                 gen_9_cmp_BSCmp_op2_3,gen_9_cmp_BSCmp_op2_2,
                 gen_9_cmp_BSCmp_op2_1,gen_9_cmp_BSCmp_op2_0}), .carryIn (
                 gen_9_cmp_BSCmp_carryIn), .sum ({gen_9_cmp_pBs_30,
                 gen_9_cmp_pBs_29,gen_9_cmp_pBs_28,gen_9_cmp_pBs_27,
                 gen_9_cmp_pBs_26,gen_9_cmp_pBs_25,gen_9_cmp_pBs_24,
                 gen_9_cmp_pBs_23,outputs_9__15,outputs_9__14,outputs_9__13,
                 outputs_9__12,outputs_9__11,outputs_9__10,outputs_9__9,
                 outputs_9__8,outputs_9__7,outputs_9__6,outputs_9__5,
                 outputs_9__4,outputs_9__3,outputs_9__2,outputs_9__1,
                 outputs_9__0}), .carryOut (\$dummy [79])) ;
    Reg_33 gen_8_cmp_pRegCmp (.D ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
           gen_8_cmp_pBs_30,gen_8_cmp_pBs_29,gen_8_cmp_pBs_28,gen_8_cmp_pBs_27,
           gen_8_cmp_pBs_26,gen_8_cmp_pBs_25,gen_8_cmp_pBs_24,gen_8_cmp_pBs_23,
           outputs_8__15,outputs_8__14,outputs_8__13,outputs_8__12,outputs_8__11
           ,outputs_8__10,outputs_8__9,outputs_8__8,outputs_8__7,outputs_8__6,
           outputs_8__5,outputs_8__4,outputs_8__3,outputs_8__2,outputs_8__1,
           outputs_8__0,gen_8_cmp_pMux_8,gen_8_cmp_pMux_7,gen_8_cmp_pMux_6,
           gen_8_cmp_pMux_5,gen_8_cmp_pMux_4,gen_8_cmp_pMux_3,nx10322}), .en (
           nx11924), .clk (nx10126), .rst (rst), .Q ({\$dummy [80],\$dummy [81],
           gen_8_cmp_pReg_30,gen_8_cmp_pReg_29,gen_8_cmp_pReg_28,
           gen_8_cmp_pReg_27,gen_8_cmp_pReg_26,gen_8_cmp_pReg_25,
           gen_8_cmp_pReg_24,gen_8_cmp_pReg_23,gen_8_cmp_pReg_22,
           gen_8_cmp_pReg_21,gen_8_cmp_pReg_20,gen_8_cmp_pReg_19,
           gen_8_cmp_pReg_18,gen_8_cmp_pReg_17,gen_8_cmp_pReg_16,
           gen_8_cmp_pReg_15,gen_8_cmp_pReg_14,gen_8_cmp_pReg_13,
           gen_8_cmp_pReg_12,gen_8_cmp_pReg_11,gen_8_cmp_pReg_10,
           gen_8_cmp_pReg_9,gen_8_cmp_pReg_8,gen_8_cmp_pReg_7,gen_8_cmp_pReg_6,
           gen_8_cmp_pReg_5,gen_8_cmp_pReg_4,gen_8_cmp_pReg_3,gen_8_cmp_pReg_2,
           gen_8_cmp_pReg_1,gen_8_cmp_pReg_0})) ;
    BinaryMux_33 gen_8_cmp_MuxCmp (.a ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_8_cmp_pReg_30,gen_8_cmp_pReg_29,gen_8_cmp_pReg_28,
                 gen_8_cmp_pReg_27,gen_8_cmp_pReg_26,gen_8_cmp_pReg_25,
                 gen_8_cmp_pReg_24,gen_8_cmp_pReg_23,gen_8_cmp_pReg_22,
                 gen_8_cmp_pReg_21,gen_8_cmp_pReg_20,gen_8_cmp_pReg_19,
                 gen_8_cmp_pReg_18,gen_8_cmp_pReg_17,gen_8_cmp_pReg_16,
                 gen_8_cmp_pReg_15,gen_8_cmp_pReg_14,gen_8_cmp_pReg_13,
                 gen_8_cmp_pReg_12,gen_8_cmp_pReg_11,gen_8_cmp_pReg_10,
                 gen_8_cmp_pReg_9,gen_8_cmp_pReg_8,gen_8_cmp_pReg_7,
                 gen_8_cmp_pReg_6,gen_8_cmp_pReg_5,gen_8_cmp_pReg_4,
                 gen_8_cmp_pReg_3,gen_8_cmp_pReg_2,gen_8_cmp_pReg_1,
                 gen_8_cmp_pReg_0}), .b ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,filter_8__7,filter_8__6
                 ,filter_8__5,filter_8__4,filter_8__3,filter_8__2,filter_8__1,
                 filter_8__0,gen_24_cmp_pInit_32}), .sel (nx11908), .f ({
                 \$dummy [82],\$dummy [83],gen_8_cmp_pMux_30,gen_8_cmp_pMux_29,
                 gen_8_cmp_pMux_28,gen_8_cmp_pMux_27,gen_8_cmp_pMux_26,
                 gen_8_cmp_pMux_25,gen_8_cmp_pMux_24,gen_8_cmp_pMux_23,
                 gen_8_cmp_pMux_22,gen_8_cmp_pMux_21,gen_8_cmp_pMux_20,
                 gen_8_cmp_pMux_19,gen_8_cmp_pMux_18,gen_8_cmp_pMux_17,
                 gen_8_cmp_pMux_16,gen_8_cmp_pMux_15,gen_8_cmp_pMux_14,
                 gen_8_cmp_pMux_13,gen_8_cmp_pMux_12,gen_8_cmp_pMux_11,
                 gen_8_cmp_pMux_10,gen_8_cmp_pMux_9,gen_8_cmp_pMux_8,
                 gen_8_cmp_pMux_7,gen_8_cmp_pMux_6,gen_8_cmp_pMux_5,
                 gen_8_cmp_pMux_4,gen_8_cmp_pMux_3,gen_8_cmp_pMux_2,
                 gen_8_cmp_pMux_1,gen_8_cmp_pMux_0})) ;
    NBitAdder_24 gen_8_cmp_BSCmp_AdderCmp (.a ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_8_cmp_pMux_30,gen_8_cmp_pMux_29,
                 gen_8_cmp_pMux_28,gen_8_cmp_pMux_27,gen_8_cmp_pMux_26,
                 gen_8_cmp_pMux_25,gen_8_cmp_pMux_24,gen_8_cmp_pMux_23,
                 gen_8_cmp_pMux_22,gen_8_cmp_pMux_21,gen_8_cmp_pMux_20,
                 gen_8_cmp_pMux_19,gen_8_cmp_pMux_18,gen_8_cmp_pMux_17,
                 gen_8_cmp_pMux_16,gen_8_cmp_pMux_15,gen_8_cmp_pMux_14,
                 gen_8_cmp_pMux_13,gen_8_cmp_pMux_12,gen_8_cmp_pMux_11,
                 gen_8_cmp_pMux_10,gen_8_cmp_pMux_9}), .b ({nx10626,nx10626,
                 nx10624,nx10632,nx10630,nx10628,nx10626,nx10624,
                 gen_8_cmp_BSCmp_op2_15,gen_8_cmp_BSCmp_op2_14,
                 gen_8_cmp_BSCmp_op2_13,gen_8_cmp_BSCmp_op2_12,
                 gen_8_cmp_BSCmp_op2_11,gen_8_cmp_BSCmp_op2_10,
                 gen_8_cmp_BSCmp_op2_9,gen_8_cmp_BSCmp_op2_8,
                 gen_8_cmp_BSCmp_op2_7,gen_8_cmp_BSCmp_op2_6,
                 gen_8_cmp_BSCmp_op2_5,gen_8_cmp_BSCmp_op2_4,
                 gen_8_cmp_BSCmp_op2_3,gen_8_cmp_BSCmp_op2_2,
                 gen_8_cmp_BSCmp_op2_1,gen_8_cmp_BSCmp_op2_0}), .carryIn (
                 gen_8_cmp_BSCmp_carryIn), .sum ({gen_8_cmp_pBs_30,
                 gen_8_cmp_pBs_29,gen_8_cmp_pBs_28,gen_8_cmp_pBs_27,
                 gen_8_cmp_pBs_26,gen_8_cmp_pBs_25,gen_8_cmp_pBs_24,
                 gen_8_cmp_pBs_23,outputs_8__15,outputs_8__14,outputs_8__13,
                 outputs_8__12,outputs_8__11,outputs_8__10,outputs_8__9,
                 outputs_8__8,outputs_8__7,outputs_8__6,outputs_8__5,
                 outputs_8__4,outputs_8__3,outputs_8__2,outputs_8__1,
                 outputs_8__0}), .carryOut (\$dummy [84])) ;
    Reg_33 gen_7_cmp_pRegCmp (.D ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
           gen_7_cmp_pBs_30,gen_7_cmp_pBs_29,gen_7_cmp_pBs_28,gen_7_cmp_pBs_27,
           gen_7_cmp_pBs_26,gen_7_cmp_pBs_25,gen_7_cmp_pBs_24,gen_7_cmp_pBs_23,
           outputs_7__15,outputs_7__14,outputs_7__13,outputs_7__12,outputs_7__11
           ,outputs_7__10,outputs_7__9,outputs_7__8,outputs_7__7,outputs_7__6,
           outputs_7__5,outputs_7__4,outputs_7__3,outputs_7__2,outputs_7__1,
           outputs_7__0,gen_7_cmp_pMux_8,gen_7_cmp_pMux_7,gen_7_cmp_pMux_6,
           gen_7_cmp_pMux_5,gen_7_cmp_pMux_4,gen_7_cmp_pMux_3,nx10334}), .en (
           nx11926), .clk (nx10126), .rst (rst), .Q ({\$dummy [85],\$dummy [86],
           gen_7_cmp_pReg_30,gen_7_cmp_pReg_29,gen_7_cmp_pReg_28,
           gen_7_cmp_pReg_27,gen_7_cmp_pReg_26,gen_7_cmp_pReg_25,
           gen_7_cmp_pReg_24,gen_7_cmp_pReg_23,gen_7_cmp_pReg_22,
           gen_7_cmp_pReg_21,gen_7_cmp_pReg_20,gen_7_cmp_pReg_19,
           gen_7_cmp_pReg_18,gen_7_cmp_pReg_17,gen_7_cmp_pReg_16,
           gen_7_cmp_pReg_15,gen_7_cmp_pReg_14,gen_7_cmp_pReg_13,
           gen_7_cmp_pReg_12,gen_7_cmp_pReg_11,gen_7_cmp_pReg_10,
           gen_7_cmp_pReg_9,gen_7_cmp_pReg_8,gen_7_cmp_pReg_7,gen_7_cmp_pReg_6,
           gen_7_cmp_pReg_5,gen_7_cmp_pReg_4,gen_7_cmp_pReg_3,gen_7_cmp_pReg_2,
           gen_7_cmp_pReg_1,gen_7_cmp_pReg_0})) ;
    BinaryMux_33 gen_7_cmp_MuxCmp (.a ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_7_cmp_pReg_30,gen_7_cmp_pReg_29,gen_7_cmp_pReg_28,
                 gen_7_cmp_pReg_27,gen_7_cmp_pReg_26,gen_7_cmp_pReg_25,
                 gen_7_cmp_pReg_24,gen_7_cmp_pReg_23,gen_7_cmp_pReg_22,
                 gen_7_cmp_pReg_21,gen_7_cmp_pReg_20,gen_7_cmp_pReg_19,
                 gen_7_cmp_pReg_18,gen_7_cmp_pReg_17,gen_7_cmp_pReg_16,
                 gen_7_cmp_pReg_15,gen_7_cmp_pReg_14,gen_7_cmp_pReg_13,
                 gen_7_cmp_pReg_12,gen_7_cmp_pReg_11,gen_7_cmp_pReg_10,
                 gen_7_cmp_pReg_9,gen_7_cmp_pReg_8,gen_7_cmp_pReg_7,
                 gen_7_cmp_pReg_6,gen_7_cmp_pReg_5,gen_7_cmp_pReg_4,
                 gen_7_cmp_pReg_3,gen_7_cmp_pReg_2,gen_7_cmp_pReg_1,
                 gen_7_cmp_pReg_0}), .b ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,filter_7__7,filter_7__6
                 ,filter_7__5,filter_7__4,filter_7__3,filter_7__2,filter_7__1,
                 filter_7__0,gen_24_cmp_pInit_32}), .sel (nx11910), .f ({
                 \$dummy [87],\$dummy [88],gen_7_cmp_pMux_30,gen_7_cmp_pMux_29,
                 gen_7_cmp_pMux_28,gen_7_cmp_pMux_27,gen_7_cmp_pMux_26,
                 gen_7_cmp_pMux_25,gen_7_cmp_pMux_24,gen_7_cmp_pMux_23,
                 gen_7_cmp_pMux_22,gen_7_cmp_pMux_21,gen_7_cmp_pMux_20,
                 gen_7_cmp_pMux_19,gen_7_cmp_pMux_18,gen_7_cmp_pMux_17,
                 gen_7_cmp_pMux_16,gen_7_cmp_pMux_15,gen_7_cmp_pMux_14,
                 gen_7_cmp_pMux_13,gen_7_cmp_pMux_12,gen_7_cmp_pMux_11,
                 gen_7_cmp_pMux_10,gen_7_cmp_pMux_9,gen_7_cmp_pMux_8,
                 gen_7_cmp_pMux_7,gen_7_cmp_pMux_6,gen_7_cmp_pMux_5,
                 gen_7_cmp_pMux_4,gen_7_cmp_pMux_3,gen_7_cmp_pMux_2,
                 gen_7_cmp_pMux_1,gen_7_cmp_pMux_0})) ;
    NBitAdder_24 gen_7_cmp_BSCmp_AdderCmp (.a ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_7_cmp_pMux_30,gen_7_cmp_pMux_29,
                 gen_7_cmp_pMux_28,gen_7_cmp_pMux_27,gen_7_cmp_pMux_26,
                 gen_7_cmp_pMux_25,gen_7_cmp_pMux_24,gen_7_cmp_pMux_23,
                 gen_7_cmp_pMux_22,gen_7_cmp_pMux_21,gen_7_cmp_pMux_20,
                 gen_7_cmp_pMux_19,gen_7_cmp_pMux_18,gen_7_cmp_pMux_17,
                 gen_7_cmp_pMux_16,gen_7_cmp_pMux_15,gen_7_cmp_pMux_14,
                 gen_7_cmp_pMux_13,gen_7_cmp_pMux_12,gen_7_cmp_pMux_11,
                 gen_7_cmp_pMux_10,gen_7_cmp_pMux_9}), .b ({nx10638,nx10638,
                 nx10636,nx10644,nx10642,nx10640,nx10638,nx10636,
                 gen_7_cmp_BSCmp_op2_15,gen_7_cmp_BSCmp_op2_14,
                 gen_7_cmp_BSCmp_op2_13,gen_7_cmp_BSCmp_op2_12,
                 gen_7_cmp_BSCmp_op2_11,gen_7_cmp_BSCmp_op2_10,
                 gen_7_cmp_BSCmp_op2_9,gen_7_cmp_BSCmp_op2_8,
                 gen_7_cmp_BSCmp_op2_7,gen_7_cmp_BSCmp_op2_6,
                 gen_7_cmp_BSCmp_op2_5,gen_7_cmp_BSCmp_op2_4,
                 gen_7_cmp_BSCmp_op2_3,gen_7_cmp_BSCmp_op2_2,
                 gen_7_cmp_BSCmp_op2_1,gen_7_cmp_BSCmp_op2_0}), .carryIn (
                 gen_7_cmp_BSCmp_carryIn), .sum ({gen_7_cmp_pBs_30,
                 gen_7_cmp_pBs_29,gen_7_cmp_pBs_28,gen_7_cmp_pBs_27,
                 gen_7_cmp_pBs_26,gen_7_cmp_pBs_25,gen_7_cmp_pBs_24,
                 gen_7_cmp_pBs_23,outputs_7__15,outputs_7__14,outputs_7__13,
                 outputs_7__12,outputs_7__11,outputs_7__10,outputs_7__9,
                 outputs_7__8,outputs_7__7,outputs_7__6,outputs_7__5,
                 outputs_7__4,outputs_7__3,outputs_7__2,outputs_7__1,
                 outputs_7__0}), .carryOut (\$dummy [89])) ;
    Reg_33 gen_6_cmp_pRegCmp (.D ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
           gen_6_cmp_pBs_30,gen_6_cmp_pBs_29,gen_6_cmp_pBs_28,gen_6_cmp_pBs_27,
           gen_6_cmp_pBs_26,gen_6_cmp_pBs_25,gen_6_cmp_pBs_24,gen_6_cmp_pBs_23,
           outputs_6__15,outputs_6__14,outputs_6__13,outputs_6__12,outputs_6__11
           ,outputs_6__10,outputs_6__9,outputs_6__8,outputs_6__7,outputs_6__6,
           outputs_6__5,outputs_6__4,outputs_6__3,outputs_6__2,outputs_6__1,
           outputs_6__0,gen_6_cmp_pMux_8,gen_6_cmp_pMux_7,gen_6_cmp_pMux_6,
           gen_6_cmp_pMux_5,gen_6_cmp_pMux_4,gen_6_cmp_pMux_3,nx10346}), .en (
           nx11926), .clk (nx10126), .rst (rst), .Q ({\$dummy [90],\$dummy [91],
           gen_6_cmp_pReg_30,gen_6_cmp_pReg_29,gen_6_cmp_pReg_28,
           gen_6_cmp_pReg_27,gen_6_cmp_pReg_26,gen_6_cmp_pReg_25,
           gen_6_cmp_pReg_24,gen_6_cmp_pReg_23,gen_6_cmp_pReg_22,
           gen_6_cmp_pReg_21,gen_6_cmp_pReg_20,gen_6_cmp_pReg_19,
           gen_6_cmp_pReg_18,gen_6_cmp_pReg_17,gen_6_cmp_pReg_16,
           gen_6_cmp_pReg_15,gen_6_cmp_pReg_14,gen_6_cmp_pReg_13,
           gen_6_cmp_pReg_12,gen_6_cmp_pReg_11,gen_6_cmp_pReg_10,
           gen_6_cmp_pReg_9,gen_6_cmp_pReg_8,gen_6_cmp_pReg_7,gen_6_cmp_pReg_6,
           gen_6_cmp_pReg_5,gen_6_cmp_pReg_4,gen_6_cmp_pReg_3,gen_6_cmp_pReg_2,
           gen_6_cmp_pReg_1,gen_6_cmp_pReg_0})) ;
    BinaryMux_33 gen_6_cmp_MuxCmp (.a ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_6_cmp_pReg_30,gen_6_cmp_pReg_29,gen_6_cmp_pReg_28,
                 gen_6_cmp_pReg_27,gen_6_cmp_pReg_26,gen_6_cmp_pReg_25,
                 gen_6_cmp_pReg_24,gen_6_cmp_pReg_23,gen_6_cmp_pReg_22,
                 gen_6_cmp_pReg_21,gen_6_cmp_pReg_20,gen_6_cmp_pReg_19,
                 gen_6_cmp_pReg_18,gen_6_cmp_pReg_17,gen_6_cmp_pReg_16,
                 gen_6_cmp_pReg_15,gen_6_cmp_pReg_14,gen_6_cmp_pReg_13,
                 gen_6_cmp_pReg_12,gen_6_cmp_pReg_11,gen_6_cmp_pReg_10,
                 gen_6_cmp_pReg_9,gen_6_cmp_pReg_8,gen_6_cmp_pReg_7,
                 gen_6_cmp_pReg_6,gen_6_cmp_pReg_5,gen_6_cmp_pReg_4,
                 gen_6_cmp_pReg_3,gen_6_cmp_pReg_2,gen_6_cmp_pReg_1,
                 gen_6_cmp_pReg_0}), .b ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,filter_6__7,filter_6__6
                 ,filter_6__5,filter_6__4,filter_6__3,filter_6__2,filter_6__1,
                 filter_6__0,gen_24_cmp_pInit_32}), .sel (nx11910), .f ({
                 \$dummy [92],\$dummy [93],gen_6_cmp_pMux_30,gen_6_cmp_pMux_29,
                 gen_6_cmp_pMux_28,gen_6_cmp_pMux_27,gen_6_cmp_pMux_26,
                 gen_6_cmp_pMux_25,gen_6_cmp_pMux_24,gen_6_cmp_pMux_23,
                 gen_6_cmp_pMux_22,gen_6_cmp_pMux_21,gen_6_cmp_pMux_20,
                 gen_6_cmp_pMux_19,gen_6_cmp_pMux_18,gen_6_cmp_pMux_17,
                 gen_6_cmp_pMux_16,gen_6_cmp_pMux_15,gen_6_cmp_pMux_14,
                 gen_6_cmp_pMux_13,gen_6_cmp_pMux_12,gen_6_cmp_pMux_11,
                 gen_6_cmp_pMux_10,gen_6_cmp_pMux_9,gen_6_cmp_pMux_8,
                 gen_6_cmp_pMux_7,gen_6_cmp_pMux_6,gen_6_cmp_pMux_5,
                 gen_6_cmp_pMux_4,gen_6_cmp_pMux_3,gen_6_cmp_pMux_2,
                 gen_6_cmp_pMux_1,gen_6_cmp_pMux_0})) ;
    NBitAdder_24 gen_6_cmp_BSCmp_AdderCmp (.a ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_6_cmp_pMux_30,gen_6_cmp_pMux_29,
                 gen_6_cmp_pMux_28,gen_6_cmp_pMux_27,gen_6_cmp_pMux_26,
                 gen_6_cmp_pMux_25,gen_6_cmp_pMux_24,gen_6_cmp_pMux_23,
                 gen_6_cmp_pMux_22,gen_6_cmp_pMux_21,gen_6_cmp_pMux_20,
                 gen_6_cmp_pMux_19,gen_6_cmp_pMux_18,gen_6_cmp_pMux_17,
                 gen_6_cmp_pMux_16,gen_6_cmp_pMux_15,gen_6_cmp_pMux_14,
                 gen_6_cmp_pMux_13,gen_6_cmp_pMux_12,gen_6_cmp_pMux_11,
                 gen_6_cmp_pMux_10,gen_6_cmp_pMux_9}), .b ({nx10650,nx10650,
                 nx10648,nx10656,nx10654,nx10652,nx10650,nx10648,
                 gen_6_cmp_BSCmp_op2_15,gen_6_cmp_BSCmp_op2_14,
                 gen_6_cmp_BSCmp_op2_13,gen_6_cmp_BSCmp_op2_12,
                 gen_6_cmp_BSCmp_op2_11,gen_6_cmp_BSCmp_op2_10,
                 gen_6_cmp_BSCmp_op2_9,gen_6_cmp_BSCmp_op2_8,
                 gen_6_cmp_BSCmp_op2_7,gen_6_cmp_BSCmp_op2_6,
                 gen_6_cmp_BSCmp_op2_5,gen_6_cmp_BSCmp_op2_4,
                 gen_6_cmp_BSCmp_op2_3,gen_6_cmp_BSCmp_op2_2,
                 gen_6_cmp_BSCmp_op2_1,gen_6_cmp_BSCmp_op2_0}), .carryIn (
                 gen_6_cmp_BSCmp_carryIn), .sum ({gen_6_cmp_pBs_30,
                 gen_6_cmp_pBs_29,gen_6_cmp_pBs_28,gen_6_cmp_pBs_27,
                 gen_6_cmp_pBs_26,gen_6_cmp_pBs_25,gen_6_cmp_pBs_24,
                 gen_6_cmp_pBs_23,outputs_6__15,outputs_6__14,outputs_6__13,
                 outputs_6__12,outputs_6__11,outputs_6__10,outputs_6__9,
                 outputs_6__8,outputs_6__7,outputs_6__6,outputs_6__5,
                 outputs_6__4,outputs_6__3,outputs_6__2,outputs_6__1,
                 outputs_6__0}), .carryOut (\$dummy [94])) ;
    Reg_33 gen_5_cmp_pRegCmp (.D ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
           gen_5_cmp_pBs_30,gen_5_cmp_pBs_29,gen_5_cmp_pBs_28,gen_5_cmp_pBs_27,
           gen_5_cmp_pBs_26,gen_5_cmp_pBs_25,gen_5_cmp_pBs_24,gen_5_cmp_pBs_23,
           outputs_5__15,outputs_5__14,outputs_5__13,outputs_5__12,outputs_5__11
           ,outputs_5__10,outputs_5__9,outputs_5__8,outputs_5__7,outputs_5__6,
           outputs_5__5,outputs_5__4,outputs_5__3,outputs_5__2,outputs_5__1,
           outputs_5__0,gen_5_cmp_pMux_8,gen_5_cmp_pMux_7,gen_5_cmp_pMux_6,
           gen_5_cmp_pMux_5,gen_5_cmp_pMux_4,gen_5_cmp_pMux_3,nx10358}), .en (
           nx11926), .clk (nx10126), .rst (rst), .Q ({\$dummy [95],\$dummy [96],
           gen_5_cmp_pReg_30,gen_5_cmp_pReg_29,gen_5_cmp_pReg_28,
           gen_5_cmp_pReg_27,gen_5_cmp_pReg_26,gen_5_cmp_pReg_25,
           gen_5_cmp_pReg_24,gen_5_cmp_pReg_23,gen_5_cmp_pReg_22,
           gen_5_cmp_pReg_21,gen_5_cmp_pReg_20,gen_5_cmp_pReg_19,
           gen_5_cmp_pReg_18,gen_5_cmp_pReg_17,gen_5_cmp_pReg_16,
           gen_5_cmp_pReg_15,gen_5_cmp_pReg_14,gen_5_cmp_pReg_13,
           gen_5_cmp_pReg_12,gen_5_cmp_pReg_11,gen_5_cmp_pReg_10,
           gen_5_cmp_pReg_9,gen_5_cmp_pReg_8,gen_5_cmp_pReg_7,gen_5_cmp_pReg_6,
           gen_5_cmp_pReg_5,gen_5_cmp_pReg_4,gen_5_cmp_pReg_3,gen_5_cmp_pReg_2,
           gen_5_cmp_pReg_1,gen_5_cmp_pReg_0})) ;
    BinaryMux_33 gen_5_cmp_MuxCmp (.a ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_5_cmp_pReg_30,gen_5_cmp_pReg_29,gen_5_cmp_pReg_28,
                 gen_5_cmp_pReg_27,gen_5_cmp_pReg_26,gen_5_cmp_pReg_25,
                 gen_5_cmp_pReg_24,gen_5_cmp_pReg_23,gen_5_cmp_pReg_22,
                 gen_5_cmp_pReg_21,gen_5_cmp_pReg_20,gen_5_cmp_pReg_19,
                 gen_5_cmp_pReg_18,gen_5_cmp_pReg_17,gen_5_cmp_pReg_16,
                 gen_5_cmp_pReg_15,gen_5_cmp_pReg_14,gen_5_cmp_pReg_13,
                 gen_5_cmp_pReg_12,gen_5_cmp_pReg_11,gen_5_cmp_pReg_10,
                 gen_5_cmp_pReg_9,gen_5_cmp_pReg_8,gen_5_cmp_pReg_7,
                 gen_5_cmp_pReg_6,gen_5_cmp_pReg_5,gen_5_cmp_pReg_4,
                 gen_5_cmp_pReg_3,gen_5_cmp_pReg_2,gen_5_cmp_pReg_1,
                 gen_5_cmp_pReg_0}), .b ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,filter_5__7,filter_5__6
                 ,filter_5__5,filter_5__4,filter_5__3,filter_5__2,filter_5__1,
                 filter_5__0,gen_24_cmp_pInit_32}), .sel (nx11910), .f ({
                 \$dummy [97],\$dummy [98],gen_5_cmp_pMux_30,gen_5_cmp_pMux_29,
                 gen_5_cmp_pMux_28,gen_5_cmp_pMux_27,gen_5_cmp_pMux_26,
                 gen_5_cmp_pMux_25,gen_5_cmp_pMux_24,gen_5_cmp_pMux_23,
                 gen_5_cmp_pMux_22,gen_5_cmp_pMux_21,gen_5_cmp_pMux_20,
                 gen_5_cmp_pMux_19,gen_5_cmp_pMux_18,gen_5_cmp_pMux_17,
                 gen_5_cmp_pMux_16,gen_5_cmp_pMux_15,gen_5_cmp_pMux_14,
                 gen_5_cmp_pMux_13,gen_5_cmp_pMux_12,gen_5_cmp_pMux_11,
                 gen_5_cmp_pMux_10,gen_5_cmp_pMux_9,gen_5_cmp_pMux_8,
                 gen_5_cmp_pMux_7,gen_5_cmp_pMux_6,gen_5_cmp_pMux_5,
                 gen_5_cmp_pMux_4,gen_5_cmp_pMux_3,gen_5_cmp_pMux_2,
                 gen_5_cmp_pMux_1,gen_5_cmp_pMux_0})) ;
    NBitAdder_24 gen_5_cmp_BSCmp_AdderCmp (.a ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_5_cmp_pMux_30,gen_5_cmp_pMux_29,
                 gen_5_cmp_pMux_28,gen_5_cmp_pMux_27,gen_5_cmp_pMux_26,
                 gen_5_cmp_pMux_25,gen_5_cmp_pMux_24,gen_5_cmp_pMux_23,
                 gen_5_cmp_pMux_22,gen_5_cmp_pMux_21,gen_5_cmp_pMux_20,
                 gen_5_cmp_pMux_19,gen_5_cmp_pMux_18,gen_5_cmp_pMux_17,
                 gen_5_cmp_pMux_16,gen_5_cmp_pMux_15,gen_5_cmp_pMux_14,
                 gen_5_cmp_pMux_13,gen_5_cmp_pMux_12,gen_5_cmp_pMux_11,
                 gen_5_cmp_pMux_10,gen_5_cmp_pMux_9}), .b ({nx10662,nx10662,
                 nx10660,nx10668,nx10666,nx10664,nx10662,nx10660,
                 gen_5_cmp_BSCmp_op2_15,gen_5_cmp_BSCmp_op2_14,
                 gen_5_cmp_BSCmp_op2_13,gen_5_cmp_BSCmp_op2_12,
                 gen_5_cmp_BSCmp_op2_11,gen_5_cmp_BSCmp_op2_10,
                 gen_5_cmp_BSCmp_op2_9,gen_5_cmp_BSCmp_op2_8,
                 gen_5_cmp_BSCmp_op2_7,gen_5_cmp_BSCmp_op2_6,
                 gen_5_cmp_BSCmp_op2_5,gen_5_cmp_BSCmp_op2_4,
                 gen_5_cmp_BSCmp_op2_3,gen_5_cmp_BSCmp_op2_2,
                 gen_5_cmp_BSCmp_op2_1,gen_5_cmp_BSCmp_op2_0}), .carryIn (
                 gen_5_cmp_BSCmp_carryIn), .sum ({gen_5_cmp_pBs_30,
                 gen_5_cmp_pBs_29,gen_5_cmp_pBs_28,gen_5_cmp_pBs_27,
                 gen_5_cmp_pBs_26,gen_5_cmp_pBs_25,gen_5_cmp_pBs_24,
                 gen_5_cmp_pBs_23,outputs_5__15,outputs_5__14,outputs_5__13,
                 outputs_5__12,outputs_5__11,outputs_5__10,outputs_5__9,
                 outputs_5__8,outputs_5__7,outputs_5__6,outputs_5__5,
                 outputs_5__4,outputs_5__3,outputs_5__2,outputs_5__1,
                 outputs_5__0}), .carryOut (\$dummy [99])) ;
    Reg_33 gen_4_cmp_pRegCmp (.D ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
           gen_4_cmp_pBs_30,gen_4_cmp_pBs_29,gen_4_cmp_pBs_28,gen_4_cmp_pBs_27,
           gen_4_cmp_pBs_26,gen_4_cmp_pBs_25,gen_4_cmp_pBs_24,gen_4_cmp_pBs_23,
           outputs_4__15,outputs_4__14,outputs_4__13,outputs_4__12,outputs_4__11
           ,outputs_4__10,outputs_4__9,outputs_4__8,outputs_4__7,outputs_4__6,
           outputs_4__5,outputs_4__4,outputs_4__3,outputs_4__2,outputs_4__1,
           outputs_4__0,gen_4_cmp_pMux_8,gen_4_cmp_pMux_7,gen_4_cmp_pMux_6,
           gen_4_cmp_pMux_5,gen_4_cmp_pMux_4,gen_4_cmp_pMux_3,nx10370}), .en (
           nx10884), .clk (nx10126), .rst (rst), .Q ({\$dummy [100],
           \$dummy [101],gen_4_cmp_pReg_30,gen_4_cmp_pReg_29,gen_4_cmp_pReg_28,
           gen_4_cmp_pReg_27,gen_4_cmp_pReg_26,gen_4_cmp_pReg_25,
           gen_4_cmp_pReg_24,gen_4_cmp_pReg_23,gen_4_cmp_pReg_22,
           gen_4_cmp_pReg_21,gen_4_cmp_pReg_20,gen_4_cmp_pReg_19,
           gen_4_cmp_pReg_18,gen_4_cmp_pReg_17,gen_4_cmp_pReg_16,
           gen_4_cmp_pReg_15,gen_4_cmp_pReg_14,gen_4_cmp_pReg_13,
           gen_4_cmp_pReg_12,gen_4_cmp_pReg_11,gen_4_cmp_pReg_10,
           gen_4_cmp_pReg_9,gen_4_cmp_pReg_8,gen_4_cmp_pReg_7,gen_4_cmp_pReg_6,
           gen_4_cmp_pReg_5,gen_4_cmp_pReg_4,gen_4_cmp_pReg_3,gen_4_cmp_pReg_2,
           gen_4_cmp_pReg_1,gen_4_cmp_pReg_0})) ;
    BinaryMux_33 gen_4_cmp_MuxCmp (.a ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_4_cmp_pReg_30,gen_4_cmp_pReg_29,gen_4_cmp_pReg_28,
                 gen_4_cmp_pReg_27,gen_4_cmp_pReg_26,gen_4_cmp_pReg_25,
                 gen_4_cmp_pReg_24,gen_4_cmp_pReg_23,gen_4_cmp_pReg_22,
                 gen_4_cmp_pReg_21,gen_4_cmp_pReg_20,gen_4_cmp_pReg_19,
                 gen_4_cmp_pReg_18,gen_4_cmp_pReg_17,gen_4_cmp_pReg_16,
                 gen_4_cmp_pReg_15,gen_4_cmp_pReg_14,gen_4_cmp_pReg_13,
                 gen_4_cmp_pReg_12,gen_4_cmp_pReg_11,gen_4_cmp_pReg_10,
                 gen_4_cmp_pReg_9,gen_4_cmp_pReg_8,gen_4_cmp_pReg_7,
                 gen_4_cmp_pReg_6,gen_4_cmp_pReg_5,gen_4_cmp_pReg_4,
                 gen_4_cmp_pReg_3,gen_4_cmp_pReg_2,gen_4_cmp_pReg_1,
                 gen_4_cmp_pReg_0}), .b ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,filter_4__7,filter_4__6
                 ,filter_4__5,filter_4__4,filter_4__3,filter_4__2,filter_4__1,
                 filter_4__0,gen_24_cmp_pInit_32}), .sel (nx11912), .f ({
                 \$dummy [102],\$dummy [103],gen_4_cmp_pMux_30,gen_4_cmp_pMux_29
                 ,gen_4_cmp_pMux_28,gen_4_cmp_pMux_27,gen_4_cmp_pMux_26,
                 gen_4_cmp_pMux_25,gen_4_cmp_pMux_24,gen_4_cmp_pMux_23,
                 gen_4_cmp_pMux_22,gen_4_cmp_pMux_21,gen_4_cmp_pMux_20,
                 gen_4_cmp_pMux_19,gen_4_cmp_pMux_18,gen_4_cmp_pMux_17,
                 gen_4_cmp_pMux_16,gen_4_cmp_pMux_15,gen_4_cmp_pMux_14,
                 gen_4_cmp_pMux_13,gen_4_cmp_pMux_12,gen_4_cmp_pMux_11,
                 gen_4_cmp_pMux_10,gen_4_cmp_pMux_9,gen_4_cmp_pMux_8,
                 gen_4_cmp_pMux_7,gen_4_cmp_pMux_6,gen_4_cmp_pMux_5,
                 gen_4_cmp_pMux_4,gen_4_cmp_pMux_3,gen_4_cmp_pMux_2,
                 gen_4_cmp_pMux_1,gen_4_cmp_pMux_0})) ;
    NBitAdder_24 gen_4_cmp_BSCmp_AdderCmp (.a ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_4_cmp_pMux_30,gen_4_cmp_pMux_29,
                 gen_4_cmp_pMux_28,gen_4_cmp_pMux_27,gen_4_cmp_pMux_26,
                 gen_4_cmp_pMux_25,gen_4_cmp_pMux_24,gen_4_cmp_pMux_23,
                 gen_4_cmp_pMux_22,gen_4_cmp_pMux_21,gen_4_cmp_pMux_20,
                 gen_4_cmp_pMux_19,gen_4_cmp_pMux_18,gen_4_cmp_pMux_17,
                 gen_4_cmp_pMux_16,gen_4_cmp_pMux_15,gen_4_cmp_pMux_14,
                 gen_4_cmp_pMux_13,gen_4_cmp_pMux_12,gen_4_cmp_pMux_11,
                 gen_4_cmp_pMux_10,gen_4_cmp_pMux_9}), .b ({nx10674,nx10674,
                 nx10672,nx10680,nx10678,nx10676,nx10674,nx10672,
                 gen_4_cmp_BSCmp_op2_15,gen_4_cmp_BSCmp_op2_14,
                 gen_4_cmp_BSCmp_op2_13,gen_4_cmp_BSCmp_op2_12,
                 gen_4_cmp_BSCmp_op2_11,gen_4_cmp_BSCmp_op2_10,
                 gen_4_cmp_BSCmp_op2_9,gen_4_cmp_BSCmp_op2_8,
                 gen_4_cmp_BSCmp_op2_7,gen_4_cmp_BSCmp_op2_6,
                 gen_4_cmp_BSCmp_op2_5,gen_4_cmp_BSCmp_op2_4,
                 gen_4_cmp_BSCmp_op2_3,gen_4_cmp_BSCmp_op2_2,
                 gen_4_cmp_BSCmp_op2_1,gen_4_cmp_BSCmp_op2_0}), .carryIn (
                 gen_4_cmp_BSCmp_carryIn), .sum ({gen_4_cmp_pBs_30,
                 gen_4_cmp_pBs_29,gen_4_cmp_pBs_28,gen_4_cmp_pBs_27,
                 gen_4_cmp_pBs_26,gen_4_cmp_pBs_25,gen_4_cmp_pBs_24,
                 gen_4_cmp_pBs_23,outputs_4__15,outputs_4__14,outputs_4__13,
                 outputs_4__12,outputs_4__11,outputs_4__10,outputs_4__9,
                 outputs_4__8,outputs_4__7,outputs_4__6,outputs_4__5,
                 outputs_4__4,outputs_4__3,outputs_4__2,outputs_4__1,
                 outputs_4__0}), .carryOut (\$dummy [104])) ;
    Reg_33 gen_3_cmp_pRegCmp (.D ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
           gen_3_cmp_pBs_30,gen_3_cmp_pBs_29,gen_3_cmp_pBs_28,gen_3_cmp_pBs_27,
           gen_3_cmp_pBs_26,gen_3_cmp_pBs_25,gen_3_cmp_pBs_24,gen_3_cmp_pBs_23,
           outputs_3__15,outputs_3__14,outputs_3__13,outputs_3__12,outputs_3__11
           ,outputs_3__10,outputs_3__9,outputs_3__8,outputs_3__7,outputs_3__6,
           outputs_3__5,outputs_3__4,outputs_3__3,outputs_3__2,outputs_3__1,
           outputs_3__0,gen_3_cmp_pMux_8,gen_3_cmp_pMux_7,gen_3_cmp_pMux_6,
           gen_3_cmp_pMux_5,gen_3_cmp_pMux_4,gen_3_cmp_pMux_3,nx10382}), .en (
           nx11928), .clk (nx10128), .rst (rst), .Q ({\$dummy [105],
           \$dummy [106],gen_3_cmp_pReg_30,gen_3_cmp_pReg_29,gen_3_cmp_pReg_28,
           gen_3_cmp_pReg_27,gen_3_cmp_pReg_26,gen_3_cmp_pReg_25,
           gen_3_cmp_pReg_24,gen_3_cmp_pReg_23,gen_3_cmp_pReg_22,
           gen_3_cmp_pReg_21,gen_3_cmp_pReg_20,gen_3_cmp_pReg_19,
           gen_3_cmp_pReg_18,gen_3_cmp_pReg_17,gen_3_cmp_pReg_16,
           gen_3_cmp_pReg_15,gen_3_cmp_pReg_14,gen_3_cmp_pReg_13,
           gen_3_cmp_pReg_12,gen_3_cmp_pReg_11,gen_3_cmp_pReg_10,
           gen_3_cmp_pReg_9,gen_3_cmp_pReg_8,gen_3_cmp_pReg_7,gen_3_cmp_pReg_6,
           gen_3_cmp_pReg_5,gen_3_cmp_pReg_4,gen_3_cmp_pReg_3,gen_3_cmp_pReg_2,
           gen_3_cmp_pReg_1,gen_3_cmp_pReg_0})) ;
    BinaryMux_33 gen_3_cmp_MuxCmp (.a ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_3_cmp_pReg_30,gen_3_cmp_pReg_29,gen_3_cmp_pReg_28,
                 gen_3_cmp_pReg_27,gen_3_cmp_pReg_26,gen_3_cmp_pReg_25,
                 gen_3_cmp_pReg_24,gen_3_cmp_pReg_23,gen_3_cmp_pReg_22,
                 gen_3_cmp_pReg_21,gen_3_cmp_pReg_20,gen_3_cmp_pReg_19,
                 gen_3_cmp_pReg_18,gen_3_cmp_pReg_17,gen_3_cmp_pReg_16,
                 gen_3_cmp_pReg_15,gen_3_cmp_pReg_14,gen_3_cmp_pReg_13,
                 gen_3_cmp_pReg_12,gen_3_cmp_pReg_11,gen_3_cmp_pReg_10,
                 gen_3_cmp_pReg_9,gen_3_cmp_pReg_8,gen_3_cmp_pReg_7,
                 gen_3_cmp_pReg_6,gen_3_cmp_pReg_5,gen_3_cmp_pReg_4,
                 gen_3_cmp_pReg_3,gen_3_cmp_pReg_2,gen_3_cmp_pReg_1,
                 gen_3_cmp_pReg_0}), .b ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,filter_3__7,filter_3__6
                 ,filter_3__5,filter_3__4,filter_3__3,filter_3__2,filter_3__1,
                 filter_3__0,gen_24_cmp_pInit_32}), .sel (nx11914), .f ({
                 \$dummy [107],\$dummy [108],gen_3_cmp_pMux_30,gen_3_cmp_pMux_29
                 ,gen_3_cmp_pMux_28,gen_3_cmp_pMux_27,gen_3_cmp_pMux_26,
                 gen_3_cmp_pMux_25,gen_3_cmp_pMux_24,gen_3_cmp_pMux_23,
                 gen_3_cmp_pMux_22,gen_3_cmp_pMux_21,gen_3_cmp_pMux_20,
                 gen_3_cmp_pMux_19,gen_3_cmp_pMux_18,gen_3_cmp_pMux_17,
                 gen_3_cmp_pMux_16,gen_3_cmp_pMux_15,gen_3_cmp_pMux_14,
                 gen_3_cmp_pMux_13,gen_3_cmp_pMux_12,gen_3_cmp_pMux_11,
                 gen_3_cmp_pMux_10,gen_3_cmp_pMux_9,gen_3_cmp_pMux_8,
                 gen_3_cmp_pMux_7,gen_3_cmp_pMux_6,gen_3_cmp_pMux_5,
                 gen_3_cmp_pMux_4,gen_3_cmp_pMux_3,gen_3_cmp_pMux_2,
                 gen_3_cmp_pMux_1,gen_3_cmp_pMux_0})) ;
    NBitAdder_24 gen_3_cmp_BSCmp_AdderCmp (.a ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_3_cmp_pMux_30,gen_3_cmp_pMux_29,
                 gen_3_cmp_pMux_28,gen_3_cmp_pMux_27,gen_3_cmp_pMux_26,
                 gen_3_cmp_pMux_25,gen_3_cmp_pMux_24,gen_3_cmp_pMux_23,
                 gen_3_cmp_pMux_22,gen_3_cmp_pMux_21,gen_3_cmp_pMux_20,
                 gen_3_cmp_pMux_19,gen_3_cmp_pMux_18,gen_3_cmp_pMux_17,
                 gen_3_cmp_pMux_16,gen_3_cmp_pMux_15,gen_3_cmp_pMux_14,
                 gen_3_cmp_pMux_13,gen_3_cmp_pMux_12,gen_3_cmp_pMux_11,
                 gen_3_cmp_pMux_10,gen_3_cmp_pMux_9}), .b ({nx10686,nx10686,
                 nx10684,nx10692,nx10690,nx10688,nx10686,nx10684,
                 gen_3_cmp_BSCmp_op2_15,gen_3_cmp_BSCmp_op2_14,
                 gen_3_cmp_BSCmp_op2_13,gen_3_cmp_BSCmp_op2_12,
                 gen_3_cmp_BSCmp_op2_11,gen_3_cmp_BSCmp_op2_10,
                 gen_3_cmp_BSCmp_op2_9,gen_3_cmp_BSCmp_op2_8,
                 gen_3_cmp_BSCmp_op2_7,gen_3_cmp_BSCmp_op2_6,
                 gen_3_cmp_BSCmp_op2_5,gen_3_cmp_BSCmp_op2_4,
                 gen_3_cmp_BSCmp_op2_3,gen_3_cmp_BSCmp_op2_2,
                 gen_3_cmp_BSCmp_op2_1,gen_3_cmp_BSCmp_op2_0}), .carryIn (
                 gen_3_cmp_BSCmp_carryIn), .sum ({gen_3_cmp_pBs_30,
                 gen_3_cmp_pBs_29,gen_3_cmp_pBs_28,gen_3_cmp_pBs_27,
                 gen_3_cmp_pBs_26,gen_3_cmp_pBs_25,gen_3_cmp_pBs_24,
                 gen_3_cmp_pBs_23,outputs_3__15,outputs_3__14,outputs_3__13,
                 outputs_3__12,outputs_3__11,outputs_3__10,outputs_3__9,
                 outputs_3__8,outputs_3__7,outputs_3__6,outputs_3__5,
                 outputs_3__4,outputs_3__3,outputs_3__2,outputs_3__1,
                 outputs_3__0}), .carryOut (\$dummy [109])) ;
    Reg_33 gen_2_cmp_pRegCmp (.D ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
           gen_2_cmp_pBs_30,gen_2_cmp_pBs_29,gen_2_cmp_pBs_28,gen_2_cmp_pBs_27,
           gen_2_cmp_pBs_26,gen_2_cmp_pBs_25,gen_2_cmp_pBs_24,gen_2_cmp_pBs_23,
           outputs_2__15,outputs_2__14,outputs_2__13,outputs_2__12,outputs_2__11
           ,outputs_2__10,outputs_2__9,outputs_2__8,outputs_2__7,outputs_2__6,
           outputs_2__5,outputs_2__4,outputs_2__3,outputs_2__2,outputs_2__1,
           outputs_2__0,gen_2_cmp_pMux_8,gen_2_cmp_pMux_7,gen_2_cmp_pMux_6,
           gen_2_cmp_pMux_5,gen_2_cmp_pMux_4,gen_2_cmp_pMux_3,nx10394}), .en (
           nx11928), .clk (nx10128), .rst (rst), .Q ({\$dummy [110],
           \$dummy [111],gen_2_cmp_pReg_30,gen_2_cmp_pReg_29,gen_2_cmp_pReg_28,
           gen_2_cmp_pReg_27,gen_2_cmp_pReg_26,gen_2_cmp_pReg_25,
           gen_2_cmp_pReg_24,gen_2_cmp_pReg_23,gen_2_cmp_pReg_22,
           gen_2_cmp_pReg_21,gen_2_cmp_pReg_20,gen_2_cmp_pReg_19,
           gen_2_cmp_pReg_18,gen_2_cmp_pReg_17,gen_2_cmp_pReg_16,
           gen_2_cmp_pReg_15,gen_2_cmp_pReg_14,gen_2_cmp_pReg_13,
           gen_2_cmp_pReg_12,gen_2_cmp_pReg_11,gen_2_cmp_pReg_10,
           gen_2_cmp_pReg_9,gen_2_cmp_pReg_8,gen_2_cmp_pReg_7,gen_2_cmp_pReg_6,
           gen_2_cmp_pReg_5,gen_2_cmp_pReg_4,gen_2_cmp_pReg_3,gen_2_cmp_pReg_2,
           gen_2_cmp_pReg_1,gen_2_cmp_pReg_0})) ;
    BinaryMux_33 gen_2_cmp_MuxCmp (.a ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_2_cmp_pReg_30,gen_2_cmp_pReg_29,gen_2_cmp_pReg_28,
                 gen_2_cmp_pReg_27,gen_2_cmp_pReg_26,gen_2_cmp_pReg_25,
                 gen_2_cmp_pReg_24,gen_2_cmp_pReg_23,gen_2_cmp_pReg_22,
                 gen_2_cmp_pReg_21,gen_2_cmp_pReg_20,gen_2_cmp_pReg_19,
                 gen_2_cmp_pReg_18,gen_2_cmp_pReg_17,gen_2_cmp_pReg_16,
                 gen_2_cmp_pReg_15,gen_2_cmp_pReg_14,gen_2_cmp_pReg_13,
                 gen_2_cmp_pReg_12,gen_2_cmp_pReg_11,gen_2_cmp_pReg_10,
                 gen_2_cmp_pReg_9,gen_2_cmp_pReg_8,gen_2_cmp_pReg_7,
                 gen_2_cmp_pReg_6,gen_2_cmp_pReg_5,gen_2_cmp_pReg_4,
                 gen_2_cmp_pReg_3,gen_2_cmp_pReg_2,gen_2_cmp_pReg_1,
                 gen_2_cmp_pReg_0}), .b ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,filter_2__7,filter_2__6
                 ,filter_2__5,filter_2__4,filter_2__3,filter_2__2,filter_2__1,
                 filter_2__0,gen_24_cmp_pInit_32}), .sel (nx11914), .f ({
                 \$dummy [112],\$dummy [113],gen_2_cmp_pMux_30,gen_2_cmp_pMux_29
                 ,gen_2_cmp_pMux_28,gen_2_cmp_pMux_27,gen_2_cmp_pMux_26,
                 gen_2_cmp_pMux_25,gen_2_cmp_pMux_24,gen_2_cmp_pMux_23,
                 gen_2_cmp_pMux_22,gen_2_cmp_pMux_21,gen_2_cmp_pMux_20,
                 gen_2_cmp_pMux_19,gen_2_cmp_pMux_18,gen_2_cmp_pMux_17,
                 gen_2_cmp_pMux_16,gen_2_cmp_pMux_15,gen_2_cmp_pMux_14,
                 gen_2_cmp_pMux_13,gen_2_cmp_pMux_12,gen_2_cmp_pMux_11,
                 gen_2_cmp_pMux_10,gen_2_cmp_pMux_9,gen_2_cmp_pMux_8,
                 gen_2_cmp_pMux_7,gen_2_cmp_pMux_6,gen_2_cmp_pMux_5,
                 gen_2_cmp_pMux_4,gen_2_cmp_pMux_3,gen_2_cmp_pMux_2,
                 gen_2_cmp_pMux_1,gen_2_cmp_pMux_0})) ;
    NBitAdder_24 gen_2_cmp_BSCmp_AdderCmp (.a ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_2_cmp_pMux_30,gen_2_cmp_pMux_29,
                 gen_2_cmp_pMux_28,gen_2_cmp_pMux_27,gen_2_cmp_pMux_26,
                 gen_2_cmp_pMux_25,gen_2_cmp_pMux_24,gen_2_cmp_pMux_23,
                 gen_2_cmp_pMux_22,gen_2_cmp_pMux_21,gen_2_cmp_pMux_20,
                 gen_2_cmp_pMux_19,gen_2_cmp_pMux_18,gen_2_cmp_pMux_17,
                 gen_2_cmp_pMux_16,gen_2_cmp_pMux_15,gen_2_cmp_pMux_14,
                 gen_2_cmp_pMux_13,gen_2_cmp_pMux_12,gen_2_cmp_pMux_11,
                 gen_2_cmp_pMux_10,gen_2_cmp_pMux_9}), .b ({nx10698,nx10698,
                 nx10696,nx10704,nx10702,nx10700,nx10698,nx10696,
                 gen_2_cmp_BSCmp_op2_15,gen_2_cmp_BSCmp_op2_14,
                 gen_2_cmp_BSCmp_op2_13,gen_2_cmp_BSCmp_op2_12,
                 gen_2_cmp_BSCmp_op2_11,gen_2_cmp_BSCmp_op2_10,
                 gen_2_cmp_BSCmp_op2_9,gen_2_cmp_BSCmp_op2_8,
                 gen_2_cmp_BSCmp_op2_7,gen_2_cmp_BSCmp_op2_6,
                 gen_2_cmp_BSCmp_op2_5,gen_2_cmp_BSCmp_op2_4,
                 gen_2_cmp_BSCmp_op2_3,gen_2_cmp_BSCmp_op2_2,
                 gen_2_cmp_BSCmp_op2_1,gen_2_cmp_BSCmp_op2_0}), .carryIn (
                 gen_2_cmp_BSCmp_carryIn), .sum ({gen_2_cmp_pBs_30,
                 gen_2_cmp_pBs_29,gen_2_cmp_pBs_28,gen_2_cmp_pBs_27,
                 gen_2_cmp_pBs_26,gen_2_cmp_pBs_25,gen_2_cmp_pBs_24,
                 gen_2_cmp_pBs_23,outputs_2__15,outputs_2__14,outputs_2__13,
                 outputs_2__12,outputs_2__11,outputs_2__10,outputs_2__9,
                 outputs_2__8,outputs_2__7,outputs_2__6,outputs_2__5,
                 outputs_2__4,outputs_2__3,outputs_2__2,outputs_2__1,
                 outputs_2__0}), .carryOut (\$dummy [114])) ;
    Reg_33 gen_1_cmp_pRegCmp (.D ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
           gen_1_cmp_pBs_30,gen_1_cmp_pBs_29,gen_1_cmp_pBs_28,gen_1_cmp_pBs_27,
           gen_1_cmp_pBs_26,gen_1_cmp_pBs_25,gen_1_cmp_pBs_24,gen_1_cmp_pBs_23,
           outputs_1__15,outputs_1__14,outputs_1__13,outputs_1__12,outputs_1__11
           ,outputs_1__10,outputs_1__9,outputs_1__8,outputs_1__7,outputs_1__6,
           outputs_1__5,outputs_1__4,outputs_1__3,outputs_1__2,outputs_1__1,
           outputs_1__0,gen_1_cmp_pMux_8,gen_1_cmp_pMux_7,gen_1_cmp_pMux_6,
           gen_1_cmp_pMux_5,gen_1_cmp_pMux_4,gen_1_cmp_pMux_3,nx10406}), .en (
           nx11928), .clk (nx10128), .rst (rst), .Q ({\$dummy [115],
           \$dummy [116],gen_1_cmp_pReg_30,gen_1_cmp_pReg_29,gen_1_cmp_pReg_28,
           gen_1_cmp_pReg_27,gen_1_cmp_pReg_26,gen_1_cmp_pReg_25,
           gen_1_cmp_pReg_24,gen_1_cmp_pReg_23,gen_1_cmp_pReg_22,
           gen_1_cmp_pReg_21,gen_1_cmp_pReg_20,gen_1_cmp_pReg_19,
           gen_1_cmp_pReg_18,gen_1_cmp_pReg_17,gen_1_cmp_pReg_16,
           gen_1_cmp_pReg_15,gen_1_cmp_pReg_14,gen_1_cmp_pReg_13,
           gen_1_cmp_pReg_12,gen_1_cmp_pReg_11,gen_1_cmp_pReg_10,
           gen_1_cmp_pReg_9,gen_1_cmp_pReg_8,gen_1_cmp_pReg_7,gen_1_cmp_pReg_6,
           gen_1_cmp_pReg_5,gen_1_cmp_pReg_4,gen_1_cmp_pReg_3,gen_1_cmp_pReg_2,
           gen_1_cmp_pReg_1,gen_1_cmp_pReg_0})) ;
    BinaryMux_33 gen_1_cmp_MuxCmp (.a ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_1_cmp_pReg_30,gen_1_cmp_pReg_29,gen_1_cmp_pReg_28,
                 gen_1_cmp_pReg_27,gen_1_cmp_pReg_26,gen_1_cmp_pReg_25,
                 gen_1_cmp_pReg_24,gen_1_cmp_pReg_23,gen_1_cmp_pReg_22,
                 gen_1_cmp_pReg_21,gen_1_cmp_pReg_20,gen_1_cmp_pReg_19,
                 gen_1_cmp_pReg_18,gen_1_cmp_pReg_17,gen_1_cmp_pReg_16,
                 gen_1_cmp_pReg_15,gen_1_cmp_pReg_14,gen_1_cmp_pReg_13,
                 gen_1_cmp_pReg_12,gen_1_cmp_pReg_11,gen_1_cmp_pReg_10,
                 gen_1_cmp_pReg_9,gen_1_cmp_pReg_8,gen_1_cmp_pReg_7,
                 gen_1_cmp_pReg_6,gen_1_cmp_pReg_5,gen_1_cmp_pReg_4,
                 gen_1_cmp_pReg_3,gen_1_cmp_pReg_2,gen_1_cmp_pReg_1,
                 gen_1_cmp_pReg_0}), .b ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,filter_1__7,filter_1__6
                 ,filter_1__5,filter_1__4,filter_1__3,filter_1__2,filter_1__1,
                 filter_1__0,gen_24_cmp_pInit_32}), .sel (nx10120), .f ({
                 \$dummy [117],\$dummy [118],gen_1_cmp_pMux_30,gen_1_cmp_pMux_29
                 ,gen_1_cmp_pMux_28,gen_1_cmp_pMux_27,gen_1_cmp_pMux_26,
                 gen_1_cmp_pMux_25,gen_1_cmp_pMux_24,gen_1_cmp_pMux_23,
                 gen_1_cmp_pMux_22,gen_1_cmp_pMux_21,gen_1_cmp_pMux_20,
                 gen_1_cmp_pMux_19,gen_1_cmp_pMux_18,gen_1_cmp_pMux_17,
                 gen_1_cmp_pMux_16,gen_1_cmp_pMux_15,gen_1_cmp_pMux_14,
                 gen_1_cmp_pMux_13,gen_1_cmp_pMux_12,gen_1_cmp_pMux_11,
                 gen_1_cmp_pMux_10,gen_1_cmp_pMux_9,gen_1_cmp_pMux_8,
                 gen_1_cmp_pMux_7,gen_1_cmp_pMux_6,gen_1_cmp_pMux_5,
                 gen_1_cmp_pMux_4,gen_1_cmp_pMux_3,gen_1_cmp_pMux_2,
                 gen_1_cmp_pMux_1,gen_1_cmp_pMux_0})) ;
    NBitAdder_24 gen_1_cmp_BSCmp_AdderCmp (.a ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_1_cmp_pMux_30,gen_1_cmp_pMux_29,
                 gen_1_cmp_pMux_28,gen_1_cmp_pMux_27,gen_1_cmp_pMux_26,
                 gen_1_cmp_pMux_25,gen_1_cmp_pMux_24,gen_1_cmp_pMux_23,
                 gen_1_cmp_pMux_22,gen_1_cmp_pMux_21,gen_1_cmp_pMux_20,
                 gen_1_cmp_pMux_19,gen_1_cmp_pMux_18,gen_1_cmp_pMux_17,
                 gen_1_cmp_pMux_16,gen_1_cmp_pMux_15,gen_1_cmp_pMux_14,
                 gen_1_cmp_pMux_13,gen_1_cmp_pMux_12,gen_1_cmp_pMux_11,
                 gen_1_cmp_pMux_10,gen_1_cmp_pMux_9}), .b ({nx10710,nx10710,
                 nx10708,nx10716,nx10714,nx10712,nx10710,nx10708,
                 gen_1_cmp_BSCmp_op2_15,gen_1_cmp_BSCmp_op2_14,
                 gen_1_cmp_BSCmp_op2_13,gen_1_cmp_BSCmp_op2_12,
                 gen_1_cmp_BSCmp_op2_11,gen_1_cmp_BSCmp_op2_10,
                 gen_1_cmp_BSCmp_op2_9,gen_1_cmp_BSCmp_op2_8,
                 gen_1_cmp_BSCmp_op2_7,gen_1_cmp_BSCmp_op2_6,
                 gen_1_cmp_BSCmp_op2_5,gen_1_cmp_BSCmp_op2_4,
                 gen_1_cmp_BSCmp_op2_3,gen_1_cmp_BSCmp_op2_2,
                 gen_1_cmp_BSCmp_op2_1,gen_1_cmp_BSCmp_op2_0}), .carryIn (
                 gen_1_cmp_BSCmp_carryIn), .sum ({gen_1_cmp_pBs_30,
                 gen_1_cmp_pBs_29,gen_1_cmp_pBs_28,gen_1_cmp_pBs_27,
                 gen_1_cmp_pBs_26,gen_1_cmp_pBs_25,gen_1_cmp_pBs_24,
                 gen_1_cmp_pBs_23,outputs_1__15,outputs_1__14,outputs_1__13,
                 outputs_1__12,outputs_1__11,outputs_1__10,outputs_1__9,
                 outputs_1__8,outputs_1__7,outputs_1__6,outputs_1__5,
                 outputs_1__4,outputs_1__3,outputs_1__2,outputs_1__1,
                 outputs_1__0}), .carryOut (\$dummy [119])) ;
    Reg_33 gen_0_cmp_pRegCmp (.D ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
           gen_0_cmp_pBs_30,gen_0_cmp_pBs_29,gen_0_cmp_pBs_28,gen_0_cmp_pBs_27,
           gen_0_cmp_pBs_26,gen_0_cmp_pBs_25,gen_0_cmp_pBs_24,gen_0_cmp_pBs_23,
           outputs_0__15,outputs_0__14,outputs_0__13,outputs_0__12,outputs_0__11
           ,outputs_0__10,outputs_0__9,outputs_0__8,outputs_0__7,outputs_0__6,
           outputs_0__5,outputs_0__4,outputs_0__3,outputs_0__2,outputs_0__1,
           outputs_0__0,gen_0_cmp_pMux_8,gen_0_cmp_pMux_7,gen_0_cmp_pMux_6,
           gen_0_cmp_pMux_5,gen_0_cmp_pMux_4,gen_0_cmp_pMux_3,nx10418}), .en (
           nx10886), .clk (nx10128), .rst (rst), .Q ({\$dummy [120],
           \$dummy [121],gen_0_cmp_pReg_30,gen_0_cmp_pReg_29,gen_0_cmp_pReg_28,
           gen_0_cmp_pReg_27,gen_0_cmp_pReg_26,gen_0_cmp_pReg_25,
           gen_0_cmp_pReg_24,gen_0_cmp_pReg_23,gen_0_cmp_pReg_22,
           gen_0_cmp_pReg_21,gen_0_cmp_pReg_20,gen_0_cmp_pReg_19,
           gen_0_cmp_pReg_18,gen_0_cmp_pReg_17,gen_0_cmp_pReg_16,
           gen_0_cmp_pReg_15,gen_0_cmp_pReg_14,gen_0_cmp_pReg_13,
           gen_0_cmp_pReg_12,gen_0_cmp_pReg_11,gen_0_cmp_pReg_10,
           gen_0_cmp_pReg_9,gen_0_cmp_pReg_8,gen_0_cmp_pReg_7,gen_0_cmp_pReg_6,
           gen_0_cmp_pReg_5,gen_0_cmp_pReg_4,gen_0_cmp_pReg_3,gen_0_cmp_pReg_2,
           gen_0_cmp_pReg_1,gen_0_cmp_pReg_0})) ;
    BinaryMux_33 gen_0_cmp_MuxCmp (.a ({gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_0_cmp_pReg_30,gen_0_cmp_pReg_29,gen_0_cmp_pReg_28,
                 gen_0_cmp_pReg_27,gen_0_cmp_pReg_26,gen_0_cmp_pReg_25,
                 gen_0_cmp_pReg_24,gen_0_cmp_pReg_23,gen_0_cmp_pReg_22,
                 gen_0_cmp_pReg_21,gen_0_cmp_pReg_20,gen_0_cmp_pReg_19,
                 gen_0_cmp_pReg_18,gen_0_cmp_pReg_17,gen_0_cmp_pReg_16,
                 gen_0_cmp_pReg_15,gen_0_cmp_pReg_14,gen_0_cmp_pReg_13,
                 gen_0_cmp_pReg_12,gen_0_cmp_pReg_11,gen_0_cmp_pReg_10,
                 gen_0_cmp_pReg_9,gen_0_cmp_pReg_8,gen_0_cmp_pReg_7,
                 gen_0_cmp_pReg_6,gen_0_cmp_pReg_5,gen_0_cmp_pReg_4,
                 gen_0_cmp_pReg_3,gen_0_cmp_pReg_2,gen_0_cmp_pReg_1,
                 gen_0_cmp_pReg_0}), .b ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_24_cmp_pInit_32,filter_0__7,filter_0__6
                 ,filter_0__5,filter_0__4,filter_0__3,filter_0__2,filter_0__1,
                 filter_0__0,gen_24_cmp_pInit_32}), .sel (nx10120), .f ({
                 \$dummy [122],\$dummy [123],gen_0_cmp_pMux_30,gen_0_cmp_pMux_29
                 ,gen_0_cmp_pMux_28,gen_0_cmp_pMux_27,gen_0_cmp_pMux_26,
                 gen_0_cmp_pMux_25,gen_0_cmp_pMux_24,gen_0_cmp_pMux_23,
                 gen_0_cmp_pMux_22,gen_0_cmp_pMux_21,gen_0_cmp_pMux_20,
                 gen_0_cmp_pMux_19,gen_0_cmp_pMux_18,gen_0_cmp_pMux_17,
                 gen_0_cmp_pMux_16,gen_0_cmp_pMux_15,gen_0_cmp_pMux_14,
                 gen_0_cmp_pMux_13,gen_0_cmp_pMux_12,gen_0_cmp_pMux_11,
                 gen_0_cmp_pMux_10,gen_0_cmp_pMux_9,gen_0_cmp_pMux_8,
                 gen_0_cmp_pMux_7,gen_0_cmp_pMux_6,gen_0_cmp_pMux_5,
                 gen_0_cmp_pMux_4,gen_0_cmp_pMux_3,gen_0_cmp_pMux_2,
                 gen_0_cmp_pMux_1,gen_0_cmp_pMux_0})) ;
    NBitAdder_24 gen_0_cmp_BSCmp_AdderCmp (.a ({gen_24_cmp_pInit_32,
                 gen_24_cmp_pInit_32,gen_0_cmp_pMux_30,gen_0_cmp_pMux_29,
                 gen_0_cmp_pMux_28,gen_0_cmp_pMux_27,gen_0_cmp_pMux_26,
                 gen_0_cmp_pMux_25,gen_0_cmp_pMux_24,gen_0_cmp_pMux_23,
                 gen_0_cmp_pMux_22,gen_0_cmp_pMux_21,gen_0_cmp_pMux_20,
                 gen_0_cmp_pMux_19,gen_0_cmp_pMux_18,gen_0_cmp_pMux_17,
                 gen_0_cmp_pMux_16,gen_0_cmp_pMux_15,gen_0_cmp_pMux_14,
                 gen_0_cmp_pMux_13,gen_0_cmp_pMux_12,gen_0_cmp_pMux_11,
                 gen_0_cmp_pMux_10,gen_0_cmp_pMux_9}), .b ({nx10722,nx10722,
                 nx10720,nx10728,nx10726,nx10724,nx10722,nx10720,
                 gen_0_cmp_BSCmp_op2_15,gen_0_cmp_BSCmp_op2_14,
                 gen_0_cmp_BSCmp_op2_13,gen_0_cmp_BSCmp_op2_12,
                 gen_0_cmp_BSCmp_op2_11,gen_0_cmp_BSCmp_op2_10,
                 gen_0_cmp_BSCmp_op2_9,gen_0_cmp_BSCmp_op2_8,
                 gen_0_cmp_BSCmp_op2_7,gen_0_cmp_BSCmp_op2_6,
                 gen_0_cmp_BSCmp_op2_5,gen_0_cmp_BSCmp_op2_4,
                 gen_0_cmp_BSCmp_op2_3,gen_0_cmp_BSCmp_op2_2,
                 gen_0_cmp_BSCmp_op2_1,gen_0_cmp_BSCmp_op2_0}), .carryIn (
                 gen_0_cmp_BSCmp_carryIn), .sum ({gen_0_cmp_pBs_30,
                 gen_0_cmp_pBs_29,gen_0_cmp_pBs_28,gen_0_cmp_pBs_27,
                 gen_0_cmp_pBs_26,gen_0_cmp_pBs_25,gen_0_cmp_pBs_24,
                 gen_0_cmp_pBs_23,outputs_0__15,outputs_0__14,outputs_0__13,
                 outputs_0__12,outputs_0__11,outputs_0__10,outputs_0__9,
                 outputs_0__8,outputs_0__7,outputs_0__6,outputs_0__5,
                 outputs_0__4,outputs_0__3,outputs_0__2,outputs_0__1,
                 outputs_0__0}), .carryOut (\$dummy [124])) ;
    nand02 ix3692 (.Y (nx3691), .A0 (nx11928), .A1 (nx3729)) ;
    dffr CounterCmp_reg_outp_3 (.Q (done), .QB (\$dummy [125]), .D (nx3691), .CLK (
         clk), .R (nx9666)) ;
    inv01 ix9667 (.Y (nx9666), .A (nx3713)) ;
    nor02_2x ix3714 (.Y (nx3713), .A0 (restartDetection), .A1 (rst)) ;
    dffr StartCaptuerCmp_reg_f (.Q (restartDetection), .QB (\$dummy [126]), .D (
         nx9650), .CLK (start), .R (nx9660)) ;
    fake_vcc ix9651 (.Y (nx9650)) ;
    inv01 ix9661 (.Y (nx9660), .A (nx3720)) ;
    nor02_2x ix3721 (.Y (nx3720), .A0 (StartCaptuerCmp_d), .A1 (rst)) ;
    dff StartCaptuerCmp_reg_d (.Q (StartCaptuerCmp_d), .QB (\$dummy [127]), .D (
        restartDetection), .CLK (nx10128)) ;
    dffr CounterCmp_reg_outp_2 (.Q (\$dummy [128]), .QB (nx3729), .D (nx3681), .CLK (
         clk), .R (nx9666)) ;
    mux21 ix3682 (.Y (nx3681), .A0 (nx3733), .A1 (nx3729), .S0 (nx11934)) ;
    nand02 ix3672 (.Y (nx3671), .A0 (nx3737), .A1 (nx3741)) ;
    nand02 ix3738 (.Y (nx3737), .A0 (CounterCmp_outp_1), .A1 (nx11934)) ;
    dffr CounterCmp_reg_outp_1 (.Q (CounterCmp_outp_1), .QB (nx3733), .D (nx3671
         ), .CLK (clk), .R (nx9666)) ;
    nand02 ix3742 (.Y (nx3741), .A0 (nx11914), .A1 (nx10886)) ;
    nor02_2x ix3698 (.Y (nx3697), .A0 (nx11938), .A1 (nx10886)) ;
    dffs_ni CounterCmp_reg_outp_0 (.Q (\$dummy [129]), .QB (nx3745), .D (nx3697)
            , .CLK (clk), .S (nx9666)) ;
    fake_gnd ix3184 (.Y (gen_24_cmp_pInit_32)) ;
    nand02 ix67 (.Y (gen_0_cmp_BSCmp_op2_1), .A0 (nx3751), .A1 (nx3771)) ;
    nor02_2x ix3752 (.Y (nx3751), .A0 (nx62), .A1 (nx58)) ;
    nor03_2x ix63 (.Y (nx62), .A0 (gen_0_cmp_mReg_0), .A1 (nx10424), .A2 (
             nx10890)) ;
    dffr gen_0_cmp_mRegCmp_reg_Q_0 (.Q (gen_0_cmp_mReg_0), .QB (nx3757), .D (
         window_0__0), .CLK (start), .R (rst)) ;
    inv01 ix3762 (.Y (nx3761), .A (gen_0_cmp_pMux_0)) ;
    nor03_2x ix59 (.Y (nx58), .A0 (nx3757), .A1 (nx10896), .A2 (nx10906)) ;
    inv02 ix3770 (.Y (nx3769), .A (gen_0_cmp_pMux_2)) ;
    nor02_2x ix3772 (.Y (nx3771), .A0 (nx48), .A1 (nx46)) ;
    nor03_2x ix49 (.Y (nx48), .A0 (nx3775), .A1 (nx10418), .A2 (nx10914)) ;
    dffr gen_0_cmp_mRegCmp_reg_Q_1 (.Q (gen_0_cmp_mReg_1), .QB (nx3775), .D (
         window_0__1), .CLK (start), .R (rst)) ;
    nor03_2x ix47 (.Y (nx46), .A0 (gen_0_cmp_mReg_1), .A1 (nx10730), .A2 (
             nx10922)) ;
    nor03_2x ix7 (.Y (nx6), .A0 (nx10424), .A1 (nx3769), .A2 (gen_0_cmp_pMux_0)
             ) ;
    nand02 ix89 (.Y (gen_0_cmp_BSCmp_op2_2), .A0 (nx3786), .A1 (nx3791)) ;
    nor02_2x ix3787 (.Y (nx3786), .A0 (nx84), .A1 (nx80)) ;
    nor03_2x ix85 (.Y (nx84), .A0 (gen_0_cmp_mReg_1), .A1 (nx10424), .A2 (
             nx10890)) ;
    nor03_2x ix81 (.Y (nx80), .A0 (nx3775), .A1 (nx10896), .A2 (nx10906)) ;
    nor02_2x ix3792 (.Y (nx3791), .A0 (nx76), .A1 (nx74)) ;
    nor03_2x ix77 (.Y (nx76), .A0 (nx3795), .A1 (nx10418), .A2 (nx10914)) ;
    dffr gen_0_cmp_mRegCmp_reg_Q_2 (.Q (gen_0_cmp_mReg_2), .QB (nx3795), .D (
         window_0__2), .CLK (start), .R (rst)) ;
    nor03_2x ix75 (.Y (nx74), .A0 (gen_0_cmp_mReg_2), .A1 (nx10730), .A2 (
             nx10922)) ;
    nand02 ix111 (.Y (gen_0_cmp_BSCmp_op2_3), .A0 (nx3801), .A1 (nx3807)) ;
    nor02_2x ix3802 (.Y (nx3801), .A0 (nx106), .A1 (nx102)) ;
    nor03_2x ix107 (.Y (nx106), .A0 (gen_0_cmp_mReg_2), .A1 (nx10424), .A2 (
             nx10890)) ;
    nor03_2x ix103 (.Y (nx102), .A0 (nx3795), .A1 (nx10896), .A2 (nx10906)) ;
    nor02_2x ix3808 (.Y (nx3807), .A0 (nx98), .A1 (nx96)) ;
    nor03_2x ix99 (.Y (nx98), .A0 (nx3810), .A1 (nx10418), .A2 (nx10914)) ;
    dffr gen_0_cmp_mRegCmp_reg_Q_3 (.Q (gen_0_cmp_mReg_3), .QB (nx3810), .D (
         window_0__3), .CLK (start), .R (rst)) ;
    nor03_2x ix97 (.Y (nx96), .A0 (gen_0_cmp_mReg_3), .A1 (nx10730), .A2 (
             nx10922)) ;
    nand02 ix133 (.Y (gen_0_cmp_BSCmp_op2_4), .A0 (nx3817), .A1 (nx3823)) ;
    nor02_2x ix3818 (.Y (nx3817), .A0 (nx128), .A1 (nx124)) ;
    nor03_2x ix129 (.Y (nx128), .A0 (gen_0_cmp_mReg_3), .A1 (nx10424), .A2 (
             nx10890)) ;
    nor03_2x ix125 (.Y (nx124), .A0 (nx3810), .A1 (nx10896), .A2 (nx10906)) ;
    nor02_2x ix3824 (.Y (nx3823), .A0 (nx120), .A1 (nx118)) ;
    nor03_2x ix121 (.Y (nx120), .A0 (nx3827), .A1 (nx10418), .A2 (nx10914)) ;
    dffr gen_0_cmp_mRegCmp_reg_Q_4 (.Q (gen_0_cmp_mReg_4), .QB (nx3827), .D (
         window_0__4), .CLK (start), .R (rst)) ;
    nor03_2x ix119 (.Y (nx118), .A0 (gen_0_cmp_mReg_4), .A1 (nx10730), .A2 (
             nx10922)) ;
    nand02 ix155 (.Y (gen_0_cmp_BSCmp_op2_5), .A0 (nx3831), .A1 (nx3837)) ;
    nor02_2x ix3832 (.Y (nx3831), .A0 (nx150), .A1 (nx146)) ;
    nor03_2x ix151 (.Y (nx150), .A0 (gen_0_cmp_mReg_4), .A1 (nx10424), .A2 (
             nx10890)) ;
    nor03_2x ix147 (.Y (nx146), .A0 (nx3827), .A1 (nx10896), .A2 (nx10906)) ;
    nor02_2x ix3838 (.Y (nx3837), .A0 (nx142), .A1 (nx140)) ;
    nor03_2x ix143 (.Y (nx142), .A0 (nx3841), .A1 (nx10420), .A2 (nx10914)) ;
    dffr gen_0_cmp_mRegCmp_reg_Q_5 (.Q (gen_0_cmp_mReg_5), .QB (nx3841), .D (
         window_0__5), .CLK (start), .R (rst)) ;
    nor03_2x ix141 (.Y (nx140), .A0 (gen_0_cmp_mReg_5), .A1 (nx10730), .A2 (
             nx10922)) ;
    nand02 ix177 (.Y (gen_0_cmp_BSCmp_op2_6), .A0 (nx3845), .A1 (nx3851)) ;
    nor02_2x ix3846 (.Y (nx3845), .A0 (nx172), .A1 (nx168)) ;
    nor03_2x ix173 (.Y (nx172), .A0 (gen_0_cmp_mReg_5), .A1 (nx10426), .A2 (
             nx10890)) ;
    nor03_2x ix169 (.Y (nx168), .A0 (nx3841), .A1 (nx10896), .A2 (nx10906)) ;
    nor02_2x ix3852 (.Y (nx3851), .A0 (nx164), .A1 (nx162)) ;
    nor03_2x ix165 (.Y (nx164), .A0 (nx3855), .A1 (nx10420), .A2 (nx10914)) ;
    dffr gen_0_cmp_mRegCmp_reg_Q_6 (.Q (gen_0_cmp_mReg_6), .QB (nx3855), .D (
         window_0__6), .CLK (start), .R (rst)) ;
    nor03_2x ix163 (.Y (nx162), .A0 (gen_0_cmp_mReg_6), .A1 (nx10730), .A2 (
             nx10922)) ;
    nand02 ix199 (.Y (gen_0_cmp_BSCmp_op2_7), .A0 (nx3861), .A1 (nx3867)) ;
    nor02_2x ix3862 (.Y (nx3861), .A0 (nx194), .A1 (nx190)) ;
    nor03_2x ix195 (.Y (nx194), .A0 (gen_0_cmp_mReg_6), .A1 (nx10426), .A2 (
             nx10892)) ;
    nor03_2x ix191 (.Y (nx190), .A0 (nx3855), .A1 (nx10898), .A2 (nx10908)) ;
    nor02_2x ix3868 (.Y (nx3867), .A0 (nx186), .A1 (nx184)) ;
    nor03_2x ix187 (.Y (nx186), .A0 (nx3870), .A1 (nx10420), .A2 (nx10916)) ;
    dffr gen_0_cmp_mRegCmp_reg_Q_7 (.Q (gen_0_cmp_mReg_7), .QB (nx3870), .D (
         window_0__7), .CLK (start), .R (rst)) ;
    nor03_2x ix185 (.Y (nx184), .A0 (gen_0_cmp_mReg_7), .A1 (nx10730), .A2 (
             nx10924)) ;
    nand02 ix221 (.Y (gen_0_cmp_BSCmp_op2_8), .A0 (nx3874), .A1 (nx3879)) ;
    nor02_2x ix3875 (.Y (nx3874), .A0 (nx216), .A1 (nx212)) ;
    nor03_2x ix217 (.Y (nx216), .A0 (gen_0_cmp_mReg_7), .A1 (nx10426), .A2 (
             nx10892)) ;
    nor03_2x ix213 (.Y (nx212), .A0 (nx3870), .A1 (nx10898), .A2 (nx10908)) ;
    nor02_2x ix3880 (.Y (nx3879), .A0 (nx208), .A1 (nx206)) ;
    nor03_2x ix209 (.Y (nx208), .A0 (nx3883), .A1 (nx10420), .A2 (nx10916)) ;
    dffr gen_0_cmp_mRegCmp_reg_Q_8 (.Q (gen_0_cmp_mReg_8), .QB (nx3883), .D (
         window_0__8), .CLK (start), .R (rst)) ;
    nor03_2x ix207 (.Y (nx206), .A0 (gen_0_cmp_mReg_8), .A1 (nx10732), .A2 (
             nx10924)) ;
    nand02 ix243 (.Y (gen_0_cmp_BSCmp_op2_9), .A0 (nx3889), .A1 (nx3895)) ;
    nor02_2x ix3890 (.Y (nx3889), .A0 (nx238), .A1 (nx234)) ;
    nor03_2x ix239 (.Y (nx238), .A0 (gen_0_cmp_mReg_8), .A1 (nx10426), .A2 (
             nx10892)) ;
    nor03_2x ix235 (.Y (nx234), .A0 (nx3883), .A1 (nx10898), .A2 (nx10908)) ;
    nor02_2x ix3896 (.Y (nx3895), .A0 (nx230), .A1 (nx228)) ;
    nor03_2x ix231 (.Y (nx230), .A0 (nx3899), .A1 (nx10420), .A2 (nx10916)) ;
    dffr gen_0_cmp_mRegCmp_reg_Q_9 (.Q (gen_0_cmp_mReg_9), .QB (nx3899), .D (
         window_0__9), .CLK (start), .R (rst)) ;
    nor03_2x ix229 (.Y (nx228), .A0 (gen_0_cmp_mReg_9), .A1 (nx10732), .A2 (
             nx10924)) ;
    nand02 ix265 (.Y (gen_0_cmp_BSCmp_op2_10), .A0 (nx3903), .A1 (nx3909)) ;
    nor02_2x ix3904 (.Y (nx3903), .A0 (nx260), .A1 (nx256)) ;
    nor03_2x ix261 (.Y (nx260), .A0 (gen_0_cmp_mReg_9), .A1 (nx10426), .A2 (
             nx10892)) ;
    nor03_2x ix257 (.Y (nx256), .A0 (nx3899), .A1 (nx10898), .A2 (nx10908)) ;
    nor02_2x ix3910 (.Y (nx3909), .A0 (nx252), .A1 (nx250)) ;
    nor03_2x ix253 (.Y (nx252), .A0 (nx3913), .A1 (nx10420), .A2 (nx10916)) ;
    dffr gen_0_cmp_mRegCmp_reg_Q_10 (.Q (gen_0_cmp_mReg_10), .QB (nx3913), .D (
         window_0__10), .CLK (start), .R (rst)) ;
    nor03_2x ix251 (.Y (nx250), .A0 (gen_0_cmp_mReg_10), .A1 (nx10732), .A2 (
             nx10924)) ;
    nand02 ix287 (.Y (gen_0_cmp_BSCmp_op2_11), .A0 (nx3919), .A1 (nx3923)) ;
    nor02_2x ix3920 (.Y (nx3919), .A0 (nx282), .A1 (nx278)) ;
    nor03_2x ix283 (.Y (nx282), .A0 (gen_0_cmp_mReg_10), .A1 (nx10426), .A2 (
             nx10892)) ;
    nor03_2x ix279 (.Y (nx278), .A0 (nx3913), .A1 (nx10898), .A2 (nx10908)) ;
    nor02_2x ix3924 (.Y (nx3923), .A0 (nx274), .A1 (nx272)) ;
    nor03_2x ix275 (.Y (nx274), .A0 (nx3927), .A1 (nx10420), .A2 (nx10916)) ;
    dffr gen_0_cmp_mRegCmp_reg_Q_11 (.Q (gen_0_cmp_mReg_11), .QB (nx3927), .D (
         window_0__11), .CLK (start), .R (rst)) ;
    nor03_2x ix273 (.Y (nx272), .A0 (gen_0_cmp_mReg_11), .A1 (nx10732), .A2 (
             nx10924)) ;
    nand02 ix309 (.Y (gen_0_cmp_BSCmp_op2_12), .A0 (nx3931), .A1 (nx3937)) ;
    nor02_2x ix3932 (.Y (nx3931), .A0 (nx304), .A1 (nx300)) ;
    nor03_2x ix305 (.Y (nx304), .A0 (gen_0_cmp_mReg_11), .A1 (nx10426), .A2 (
             nx10892)) ;
    nor03_2x ix301 (.Y (nx300), .A0 (nx3927), .A1 (nx10898), .A2 (nx10908)) ;
    nor02_2x ix3938 (.Y (nx3937), .A0 (nx296), .A1 (nx294)) ;
    nor03_2x ix297 (.Y (nx296), .A0 (nx3941), .A1 (nx10422), .A2 (nx10916)) ;
    dffr gen_0_cmp_mRegCmp_reg_Q_12 (.Q (gen_0_cmp_mReg_12), .QB (nx3941), .D (
         window_0__12), .CLK (start), .R (rst)) ;
    nor03_2x ix295 (.Y (nx294), .A0 (gen_0_cmp_mReg_12), .A1 (nx10732), .A2 (
             nx10924)) ;
    nand02 ix331 (.Y (gen_0_cmp_BSCmp_op2_13), .A0 (nx3945), .A1 (nx3951)) ;
    nor02_2x ix3946 (.Y (nx3945), .A0 (nx326), .A1 (nx322)) ;
    nor03_2x ix327 (.Y (nx326), .A0 (gen_0_cmp_mReg_12), .A1 (nx10428), .A2 (
             nx10894)) ;
    nor03_2x ix323 (.Y (nx322), .A0 (nx3941), .A1 (nx10898), .A2 (nx10910)) ;
    nor02_2x ix3952 (.Y (nx3951), .A0 (nx318), .A1 (nx316)) ;
    nor03_2x ix319 (.Y (nx318), .A0 (nx3954), .A1 (nx10422), .A2 (nx10918)) ;
    dffr gen_0_cmp_mRegCmp_reg_Q_13 (.Q (gen_0_cmp_mReg_13), .QB (nx3954), .D (
         window_0__13), .CLK (start), .R (rst)) ;
    nor03_2x ix317 (.Y (nx316), .A0 (gen_0_cmp_mReg_13), .A1 (nx10732), .A2 (
             nx10926)) ;
    nand02 ix353 (.Y (gen_0_cmp_BSCmp_op2_14), .A0 (nx3961), .A1 (nx3967)) ;
    nor02_2x ix3962 (.Y (nx3961), .A0 (nx348), .A1 (nx344)) ;
    nor03_2x ix349 (.Y (nx348), .A0 (gen_0_cmp_mReg_13), .A1 (nx10428), .A2 (
             nx10894)) ;
    nor03_2x ix345 (.Y (nx344), .A0 (nx3954), .A1 (nx10900), .A2 (nx10910)) ;
    nor02_2x ix3968 (.Y (nx3967), .A0 (nx340), .A1 (nx338)) ;
    nor03_2x ix341 (.Y (nx340), .A0 (nx3971), .A1 (nx10422), .A2 (nx10918)) ;
    dffr gen_0_cmp_mRegCmp_reg_Q_14 (.Q (gen_0_cmp_mReg_14), .QB (nx3971), .D (
         window_0__14), .CLK (start), .R (rst)) ;
    nor03_2x ix339 (.Y (nx338), .A0 (gen_0_cmp_mReg_14), .A1 (nx10732), .A2 (
             nx10926)) ;
    nand02 ix375 (.Y (gen_0_cmp_BSCmp_op2_15), .A0 (nx3975), .A1 (nx3981)) ;
    nor02_2x ix3976 (.Y (nx3975), .A0 (nx370), .A1 (nx366)) ;
    nor03_2x ix371 (.Y (nx370), .A0 (gen_0_cmp_mReg_14), .A1 (nx10428), .A2 (
             nx10894)) ;
    nor03_2x ix367 (.Y (nx366), .A0 (nx3971), .A1 (nx10900), .A2 (nx10910)) ;
    nor02_2x ix3982 (.Y (nx3981), .A0 (nx362), .A1 (nx360)) ;
    nor03_2x ix363 (.Y (nx362), .A0 (nx3985), .A1 (nx10422), .A2 (nx10918)) ;
    dffr gen_0_cmp_mRegCmp_reg_Q_15 (.Q (gen_0_cmp_mReg_15), .QB (nx3985), .D (
         window_0__15), .CLK (start), .R (rst)) ;
    nor03_2x ix361 (.Y (nx360), .A0 (gen_0_cmp_mReg_15), .A1 (nx10734), .A2 (
             nx10926)) ;
    nand02 ix385 (.Y (gen_0_cmp_BSCmp_op2_16), .A0 (nx3989), .A1 (nx3981)) ;
    nor02_2x ix3990 (.Y (nx3989), .A0 (nx380), .A1 (nx376)) ;
    nor03_2x ix381 (.Y (nx380), .A0 (gen_0_cmp_mReg_15), .A1 (nx10428), .A2 (
             nx10894)) ;
    nor03_2x ix377 (.Y (nx376), .A0 (nx3985), .A1 (nx10900), .A2 (nx10910)) ;
    nand02 ix453 (.Y (gen_1_cmp_BSCmp_op2_1), .A0 (nx3996), .A1 (nx4015)) ;
    nor02_2x ix3997 (.Y (nx3996), .A0 (nx448), .A1 (nx444)) ;
    nor03_2x ix449 (.Y (nx448), .A0 (gen_1_cmp_mReg_0), .A1 (nx10412), .A2 (
             nx10930)) ;
    dffr gen_1_cmp_mRegCmp_reg_Q_0 (.Q (gen_1_cmp_mReg_0), .QB (nx4001), .D (
         window_1__0), .CLK (start), .R (rst)) ;
    inv01 ix4006 (.Y (nx4005), .A (gen_1_cmp_pMux_0)) ;
    nor03_2x ix445 (.Y (nx444), .A0 (nx4001), .A1 (nx10936), .A2 (nx10946)) ;
    inv02 ix4014 (.Y (nx4013), .A (gen_1_cmp_pMux_2)) ;
    nor02_2x ix4016 (.Y (nx4015), .A0 (nx434), .A1 (nx432)) ;
    nor03_2x ix435 (.Y (nx434), .A0 (nx4018), .A1 (nx10406), .A2 (nx10954)) ;
    dffr gen_1_cmp_mRegCmp_reg_Q_1 (.Q (gen_1_cmp_mReg_1), .QB (nx4018), .D (
         window_1__1), .CLK (start), .R (rst)) ;
    nor03_2x ix433 (.Y (nx432), .A0 (gen_1_cmp_mReg_1), .A1 (nx10736), .A2 (
             nx10962)) ;
    nor03_2x ix393 (.Y (nx392), .A0 (nx10412), .A1 (nx4013), .A2 (
             gen_1_cmp_pMux_0)) ;
    nand02 ix475 (.Y (gen_1_cmp_BSCmp_op2_2), .A0 (nx4031), .A1 (nx4037)) ;
    nor02_2x ix4032 (.Y (nx4031), .A0 (nx470), .A1 (nx466)) ;
    nor03_2x ix471 (.Y (nx470), .A0 (gen_1_cmp_mReg_1), .A1 (nx10412), .A2 (
             nx10930)) ;
    nor03_2x ix467 (.Y (nx466), .A0 (nx4018), .A1 (nx10936), .A2 (nx10946)) ;
    nor02_2x ix4038 (.Y (nx4037), .A0 (nx462), .A1 (nx460)) ;
    nor03_2x ix463 (.Y (nx462), .A0 (nx4040), .A1 (nx10406), .A2 (nx10954)) ;
    dffr gen_1_cmp_mRegCmp_reg_Q_2 (.Q (gen_1_cmp_mReg_2), .QB (nx4040), .D (
         window_1__2), .CLK (start), .R (rst)) ;
    nor03_2x ix461 (.Y (nx460), .A0 (gen_1_cmp_mReg_2), .A1 (nx10736), .A2 (
             nx10962)) ;
    nand02 ix497 (.Y (gen_1_cmp_BSCmp_op2_3), .A0 (nx4045), .A1 (nx4051)) ;
    nor02_2x ix4046 (.Y (nx4045), .A0 (nx492), .A1 (nx488)) ;
    nor03_2x ix493 (.Y (nx492), .A0 (gen_1_cmp_mReg_2), .A1 (nx10412), .A2 (
             nx10930)) ;
    nor03_2x ix489 (.Y (nx488), .A0 (nx4040), .A1 (nx10936), .A2 (nx10946)) ;
    nor02_2x ix4052 (.Y (nx4051), .A0 (nx484), .A1 (nx482)) ;
    nor03_2x ix485 (.Y (nx484), .A0 (nx4055), .A1 (nx10406), .A2 (nx10954)) ;
    dffr gen_1_cmp_mRegCmp_reg_Q_3 (.Q (gen_1_cmp_mReg_3), .QB (nx4055), .D (
         window_1__3), .CLK (start), .R (rst)) ;
    nor03_2x ix483 (.Y (nx482), .A0 (gen_1_cmp_mReg_3), .A1 (nx10736), .A2 (
             nx10962)) ;
    nand02 ix519 (.Y (gen_1_cmp_BSCmp_op2_4), .A0 (nx4061), .A1 (nx4065)) ;
    nor02_2x ix4062 (.Y (nx4061), .A0 (nx514), .A1 (nx510)) ;
    nor03_2x ix515 (.Y (nx514), .A0 (gen_1_cmp_mReg_3), .A1 (nx10412), .A2 (
             nx10930)) ;
    nor03_2x ix511 (.Y (nx510), .A0 (nx4055), .A1 (nx10936), .A2 (nx10946)) ;
    nor02_2x ix4066 (.Y (nx4065), .A0 (nx506), .A1 (nx504)) ;
    nor03_2x ix507 (.Y (nx506), .A0 (nx4069), .A1 (nx10406), .A2 (nx10954)) ;
    dffr gen_1_cmp_mRegCmp_reg_Q_4 (.Q (gen_1_cmp_mReg_4), .QB (nx4069), .D (
         window_1__4), .CLK (start), .R (rst)) ;
    nor03_2x ix505 (.Y (nx504), .A0 (gen_1_cmp_mReg_4), .A1 (nx10736), .A2 (
             nx10962)) ;
    nand02 ix541 (.Y (gen_1_cmp_BSCmp_op2_5), .A0 (nx4075), .A1 (nx4081)) ;
    nor02_2x ix4076 (.Y (nx4075), .A0 (nx536), .A1 (nx532)) ;
    nor03_2x ix537 (.Y (nx536), .A0 (gen_1_cmp_mReg_4), .A1 (nx10412), .A2 (
             nx10930)) ;
    nor03_2x ix533 (.Y (nx532), .A0 (nx4069), .A1 (nx10936), .A2 (nx10946)) ;
    nor02_2x ix4082 (.Y (nx4081), .A0 (nx528), .A1 (nx526)) ;
    nor03_2x ix529 (.Y (nx528), .A0 (nx4084), .A1 (nx10408), .A2 (nx10954)) ;
    dffr gen_1_cmp_mRegCmp_reg_Q_5 (.Q (gen_1_cmp_mReg_5), .QB (nx4084), .D (
         window_1__5), .CLK (start), .R (rst)) ;
    nor03_2x ix527 (.Y (nx526), .A0 (gen_1_cmp_mReg_5), .A1 (nx10736), .A2 (
             nx10962)) ;
    nand02 ix563 (.Y (gen_1_cmp_BSCmp_op2_6), .A0 (nx4089), .A1 (nx4095)) ;
    nor02_2x ix4090 (.Y (nx4089), .A0 (nx558), .A1 (nx554)) ;
    nor03_2x ix559 (.Y (nx558), .A0 (gen_1_cmp_mReg_5), .A1 (nx10414), .A2 (
             nx10930)) ;
    nor03_2x ix555 (.Y (nx554), .A0 (nx4084), .A1 (nx10936), .A2 (nx10946)) ;
    nor02_2x ix4096 (.Y (nx4095), .A0 (nx550), .A1 (nx548)) ;
    nor03_2x ix551 (.Y (nx550), .A0 (nx4099), .A1 (nx10408), .A2 (nx10954)) ;
    dffr gen_1_cmp_mRegCmp_reg_Q_6 (.Q (gen_1_cmp_mReg_6), .QB (nx4099), .D (
         window_1__6), .CLK (start), .R (rst)) ;
    nor03_2x ix549 (.Y (nx548), .A0 (gen_1_cmp_mReg_6), .A1 (nx10736), .A2 (
             nx10962)) ;
    nand02 ix585 (.Y (gen_1_cmp_BSCmp_op2_7), .A0 (nx4105), .A1 (nx4109)) ;
    nor02_2x ix4106 (.Y (nx4105), .A0 (nx580), .A1 (nx576)) ;
    nor03_2x ix581 (.Y (nx580), .A0 (gen_1_cmp_mReg_6), .A1 (nx10414), .A2 (
             nx10932)) ;
    nor03_2x ix577 (.Y (nx576), .A0 (nx4099), .A1 (nx10938), .A2 (nx10948)) ;
    nor02_2x ix4110 (.Y (nx4109), .A0 (nx572), .A1 (nx570)) ;
    nor03_2x ix573 (.Y (nx572), .A0 (nx4113), .A1 (nx10408), .A2 (nx10956)) ;
    dffr gen_1_cmp_mRegCmp_reg_Q_7 (.Q (gen_1_cmp_mReg_7), .QB (nx4113), .D (
         window_1__7), .CLK (start), .R (rst)) ;
    nor03_2x ix571 (.Y (nx570), .A0 (gen_1_cmp_mReg_7), .A1 (nx10736), .A2 (
             nx10964)) ;
    nand02 ix607 (.Y (gen_1_cmp_BSCmp_op2_8), .A0 (nx4119), .A1 (nx4125)) ;
    nor02_2x ix4120 (.Y (nx4119), .A0 (nx602), .A1 (nx598)) ;
    nor03_2x ix603 (.Y (nx602), .A0 (gen_1_cmp_mReg_7), .A1 (nx10414), .A2 (
             nx10932)) ;
    nor03_2x ix599 (.Y (nx598), .A0 (nx4113), .A1 (nx10938), .A2 (nx10948)) ;
    nor02_2x ix4126 (.Y (nx4125), .A0 (nx594), .A1 (nx592)) ;
    nor03_2x ix595 (.Y (nx594), .A0 (nx4128), .A1 (nx10408), .A2 (nx10956)) ;
    dffr gen_1_cmp_mRegCmp_reg_Q_8 (.Q (gen_1_cmp_mReg_8), .QB (nx4128), .D (
         window_1__8), .CLK (start), .R (rst)) ;
    nor03_2x ix593 (.Y (nx592), .A0 (gen_1_cmp_mReg_8), .A1 (nx10738), .A2 (
             nx10964)) ;
    nand02 ix629 (.Y (gen_1_cmp_BSCmp_op2_9), .A0 (nx4133), .A1 (nx4139)) ;
    nor02_2x ix4134 (.Y (nx4133), .A0 (nx624), .A1 (nx620)) ;
    nor03_2x ix625 (.Y (nx624), .A0 (gen_1_cmp_mReg_8), .A1 (nx10414), .A2 (
             nx10932)) ;
    nor03_2x ix621 (.Y (nx620), .A0 (nx4128), .A1 (nx10938), .A2 (nx10948)) ;
    nor02_2x ix4140 (.Y (nx4139), .A0 (nx616), .A1 (nx614)) ;
    nor03_2x ix617 (.Y (nx616), .A0 (nx4143), .A1 (nx10408), .A2 (nx10956)) ;
    dffr gen_1_cmp_mRegCmp_reg_Q_9 (.Q (gen_1_cmp_mReg_9), .QB (nx4143), .D (
         window_1__9), .CLK (start), .R (rst)) ;
    nor03_2x ix615 (.Y (nx614), .A0 (gen_1_cmp_mReg_9), .A1 (nx10738), .A2 (
             nx10964)) ;
    nand02 ix651 (.Y (gen_1_cmp_BSCmp_op2_10), .A0 (nx4149), .A1 (nx4153)) ;
    nor02_2x ix4150 (.Y (nx4149), .A0 (nx646), .A1 (nx642)) ;
    nor03_2x ix647 (.Y (nx646), .A0 (gen_1_cmp_mReg_9), .A1 (nx10414), .A2 (
             nx10932)) ;
    nor03_2x ix643 (.Y (nx642), .A0 (nx4143), .A1 (nx10938), .A2 (nx10948)) ;
    nor02_2x ix4154 (.Y (nx4153), .A0 (nx638), .A1 (nx636)) ;
    nor03_2x ix639 (.Y (nx638), .A0 (nx4157), .A1 (nx10408), .A2 (nx10956)) ;
    dffr gen_1_cmp_mRegCmp_reg_Q_10 (.Q (gen_1_cmp_mReg_10), .QB (nx4157), .D (
         window_1__10), .CLK (start), .R (rst)) ;
    nor03_2x ix637 (.Y (nx636), .A0 (gen_1_cmp_mReg_10), .A1 (nx10738), .A2 (
             nx10964)) ;
    nand02 ix673 (.Y (gen_1_cmp_BSCmp_op2_11), .A0 (nx4163), .A1 (nx4169)) ;
    nor02_2x ix4164 (.Y (nx4163), .A0 (nx668), .A1 (nx664)) ;
    nor03_2x ix669 (.Y (nx668), .A0 (gen_1_cmp_mReg_10), .A1 (nx10414), .A2 (
             nx10932)) ;
    nor03_2x ix665 (.Y (nx664), .A0 (nx4157), .A1 (nx10938), .A2 (nx10948)) ;
    nor02_2x ix4170 (.Y (nx4169), .A0 (nx660), .A1 (nx658)) ;
    nor03_2x ix661 (.Y (nx660), .A0 (nx4172), .A1 (nx10408), .A2 (nx10956)) ;
    dffr gen_1_cmp_mRegCmp_reg_Q_11 (.Q (gen_1_cmp_mReg_11), .QB (nx4172), .D (
         window_1__11), .CLK (start), .R (rst)) ;
    nor03_2x ix659 (.Y (nx658), .A0 (gen_1_cmp_mReg_11), .A1 (nx10738), .A2 (
             nx10964)) ;
    nand02 ix695 (.Y (gen_1_cmp_BSCmp_op2_12), .A0 (nx4177), .A1 (nx4183)) ;
    nor02_2x ix4178 (.Y (nx4177), .A0 (nx690), .A1 (nx686)) ;
    nor03_2x ix691 (.Y (nx690), .A0 (gen_1_cmp_mReg_11), .A1 (nx10414), .A2 (
             nx10932)) ;
    nor03_2x ix687 (.Y (nx686), .A0 (nx4172), .A1 (nx10938), .A2 (nx10948)) ;
    nor02_2x ix4184 (.Y (nx4183), .A0 (nx682), .A1 (nx680)) ;
    nor03_2x ix683 (.Y (nx682), .A0 (nx4187), .A1 (nx10410), .A2 (nx10956)) ;
    dffr gen_1_cmp_mRegCmp_reg_Q_12 (.Q (gen_1_cmp_mReg_12), .QB (nx4187), .D (
         window_1__12), .CLK (start), .R (rst)) ;
    nor03_2x ix681 (.Y (nx680), .A0 (gen_1_cmp_mReg_12), .A1 (nx10738), .A2 (
             nx10964)) ;
    nand02 ix717 (.Y (gen_1_cmp_BSCmp_op2_13), .A0 (nx4193), .A1 (nx4197)) ;
    nor02_2x ix4194 (.Y (nx4193), .A0 (nx712), .A1 (nx708)) ;
    nor03_2x ix713 (.Y (nx712), .A0 (gen_1_cmp_mReg_12), .A1 (nx10416), .A2 (
             nx10934)) ;
    nor03_2x ix709 (.Y (nx708), .A0 (nx4187), .A1 (nx10938), .A2 (nx10950)) ;
    nor02_2x ix4198 (.Y (nx4197), .A0 (nx704), .A1 (nx702)) ;
    nor03_2x ix705 (.Y (nx704), .A0 (nx4201), .A1 (nx10410), .A2 (nx10958)) ;
    dffr gen_1_cmp_mRegCmp_reg_Q_13 (.Q (gen_1_cmp_mReg_13), .QB (nx4201), .D (
         window_1__13), .CLK (start), .R (rst)) ;
    nor03_2x ix703 (.Y (nx702), .A0 (gen_1_cmp_mReg_13), .A1 (nx10738), .A2 (
             nx10966)) ;
    nand02 ix739 (.Y (gen_1_cmp_BSCmp_op2_14), .A0 (nx4207), .A1 (nx4213)) ;
    nor02_2x ix4208 (.Y (nx4207), .A0 (nx734), .A1 (nx730)) ;
    nor03_2x ix735 (.Y (nx734), .A0 (gen_1_cmp_mReg_13), .A1 (nx10416), .A2 (
             nx10934)) ;
    nor03_2x ix731 (.Y (nx730), .A0 (nx4201), .A1 (nx10940), .A2 (nx10950)) ;
    nor02_2x ix4214 (.Y (nx4213), .A0 (nx726), .A1 (nx724)) ;
    nor03_2x ix727 (.Y (nx726), .A0 (nx4216), .A1 (nx10410), .A2 (nx10958)) ;
    dffr gen_1_cmp_mRegCmp_reg_Q_14 (.Q (gen_1_cmp_mReg_14), .QB (nx4216), .D (
         window_1__14), .CLK (start), .R (rst)) ;
    nor03_2x ix725 (.Y (nx724), .A0 (gen_1_cmp_mReg_14), .A1 (nx10738), .A2 (
             nx10966)) ;
    nand02 ix761 (.Y (gen_1_cmp_BSCmp_op2_15), .A0 (nx4221), .A1 (nx4227)) ;
    nor02_2x ix4222 (.Y (nx4221), .A0 (nx756), .A1 (nx752)) ;
    nor03_2x ix757 (.Y (nx756), .A0 (gen_1_cmp_mReg_14), .A1 (nx10416), .A2 (
             nx10934)) ;
    nor03_2x ix753 (.Y (nx752), .A0 (nx4216), .A1 (nx10940), .A2 (nx10950)) ;
    nor02_2x ix4228 (.Y (nx4227), .A0 (nx748), .A1 (nx746)) ;
    nor03_2x ix749 (.Y (nx748), .A0 (nx4231), .A1 (nx10410), .A2 (nx10958)) ;
    dffr gen_1_cmp_mRegCmp_reg_Q_15 (.Q (gen_1_cmp_mReg_15), .QB (nx4231), .D (
         window_1__15), .CLK (start), .R (rst)) ;
    nor03_2x ix747 (.Y (nx746), .A0 (gen_1_cmp_mReg_15), .A1 (nx10740), .A2 (
             nx10966)) ;
    nand02 ix771 (.Y (gen_1_cmp_BSCmp_op2_16), .A0 (nx4237), .A1 (nx4227)) ;
    nor02_2x ix4238 (.Y (nx4237), .A0 (nx766), .A1 (nx762)) ;
    nor03_2x ix767 (.Y (nx766), .A0 (gen_1_cmp_mReg_15), .A1 (nx10416), .A2 (
             nx10934)) ;
    nor03_2x ix763 (.Y (nx762), .A0 (nx4231), .A1 (nx10940), .A2 (nx10950)) ;
    nand02 ix839 (.Y (gen_2_cmp_BSCmp_op2_1), .A0 (nx4243), .A1 (nx4263)) ;
    nor02_2x ix4244 (.Y (nx4243), .A0 (nx834), .A1 (nx830)) ;
    nor03_2x ix835 (.Y (nx834), .A0 (gen_2_cmp_mReg_0), .A1 (nx10400), .A2 (
             nx10970)) ;
    dffr gen_2_cmp_mRegCmp_reg_Q_0 (.Q (gen_2_cmp_mReg_0), .QB (nx4249), .D (
         window_2__0), .CLK (start), .R (rst)) ;
    inv01 ix4254 (.Y (nx4253), .A (gen_2_cmp_pMux_0)) ;
    nor03_2x ix831 (.Y (nx830), .A0 (nx4249), .A1 (nx10976), .A2 (nx10986)) ;
    inv02 ix4261 (.Y (nx4260), .A (gen_2_cmp_pMux_2)) ;
    nor02_2x ix4264 (.Y (nx4263), .A0 (nx820), .A1 (nx818)) ;
    nor03_2x ix821 (.Y (nx820), .A0 (nx4267), .A1 (nx10394), .A2 (nx10994)) ;
    dffr gen_2_cmp_mRegCmp_reg_Q_1 (.Q (gen_2_cmp_mReg_1), .QB (nx4267), .D (
         window_2__1), .CLK (start), .R (rst)) ;
    nor03_2x ix819 (.Y (nx818), .A0 (gen_2_cmp_mReg_1), .A1 (nx10742), .A2 (
             nx11002)) ;
    nor03_2x ix779 (.Y (nx778), .A0 (nx10400), .A1 (nx4260), .A2 (
             gen_2_cmp_pMux_0)) ;
    nand02 ix861 (.Y (gen_2_cmp_BSCmp_op2_2), .A0 (nx4279), .A1 (nx4285)) ;
    nor02_2x ix4280 (.Y (nx4279), .A0 (nx856), .A1 (nx852)) ;
    nor03_2x ix857 (.Y (nx856), .A0 (gen_2_cmp_mReg_1), .A1 (nx10400), .A2 (
             nx10970)) ;
    nor03_2x ix853 (.Y (nx852), .A0 (nx4267), .A1 (nx10976), .A2 (nx10986)) ;
    nor02_2x ix4286 (.Y (nx4285), .A0 (nx848), .A1 (nx846)) ;
    nor03_2x ix849 (.Y (nx848), .A0 (nx4288), .A1 (nx10394), .A2 (nx10994)) ;
    dffr gen_2_cmp_mRegCmp_reg_Q_2 (.Q (gen_2_cmp_mReg_2), .QB (nx4288), .D (
         window_2__2), .CLK (start), .R (rst)) ;
    nor03_2x ix847 (.Y (nx846), .A0 (gen_2_cmp_mReg_2), .A1 (nx10742), .A2 (
             nx11002)) ;
    nand02 ix883 (.Y (gen_2_cmp_BSCmp_op2_3), .A0 (nx4293), .A1 (nx4299)) ;
    nor02_2x ix4294 (.Y (nx4293), .A0 (nx878), .A1 (nx874)) ;
    nor03_2x ix879 (.Y (nx878), .A0 (gen_2_cmp_mReg_2), .A1 (nx10400), .A2 (
             nx10970)) ;
    nor03_2x ix875 (.Y (nx874), .A0 (nx4288), .A1 (nx10976), .A2 (nx10986)) ;
    nor02_2x ix4300 (.Y (nx4299), .A0 (nx870), .A1 (nx868)) ;
    nor03_2x ix871 (.Y (nx870), .A0 (nx4303), .A1 (nx10394), .A2 (nx10994)) ;
    dffr gen_2_cmp_mRegCmp_reg_Q_3 (.Q (gen_2_cmp_mReg_3), .QB (nx4303), .D (
         window_2__3), .CLK (start), .R (rst)) ;
    nor03_2x ix869 (.Y (nx868), .A0 (gen_2_cmp_mReg_3), .A1 (nx10742), .A2 (
             nx11002)) ;
    nand02 ix905 (.Y (gen_2_cmp_BSCmp_op2_4), .A0 (nx4309), .A1 (nx4315)) ;
    nor02_2x ix4310 (.Y (nx4309), .A0 (nx900), .A1 (nx896)) ;
    nor03_2x ix901 (.Y (nx900), .A0 (gen_2_cmp_mReg_3), .A1 (nx10400), .A2 (
             nx10970)) ;
    nor03_2x ix897 (.Y (nx896), .A0 (nx4303), .A1 (nx10976), .A2 (nx10986)) ;
    nor02_2x ix4316 (.Y (nx4315), .A0 (nx892), .A1 (nx890)) ;
    nor03_2x ix893 (.Y (nx892), .A0 (nx4318), .A1 (nx10394), .A2 (nx10994)) ;
    dffr gen_2_cmp_mRegCmp_reg_Q_4 (.Q (gen_2_cmp_mReg_4), .QB (nx4318), .D (
         window_2__4), .CLK (start), .R (rst)) ;
    nor03_2x ix891 (.Y (nx890), .A0 (gen_2_cmp_mReg_4), .A1 (nx10742), .A2 (
             nx11002)) ;
    nand02 ix927 (.Y (gen_2_cmp_BSCmp_op2_5), .A0 (nx4325), .A1 (nx4331)) ;
    nor02_2x ix4326 (.Y (nx4325), .A0 (nx922), .A1 (nx918)) ;
    nor03_2x ix923 (.Y (nx922), .A0 (gen_2_cmp_mReg_4), .A1 (nx10400), .A2 (
             nx10970)) ;
    nor03_2x ix919 (.Y (nx918), .A0 (nx4318), .A1 (nx10976), .A2 (nx10986)) ;
    nor02_2x ix4332 (.Y (nx4331), .A0 (nx914), .A1 (nx912)) ;
    nor03_2x ix915 (.Y (nx914), .A0 (nx4335), .A1 (nx10396), .A2 (nx10994)) ;
    dffr gen_2_cmp_mRegCmp_reg_Q_5 (.Q (gen_2_cmp_mReg_5), .QB (nx4335), .D (
         window_2__5), .CLK (start), .R (rst)) ;
    nor03_2x ix913 (.Y (nx912), .A0 (gen_2_cmp_mReg_5), .A1 (nx10742), .A2 (
             nx11002)) ;
    nand02 ix949 (.Y (gen_2_cmp_BSCmp_op2_6), .A0 (nx4339), .A1 (nx4345)) ;
    nor02_2x ix4340 (.Y (nx4339), .A0 (nx944), .A1 (nx940)) ;
    nor03_2x ix945 (.Y (nx944), .A0 (gen_2_cmp_mReg_5), .A1 (nx10402), .A2 (
             nx10970)) ;
    nor03_2x ix941 (.Y (nx940), .A0 (nx4335), .A1 (nx10976), .A2 (nx10986)) ;
    nor02_2x ix4346 (.Y (nx4345), .A0 (nx936), .A1 (nx934)) ;
    nor03_2x ix937 (.Y (nx936), .A0 (nx4349), .A1 (nx10396), .A2 (nx10994)) ;
    dffr gen_2_cmp_mRegCmp_reg_Q_6 (.Q (gen_2_cmp_mReg_6), .QB (nx4349), .D (
         window_2__6), .CLK (start), .R (rst)) ;
    nor03_2x ix935 (.Y (nx934), .A0 (gen_2_cmp_mReg_6), .A1 (nx10742), .A2 (
             nx11002)) ;
    nand02 ix971 (.Y (gen_2_cmp_BSCmp_op2_7), .A0 (nx4353), .A1 (nx4359)) ;
    nor02_2x ix4354 (.Y (nx4353), .A0 (nx966), .A1 (nx962)) ;
    nor03_2x ix967 (.Y (nx966), .A0 (gen_2_cmp_mReg_6), .A1 (nx10402), .A2 (
             nx10972)) ;
    nor03_2x ix963 (.Y (nx962), .A0 (nx4349), .A1 (nx10978), .A2 (nx10988)) ;
    nor02_2x ix4360 (.Y (nx4359), .A0 (nx958), .A1 (nx956)) ;
    nor03_2x ix959 (.Y (nx958), .A0 (nx4362), .A1 (nx10396), .A2 (nx10996)) ;
    dffr gen_2_cmp_mRegCmp_reg_Q_7 (.Q (gen_2_cmp_mReg_7), .QB (nx4362), .D (
         window_2__7), .CLK (start), .R (rst)) ;
    nor03_2x ix957 (.Y (nx956), .A0 (gen_2_cmp_mReg_7), .A1 (nx10742), .A2 (
             nx11004)) ;
    nand02 ix993 (.Y (gen_2_cmp_BSCmp_op2_8), .A0 (nx4369), .A1 (nx4375)) ;
    nor02_2x ix4370 (.Y (nx4369), .A0 (nx988), .A1 (nx984)) ;
    nor03_2x ix989 (.Y (nx988), .A0 (gen_2_cmp_mReg_7), .A1 (nx10402), .A2 (
             nx10972)) ;
    nor03_2x ix985 (.Y (nx984), .A0 (nx4362), .A1 (nx10978), .A2 (nx10988)) ;
    nor02_2x ix4376 (.Y (nx4375), .A0 (nx980), .A1 (nx978)) ;
    nor03_2x ix981 (.Y (nx980), .A0 (nx4379), .A1 (nx10396), .A2 (nx10996)) ;
    dffr gen_2_cmp_mRegCmp_reg_Q_8 (.Q (gen_2_cmp_mReg_8), .QB (nx4379), .D (
         window_2__8), .CLK (start), .R (rst)) ;
    nor03_2x ix979 (.Y (nx978), .A0 (gen_2_cmp_mReg_8), .A1 (nx10744), .A2 (
             nx11004)) ;
    nand02 ix1015 (.Y (gen_2_cmp_BSCmp_op2_9), .A0 (nx4383), .A1 (nx4389)) ;
    nor02_2x ix4384 (.Y (nx4383), .A0 (nx1010), .A1 (nx1006)) ;
    nor03_2x ix1011 (.Y (nx1010), .A0 (gen_2_cmp_mReg_8), .A1 (nx10402), .A2 (
             nx10972)) ;
    nor03_2x ix1007 (.Y (nx1006), .A0 (nx4379), .A1 (nx10978), .A2 (nx10988)) ;
    nor02_2x ix4390 (.Y (nx4389), .A0 (nx1002), .A1 (nx1000)) ;
    nor03_2x ix1003 (.Y (nx1002), .A0 (nx4393), .A1 (nx10396), .A2 (nx10996)) ;
    dffr gen_2_cmp_mRegCmp_reg_Q_9 (.Q (gen_2_cmp_mReg_9), .QB (nx4393), .D (
         window_2__9), .CLK (start), .R (rst)) ;
    nor03_2x ix1001 (.Y (nx1000), .A0 (gen_2_cmp_mReg_9), .A1 (nx10744), .A2 (
             nx11004)) ;
    nand02 ix1037 (.Y (gen_2_cmp_BSCmp_op2_10), .A0 (nx4397), .A1 (nx4403)) ;
    nor02_2x ix4398 (.Y (nx4397), .A0 (nx1032), .A1 (nx1028)) ;
    nor03_2x ix1033 (.Y (nx1032), .A0 (gen_2_cmp_mReg_9), .A1 (nx10402), .A2 (
             nx10972)) ;
    nor03_2x ix1029 (.Y (nx1028), .A0 (nx4393), .A1 (nx10978), .A2 (nx10988)) ;
    nor02_2x ix4404 (.Y (nx4403), .A0 (nx1024), .A1 (nx1022)) ;
    nor03_2x ix1025 (.Y (nx1024), .A0 (nx4406), .A1 (nx10396), .A2 (nx10996)) ;
    dffr gen_2_cmp_mRegCmp_reg_Q_10 (.Q (gen_2_cmp_mReg_10), .QB (nx4406), .D (
         window_2__10), .CLK (start), .R (rst)) ;
    nor03_2x ix1023 (.Y (nx1022), .A0 (gen_2_cmp_mReg_10), .A1 (nx10744), .A2 (
             nx11004)) ;
    nand02 ix1059 (.Y (gen_2_cmp_BSCmp_op2_11), .A0 (nx4413), .A1 (nx4419)) ;
    nor02_2x ix4414 (.Y (nx4413), .A0 (nx1054), .A1 (nx1050)) ;
    nor03_2x ix1055 (.Y (nx1054), .A0 (gen_2_cmp_mReg_10), .A1 (nx10402), .A2 (
             nx10972)) ;
    nor03_2x ix1051 (.Y (nx1050), .A0 (nx4406), .A1 (nx10978), .A2 (nx10988)) ;
    nor02_2x ix4420 (.Y (nx4419), .A0 (nx1046), .A1 (nx1044)) ;
    nor03_2x ix1047 (.Y (nx1046), .A0 (nx4423), .A1 (nx10396), .A2 (nx10996)) ;
    dffr gen_2_cmp_mRegCmp_reg_Q_11 (.Q (gen_2_cmp_mReg_11), .QB (nx4423), .D (
         window_2__11), .CLK (start), .R (rst)) ;
    nor03_2x ix1045 (.Y (nx1044), .A0 (gen_2_cmp_mReg_11), .A1 (nx10744), .A2 (
             nx11004)) ;
    nand02 ix1081 (.Y (gen_2_cmp_BSCmp_op2_12), .A0 (nx4427), .A1 (nx4433)) ;
    nor02_2x ix4428 (.Y (nx4427), .A0 (nx1076), .A1 (nx1072)) ;
    nor03_2x ix1077 (.Y (nx1076), .A0 (gen_2_cmp_mReg_11), .A1 (nx10402), .A2 (
             nx10972)) ;
    nor03_2x ix1073 (.Y (nx1072), .A0 (nx4423), .A1 (nx10978), .A2 (nx10988)) ;
    nor02_2x ix4434 (.Y (nx4433), .A0 (nx1068), .A1 (nx1066)) ;
    nor03_2x ix1069 (.Y (nx1068), .A0 (nx4437), .A1 (nx10398), .A2 (nx10996)) ;
    dffr gen_2_cmp_mRegCmp_reg_Q_12 (.Q (gen_2_cmp_mReg_12), .QB (nx4437), .D (
         window_2__12), .CLK (start), .R (rst)) ;
    nor03_2x ix1067 (.Y (nx1066), .A0 (gen_2_cmp_mReg_12), .A1 (nx10744), .A2 (
             nx11004)) ;
    nand02 ix1103 (.Y (gen_2_cmp_BSCmp_op2_13), .A0 (nx4441), .A1 (nx4447)) ;
    nor02_2x ix4442 (.Y (nx4441), .A0 (nx1098), .A1 (nx1094)) ;
    nor03_2x ix1099 (.Y (nx1098), .A0 (gen_2_cmp_mReg_12), .A1 (nx10404), .A2 (
             nx10974)) ;
    nor03_2x ix1095 (.Y (nx1094), .A0 (nx4437), .A1 (nx10978), .A2 (nx10990)) ;
    nor02_2x ix4448 (.Y (nx4447), .A0 (nx1090), .A1 (nx1088)) ;
    nor03_2x ix1091 (.Y (nx1090), .A0 (nx4450), .A1 (nx10398), .A2 (nx10998)) ;
    dffr gen_2_cmp_mRegCmp_reg_Q_13 (.Q (gen_2_cmp_mReg_13), .QB (nx4450), .D (
         window_2__13), .CLK (start), .R (rst)) ;
    nor03_2x ix1089 (.Y (nx1088), .A0 (gen_2_cmp_mReg_13), .A1 (nx10744), .A2 (
             nx11006)) ;
    nand02 ix1125 (.Y (gen_2_cmp_BSCmp_op2_14), .A0 (nx4457), .A1 (nx4463)) ;
    nor02_2x ix4458 (.Y (nx4457), .A0 (nx1120), .A1 (nx1116)) ;
    nor03_2x ix1121 (.Y (nx1120), .A0 (gen_2_cmp_mReg_13), .A1 (nx10404), .A2 (
             nx10974)) ;
    nor03_2x ix1117 (.Y (nx1116), .A0 (nx4450), .A1 (nx10980), .A2 (nx10990)) ;
    nor02_2x ix4464 (.Y (nx4463), .A0 (nx1112), .A1 (nx1110)) ;
    nor03_2x ix1113 (.Y (nx1112), .A0 (nx4467), .A1 (nx10398), .A2 (nx10998)) ;
    dffr gen_2_cmp_mRegCmp_reg_Q_14 (.Q (gen_2_cmp_mReg_14), .QB (nx4467), .D (
         window_2__14), .CLK (start), .R (rst)) ;
    nor03_2x ix1111 (.Y (nx1110), .A0 (gen_2_cmp_mReg_14), .A1 (nx10744), .A2 (
             nx11006)) ;
    nand02 ix1147 (.Y (gen_2_cmp_BSCmp_op2_15), .A0 (nx4471), .A1 (nx4477)) ;
    nor02_2x ix4472 (.Y (nx4471), .A0 (nx1142), .A1 (nx1138)) ;
    nor03_2x ix1143 (.Y (nx1142), .A0 (gen_2_cmp_mReg_14), .A1 (nx10404), .A2 (
             nx10974)) ;
    nor03_2x ix1139 (.Y (nx1138), .A0 (nx4467), .A1 (nx10980), .A2 (nx10990)) ;
    nor02_2x ix4478 (.Y (nx4477), .A0 (nx1134), .A1 (nx1132)) ;
    nor03_2x ix1135 (.Y (nx1134), .A0 (nx4481), .A1 (nx10398), .A2 (nx10998)) ;
    dffr gen_2_cmp_mRegCmp_reg_Q_15 (.Q (gen_2_cmp_mReg_15), .QB (nx4481), .D (
         window_2__15), .CLK (start), .R (rst)) ;
    nor03_2x ix1133 (.Y (nx1132), .A0 (gen_2_cmp_mReg_15), .A1 (nx10746), .A2 (
             nx11006)) ;
    nand02 ix1157 (.Y (gen_2_cmp_BSCmp_op2_16), .A0 (nx4485), .A1 (nx4477)) ;
    nor02_2x ix4486 (.Y (nx4485), .A0 (nx1152), .A1 (nx1148)) ;
    nor03_2x ix1153 (.Y (nx1152), .A0 (gen_2_cmp_mReg_15), .A1 (nx10404), .A2 (
             nx10974)) ;
    nor03_2x ix1149 (.Y (nx1148), .A0 (nx4481), .A1 (nx10980), .A2 (nx10990)) ;
    nand02 ix1225 (.Y (gen_3_cmp_BSCmp_op2_1), .A0 (nx4492), .A1 (nx4511)) ;
    nor02_2x ix4493 (.Y (nx4492), .A0 (nx1220), .A1 (nx1216)) ;
    nor03_2x ix1221 (.Y (nx1220), .A0 (gen_3_cmp_mReg_0), .A1 (nx10388), .A2 (
             nx11010)) ;
    dffr gen_3_cmp_mRegCmp_reg_Q_0 (.Q (gen_3_cmp_mReg_0), .QB (nx4497), .D (
         window_3__0), .CLK (start), .R (rst)) ;
    inv01 ix4502 (.Y (nx4501), .A (gen_3_cmp_pMux_0)) ;
    nor03_2x ix1217 (.Y (nx1216), .A0 (nx4497), .A1 (nx11016), .A2 (nx11026)) ;
    inv02 ix4510 (.Y (nx4509), .A (gen_3_cmp_pMux_2)) ;
    nor02_2x ix4512 (.Y (nx4511), .A0 (nx1206), .A1 (nx1204)) ;
    nor03_2x ix1207 (.Y (nx1206), .A0 (nx4514), .A1 (nx10382), .A2 (nx11034)) ;
    dffr gen_3_cmp_mRegCmp_reg_Q_1 (.Q (gen_3_cmp_mReg_1), .QB (nx4514), .D (
         window_3__1), .CLK (start), .R (rst)) ;
    nor03_2x ix1205 (.Y (nx1204), .A0 (gen_3_cmp_mReg_1), .A1 (nx10748), .A2 (
             nx11042)) ;
    nor03_2x ix1165 (.Y (nx1164), .A0 (nx10388), .A1 (nx4509), .A2 (
             gen_3_cmp_pMux_0)) ;
    nand02 ix1247 (.Y (gen_3_cmp_BSCmp_op2_2), .A0 (nx4527), .A1 (nx4533)) ;
    nor02_2x ix4528 (.Y (nx4527), .A0 (nx1242), .A1 (nx1238)) ;
    nor03_2x ix1243 (.Y (nx1242), .A0 (gen_3_cmp_mReg_1), .A1 (nx10388), .A2 (
             nx11010)) ;
    nor03_2x ix1239 (.Y (nx1238), .A0 (nx4514), .A1 (nx11016), .A2 (nx11026)) ;
    nor02_2x ix4534 (.Y (nx4533), .A0 (nx1234), .A1 (nx1232)) ;
    nor03_2x ix1235 (.Y (nx1234), .A0 (nx4536), .A1 (nx10382), .A2 (nx11034)) ;
    dffr gen_3_cmp_mRegCmp_reg_Q_2 (.Q (gen_3_cmp_mReg_2), .QB (nx4536), .D (
         window_3__2), .CLK (start), .R (rst)) ;
    nor03_2x ix1233 (.Y (nx1232), .A0 (gen_3_cmp_mReg_2), .A1 (nx10748), .A2 (
             nx11042)) ;
    nand02 ix1269 (.Y (gen_3_cmp_BSCmp_op2_3), .A0 (nx4541), .A1 (nx4547)) ;
    nor02_2x ix4542 (.Y (nx4541), .A0 (nx1264), .A1 (nx1260)) ;
    nor03_2x ix1265 (.Y (nx1264), .A0 (gen_3_cmp_mReg_2), .A1 (nx10388), .A2 (
             nx11010)) ;
    nor03_2x ix1261 (.Y (nx1260), .A0 (nx4536), .A1 (nx11016), .A2 (nx11026)) ;
    nor02_2x ix4548 (.Y (nx4547), .A0 (nx1256), .A1 (nx1254)) ;
    nor03_2x ix1257 (.Y (nx1256), .A0 (nx4551), .A1 (nx10382), .A2 (nx11034)) ;
    dffr gen_3_cmp_mRegCmp_reg_Q_3 (.Q (gen_3_cmp_mReg_3), .QB (nx4551), .D (
         window_3__3), .CLK (start), .R (rst)) ;
    nor03_2x ix1255 (.Y (nx1254), .A0 (gen_3_cmp_mReg_3), .A1 (nx10748), .A2 (
             nx11042)) ;
    nand02 ix1291 (.Y (gen_3_cmp_BSCmp_op2_4), .A0 (nx4557), .A1 (nx4561)) ;
    nor02_2x ix4558 (.Y (nx4557), .A0 (nx1286), .A1 (nx1282)) ;
    nor03_2x ix1287 (.Y (nx1286), .A0 (gen_3_cmp_mReg_3), .A1 (nx10388), .A2 (
             nx11010)) ;
    nor03_2x ix1283 (.Y (nx1282), .A0 (nx4551), .A1 (nx11016), .A2 (nx11026)) ;
    nor02_2x ix4562 (.Y (nx4561), .A0 (nx1278), .A1 (nx1276)) ;
    nor03_2x ix1279 (.Y (nx1278), .A0 (nx4565), .A1 (nx10382), .A2 (nx11034)) ;
    dffr gen_3_cmp_mRegCmp_reg_Q_4 (.Q (gen_3_cmp_mReg_4), .QB (nx4565), .D (
         window_3__4), .CLK (start), .R (rst)) ;
    nor03_2x ix1277 (.Y (nx1276), .A0 (gen_3_cmp_mReg_4), .A1 (nx10748), .A2 (
             nx11042)) ;
    nand02 ix1313 (.Y (gen_3_cmp_BSCmp_op2_5), .A0 (nx4571), .A1 (nx4577)) ;
    nor02_2x ix4572 (.Y (nx4571), .A0 (nx1308), .A1 (nx1304)) ;
    nor03_2x ix1309 (.Y (nx1308), .A0 (gen_3_cmp_mReg_4), .A1 (nx10388), .A2 (
             nx11010)) ;
    nor03_2x ix1305 (.Y (nx1304), .A0 (nx4565), .A1 (nx11016), .A2 (nx11026)) ;
    nor02_2x ix4578 (.Y (nx4577), .A0 (nx1300), .A1 (nx1298)) ;
    nor03_2x ix1301 (.Y (nx1300), .A0 (nx4580), .A1 (nx10384), .A2 (nx11034)) ;
    dffr gen_3_cmp_mRegCmp_reg_Q_5 (.Q (gen_3_cmp_mReg_5), .QB (nx4580), .D (
         window_3__5), .CLK (start), .R (rst)) ;
    nor03_2x ix1299 (.Y (nx1298), .A0 (gen_3_cmp_mReg_5), .A1 (nx10748), .A2 (
             nx11042)) ;
    nand02 ix1335 (.Y (gen_3_cmp_BSCmp_op2_6), .A0 (nx4585), .A1 (nx4591)) ;
    nor02_2x ix4586 (.Y (nx4585), .A0 (nx1330), .A1 (nx1326)) ;
    nor03_2x ix1331 (.Y (nx1330), .A0 (gen_3_cmp_mReg_5), .A1 (nx10390), .A2 (
             nx11010)) ;
    nor03_2x ix1327 (.Y (nx1326), .A0 (nx4580), .A1 (nx11016), .A2 (nx11026)) ;
    nor02_2x ix4592 (.Y (nx4591), .A0 (nx1322), .A1 (nx1320)) ;
    nor03_2x ix1323 (.Y (nx1322), .A0 (nx4595), .A1 (nx10384), .A2 (nx11034)) ;
    dffr gen_3_cmp_mRegCmp_reg_Q_6 (.Q (gen_3_cmp_mReg_6), .QB (nx4595), .D (
         window_3__6), .CLK (start), .R (rst)) ;
    nor03_2x ix1321 (.Y (nx1320), .A0 (gen_3_cmp_mReg_6), .A1 (nx10748), .A2 (
             nx11042)) ;
    nand02 ix1357 (.Y (gen_3_cmp_BSCmp_op2_7), .A0 (nx4601), .A1 (nx4605)) ;
    nor02_2x ix4602 (.Y (nx4601), .A0 (nx1352), .A1 (nx1348)) ;
    nor03_2x ix1353 (.Y (nx1352), .A0 (gen_3_cmp_mReg_6), .A1 (nx10390), .A2 (
             nx11012)) ;
    nor03_2x ix1349 (.Y (nx1348), .A0 (nx4595), .A1 (nx11018), .A2 (nx11028)) ;
    nor02_2x ix4606 (.Y (nx4605), .A0 (nx1344), .A1 (nx1342)) ;
    nor03_2x ix1345 (.Y (nx1344), .A0 (nx4609), .A1 (nx10384), .A2 (nx11036)) ;
    dffr gen_3_cmp_mRegCmp_reg_Q_7 (.Q (gen_3_cmp_mReg_7), .QB (nx4609), .D (
         window_3__7), .CLK (start), .R (rst)) ;
    nor03_2x ix1343 (.Y (nx1342), .A0 (gen_3_cmp_mReg_7), .A1 (nx10748), .A2 (
             nx11044)) ;
    nand02 ix1379 (.Y (gen_3_cmp_BSCmp_op2_8), .A0 (nx4615), .A1 (nx4621)) ;
    nor02_2x ix4616 (.Y (nx4615), .A0 (nx1374), .A1 (nx1370)) ;
    nor03_2x ix1375 (.Y (nx1374), .A0 (gen_3_cmp_mReg_7), .A1 (nx10390), .A2 (
             nx11012)) ;
    nor03_2x ix1371 (.Y (nx1370), .A0 (nx4609), .A1 (nx11018), .A2 (nx11028)) ;
    nor02_2x ix4622 (.Y (nx4621), .A0 (nx1366), .A1 (nx1364)) ;
    nor03_2x ix1367 (.Y (nx1366), .A0 (nx4625), .A1 (nx10384), .A2 (nx11036)) ;
    dffr gen_3_cmp_mRegCmp_reg_Q_8 (.Q (gen_3_cmp_mReg_8), .QB (nx4625), .D (
         window_3__8), .CLK (start), .R (rst)) ;
    nor03_2x ix1365 (.Y (nx1364), .A0 (gen_3_cmp_mReg_8), .A1 (nx10750), .A2 (
             nx11044)) ;
    nand02 ix1401 (.Y (gen_3_cmp_BSCmp_op2_9), .A0 (nx4631), .A1 (nx4637)) ;
    nor02_2x ix4632 (.Y (nx4631), .A0 (nx1396), .A1 (nx1392)) ;
    nor03_2x ix1397 (.Y (nx1396), .A0 (gen_3_cmp_mReg_8), .A1 (nx10390), .A2 (
             nx11012)) ;
    nor03_2x ix1393 (.Y (nx1392), .A0 (nx4625), .A1 (nx11018), .A2 (nx11028)) ;
    nor02_2x ix4638 (.Y (nx4637), .A0 (nx1388), .A1 (nx1386)) ;
    nor03_2x ix1389 (.Y (nx1388), .A0 (nx4641), .A1 (nx10384), .A2 (nx11036)) ;
    dffr gen_3_cmp_mRegCmp_reg_Q_9 (.Q (gen_3_cmp_mReg_9), .QB (nx4641), .D (
         window_3__9), .CLK (start), .R (rst)) ;
    nor03_2x ix1387 (.Y (nx1386), .A0 (gen_3_cmp_mReg_9), .A1 (nx10750), .A2 (
             nx11044)) ;
    nand02 ix1423 (.Y (gen_3_cmp_BSCmp_op2_10), .A0 (nx4645), .A1 (nx4649)) ;
    nor02_2x ix4646 (.Y (nx4645), .A0 (nx1418), .A1 (nx1414)) ;
    nor03_2x ix1419 (.Y (nx1418), .A0 (gen_3_cmp_mReg_9), .A1 (nx10390), .A2 (
             nx11012)) ;
    nor03_2x ix1415 (.Y (nx1414), .A0 (nx4641), .A1 (nx11018), .A2 (nx11028)) ;
    nor02_2x ix4650 (.Y (nx4649), .A0 (nx1410), .A1 (nx1408)) ;
    nor03_2x ix1411 (.Y (nx1410), .A0 (nx4653), .A1 (nx10384), .A2 (nx11036)) ;
    dffr gen_3_cmp_mRegCmp_reg_Q_10 (.Q (gen_3_cmp_mReg_10), .QB (nx4653), .D (
         window_3__10), .CLK (start), .R (rst)) ;
    nor03_2x ix1409 (.Y (nx1408), .A0 (gen_3_cmp_mReg_10), .A1 (nx10750), .A2 (
             nx11044)) ;
    nand02 ix1445 (.Y (gen_3_cmp_BSCmp_op2_11), .A0 (nx4659), .A1 (nx4665)) ;
    nor02_2x ix4660 (.Y (nx4659), .A0 (nx1440), .A1 (nx1436)) ;
    nor03_2x ix1441 (.Y (nx1440), .A0 (gen_3_cmp_mReg_10), .A1 (nx10390), .A2 (
             nx11012)) ;
    nor03_2x ix1437 (.Y (nx1436), .A0 (nx4653), .A1 (nx11018), .A2 (nx11028)) ;
    nor02_2x ix4666 (.Y (nx4665), .A0 (nx1432), .A1 (nx1430)) ;
    nor03_2x ix1433 (.Y (nx1432), .A0 (nx4669), .A1 (nx10384), .A2 (nx11036)) ;
    dffr gen_3_cmp_mRegCmp_reg_Q_11 (.Q (gen_3_cmp_mReg_11), .QB (nx4669), .D (
         window_3__11), .CLK (start), .R (rst)) ;
    nor03_2x ix1431 (.Y (nx1430), .A0 (gen_3_cmp_mReg_11), .A1 (nx10750), .A2 (
             nx11044)) ;
    nand02 ix1467 (.Y (gen_3_cmp_BSCmp_op2_12), .A0 (nx4674), .A1 (nx4679)) ;
    nor02_2x ix4675 (.Y (nx4674), .A0 (nx1462), .A1 (nx1458)) ;
    nor03_2x ix1463 (.Y (nx1462), .A0 (gen_3_cmp_mReg_11), .A1 (nx10390), .A2 (
             nx11012)) ;
    nor03_2x ix1459 (.Y (nx1458), .A0 (nx4669), .A1 (nx11018), .A2 (nx11028)) ;
    nor02_2x ix4680 (.Y (nx4679), .A0 (nx1454), .A1 (nx1452)) ;
    nor03_2x ix1455 (.Y (nx1454), .A0 (nx4683), .A1 (nx10386), .A2 (nx11036)) ;
    dffr gen_3_cmp_mRegCmp_reg_Q_12 (.Q (gen_3_cmp_mReg_12), .QB (nx4683), .D (
         window_3__12), .CLK (start), .R (rst)) ;
    nor03_2x ix1453 (.Y (nx1452), .A0 (gen_3_cmp_mReg_12), .A1 (nx10750), .A2 (
             nx11044)) ;
    nand02 ix1489 (.Y (gen_3_cmp_BSCmp_op2_13), .A0 (nx4687), .A1 (nx4693)) ;
    nor02_2x ix4688 (.Y (nx4687), .A0 (nx1484), .A1 (nx1480)) ;
    nor03_2x ix1485 (.Y (nx1484), .A0 (gen_3_cmp_mReg_12), .A1 (nx10392), .A2 (
             nx11014)) ;
    nor03_2x ix1481 (.Y (nx1480), .A0 (nx4683), .A1 (nx11018), .A2 (nx11030)) ;
    nor02_2x ix4694 (.Y (nx4693), .A0 (nx1476), .A1 (nx1474)) ;
    nor03_2x ix1477 (.Y (nx1476), .A0 (nx4697), .A1 (nx10386), .A2 (nx11038)) ;
    dffr gen_3_cmp_mRegCmp_reg_Q_13 (.Q (gen_3_cmp_mReg_13), .QB (nx4697), .D (
         window_3__13), .CLK (start), .R (rst)) ;
    nor03_2x ix1475 (.Y (nx1474), .A0 (gen_3_cmp_mReg_13), .A1 (nx10750), .A2 (
             nx11046)) ;
    nand02 ix1511 (.Y (gen_3_cmp_BSCmp_op2_14), .A0 (nx4702), .A1 (nx4707)) ;
    nor02_2x ix4703 (.Y (nx4702), .A0 (nx1506), .A1 (nx1502)) ;
    nor03_2x ix1507 (.Y (nx1506), .A0 (gen_3_cmp_mReg_13), .A1 (nx10392), .A2 (
             nx11014)) ;
    nor03_2x ix1503 (.Y (nx1502), .A0 (nx4697), .A1 (nx11020), .A2 (nx11030)) ;
    nor02_2x ix4708 (.Y (nx4707), .A0 (nx1498), .A1 (nx1496)) ;
    nor03_2x ix1499 (.Y (nx1498), .A0 (nx4711), .A1 (nx10386), .A2 (nx11038)) ;
    dffr gen_3_cmp_mRegCmp_reg_Q_14 (.Q (gen_3_cmp_mReg_14), .QB (nx4711), .D (
         window_3__14), .CLK (start), .R (rst)) ;
    nor03_2x ix1497 (.Y (nx1496), .A0 (gen_3_cmp_mReg_14), .A1 (nx10750), .A2 (
             nx11046)) ;
    nand02 ix1533 (.Y (gen_3_cmp_BSCmp_op2_15), .A0 (nx4717), .A1 (nx4723)) ;
    nor02_2x ix4718 (.Y (nx4717), .A0 (nx1528), .A1 (nx1524)) ;
    nor03_2x ix1529 (.Y (nx1528), .A0 (gen_3_cmp_mReg_14), .A1 (nx10392), .A2 (
             nx11014)) ;
    nor03_2x ix1525 (.Y (nx1524), .A0 (nx4711), .A1 (nx11020), .A2 (nx11030)) ;
    nor02_2x ix4724 (.Y (nx4723), .A0 (nx1520), .A1 (nx1518)) ;
    nor03_2x ix1521 (.Y (nx1520), .A0 (nx4726), .A1 (nx10386), .A2 (nx11038)) ;
    dffr gen_3_cmp_mRegCmp_reg_Q_15 (.Q (gen_3_cmp_mReg_15), .QB (nx4726), .D (
         window_3__15), .CLK (start), .R (rst)) ;
    nor03_2x ix1519 (.Y (nx1518), .A0 (gen_3_cmp_mReg_15), .A1 (nx10752), .A2 (
             nx11046)) ;
    nand02 ix1543 (.Y (gen_3_cmp_BSCmp_op2_16), .A0 (nx4733), .A1 (nx4723)) ;
    nor02_2x ix4734 (.Y (nx4733), .A0 (nx1538), .A1 (nx1534)) ;
    nor03_2x ix1539 (.Y (nx1538), .A0 (gen_3_cmp_mReg_15), .A1 (nx10392), .A2 (
             nx11014)) ;
    nor03_2x ix1535 (.Y (nx1534), .A0 (nx4726), .A1 (nx11020), .A2 (nx11030)) ;
    nand02 ix1611 (.Y (gen_4_cmp_BSCmp_op2_1), .A0 (nx4739), .A1 (nx4759)) ;
    nor02_2x ix4740 (.Y (nx4739), .A0 (nx1606), .A1 (nx1602)) ;
    nor03_2x ix1607 (.Y (nx1606), .A0 (gen_4_cmp_mReg_0), .A1 (nx10376), .A2 (
             nx11050)) ;
    dffr gen_4_cmp_mRegCmp_reg_Q_0 (.Q (gen_4_cmp_mReg_0), .QB (nx4745), .D (
         window_4__0), .CLK (start), .R (rst)) ;
    inv01 ix4750 (.Y (nx4748), .A (gen_4_cmp_pMux_0)) ;
    nor03_2x ix1603 (.Y (nx1602), .A0 (nx4745), .A1 (nx11056), .A2 (nx11066)) ;
    inv02 ix4758 (.Y (nx4757), .A (gen_4_cmp_pMux_2)) ;
    nor02_2x ix4760 (.Y (nx4759), .A0 (nx1592), .A1 (nx1590)) ;
    nor03_2x ix1593 (.Y (nx1592), .A0 (nx4763), .A1 (nx10370), .A2 (nx11074)) ;
    dffr gen_4_cmp_mRegCmp_reg_Q_1 (.Q (gen_4_cmp_mReg_1), .QB (nx4763), .D (
         window_4__1), .CLK (start), .R (rst)) ;
    nor03_2x ix1591 (.Y (nx1590), .A0 (gen_4_cmp_mReg_1), .A1 (nx10754), .A2 (
             nx11082)) ;
    nor03_2x ix1551 (.Y (nx1550), .A0 (nx10376), .A1 (nx4757), .A2 (
             gen_4_cmp_pMux_0)) ;
    nand02 ix1633 (.Y (gen_4_cmp_BSCmp_op2_2), .A0 (nx4773), .A1 (nx4779)) ;
    nor02_2x ix4774 (.Y (nx4773), .A0 (nx1628), .A1 (nx1624)) ;
    nor03_2x ix1629 (.Y (nx1628), .A0 (gen_4_cmp_mReg_1), .A1 (nx10376), .A2 (
             nx11050)) ;
    nor03_2x ix1625 (.Y (nx1624), .A0 (nx4763), .A1 (nx11056), .A2 (nx11066)) ;
    nor02_2x ix4780 (.Y (nx4779), .A0 (nx1620), .A1 (nx1618)) ;
    nor03_2x ix1621 (.Y (nx1620), .A0 (nx4783), .A1 (nx10370), .A2 (nx11074)) ;
    dffr gen_4_cmp_mRegCmp_reg_Q_2 (.Q (gen_4_cmp_mReg_2), .QB (nx4783), .D (
         window_4__2), .CLK (start), .R (rst)) ;
    nor03_2x ix1619 (.Y (nx1618), .A0 (gen_4_cmp_mReg_2), .A1 (nx10754), .A2 (
             nx11082)) ;
    nand02 ix1655 (.Y (gen_4_cmp_BSCmp_op2_3), .A0 (nx4789), .A1 (nx4793)) ;
    nor02_2x ix4790 (.Y (nx4789), .A0 (nx1650), .A1 (nx1646)) ;
    nor03_2x ix1651 (.Y (nx1650), .A0 (gen_4_cmp_mReg_2), .A1 (nx10376), .A2 (
             nx11050)) ;
    nor03_2x ix1647 (.Y (nx1646), .A0 (nx4783), .A1 (nx11056), .A2 (nx11066)) ;
    nor02_2x ix4794 (.Y (nx4793), .A0 (nx1642), .A1 (nx1640)) ;
    nor03_2x ix1643 (.Y (nx1642), .A0 (nx4797), .A1 (nx10370), .A2 (nx11074)) ;
    dffr gen_4_cmp_mRegCmp_reg_Q_3 (.Q (gen_4_cmp_mReg_3), .QB (nx4797), .D (
         window_4__3), .CLK (start), .R (rst)) ;
    nor03_2x ix1641 (.Y (nx1640), .A0 (gen_4_cmp_mReg_3), .A1 (nx10754), .A2 (
             nx11082)) ;
    nand02 ix1677 (.Y (gen_4_cmp_BSCmp_op2_4), .A0 (nx4803), .A1 (nx4809)) ;
    nor02_2x ix4804 (.Y (nx4803), .A0 (nx1672), .A1 (nx1668)) ;
    nor03_2x ix1673 (.Y (nx1672), .A0 (gen_4_cmp_mReg_3), .A1 (nx10376), .A2 (
             nx11050)) ;
    nor03_2x ix1669 (.Y (nx1668), .A0 (nx4797), .A1 (nx11056), .A2 (nx11066)) ;
    nor02_2x ix4810 (.Y (nx4809), .A0 (nx1664), .A1 (nx1662)) ;
    nor03_2x ix1665 (.Y (nx1664), .A0 (nx4812), .A1 (nx10370), .A2 (nx11074)) ;
    dffr gen_4_cmp_mRegCmp_reg_Q_4 (.Q (gen_4_cmp_mReg_4), .QB (nx4812), .D (
         window_4__4), .CLK (start), .R (rst)) ;
    nor03_2x ix1663 (.Y (nx1662), .A0 (gen_4_cmp_mReg_4), .A1 (nx10754), .A2 (
             nx11082)) ;
    nand02 ix1699 (.Y (gen_4_cmp_BSCmp_op2_5), .A0 (nx4817), .A1 (nx4823)) ;
    nor02_2x ix4818 (.Y (nx4817), .A0 (nx1694), .A1 (nx1690)) ;
    nor03_2x ix1695 (.Y (nx1694), .A0 (gen_4_cmp_mReg_4), .A1 (nx10376), .A2 (
             nx11050)) ;
    nor03_2x ix1691 (.Y (nx1690), .A0 (nx4812), .A1 (nx11056), .A2 (nx11066)) ;
    nor02_2x ix4824 (.Y (nx4823), .A0 (nx1686), .A1 (nx1684)) ;
    nor03_2x ix1687 (.Y (nx1686), .A0 (nx4827), .A1 (nx10372), .A2 (nx11074)) ;
    dffr gen_4_cmp_mRegCmp_reg_Q_5 (.Q (gen_4_cmp_mReg_5), .QB (nx4827), .D (
         window_4__5), .CLK (start), .R (rst)) ;
    nor03_2x ix1685 (.Y (nx1684), .A0 (gen_4_cmp_mReg_5), .A1 (nx10754), .A2 (
             nx11082)) ;
    nand02 ix1721 (.Y (gen_4_cmp_BSCmp_op2_6), .A0 (nx4833), .A1 (nx4837)) ;
    nor02_2x ix4834 (.Y (nx4833), .A0 (nx1716), .A1 (nx1712)) ;
    nor03_2x ix1717 (.Y (nx1716), .A0 (gen_4_cmp_mReg_5), .A1 (nx10378), .A2 (
             nx11050)) ;
    nor03_2x ix1713 (.Y (nx1712), .A0 (nx4827), .A1 (nx11056), .A2 (nx11066)) ;
    nor02_2x ix4838 (.Y (nx4837), .A0 (nx1708), .A1 (nx1706)) ;
    nor03_2x ix1709 (.Y (nx1708), .A0 (nx4841), .A1 (nx10372), .A2 (nx11074)) ;
    dffr gen_4_cmp_mRegCmp_reg_Q_6 (.Q (gen_4_cmp_mReg_6), .QB (nx4841), .D (
         window_4__6), .CLK (start), .R (rst)) ;
    nor03_2x ix1707 (.Y (nx1706), .A0 (gen_4_cmp_mReg_6), .A1 (nx10754), .A2 (
             nx11082)) ;
    nand02 ix1743 (.Y (gen_4_cmp_BSCmp_op2_7), .A0 (nx4847), .A1 (nx4853)) ;
    nor02_2x ix4848 (.Y (nx4847), .A0 (nx1738), .A1 (nx1734)) ;
    nor03_2x ix1739 (.Y (nx1738), .A0 (gen_4_cmp_mReg_6), .A1 (nx10378), .A2 (
             nx11052)) ;
    nor03_2x ix1735 (.Y (nx1734), .A0 (nx4841), .A1 (nx11058), .A2 (nx11068)) ;
    nor02_2x ix4854 (.Y (nx4853), .A0 (nx1730), .A1 (nx1728)) ;
    nor03_2x ix1731 (.Y (nx1730), .A0 (nx4856), .A1 (nx10372), .A2 (nx11076)) ;
    dffr gen_4_cmp_mRegCmp_reg_Q_7 (.Q (gen_4_cmp_mReg_7), .QB (nx4856), .D (
         window_4__7), .CLK (start), .R (rst)) ;
    nor03_2x ix1729 (.Y (nx1728), .A0 (gen_4_cmp_mReg_7), .A1 (nx10754), .A2 (
             nx11084)) ;
    nand02 ix1765 (.Y (gen_4_cmp_BSCmp_op2_8), .A0 (nx4861), .A1 (nx4867)) ;
    nor02_2x ix4862 (.Y (nx4861), .A0 (nx1760), .A1 (nx1756)) ;
    nor03_2x ix1761 (.Y (nx1760), .A0 (gen_4_cmp_mReg_7), .A1 (nx10378), .A2 (
             nx11052)) ;
    nor03_2x ix1757 (.Y (nx1756), .A0 (nx4856), .A1 (nx11058), .A2 (nx11068)) ;
    nor02_2x ix4868 (.Y (nx4867), .A0 (nx1752), .A1 (nx1750)) ;
    nor03_2x ix1753 (.Y (nx1752), .A0 (nx4871), .A1 (nx10372), .A2 (nx11076)) ;
    dffr gen_4_cmp_mRegCmp_reg_Q_8 (.Q (gen_4_cmp_mReg_8), .QB (nx4871), .D (
         window_4__8), .CLK (start), .R (rst)) ;
    nor03_2x ix1751 (.Y (nx1750), .A0 (gen_4_cmp_mReg_8), .A1 (nx10756), .A2 (
             nx11084)) ;
    nand02 ix1787 (.Y (gen_4_cmp_BSCmp_op2_9), .A0 (nx4877), .A1 (nx4881)) ;
    nor02_2x ix4878 (.Y (nx4877), .A0 (nx1782), .A1 (nx1778)) ;
    nor03_2x ix1783 (.Y (nx1782), .A0 (gen_4_cmp_mReg_8), .A1 (nx10378), .A2 (
             nx11052)) ;
    nor03_2x ix1779 (.Y (nx1778), .A0 (nx4871), .A1 (nx11058), .A2 (nx11068)) ;
    nor02_2x ix4882 (.Y (nx4881), .A0 (nx1774), .A1 (nx1772)) ;
    nor03_2x ix1775 (.Y (nx1774), .A0 (nx4885), .A1 (nx10372), .A2 (nx11076)) ;
    dffr gen_4_cmp_mRegCmp_reg_Q_9 (.Q (gen_4_cmp_mReg_9), .QB (nx4885), .D (
         window_4__9), .CLK (start), .R (rst)) ;
    nor03_2x ix1773 (.Y (nx1772), .A0 (gen_4_cmp_mReg_9), .A1 (nx10756), .A2 (
             nx11084)) ;
    nand02 ix1809 (.Y (gen_4_cmp_BSCmp_op2_10), .A0 (nx4891), .A1 (nx4897)) ;
    nor02_2x ix4892 (.Y (nx4891), .A0 (nx1804), .A1 (nx1800)) ;
    nor03_2x ix1805 (.Y (nx1804), .A0 (gen_4_cmp_mReg_9), .A1 (nx10378), .A2 (
             nx11052)) ;
    nor03_2x ix1801 (.Y (nx1800), .A0 (nx4885), .A1 (nx11058), .A2 (nx11068)) ;
    nor02_2x ix4898 (.Y (nx4897), .A0 (nx1796), .A1 (nx1794)) ;
    nor03_2x ix1797 (.Y (nx1796), .A0 (nx4900), .A1 (nx10372), .A2 (nx11076)) ;
    dffr gen_4_cmp_mRegCmp_reg_Q_10 (.Q (gen_4_cmp_mReg_10), .QB (nx4900), .D (
         window_4__10), .CLK (start), .R (rst)) ;
    nor03_2x ix1795 (.Y (nx1794), .A0 (gen_4_cmp_mReg_10), .A1 (nx10756), .A2 (
             nx11084)) ;
    nand02 ix1831 (.Y (gen_4_cmp_BSCmp_op2_11), .A0 (nx4905), .A1 (nx4911)) ;
    nor02_2x ix4906 (.Y (nx4905), .A0 (nx1826), .A1 (nx1822)) ;
    nor03_2x ix1827 (.Y (nx1826), .A0 (gen_4_cmp_mReg_10), .A1 (nx10378), .A2 (
             nx11052)) ;
    nor03_2x ix1823 (.Y (nx1822), .A0 (nx4900), .A1 (nx11058), .A2 (nx11068)) ;
    nor02_2x ix4912 (.Y (nx4911), .A0 (nx1818), .A1 (nx1816)) ;
    nor03_2x ix1819 (.Y (nx1818), .A0 (nx4915), .A1 (nx10372), .A2 (nx11076)) ;
    dffr gen_4_cmp_mRegCmp_reg_Q_11 (.Q (gen_4_cmp_mReg_11), .QB (nx4915), .D (
         window_4__11), .CLK (start), .R (rst)) ;
    nor03_2x ix1817 (.Y (nx1816), .A0 (gen_4_cmp_mReg_11), .A1 (nx10756), .A2 (
             nx11084)) ;
    nand02 ix1853 (.Y (gen_4_cmp_BSCmp_op2_12), .A0 (nx4921), .A1 (nx4925)) ;
    nor02_2x ix4922 (.Y (nx4921), .A0 (nx1848), .A1 (nx1844)) ;
    nor03_2x ix1849 (.Y (nx1848), .A0 (gen_4_cmp_mReg_11), .A1 (nx10378), .A2 (
             nx11052)) ;
    nor03_2x ix1845 (.Y (nx1844), .A0 (nx4915), .A1 (nx11058), .A2 (nx11068)) ;
    nor02_2x ix4926 (.Y (nx4925), .A0 (nx1840), .A1 (nx1838)) ;
    nor03_2x ix1841 (.Y (nx1840), .A0 (nx4929), .A1 (nx10374), .A2 (nx11076)) ;
    dffr gen_4_cmp_mRegCmp_reg_Q_12 (.Q (gen_4_cmp_mReg_12), .QB (nx4929), .D (
         window_4__12), .CLK (start), .R (rst)) ;
    nor03_2x ix1839 (.Y (nx1838), .A0 (gen_4_cmp_mReg_12), .A1 (nx10756), .A2 (
             nx11084)) ;
    nand02 ix1875 (.Y (gen_4_cmp_BSCmp_op2_13), .A0 (nx4935), .A1 (nx4941)) ;
    nor02_2x ix4936 (.Y (nx4935), .A0 (nx1870), .A1 (nx1866)) ;
    nor03_2x ix1871 (.Y (nx1870), .A0 (gen_4_cmp_mReg_12), .A1 (nx10380), .A2 (
             nx11054)) ;
    nor03_2x ix1867 (.Y (nx1866), .A0 (nx4929), .A1 (nx11058), .A2 (nx11070)) ;
    nor02_2x ix4942 (.Y (nx4941), .A0 (nx1862), .A1 (nx1860)) ;
    nor03_2x ix1863 (.Y (nx1862), .A0 (nx4944), .A1 (nx10374), .A2 (nx11078)) ;
    dffr gen_4_cmp_mRegCmp_reg_Q_13 (.Q (gen_4_cmp_mReg_13), .QB (nx4944), .D (
         window_4__13), .CLK (start), .R (rst)) ;
    nor03_2x ix1861 (.Y (nx1860), .A0 (gen_4_cmp_mReg_13), .A1 (nx10756), .A2 (
             nx11086)) ;
    nand02 ix1897 (.Y (gen_4_cmp_BSCmp_op2_14), .A0 (nx4949), .A1 (nx4955)) ;
    nor02_2x ix4950 (.Y (nx4949), .A0 (nx1892), .A1 (nx1888)) ;
    nor03_2x ix1893 (.Y (nx1892), .A0 (gen_4_cmp_mReg_13), .A1 (nx10380), .A2 (
             nx11054)) ;
    nor03_2x ix1889 (.Y (nx1888), .A0 (nx4944), .A1 (nx11060), .A2 (nx11070)) ;
    nor02_2x ix4956 (.Y (nx4955), .A0 (nx1884), .A1 (nx1882)) ;
    nor03_2x ix1885 (.Y (nx1884), .A0 (nx4959), .A1 (nx10374), .A2 (nx11078)) ;
    dffr gen_4_cmp_mRegCmp_reg_Q_14 (.Q (gen_4_cmp_mReg_14), .QB (nx4959), .D (
         window_4__14), .CLK (start), .R (rst)) ;
    nor03_2x ix1883 (.Y (nx1882), .A0 (gen_4_cmp_mReg_14), .A1 (nx10756), .A2 (
             nx11086)) ;
    nand02 ix1919 (.Y (gen_4_cmp_BSCmp_op2_15), .A0 (nx4965), .A1 (nx4969)) ;
    nor02_2x ix4966 (.Y (nx4965), .A0 (nx1914), .A1 (nx1910)) ;
    nor03_2x ix1915 (.Y (nx1914), .A0 (gen_4_cmp_mReg_14), .A1 (nx10380), .A2 (
             nx11054)) ;
    nor03_2x ix1911 (.Y (nx1910), .A0 (nx4959), .A1 (nx11060), .A2 (nx11070)) ;
    nor02_2x ix4970 (.Y (nx4969), .A0 (nx1906), .A1 (nx1904)) ;
    nor03_2x ix1907 (.Y (nx1906), .A0 (nx4973), .A1 (nx10374), .A2 (nx11078)) ;
    dffr gen_4_cmp_mRegCmp_reg_Q_15 (.Q (gen_4_cmp_mReg_15), .QB (nx4973), .D (
         window_4__15), .CLK (start), .R (rst)) ;
    nor03_2x ix1905 (.Y (nx1904), .A0 (gen_4_cmp_mReg_15), .A1 (nx10758), .A2 (
             nx11086)) ;
    nand02 ix1929 (.Y (gen_4_cmp_BSCmp_op2_16), .A0 (nx4979), .A1 (nx4969)) ;
    nor02_2x ix4980 (.Y (nx4979), .A0 (nx1924), .A1 (nx1920)) ;
    nor03_2x ix1925 (.Y (nx1924), .A0 (gen_4_cmp_mReg_15), .A1 (nx10380), .A2 (
             nx11054)) ;
    nor03_2x ix1921 (.Y (nx1920), .A0 (nx4973), .A1 (nx11060), .A2 (nx11070)) ;
    nand02 ix1997 (.Y (gen_5_cmp_BSCmp_op2_1), .A0 (nx4987), .A1 (nx5005)) ;
    nor02_2x ix4988 (.Y (nx4987), .A0 (nx1992), .A1 (nx1988)) ;
    nor03_2x ix1993 (.Y (nx1992), .A0 (gen_5_cmp_mReg_0), .A1 (nx10364), .A2 (
             nx11090)) ;
    dffr gen_5_cmp_mRegCmp_reg_Q_0 (.Q (gen_5_cmp_mReg_0), .QB (nx4991), .D (
         window_5__0), .CLK (start), .R (rst)) ;
    inv01 ix4996 (.Y (nx4995), .A (gen_5_cmp_pMux_0)) ;
    nor03_2x ix1989 (.Y (nx1988), .A0 (nx4991), .A1 (nx11096), .A2 (nx11106)) ;
    inv02 ix5004 (.Y (nx5003), .A (gen_5_cmp_pMux_2)) ;
    nor02_2x ix5006 (.Y (nx5005), .A0 (nx1978), .A1 (nx1976)) ;
    nor03_2x ix1979 (.Y (nx1978), .A0 (nx5009), .A1 (nx10358), .A2 (nx11114)) ;
    dffr gen_5_cmp_mRegCmp_reg_Q_1 (.Q (gen_5_cmp_mReg_1), .QB (nx5009), .D (
         window_5__1), .CLK (start), .R (rst)) ;
    nor03_2x ix1977 (.Y (nx1976), .A0 (gen_5_cmp_mReg_1), .A1 (nx10760), .A2 (
             nx11122)) ;
    nor03_2x ix1937 (.Y (nx1936), .A0 (nx10364), .A1 (nx5003), .A2 (
             gen_5_cmp_pMux_0)) ;
    nand02 ix2019 (.Y (gen_5_cmp_BSCmp_op2_2), .A0 (nx5021), .A1 (nx5027)) ;
    nor02_2x ix5022 (.Y (nx5021), .A0 (nx2014), .A1 (nx2010)) ;
    nor03_2x ix2015 (.Y (nx2014), .A0 (gen_5_cmp_mReg_1), .A1 (nx10364), .A2 (
             nx11090)) ;
    nor03_2x ix2011 (.Y (nx2010), .A0 (nx5009), .A1 (nx11096), .A2 (nx11106)) ;
    nor02_2x ix5028 (.Y (nx5027), .A0 (nx2006), .A1 (nx2004)) ;
    nor03_2x ix2007 (.Y (nx2006), .A0 (nx5030), .A1 (nx10358), .A2 (nx11114)) ;
    dffr gen_5_cmp_mRegCmp_reg_Q_2 (.Q (gen_5_cmp_mReg_2), .QB (nx5030), .D (
         window_5__2), .CLK (start), .R (rst)) ;
    nor03_2x ix2005 (.Y (nx2004), .A0 (gen_5_cmp_mReg_2), .A1 (nx10760), .A2 (
             nx11122)) ;
    nand02 ix2041 (.Y (gen_5_cmp_BSCmp_op2_3), .A0 (nx5035), .A1 (nx5041)) ;
    nor02_2x ix5036 (.Y (nx5035), .A0 (nx2036), .A1 (nx2032)) ;
    nor03_2x ix2037 (.Y (nx2036), .A0 (gen_5_cmp_mReg_2), .A1 (nx10364), .A2 (
             nx11090)) ;
    nor03_2x ix2033 (.Y (nx2032), .A0 (nx5030), .A1 (nx11096), .A2 (nx11106)) ;
    nor02_2x ix5042 (.Y (nx5041), .A0 (nx2028), .A1 (nx2026)) ;
    nor03_2x ix2029 (.Y (nx2028), .A0 (nx5045), .A1 (nx10358), .A2 (nx11114)) ;
    dffr gen_5_cmp_mRegCmp_reg_Q_3 (.Q (gen_5_cmp_mReg_3), .QB (nx5045), .D (
         window_5__3), .CLK (start), .R (rst)) ;
    nor03_2x ix2027 (.Y (nx2026), .A0 (gen_5_cmp_mReg_3), .A1 (nx10760), .A2 (
             nx11122)) ;
    nand02 ix2063 (.Y (gen_5_cmp_BSCmp_op2_4), .A0 (nx5051), .A1 (nx5057)) ;
    nor02_2x ix5052 (.Y (nx5051), .A0 (nx2058), .A1 (nx2054)) ;
    nor03_2x ix2059 (.Y (nx2058), .A0 (gen_5_cmp_mReg_3), .A1 (nx10364), .A2 (
             nx11090)) ;
    nor03_2x ix2055 (.Y (nx2054), .A0 (nx5045), .A1 (nx11096), .A2 (nx11106)) ;
    nor02_2x ix5058 (.Y (nx5057), .A0 (nx2050), .A1 (nx2048)) ;
    nor03_2x ix2051 (.Y (nx2050), .A0 (nx5060), .A1 (nx10358), .A2 (nx11114)) ;
    dffr gen_5_cmp_mRegCmp_reg_Q_4 (.Q (gen_5_cmp_mReg_4), .QB (nx5060), .D (
         window_5__4), .CLK (start), .R (rst)) ;
    nor03_2x ix2049 (.Y (nx2048), .A0 (gen_5_cmp_mReg_4), .A1 (nx10760), .A2 (
             nx11122)) ;
    nand02 ix2085 (.Y (gen_5_cmp_BSCmp_op2_5), .A0 (nx5065), .A1 (nx5071)) ;
    nor02_2x ix5066 (.Y (nx5065), .A0 (nx2080), .A1 (nx2076)) ;
    nor03_2x ix2081 (.Y (nx2080), .A0 (gen_5_cmp_mReg_4), .A1 (nx10364), .A2 (
             nx11090)) ;
    nor03_2x ix2077 (.Y (nx2076), .A0 (nx5060), .A1 (nx11096), .A2 (nx11106)) ;
    nor02_2x ix5072 (.Y (nx5071), .A0 (nx2072), .A1 (nx2070)) ;
    nor03_2x ix2073 (.Y (nx2072), .A0 (nx5075), .A1 (nx10360), .A2 (nx11114)) ;
    dffr gen_5_cmp_mRegCmp_reg_Q_5 (.Q (gen_5_cmp_mReg_5), .QB (nx5075), .D (
         window_5__5), .CLK (start), .R (rst)) ;
    nor03_2x ix2071 (.Y (nx2070), .A0 (gen_5_cmp_mReg_5), .A1 (nx10760), .A2 (
             nx11122)) ;
    nand02 ix2107 (.Y (gen_5_cmp_BSCmp_op2_6), .A0 (nx5081), .A1 (nx5087)) ;
    nor02_2x ix5082 (.Y (nx5081), .A0 (nx2102), .A1 (nx2098)) ;
    nor03_2x ix2103 (.Y (nx2102), .A0 (gen_5_cmp_mReg_5), .A1 (nx10366), .A2 (
             nx11090)) ;
    nor03_2x ix2099 (.Y (nx2098), .A0 (nx5075), .A1 (nx11096), .A2 (nx11106)) ;
    nor02_2x ix5088 (.Y (nx5087), .A0 (nx2094), .A1 (nx2092)) ;
    nor03_2x ix2095 (.Y (nx2094), .A0 (nx5090), .A1 (nx10360), .A2 (nx11114)) ;
    dffr gen_5_cmp_mRegCmp_reg_Q_6 (.Q (gen_5_cmp_mReg_6), .QB (nx5090), .D (
         window_5__6), .CLK (start), .R (rst)) ;
    nor03_2x ix2093 (.Y (nx2092), .A0 (gen_5_cmp_mReg_6), .A1 (nx10760), .A2 (
             nx11122)) ;
    nand02 ix2129 (.Y (gen_5_cmp_BSCmp_op2_7), .A0 (nx5097), .A1 (nx5103)) ;
    nor02_2x ix5098 (.Y (nx5097), .A0 (nx2124), .A1 (nx2120)) ;
    nor03_2x ix2125 (.Y (nx2124), .A0 (gen_5_cmp_mReg_6), .A1 (nx10366), .A2 (
             nx11092)) ;
    nor03_2x ix2121 (.Y (nx2120), .A0 (nx5090), .A1 (nx11098), .A2 (nx11108)) ;
    nor02_2x ix5104 (.Y (nx5103), .A0 (nx2116), .A1 (nx2114)) ;
    nor03_2x ix2117 (.Y (nx2116), .A0 (nx5107), .A1 (nx10360), .A2 (nx11116)) ;
    dffr gen_5_cmp_mRegCmp_reg_Q_7 (.Q (gen_5_cmp_mReg_7), .QB (nx5107), .D (
         window_5__7), .CLK (start), .R (rst)) ;
    nor03_2x ix2115 (.Y (nx2114), .A0 (gen_5_cmp_mReg_7), .A1 (nx10760), .A2 (
             nx11124)) ;
    nand02 ix2151 (.Y (gen_5_cmp_BSCmp_op2_8), .A0 (nx5111), .A1 (nx5117)) ;
    nor02_2x ix5112 (.Y (nx5111), .A0 (nx2146), .A1 (nx2142)) ;
    nor03_2x ix2147 (.Y (nx2146), .A0 (gen_5_cmp_mReg_7), .A1 (nx10366), .A2 (
             nx11092)) ;
    nor03_2x ix2143 (.Y (nx2142), .A0 (nx5107), .A1 (nx11098), .A2 (nx11108)) ;
    nor02_2x ix5118 (.Y (nx5117), .A0 (nx2138), .A1 (nx2136)) ;
    nor03_2x ix2139 (.Y (nx2138), .A0 (nx5121), .A1 (nx10360), .A2 (nx11116)) ;
    dffr gen_5_cmp_mRegCmp_reg_Q_8 (.Q (gen_5_cmp_mReg_8), .QB (nx5121), .D (
         window_5__8), .CLK (start), .R (rst)) ;
    nor03_2x ix2137 (.Y (nx2136), .A0 (gen_5_cmp_mReg_8), .A1 (nx10762), .A2 (
             nx11124)) ;
    nand02 ix2173 (.Y (gen_5_cmp_BSCmp_op2_9), .A0 (nx5125), .A1 (nx5131)) ;
    nor02_2x ix5126 (.Y (nx5125), .A0 (nx2168), .A1 (nx2164)) ;
    nor03_2x ix2169 (.Y (nx2168), .A0 (gen_5_cmp_mReg_8), .A1 (nx10366), .A2 (
             nx11092)) ;
    nor03_2x ix2165 (.Y (nx2164), .A0 (nx5121), .A1 (nx11098), .A2 (nx11108)) ;
    nor02_2x ix5132 (.Y (nx5131), .A0 (nx2160), .A1 (nx2158)) ;
    nor03_2x ix2161 (.Y (nx2160), .A0 (nx5134), .A1 (nx10360), .A2 (nx11116)) ;
    dffr gen_5_cmp_mRegCmp_reg_Q_9 (.Q (gen_5_cmp_mReg_9), .QB (nx5134), .D (
         window_5__9), .CLK (start), .R (rst)) ;
    nor03_2x ix2159 (.Y (nx2158), .A0 (gen_5_cmp_mReg_9), .A1 (nx10762), .A2 (
             nx11124)) ;
    nand02 ix2195 (.Y (gen_5_cmp_BSCmp_op2_10), .A0 (nx5141), .A1 (nx5147)) ;
    nor02_2x ix5142 (.Y (nx5141), .A0 (nx2190), .A1 (nx2186)) ;
    nor03_2x ix2191 (.Y (nx2190), .A0 (gen_5_cmp_mReg_9), .A1 (nx10366), .A2 (
             nx11092)) ;
    nor03_2x ix2187 (.Y (nx2186), .A0 (nx5134), .A1 (nx11098), .A2 (nx11108)) ;
    nor02_2x ix5148 (.Y (nx5147), .A0 (nx2182), .A1 (nx2180)) ;
    nor03_2x ix2183 (.Y (nx2182), .A0 (nx5151), .A1 (nx10360), .A2 (nx11116)) ;
    dffr gen_5_cmp_mRegCmp_reg_Q_10 (.Q (gen_5_cmp_mReg_10), .QB (nx5151), .D (
         window_5__10), .CLK (start), .R (rst)) ;
    nor03_2x ix2181 (.Y (nx2180), .A0 (gen_5_cmp_mReg_10), .A1 (nx10762), .A2 (
             nx11124)) ;
    nand02 ix2217 (.Y (gen_5_cmp_BSCmp_op2_11), .A0 (nx5155), .A1 (nx5161)) ;
    nor02_2x ix5156 (.Y (nx5155), .A0 (nx2212), .A1 (nx2208)) ;
    nor03_2x ix2213 (.Y (nx2212), .A0 (gen_5_cmp_mReg_10), .A1 (nx10366), .A2 (
             nx11092)) ;
    nor03_2x ix2209 (.Y (nx2208), .A0 (nx5151), .A1 (nx11098), .A2 (nx11108)) ;
    nor02_2x ix5162 (.Y (nx5161), .A0 (nx2204), .A1 (nx2202)) ;
    nor03_2x ix2205 (.Y (nx2204), .A0 (nx5165), .A1 (nx10360), .A2 (nx11116)) ;
    dffr gen_5_cmp_mRegCmp_reg_Q_11 (.Q (gen_5_cmp_mReg_11), .QB (nx5165), .D (
         window_5__11), .CLK (start), .R (rst)) ;
    nor03_2x ix2203 (.Y (nx2202), .A0 (gen_5_cmp_mReg_11), .A1 (nx10762), .A2 (
             nx11124)) ;
    nand02 ix2239 (.Y (gen_5_cmp_BSCmp_op2_12), .A0 (nx5169), .A1 (nx5175)) ;
    nor02_2x ix5170 (.Y (nx5169), .A0 (nx2234), .A1 (nx2230)) ;
    nor03_2x ix2235 (.Y (nx2234), .A0 (gen_5_cmp_mReg_11), .A1 (nx10366), .A2 (
             nx11092)) ;
    nor03_2x ix2231 (.Y (nx2230), .A0 (nx5165), .A1 (nx11098), .A2 (nx11108)) ;
    nor02_2x ix5176 (.Y (nx5175), .A0 (nx2226), .A1 (nx2224)) ;
    nor03_2x ix2227 (.Y (nx2226), .A0 (nx5178), .A1 (nx10362), .A2 (nx11116)) ;
    dffr gen_5_cmp_mRegCmp_reg_Q_12 (.Q (gen_5_cmp_mReg_12), .QB (nx5178), .D (
         window_5__12), .CLK (start), .R (rst)) ;
    nor03_2x ix2225 (.Y (nx2224), .A0 (gen_5_cmp_mReg_12), .A1 (nx10762), .A2 (
             nx11124)) ;
    nand02 ix2261 (.Y (gen_5_cmp_BSCmp_op2_13), .A0 (nx5185), .A1 (nx5191)) ;
    nor02_2x ix5186 (.Y (nx5185), .A0 (nx2256), .A1 (nx2252)) ;
    nor03_2x ix2257 (.Y (nx2256), .A0 (gen_5_cmp_mReg_12), .A1 (nx10368), .A2 (
             nx11094)) ;
    nor03_2x ix2253 (.Y (nx2252), .A0 (nx5178), .A1 (nx11098), .A2 (nx11110)) ;
    nor02_2x ix5192 (.Y (nx5191), .A0 (nx2248), .A1 (nx2246)) ;
    nor03_2x ix2249 (.Y (nx2248), .A0 (nx5195), .A1 (nx10362), .A2 (nx11118)) ;
    dffr gen_5_cmp_mRegCmp_reg_Q_13 (.Q (gen_5_cmp_mReg_13), .QB (nx5195), .D (
         window_5__13), .CLK (start), .R (rst)) ;
    nor03_2x ix2247 (.Y (nx2246), .A0 (gen_5_cmp_mReg_13), .A1 (nx10762), .A2 (
             nx11126)) ;
    nand02 ix2283 (.Y (gen_5_cmp_BSCmp_op2_14), .A0 (nx5199), .A1 (nx5205)) ;
    nor02_2x ix5200 (.Y (nx5199), .A0 (nx2278), .A1 (nx2274)) ;
    nor03_2x ix2279 (.Y (nx2278), .A0 (gen_5_cmp_mReg_13), .A1 (nx10368), .A2 (
             nx11094)) ;
    nor03_2x ix2275 (.Y (nx2274), .A0 (nx5195), .A1 (nx11100), .A2 (nx11110)) ;
    nor02_2x ix5206 (.Y (nx5205), .A0 (nx2270), .A1 (nx2268)) ;
    nor03_2x ix2271 (.Y (nx2270), .A0 (nx5209), .A1 (nx10362), .A2 (nx11118)) ;
    dffr gen_5_cmp_mRegCmp_reg_Q_14 (.Q (gen_5_cmp_mReg_14), .QB (nx5209), .D (
         window_5__14), .CLK (start), .R (rst)) ;
    nor03_2x ix2269 (.Y (nx2268), .A0 (gen_5_cmp_mReg_14), .A1 (nx10762), .A2 (
             nx11126)) ;
    nand02 ix2305 (.Y (gen_5_cmp_BSCmp_op2_15), .A0 (nx5213), .A1 (nx5219)) ;
    nor02_2x ix5214 (.Y (nx5213), .A0 (nx2300), .A1 (nx2296)) ;
    nor03_2x ix2301 (.Y (nx2300), .A0 (gen_5_cmp_mReg_14), .A1 (nx10368), .A2 (
             nx11094)) ;
    nor03_2x ix2297 (.Y (nx2296), .A0 (nx5209), .A1 (nx11100), .A2 (nx11110)) ;
    nor02_2x ix5220 (.Y (nx5219), .A0 (nx2292), .A1 (nx2290)) ;
    nor03_2x ix2293 (.Y (nx2292), .A0 (nx5222), .A1 (nx10362), .A2 (nx11118)) ;
    dffr gen_5_cmp_mRegCmp_reg_Q_15 (.Q (gen_5_cmp_mReg_15), .QB (nx5222), .D (
         window_5__15), .CLK (start), .R (rst)) ;
    nor03_2x ix2291 (.Y (nx2290), .A0 (gen_5_cmp_mReg_15), .A1 (nx10764), .A2 (
             nx11126)) ;
    nand02 ix2315 (.Y (gen_5_cmp_BSCmp_op2_16), .A0 (nx5229), .A1 (nx5219)) ;
    nor02_2x ix5230 (.Y (nx5229), .A0 (nx2310), .A1 (nx2306)) ;
    nor03_2x ix2311 (.Y (nx2310), .A0 (gen_5_cmp_mReg_15), .A1 (nx10368), .A2 (
             nx11094)) ;
    nor03_2x ix2307 (.Y (nx2306), .A0 (nx5222), .A1 (nx11100), .A2 (nx11110)) ;
    nand02 ix2383 (.Y (gen_6_cmp_BSCmp_op2_1), .A0 (nx5235), .A1 (nx5255)) ;
    nor02_2x ix5236 (.Y (nx5235), .A0 (nx2378), .A1 (nx2374)) ;
    nor03_2x ix2379 (.Y (nx2378), .A0 (gen_6_cmp_mReg_0), .A1 (nx10352), .A2 (
             nx11130)) ;
    dffr gen_6_cmp_mRegCmp_reg_Q_0 (.Q (gen_6_cmp_mReg_0), .QB (nx5241), .D (
         window_6__0), .CLK (start), .R (rst)) ;
    inv01 ix5246 (.Y (nx5244), .A (gen_6_cmp_pMux_0)) ;
    nor03_2x ix2375 (.Y (nx2374), .A0 (nx5241), .A1 (nx11136), .A2 (nx11146)) ;
    inv02 ix5254 (.Y (nx5253), .A (gen_6_cmp_pMux_2)) ;
    nor02_2x ix5256 (.Y (nx5255), .A0 (nx2364), .A1 (nx2362)) ;
    nor03_2x ix2365 (.Y (nx2364), .A0 (nx5259), .A1 (nx10346), .A2 (nx11154)) ;
    dffr gen_6_cmp_mRegCmp_reg_Q_1 (.Q (gen_6_cmp_mReg_1), .QB (nx5259), .D (
         window_6__1), .CLK (start), .R (rst)) ;
    nor03_2x ix2363 (.Y (nx2362), .A0 (gen_6_cmp_mReg_1), .A1 (nx10766), .A2 (
             nx11162)) ;
    nor03_2x ix2323 (.Y (nx2322), .A0 (nx10352), .A1 (nx5253), .A2 (
             gen_6_cmp_pMux_0)) ;
    nand02 ix2405 (.Y (gen_6_cmp_BSCmp_op2_2), .A0 (nx5269), .A1 (nx5275)) ;
    nor02_2x ix5270 (.Y (nx5269), .A0 (nx2400), .A1 (nx2396)) ;
    nor03_2x ix2401 (.Y (nx2400), .A0 (gen_6_cmp_mReg_1), .A1 (nx10352), .A2 (
             nx11130)) ;
    nor03_2x ix2397 (.Y (nx2396), .A0 (nx5259), .A1 (nx11136), .A2 (nx11146)) ;
    nor02_2x ix5276 (.Y (nx5275), .A0 (nx2392), .A1 (nx2390)) ;
    nor03_2x ix2393 (.Y (nx2392), .A0 (nx5279), .A1 (nx10346), .A2 (nx11154)) ;
    dffr gen_6_cmp_mRegCmp_reg_Q_2 (.Q (gen_6_cmp_mReg_2), .QB (nx5279), .D (
         window_6__2), .CLK (start), .R (rst)) ;
    nor03_2x ix2391 (.Y (nx2390), .A0 (gen_6_cmp_mReg_2), .A1 (nx10766), .A2 (
             nx11162)) ;
    nand02 ix2427 (.Y (gen_6_cmp_BSCmp_op2_3), .A0 (nx5285), .A1 (nx5289)) ;
    nor02_2x ix5286 (.Y (nx5285), .A0 (nx2422), .A1 (nx2418)) ;
    nor03_2x ix2423 (.Y (nx2422), .A0 (gen_6_cmp_mReg_2), .A1 (nx10352), .A2 (
             nx11130)) ;
    nor03_2x ix2419 (.Y (nx2418), .A0 (nx5279), .A1 (nx11136), .A2 (nx11146)) ;
    nor02_2x ix5290 (.Y (nx5289), .A0 (nx2414), .A1 (nx2412)) ;
    nor03_2x ix2415 (.Y (nx2414), .A0 (nx5293), .A1 (nx10346), .A2 (nx11154)) ;
    dffr gen_6_cmp_mRegCmp_reg_Q_3 (.Q (gen_6_cmp_mReg_3), .QB (nx5293), .D (
         window_6__3), .CLK (start), .R (rst)) ;
    nor03_2x ix2413 (.Y (nx2412), .A0 (gen_6_cmp_mReg_3), .A1 (nx10766), .A2 (
             nx11162)) ;
    nand02 ix2449 (.Y (gen_6_cmp_BSCmp_op2_4), .A0 (nx5299), .A1 (nx5305)) ;
    nor02_2x ix5300 (.Y (nx5299), .A0 (nx2444), .A1 (nx2440)) ;
    nor03_2x ix2445 (.Y (nx2444), .A0 (gen_6_cmp_mReg_3), .A1 (nx10352), .A2 (
             nx11130)) ;
    nor03_2x ix2441 (.Y (nx2440), .A0 (nx5293), .A1 (nx11136), .A2 (nx11146)) ;
    nor02_2x ix5306 (.Y (nx5305), .A0 (nx2436), .A1 (nx2434)) ;
    nor03_2x ix2437 (.Y (nx2436), .A0 (nx5308), .A1 (nx10346), .A2 (nx11154)) ;
    dffr gen_6_cmp_mRegCmp_reg_Q_4 (.Q (gen_6_cmp_mReg_4), .QB (nx5308), .D (
         window_6__4), .CLK (start), .R (rst)) ;
    nor03_2x ix2435 (.Y (nx2434), .A0 (gen_6_cmp_mReg_4), .A1 (nx10766), .A2 (
             nx11162)) ;
    nand02 ix2471 (.Y (gen_6_cmp_BSCmp_op2_5), .A0 (nx5313), .A1 (nx5319)) ;
    nor02_2x ix5314 (.Y (nx5313), .A0 (nx2466), .A1 (nx2462)) ;
    nor03_2x ix2467 (.Y (nx2466), .A0 (gen_6_cmp_mReg_4), .A1 (nx10352), .A2 (
             nx11130)) ;
    nor03_2x ix2463 (.Y (nx2462), .A0 (nx5308), .A1 (nx11136), .A2 (nx11146)) ;
    nor02_2x ix5320 (.Y (nx5319), .A0 (nx2458), .A1 (nx2456)) ;
    nor03_2x ix2459 (.Y (nx2458), .A0 (nx5323), .A1 (nx10348), .A2 (nx11154)) ;
    dffr gen_6_cmp_mRegCmp_reg_Q_5 (.Q (gen_6_cmp_mReg_5), .QB (nx5323), .D (
         window_6__5), .CLK (start), .R (rst)) ;
    nor03_2x ix2457 (.Y (nx2456), .A0 (gen_6_cmp_mReg_5), .A1 (nx10766), .A2 (
             nx11162)) ;
    nand02 ix2493 (.Y (gen_6_cmp_BSCmp_op2_6), .A0 (nx5329), .A1 (nx5333)) ;
    nor02_2x ix5330 (.Y (nx5329), .A0 (nx2488), .A1 (nx2484)) ;
    nor03_2x ix2489 (.Y (nx2488), .A0 (gen_6_cmp_mReg_5), .A1 (nx10354), .A2 (
             nx11130)) ;
    nor03_2x ix2485 (.Y (nx2484), .A0 (nx5323), .A1 (nx11136), .A2 (nx11146)) ;
    nor02_2x ix5334 (.Y (nx5333), .A0 (nx2480), .A1 (nx2478)) ;
    nor03_2x ix2481 (.Y (nx2480), .A0 (nx5337), .A1 (nx10348), .A2 (nx11154)) ;
    dffr gen_6_cmp_mRegCmp_reg_Q_6 (.Q (gen_6_cmp_mReg_6), .QB (nx5337), .D (
         window_6__6), .CLK (start), .R (rst)) ;
    nor03_2x ix2479 (.Y (nx2478), .A0 (gen_6_cmp_mReg_6), .A1 (nx10766), .A2 (
             nx11162)) ;
    nand02 ix2515 (.Y (gen_6_cmp_BSCmp_op2_7), .A0 (nx5343), .A1 (nx5349)) ;
    nor02_2x ix5344 (.Y (nx5343), .A0 (nx2510), .A1 (nx2506)) ;
    nor03_2x ix2511 (.Y (nx2510), .A0 (gen_6_cmp_mReg_6), .A1 (nx10354), .A2 (
             nx11132)) ;
    nor03_2x ix2507 (.Y (nx2506), .A0 (nx5337), .A1 (nx11138), .A2 (nx11148)) ;
    nor02_2x ix5350 (.Y (nx5349), .A0 (nx2502), .A1 (nx2500)) ;
    nor03_2x ix2503 (.Y (nx2502), .A0 (nx5352), .A1 (nx10348), .A2 (nx11156)) ;
    dffr gen_6_cmp_mRegCmp_reg_Q_7 (.Q (gen_6_cmp_mReg_7), .QB (nx5352), .D (
         window_6__7), .CLK (start), .R (rst)) ;
    nor03_2x ix2501 (.Y (nx2500), .A0 (gen_6_cmp_mReg_7), .A1 (nx10766), .A2 (
             nx11164)) ;
    nand02 ix2537 (.Y (gen_6_cmp_BSCmp_op2_8), .A0 (nx5357), .A1 (nx5363)) ;
    nor02_2x ix5358 (.Y (nx5357), .A0 (nx2532), .A1 (nx2528)) ;
    nor03_2x ix2533 (.Y (nx2532), .A0 (gen_6_cmp_mReg_7), .A1 (nx10354), .A2 (
             nx11132)) ;
    nor03_2x ix2529 (.Y (nx2528), .A0 (nx5352), .A1 (nx11138), .A2 (nx11148)) ;
    nor02_2x ix5364 (.Y (nx5363), .A0 (nx2524), .A1 (nx2522)) ;
    nor03_2x ix2525 (.Y (nx2524), .A0 (nx5367), .A1 (nx10348), .A2 (nx11156)) ;
    dffr gen_6_cmp_mRegCmp_reg_Q_8 (.Q (gen_6_cmp_mReg_8), .QB (nx5367), .D (
         window_6__8), .CLK (start), .R (rst)) ;
    nor03_2x ix2523 (.Y (nx2522), .A0 (gen_6_cmp_mReg_8), .A1 (nx10768), .A2 (
             nx11164)) ;
    nand02 ix2559 (.Y (gen_6_cmp_BSCmp_op2_9), .A0 (nx5373), .A1 (nx5377)) ;
    nor02_2x ix5374 (.Y (nx5373), .A0 (nx2554), .A1 (nx2550)) ;
    nor03_2x ix2555 (.Y (nx2554), .A0 (gen_6_cmp_mReg_8), .A1 (nx10354), .A2 (
             nx11132)) ;
    nor03_2x ix2551 (.Y (nx2550), .A0 (nx5367), .A1 (nx11138), .A2 (nx11148)) ;
    nor02_2x ix5378 (.Y (nx5377), .A0 (nx2546), .A1 (nx2544)) ;
    nor03_2x ix2547 (.Y (nx2546), .A0 (nx5381), .A1 (nx10348), .A2 (nx11156)) ;
    dffr gen_6_cmp_mRegCmp_reg_Q_9 (.Q (gen_6_cmp_mReg_9), .QB (nx5381), .D (
         window_6__9), .CLK (start), .R (rst)) ;
    nor03_2x ix2545 (.Y (nx2544), .A0 (gen_6_cmp_mReg_9), .A1 (nx10768), .A2 (
             nx11164)) ;
    nand02 ix2581 (.Y (gen_6_cmp_BSCmp_op2_10), .A0 (nx5387), .A1 (nx5393)) ;
    nor02_2x ix5388 (.Y (nx5387), .A0 (nx2576), .A1 (nx2572)) ;
    nor03_2x ix2577 (.Y (nx2576), .A0 (gen_6_cmp_mReg_9), .A1 (nx10354), .A2 (
             nx11132)) ;
    nor03_2x ix2573 (.Y (nx2572), .A0 (nx5381), .A1 (nx11138), .A2 (nx11148)) ;
    nor02_2x ix5394 (.Y (nx5393), .A0 (nx2568), .A1 (nx2566)) ;
    nor03_2x ix2569 (.Y (nx2568), .A0 (nx5397), .A1 (nx10348), .A2 (nx11156)) ;
    dffr gen_6_cmp_mRegCmp_reg_Q_10 (.Q (gen_6_cmp_mReg_10), .QB (nx5397), .D (
         window_6__10), .CLK (start), .R (rst)) ;
    nor03_2x ix2567 (.Y (nx2566), .A0 (gen_6_cmp_mReg_10), .A1 (nx10768), .A2 (
             nx11164)) ;
    nand02 ix2603 (.Y (gen_6_cmp_BSCmp_op2_11), .A0 (nx5403), .A1 (nx5409)) ;
    nor02_2x ix5404 (.Y (nx5403), .A0 (nx2598), .A1 (nx2594)) ;
    nor03_2x ix2599 (.Y (nx2598), .A0 (gen_6_cmp_mReg_10), .A1 (nx10354), .A2 (
             nx11132)) ;
    nor03_2x ix2595 (.Y (nx2594), .A0 (nx5397), .A1 (nx11138), .A2 (nx11148)) ;
    nor02_2x ix5410 (.Y (nx5409), .A0 (nx2590), .A1 (nx2588)) ;
    nor03_2x ix2591 (.Y (nx2590), .A0 (nx5413), .A1 (nx10348), .A2 (nx11156)) ;
    dffr gen_6_cmp_mRegCmp_reg_Q_11 (.Q (gen_6_cmp_mReg_11), .QB (nx5413), .D (
         window_6__11), .CLK (start), .R (rst)) ;
    nor03_2x ix2589 (.Y (nx2588), .A0 (gen_6_cmp_mReg_11), .A1 (nx10768), .A2 (
             nx11164)) ;
    nand02 ix2625 (.Y (gen_6_cmp_BSCmp_op2_12), .A0 (nx5417), .A1 (nx5421)) ;
    nor02_2x ix5418 (.Y (nx5417), .A0 (nx2620), .A1 (nx2616)) ;
    nor03_2x ix2621 (.Y (nx2620), .A0 (gen_6_cmp_mReg_11), .A1 (nx10354), .A2 (
             nx11132)) ;
    nor03_2x ix2617 (.Y (nx2616), .A0 (nx5413), .A1 (nx11138), .A2 (nx11148)) ;
    nor02_2x ix5422 (.Y (nx5421), .A0 (nx2612), .A1 (nx2610)) ;
    nor03_2x ix2613 (.Y (nx2612), .A0 (nx5425), .A1 (nx10350), .A2 (nx11156)) ;
    dffr gen_6_cmp_mRegCmp_reg_Q_12 (.Q (gen_6_cmp_mReg_12), .QB (nx5425), .D (
         window_6__12), .CLK (start), .R (rst)) ;
    nor03_2x ix2611 (.Y (nx2610), .A0 (gen_6_cmp_mReg_12), .A1 (nx10768), .A2 (
             nx11164)) ;
    nand02 ix2647 (.Y (gen_6_cmp_BSCmp_op2_13), .A0 (nx5431), .A1 (nx5437)) ;
    nor02_2x ix5432 (.Y (nx5431), .A0 (nx2642), .A1 (nx2638)) ;
    nor03_2x ix2643 (.Y (nx2642), .A0 (gen_6_cmp_mReg_12), .A1 (nx10356), .A2 (
             nx11134)) ;
    nor03_2x ix2639 (.Y (nx2638), .A0 (nx5425), .A1 (nx11138), .A2 (nx11150)) ;
    nor02_2x ix5438 (.Y (nx5437), .A0 (nx2634), .A1 (nx2632)) ;
    nor03_2x ix2635 (.Y (nx2634), .A0 (nx5441), .A1 (nx10350), .A2 (nx11158)) ;
    dffr gen_6_cmp_mRegCmp_reg_Q_13 (.Q (gen_6_cmp_mReg_13), .QB (nx5441), .D (
         window_6__13), .CLK (start), .R (rst)) ;
    nor03_2x ix2633 (.Y (nx2632), .A0 (gen_6_cmp_mReg_13), .A1 (nx10768), .A2 (
             nx11166)) ;
    nand02 ix2669 (.Y (gen_6_cmp_BSCmp_op2_14), .A0 (nx5446), .A1 (nx5451)) ;
    nor02_2x ix5447 (.Y (nx5446), .A0 (nx2664), .A1 (nx2660)) ;
    nor03_2x ix2665 (.Y (nx2664), .A0 (gen_6_cmp_mReg_13), .A1 (nx10356), .A2 (
             nx11134)) ;
    nor03_2x ix2661 (.Y (nx2660), .A0 (nx5441), .A1 (nx11140), .A2 (nx11150)) ;
    nor02_2x ix5452 (.Y (nx5451), .A0 (nx2656), .A1 (nx2654)) ;
    nor03_2x ix2657 (.Y (nx2656), .A0 (nx5455), .A1 (nx10350), .A2 (nx11158)) ;
    dffr gen_6_cmp_mRegCmp_reg_Q_14 (.Q (gen_6_cmp_mReg_14), .QB (nx5455), .D (
         window_6__14), .CLK (start), .R (rst)) ;
    nor03_2x ix2655 (.Y (nx2654), .A0 (gen_6_cmp_mReg_14), .A1 (nx10768), .A2 (
             nx11166)) ;
    nand02 ix2691 (.Y (gen_6_cmp_BSCmp_op2_15), .A0 (nx5459), .A1 (nx5465)) ;
    nor02_2x ix5460 (.Y (nx5459), .A0 (nx2686), .A1 (nx2682)) ;
    nor03_2x ix2687 (.Y (nx2686), .A0 (gen_6_cmp_mReg_14), .A1 (nx10356), .A2 (
             nx11134)) ;
    nor03_2x ix2683 (.Y (nx2682), .A0 (nx5455), .A1 (nx11140), .A2 (nx11150)) ;
    nor02_2x ix5466 (.Y (nx5465), .A0 (nx2678), .A1 (nx2676)) ;
    nor03_2x ix2679 (.Y (nx2678), .A0 (nx5469), .A1 (nx10350), .A2 (nx11158)) ;
    dffr gen_6_cmp_mRegCmp_reg_Q_15 (.Q (gen_6_cmp_mReg_15), .QB (nx5469), .D (
         window_6__15), .CLK (start), .R (rst)) ;
    nor03_2x ix2677 (.Y (nx2676), .A0 (gen_6_cmp_mReg_15), .A1 (nx10770), .A2 (
             nx11166)) ;
    nand02 ix2701 (.Y (gen_6_cmp_BSCmp_op2_16), .A0 (nx5474), .A1 (nx5465)) ;
    nor02_2x ix5475 (.Y (nx5474), .A0 (nx2696), .A1 (nx2692)) ;
    nor03_2x ix2697 (.Y (nx2696), .A0 (gen_6_cmp_mReg_15), .A1 (nx10356), .A2 (
             nx11134)) ;
    nor03_2x ix2693 (.Y (nx2692), .A0 (nx5469), .A1 (nx11140), .A2 (nx11150)) ;
    nand02 ix2769 (.Y (gen_7_cmp_BSCmp_op2_1), .A0 (nx5481), .A1 (nx5501)) ;
    nor02_2x ix5482 (.Y (nx5481), .A0 (nx2764), .A1 (nx2760)) ;
    nor03_2x ix2765 (.Y (nx2764), .A0 (gen_7_cmp_mReg_0), .A1 (nx10340), .A2 (
             nx11170)) ;
    dffr gen_7_cmp_mRegCmp_reg_Q_0 (.Q (gen_7_cmp_mReg_0), .QB (nx5487), .D (
         window_7__0), .CLK (start), .R (rst)) ;
    inv01 ix5492 (.Y (nx5491), .A (gen_7_cmp_pMux_0)) ;
    nor03_2x ix2761 (.Y (nx2760), .A0 (nx5487), .A1 (nx11176), .A2 (nx11186)) ;
    inv02 ix5500 (.Y (nx5499), .A (gen_7_cmp_pMux_2)) ;
    nor02_2x ix5502 (.Y (nx5501), .A0 (nx2750), .A1 (nx2748)) ;
    nor03_2x ix2751 (.Y (nx2750), .A0 (nx5505), .A1 (nx10334), .A2 (nx11194)) ;
    dffr gen_7_cmp_mRegCmp_reg_Q_1 (.Q (gen_7_cmp_mReg_1), .QB (nx5505), .D (
         window_7__1), .CLK (start), .R (rst)) ;
    nor03_2x ix2749 (.Y (nx2748), .A0 (gen_7_cmp_mReg_1), .A1 (nx10772), .A2 (
             nx11202)) ;
    nor03_2x ix2709 (.Y (nx2708), .A0 (nx10340), .A1 (nx5499), .A2 (
             gen_7_cmp_pMux_0)) ;
    nand02 ix2791 (.Y (gen_7_cmp_BSCmp_op2_2), .A0 (nx5515), .A1 (nx5519)) ;
    nor02_2x ix5516 (.Y (nx5515), .A0 (nx2786), .A1 (nx2782)) ;
    nor03_2x ix2787 (.Y (nx2786), .A0 (gen_7_cmp_mReg_1), .A1 (nx10340), .A2 (
             nx11170)) ;
    nor03_2x ix2783 (.Y (nx2782), .A0 (nx5505), .A1 (nx11176), .A2 (nx11186)) ;
    nor02_2x ix5520 (.Y (nx5519), .A0 (nx2778), .A1 (nx2776)) ;
    nor03_2x ix2779 (.Y (nx2778), .A0 (nx5523), .A1 (nx10334), .A2 (nx11194)) ;
    dffr gen_7_cmp_mRegCmp_reg_Q_2 (.Q (gen_7_cmp_mReg_2), .QB (nx5523), .D (
         window_7__2), .CLK (start), .R (rst)) ;
    nor03_2x ix2777 (.Y (nx2776), .A0 (gen_7_cmp_mReg_2), .A1 (nx10772), .A2 (
             nx11202)) ;
    nand02 ix2813 (.Y (gen_7_cmp_BSCmp_op2_3), .A0 (nx5529), .A1 (nx5533)) ;
    nor02_2x ix5530 (.Y (nx5529), .A0 (nx2808), .A1 (nx2804)) ;
    nor03_2x ix2809 (.Y (nx2808), .A0 (gen_7_cmp_mReg_2), .A1 (nx10340), .A2 (
             nx11170)) ;
    nor03_2x ix2805 (.Y (nx2804), .A0 (nx5523), .A1 (nx11176), .A2 (nx11186)) ;
    nor02_2x ix5534 (.Y (nx5533), .A0 (nx2800), .A1 (nx2798)) ;
    nor03_2x ix2801 (.Y (nx2800), .A0 (nx5537), .A1 (nx10334), .A2 (nx11194)) ;
    dffr gen_7_cmp_mRegCmp_reg_Q_3 (.Q (gen_7_cmp_mReg_3), .QB (nx5537), .D (
         window_7__3), .CLK (start), .R (rst)) ;
    nor03_2x ix2799 (.Y (nx2798), .A0 (gen_7_cmp_mReg_3), .A1 (nx10772), .A2 (
             nx11202)) ;
    nand02 ix2835 (.Y (gen_7_cmp_BSCmp_op2_4), .A0 (nx5541), .A1 (nx5547)) ;
    nor02_2x ix5542 (.Y (nx5541), .A0 (nx2830), .A1 (nx2826)) ;
    nor03_2x ix2831 (.Y (nx2830), .A0 (gen_7_cmp_mReg_3), .A1 (nx10340), .A2 (
             nx11170)) ;
    nor03_2x ix2827 (.Y (nx2826), .A0 (nx5537), .A1 (nx11176), .A2 (nx11186)) ;
    nor02_2x ix5548 (.Y (nx5547), .A0 (nx2822), .A1 (nx2820)) ;
    nor03_2x ix2823 (.Y (nx2822), .A0 (nx5551), .A1 (nx10334), .A2 (nx11194)) ;
    dffr gen_7_cmp_mRegCmp_reg_Q_4 (.Q (gen_7_cmp_mReg_4), .QB (nx5551), .D (
         window_7__4), .CLK (start), .R (rst)) ;
    nor03_2x ix2821 (.Y (nx2820), .A0 (gen_7_cmp_mReg_4), .A1 (nx10772), .A2 (
             nx11202)) ;
    nand02 ix2857 (.Y (gen_7_cmp_BSCmp_op2_5), .A0 (nx5555), .A1 (nx5561)) ;
    nor02_2x ix5556 (.Y (nx5555), .A0 (nx2852), .A1 (nx2848)) ;
    nor03_2x ix2853 (.Y (nx2852), .A0 (gen_7_cmp_mReg_4), .A1 (nx10340), .A2 (
             nx11170)) ;
    nor03_2x ix2849 (.Y (nx2848), .A0 (nx5551), .A1 (nx11176), .A2 (nx11186)) ;
    nor02_2x ix5562 (.Y (nx5561), .A0 (nx2844), .A1 (nx2842)) ;
    nor03_2x ix2845 (.Y (nx2844), .A0 (nx5564), .A1 (nx10336), .A2 (nx11194)) ;
    dffr gen_7_cmp_mRegCmp_reg_Q_5 (.Q (gen_7_cmp_mReg_5), .QB (nx5564), .D (
         window_7__5), .CLK (start), .R (rst)) ;
    nor03_2x ix2843 (.Y (nx2842), .A0 (gen_7_cmp_mReg_5), .A1 (nx10772), .A2 (
             nx11202)) ;
    nand02 ix2879 (.Y (gen_7_cmp_BSCmp_op2_6), .A0 (nx5571), .A1 (nx5577)) ;
    nor02_2x ix5572 (.Y (nx5571), .A0 (nx2874), .A1 (nx2870)) ;
    nor03_2x ix2875 (.Y (nx2874), .A0 (gen_7_cmp_mReg_5), .A1 (nx10342), .A2 (
             nx11170)) ;
    nor03_2x ix2871 (.Y (nx2870), .A0 (nx5564), .A1 (nx11176), .A2 (nx11186)) ;
    nor02_2x ix5578 (.Y (nx5577), .A0 (nx2866), .A1 (nx2864)) ;
    nor03_2x ix2867 (.Y (nx2866), .A0 (nx5581), .A1 (nx10336), .A2 (nx11194)) ;
    dffr gen_7_cmp_mRegCmp_reg_Q_6 (.Q (gen_7_cmp_mReg_6), .QB (nx5581), .D (
         window_7__6), .CLK (start), .R (rst)) ;
    nor03_2x ix2865 (.Y (nx2864), .A0 (gen_7_cmp_mReg_6), .A1 (nx10772), .A2 (
             nx11202)) ;
    nand02 ix2901 (.Y (gen_7_cmp_BSCmp_op2_7), .A0 (nx5585), .A1 (nx5591)) ;
    nor02_2x ix5586 (.Y (nx5585), .A0 (nx2896), .A1 (nx2892)) ;
    nor03_2x ix2897 (.Y (nx2896), .A0 (gen_7_cmp_mReg_6), .A1 (nx10342), .A2 (
             nx11172)) ;
    nor03_2x ix2893 (.Y (nx2892), .A0 (nx5581), .A1 (nx11178), .A2 (nx11188)) ;
    nor02_2x ix5592 (.Y (nx5591), .A0 (nx2888), .A1 (nx2886)) ;
    nor03_2x ix2889 (.Y (nx2888), .A0 (nx5595), .A1 (nx10336), .A2 (nx11196)) ;
    dffr gen_7_cmp_mRegCmp_reg_Q_7 (.Q (gen_7_cmp_mReg_7), .QB (nx5595), .D (
         window_7__7), .CLK (start), .R (rst)) ;
    nor03_2x ix2887 (.Y (nx2886), .A0 (gen_7_cmp_mReg_7), .A1 (nx10772), .A2 (
             nx11204)) ;
    nand02 ix2923 (.Y (gen_7_cmp_BSCmp_op2_8), .A0 (nx5599), .A1 (nx5605)) ;
    nor02_2x ix5600 (.Y (nx5599), .A0 (nx2918), .A1 (nx2914)) ;
    nor03_2x ix2919 (.Y (nx2918), .A0 (gen_7_cmp_mReg_7), .A1 (nx10342), .A2 (
             nx11172)) ;
    nor03_2x ix2915 (.Y (nx2914), .A0 (nx5595), .A1 (nx11178), .A2 (nx11188)) ;
    nor02_2x ix5606 (.Y (nx5605), .A0 (nx2910), .A1 (nx2908)) ;
    nor03_2x ix2911 (.Y (nx2910), .A0 (nx5608), .A1 (nx10336), .A2 (nx11196)) ;
    dffr gen_7_cmp_mRegCmp_reg_Q_8 (.Q (gen_7_cmp_mReg_8), .QB (nx5608), .D (
         window_7__8), .CLK (start), .R (rst)) ;
    nor03_2x ix2909 (.Y (nx2908), .A0 (gen_7_cmp_mReg_8), .A1 (nx10774), .A2 (
             nx11204)) ;
    nand02 ix2945 (.Y (gen_7_cmp_BSCmp_op2_9), .A0 (nx5615), .A1 (nx5621)) ;
    nor02_2x ix5616 (.Y (nx5615), .A0 (nx2940), .A1 (nx2936)) ;
    nor03_2x ix2941 (.Y (nx2940), .A0 (gen_7_cmp_mReg_8), .A1 (nx10342), .A2 (
             nx11172)) ;
    nor03_2x ix2937 (.Y (nx2936), .A0 (nx5608), .A1 (nx11178), .A2 (nx11188)) ;
    nor02_2x ix5622 (.Y (nx5621), .A0 (nx2932), .A1 (nx2930)) ;
    nor03_2x ix2933 (.Y (nx2932), .A0 (nx5625), .A1 (nx10336), .A2 (nx11196)) ;
    dffr gen_7_cmp_mRegCmp_reg_Q_9 (.Q (gen_7_cmp_mReg_9), .QB (nx5625), .D (
         window_7__9), .CLK (start), .R (rst)) ;
    nor03_2x ix2931 (.Y (nx2930), .A0 (gen_7_cmp_mReg_9), .A1 (nx10774), .A2 (
             nx11204)) ;
    nand02 ix2967 (.Y (gen_7_cmp_BSCmp_op2_10), .A0 (nx5629), .A1 (nx5635)) ;
    nor02_2x ix5630 (.Y (nx5629), .A0 (nx2962), .A1 (nx2958)) ;
    nor03_2x ix2963 (.Y (nx2962), .A0 (gen_7_cmp_mReg_9), .A1 (nx10342), .A2 (
             nx11172)) ;
    nor03_2x ix2959 (.Y (nx2958), .A0 (nx5625), .A1 (nx11178), .A2 (nx11188)) ;
    nor02_2x ix5636 (.Y (nx5635), .A0 (nx2954), .A1 (nx2952)) ;
    nor03_2x ix2955 (.Y (nx2954), .A0 (nx5639), .A1 (nx10336), .A2 (nx11196)) ;
    dffr gen_7_cmp_mRegCmp_reg_Q_10 (.Q (gen_7_cmp_mReg_10), .QB (nx5639), .D (
         window_7__10), .CLK (start), .R (rst)) ;
    nor03_2x ix2953 (.Y (nx2952), .A0 (gen_7_cmp_mReg_10), .A1 (nx10774), .A2 (
             nx11204)) ;
    nand02 ix2989 (.Y (gen_7_cmp_BSCmp_op2_11), .A0 (nx5643), .A1 (nx5649)) ;
    nor02_2x ix5644 (.Y (nx5643), .A0 (nx2984), .A1 (nx2980)) ;
    nor03_2x ix2985 (.Y (nx2984), .A0 (gen_7_cmp_mReg_10), .A1 (nx10342), .A2 (
             nx11172)) ;
    nor03_2x ix2981 (.Y (nx2980), .A0 (nx5639), .A1 (nx11178), .A2 (nx11188)) ;
    nor02_2x ix5650 (.Y (nx5649), .A0 (nx2976), .A1 (nx2974)) ;
    nor03_2x ix2977 (.Y (nx2976), .A0 (nx5652), .A1 (nx10336), .A2 (nx11196)) ;
    dffr gen_7_cmp_mRegCmp_reg_Q_11 (.Q (gen_7_cmp_mReg_11), .QB (nx5652), .D (
         window_7__11), .CLK (start), .R (rst)) ;
    nor03_2x ix2975 (.Y (nx2974), .A0 (gen_7_cmp_mReg_11), .A1 (nx10774), .A2 (
             nx11204)) ;
    nand02 ix3011 (.Y (gen_7_cmp_BSCmp_op2_12), .A0 (nx5659), .A1 (nx5665)) ;
    nor02_2x ix5660 (.Y (nx5659), .A0 (nx3006), .A1 (nx3002)) ;
    nor03_2x ix3007 (.Y (nx3006), .A0 (gen_7_cmp_mReg_11), .A1 (nx10342), .A2 (
             nx11172)) ;
    nor03_2x ix3003 (.Y (nx3002), .A0 (nx5652), .A1 (nx11178), .A2 (nx11188)) ;
    nor02_2x ix5666 (.Y (nx5665), .A0 (nx2998), .A1 (nx2996)) ;
    nor03_2x ix2999 (.Y (nx2998), .A0 (nx5669), .A1 (nx10338), .A2 (nx11196)) ;
    dffr gen_7_cmp_mRegCmp_reg_Q_12 (.Q (gen_7_cmp_mReg_12), .QB (nx5669), .D (
         window_7__12), .CLK (start), .R (rst)) ;
    nor03_2x ix2997 (.Y (nx2996), .A0 (gen_7_cmp_mReg_12), .A1 (nx10774), .A2 (
             nx11204)) ;
    nand02 ix3033 (.Y (gen_7_cmp_BSCmp_op2_13), .A0 (nx5673), .A1 (nx5679)) ;
    nor02_2x ix5674 (.Y (nx5673), .A0 (nx3028), .A1 (nx3024)) ;
    nor03_2x ix3029 (.Y (nx3028), .A0 (gen_7_cmp_mReg_12), .A1 (nx10344), .A2 (
             nx11174)) ;
    nor03_2x ix3025 (.Y (nx3024), .A0 (nx5669), .A1 (nx11178), .A2 (nx11190)) ;
    nor02_2x ix5680 (.Y (nx5679), .A0 (nx3020), .A1 (nx3018)) ;
    nor03_2x ix3021 (.Y (nx3020), .A0 (nx5683), .A1 (nx10338), .A2 (nx11198)) ;
    dffr gen_7_cmp_mRegCmp_reg_Q_13 (.Q (gen_7_cmp_mReg_13), .QB (nx5683), .D (
         window_7__13), .CLK (start), .R (rst)) ;
    nor03_2x ix3019 (.Y (nx3018), .A0 (gen_7_cmp_mReg_13), .A1 (nx10774), .A2 (
             nx11206)) ;
    nand02 ix3055 (.Y (gen_7_cmp_BSCmp_op2_14), .A0 (nx5687), .A1 (nx5693)) ;
    nor02_2x ix5688 (.Y (nx5687), .A0 (nx3050), .A1 (nx3046)) ;
    nor03_2x ix3051 (.Y (nx3050), .A0 (gen_7_cmp_mReg_13), .A1 (nx10344), .A2 (
             nx11174)) ;
    nor03_2x ix3047 (.Y (nx3046), .A0 (nx5683), .A1 (nx11180), .A2 (nx11190)) ;
    nor02_2x ix5694 (.Y (nx5693), .A0 (nx3042), .A1 (nx3040)) ;
    nor03_2x ix3043 (.Y (nx3042), .A0 (nx5696), .A1 (nx10338), .A2 (nx11198)) ;
    dffr gen_7_cmp_mRegCmp_reg_Q_14 (.Q (gen_7_cmp_mReg_14), .QB (nx5696), .D (
         window_7__14), .CLK (start), .R (rst)) ;
    nor03_2x ix3041 (.Y (nx3040), .A0 (gen_7_cmp_mReg_14), .A1 (nx10774), .A2 (
             nx11206)) ;
    nand02 ix3077 (.Y (gen_7_cmp_BSCmp_op2_15), .A0 (nx5703), .A1 (nx5709)) ;
    nor02_2x ix5704 (.Y (nx5703), .A0 (nx3072), .A1 (nx3068)) ;
    nor03_2x ix3073 (.Y (nx3072), .A0 (gen_7_cmp_mReg_14), .A1 (nx10344), .A2 (
             nx11174)) ;
    nor03_2x ix3069 (.Y (nx3068), .A0 (nx5696), .A1 (nx11180), .A2 (nx11190)) ;
    nor02_2x ix5710 (.Y (nx5709), .A0 (nx3064), .A1 (nx3062)) ;
    nor03_2x ix3065 (.Y (nx3064), .A0 (nx5713), .A1 (nx10338), .A2 (nx11198)) ;
    dffr gen_7_cmp_mRegCmp_reg_Q_15 (.Q (gen_7_cmp_mReg_15), .QB (nx5713), .D (
         window_7__15), .CLK (start), .R (rst)) ;
    nor03_2x ix3063 (.Y (nx3062), .A0 (gen_7_cmp_mReg_15), .A1 (nx10776), .A2 (
             nx11206)) ;
    nand02 ix3087 (.Y (gen_7_cmp_BSCmp_op2_16), .A0 (nx5717), .A1 (nx5709)) ;
    nor02_2x ix5718 (.Y (nx5717), .A0 (nx3082), .A1 (nx3078)) ;
    nor03_2x ix3083 (.Y (nx3082), .A0 (gen_7_cmp_mReg_15), .A1 (nx10344), .A2 (
             nx11174)) ;
    nor03_2x ix3079 (.Y (nx3078), .A0 (nx5713), .A1 (nx11180), .A2 (nx11190)) ;
    nand02 ix3155 (.Y (gen_8_cmp_BSCmp_op2_1), .A0 (nx5725), .A1 (nx5745)) ;
    nor02_2x ix5726 (.Y (nx5725), .A0 (nx3150), .A1 (nx3146)) ;
    nor03_2x ix3151 (.Y (nx3150), .A0 (gen_8_cmp_mReg_0), .A1 (nx10328), .A2 (
             nx11210)) ;
    dffr gen_8_cmp_mRegCmp_reg_Q_0 (.Q (gen_8_cmp_mReg_0), .QB (nx5731), .D (
         window_8__0), .CLK (start), .R (rst)) ;
    inv01 ix5736 (.Y (nx5735), .A (gen_8_cmp_pMux_0)) ;
    nor03_2x ix3147 (.Y (nx3146), .A0 (nx5731), .A1 (nx11216), .A2 (nx11226)) ;
    inv02 ix5744 (.Y (nx5743), .A (gen_8_cmp_pMux_2)) ;
    nor02_2x ix5746 (.Y (nx5745), .A0 (nx3136), .A1 (nx3134)) ;
    nor03_2x ix3137 (.Y (nx3136), .A0 (nx5749), .A1 (nx10322), .A2 (nx11234)) ;
    dffr gen_8_cmp_mRegCmp_reg_Q_1 (.Q (gen_8_cmp_mReg_1), .QB (nx5749), .D (
         window_8__1), .CLK (start), .R (rst)) ;
    nor03_2x ix3135 (.Y (nx3134), .A0 (gen_8_cmp_mReg_1), .A1 (nx10778), .A2 (
             nx11242)) ;
    nor03_2x ix3095 (.Y (nx3094), .A0 (nx10328), .A1 (nx5743), .A2 (
             gen_8_cmp_pMux_0)) ;
    nand02 ix3177 (.Y (gen_8_cmp_BSCmp_op2_2), .A0 (nx5760), .A1 (nx5765)) ;
    nor02_2x ix5761 (.Y (nx5760), .A0 (nx3172), .A1 (nx3168)) ;
    nor03_2x ix3173 (.Y (nx3172), .A0 (gen_8_cmp_mReg_1), .A1 (nx10328), .A2 (
             nx11210)) ;
    nor03_2x ix3169 (.Y (nx3168), .A0 (nx5749), .A1 (nx11216), .A2 (nx11226)) ;
    nor02_2x ix5766 (.Y (nx5765), .A0 (nx3164), .A1 (nx3162)) ;
    nor03_2x ix3165 (.Y (nx3164), .A0 (nx5769), .A1 (nx10322), .A2 (nx11234)) ;
    dffr gen_8_cmp_mRegCmp_reg_Q_2 (.Q (gen_8_cmp_mReg_2), .QB (nx5769), .D (
         window_8__2), .CLK (start), .R (rst)) ;
    nor03_2x ix3163 (.Y (nx3162), .A0 (gen_8_cmp_mReg_2), .A1 (nx10778), .A2 (
             nx11242)) ;
    nand02 ix3199 (.Y (gen_8_cmp_BSCmp_op2_3), .A0 (nx5775), .A1 (nx5781)) ;
    nor02_2x ix5776 (.Y (nx5775), .A0 (nx3194), .A1 (nx3190)) ;
    nor03_2x ix3195 (.Y (nx3194), .A0 (gen_8_cmp_mReg_2), .A1 (nx10328), .A2 (
             nx11210)) ;
    nor03_2x ix3191 (.Y (nx3190), .A0 (nx5769), .A1 (nx11216), .A2 (nx11226)) ;
    nor02_2x ix5782 (.Y (nx5781), .A0 (nx3186), .A1 (nx3184)) ;
    nor03_2x ix3187 (.Y (nx3186), .A0 (nx5785), .A1 (nx10322), .A2 (nx11234)) ;
    dffr gen_8_cmp_mRegCmp_reg_Q_3 (.Q (gen_8_cmp_mReg_3), .QB (nx5785), .D (
         window_8__3), .CLK (start), .R (rst)) ;
    nor03_2x ix3185 (.Y (nx3184), .A0 (gen_8_cmp_mReg_3), .A1 (nx10778), .A2 (
             nx11242)) ;
    nand02 ix3221 (.Y (gen_8_cmp_BSCmp_op2_4), .A0 (nx5791), .A1 (nx5797)) ;
    nor02_2x ix5792 (.Y (nx5791), .A0 (nx3216), .A1 (nx3212)) ;
    nor03_2x ix3217 (.Y (nx3216), .A0 (gen_8_cmp_mReg_3), .A1 (nx10328), .A2 (
             nx11210)) ;
    nor03_2x ix3213 (.Y (nx3212), .A0 (nx5785), .A1 (nx11216), .A2 (nx11226)) ;
    nor02_2x ix5798 (.Y (nx5797), .A0 (nx3208), .A1 (nx3206)) ;
    nor03_2x ix3209 (.Y (nx3208), .A0 (nx5800), .A1 (nx10322), .A2 (nx11234)) ;
    dffr gen_8_cmp_mRegCmp_reg_Q_4 (.Q (gen_8_cmp_mReg_4), .QB (nx5800), .D (
         window_8__4), .CLK (start), .R (rst)) ;
    nor03_2x ix3207 (.Y (nx3206), .A0 (gen_8_cmp_mReg_4), .A1 (nx10778), .A2 (
             nx11242)) ;
    nand02 ix3243 (.Y (gen_8_cmp_BSCmp_op2_5), .A0 (nx5804), .A1 (nx5809)) ;
    nor02_2x ix5805 (.Y (nx5804), .A0 (nx3238), .A1 (nx3234)) ;
    nor03_2x ix3239 (.Y (nx3238), .A0 (gen_8_cmp_mReg_4), .A1 (nx10328), .A2 (
             nx11210)) ;
    nor03_2x ix3235 (.Y (nx3234), .A0 (nx5800), .A1 (nx11216), .A2 (nx11226)) ;
    nor02_2x ix5810 (.Y (nx5809), .A0 (nx3230), .A1 (nx3228)) ;
    nor03_2x ix3231 (.Y (nx3230), .A0 (nx5813), .A1 (nx10324), .A2 (nx11234)) ;
    dffr gen_8_cmp_mRegCmp_reg_Q_5 (.Q (gen_8_cmp_mReg_5), .QB (nx5813), .D (
         window_8__5), .CLK (start), .R (rst)) ;
    nor03_2x ix3229 (.Y (nx3228), .A0 (gen_8_cmp_mReg_5), .A1 (nx10778), .A2 (
             nx11242)) ;
    nand02 ix3265 (.Y (gen_8_cmp_BSCmp_op2_6), .A0 (nx5819), .A1 (nx5825)) ;
    nor02_2x ix5820 (.Y (nx5819), .A0 (nx3260), .A1 (nx3256)) ;
    nor03_2x ix3261 (.Y (nx3260), .A0 (gen_8_cmp_mReg_5), .A1 (nx10330), .A2 (
             nx11210)) ;
    nor03_2x ix3257 (.Y (nx3256), .A0 (nx5813), .A1 (nx11216), .A2 (nx11226)) ;
    nor02_2x ix5826 (.Y (nx5825), .A0 (nx3252), .A1 (nx3250)) ;
    nor03_2x ix3253 (.Y (nx3252), .A0 (nx5829), .A1 (nx10324), .A2 (nx11234)) ;
    dffr gen_8_cmp_mRegCmp_reg_Q_6 (.Q (gen_8_cmp_mReg_6), .QB (nx5829), .D (
         window_8__6), .CLK (start), .R (rst)) ;
    nor03_2x ix3251 (.Y (nx3250), .A0 (gen_8_cmp_mReg_6), .A1 (nx10778), .A2 (
             nx11242)) ;
    nand02 ix3287 (.Y (gen_8_cmp_BSCmp_op2_7), .A0 (nx5833), .A1 (nx5839)) ;
    nor02_2x ix5834 (.Y (nx5833), .A0 (nx3282), .A1 (nx3278)) ;
    nor03_2x ix3283 (.Y (nx3282), .A0 (gen_8_cmp_mReg_6), .A1 (nx10330), .A2 (
             nx11212)) ;
    nor03_2x ix3279 (.Y (nx3278), .A0 (nx5829), .A1 (nx11218), .A2 (nx11228)) ;
    nor02_2x ix5840 (.Y (nx5839), .A0 (nx3274), .A1 (nx3272)) ;
    nor03_2x ix3275 (.Y (nx3274), .A0 (nx5843), .A1 (nx10324), .A2 (nx11236)) ;
    dffr gen_8_cmp_mRegCmp_reg_Q_7 (.Q (gen_8_cmp_mReg_7), .QB (nx5843), .D (
         window_8__7), .CLK (start), .R (rst)) ;
    nor03_2x ix3273 (.Y (nx3272), .A0 (gen_8_cmp_mReg_7), .A1 (nx10778), .A2 (
             nx11244)) ;
    nand02 ix3309 (.Y (gen_8_cmp_BSCmp_op2_8), .A0 (nx5849), .A1 (nx5853)) ;
    nor02_2x ix5850 (.Y (nx5849), .A0 (nx3304), .A1 (nx3300)) ;
    nor03_2x ix3305 (.Y (nx3304), .A0 (gen_8_cmp_mReg_7), .A1 (nx10330), .A2 (
             nx11212)) ;
    nor03_2x ix3301 (.Y (nx3300), .A0 (nx5843), .A1 (nx11218), .A2 (nx11228)) ;
    nor02_2x ix5854 (.Y (nx5853), .A0 (nx3296), .A1 (nx3294)) ;
    nor03_2x ix3297 (.Y (nx3296), .A0 (nx5857), .A1 (nx10324), .A2 (nx11236)) ;
    dffr gen_8_cmp_mRegCmp_reg_Q_8 (.Q (gen_8_cmp_mReg_8), .QB (nx5857), .D (
         window_8__8), .CLK (start), .R (rst)) ;
    nor03_2x ix3295 (.Y (nx3294), .A0 (gen_8_cmp_mReg_8), .A1 (nx10780), .A2 (
             nx11244)) ;
    nand02 ix3331 (.Y (gen_8_cmp_BSCmp_op2_9), .A0 (nx5861), .A1 (nx5867)) ;
    nor02_2x ix5862 (.Y (nx5861), .A0 (nx3326), .A1 (nx3322)) ;
    nor03_2x ix3327 (.Y (nx3326), .A0 (gen_8_cmp_mReg_8), .A1 (nx10330), .A2 (
             nx11212)) ;
    nor03_2x ix3323 (.Y (nx3322), .A0 (nx5857), .A1 (nx11218), .A2 (nx11228)) ;
    nor02_2x ix5868 (.Y (nx5867), .A0 (nx3318), .A1 (nx3316)) ;
    nor03_2x ix3319 (.Y (nx3318), .A0 (nx5871), .A1 (nx10324), .A2 (nx11236)) ;
    dffr gen_8_cmp_mRegCmp_reg_Q_9 (.Q (gen_8_cmp_mReg_9), .QB (nx5871), .D (
         window_8__9), .CLK (start), .R (rst)) ;
    nor03_2x ix3317 (.Y (nx3316), .A0 (gen_8_cmp_mReg_9), .A1 (nx10780), .A2 (
             nx11244)) ;
    nand02 ix3353 (.Y (gen_8_cmp_BSCmp_op2_10), .A0 (nx5875), .A1 (nx5881)) ;
    nor02_2x ix5876 (.Y (nx5875), .A0 (nx3348), .A1 (nx3344)) ;
    nor03_2x ix3349 (.Y (nx3348), .A0 (gen_8_cmp_mReg_9), .A1 (nx10330), .A2 (
             nx11212)) ;
    nor03_2x ix3345 (.Y (nx3344), .A0 (nx5871), .A1 (nx11218), .A2 (nx11228)) ;
    nor02_2x ix5882 (.Y (nx5881), .A0 (nx3340), .A1 (nx3338)) ;
    nor03_2x ix3341 (.Y (nx3340), .A0 (nx5884), .A1 (nx10324), .A2 (nx11236)) ;
    dffr gen_8_cmp_mRegCmp_reg_Q_10 (.Q (gen_8_cmp_mReg_10), .QB (nx5884), .D (
         window_8__10), .CLK (start), .R (rst)) ;
    nor03_2x ix3339 (.Y (nx3338), .A0 (gen_8_cmp_mReg_10), .A1 (nx10780), .A2 (
             nx11244)) ;
    nand02 ix3375 (.Y (gen_8_cmp_BSCmp_op2_11), .A0 (nx5891), .A1 (nx5897)) ;
    nor02_2x ix5892 (.Y (nx5891), .A0 (nx3370), .A1 (nx3366)) ;
    nor03_2x ix3371 (.Y (nx3370), .A0 (gen_8_cmp_mReg_10), .A1 (nx10330), .A2 (
             nx11212)) ;
    nor03_2x ix3367 (.Y (nx3366), .A0 (nx5884), .A1 (nx11218), .A2 (nx11228)) ;
    nor02_2x ix5898 (.Y (nx5897), .A0 (nx3362), .A1 (nx3360)) ;
    nor03_2x ix3363 (.Y (nx3362), .A0 (nx5901), .A1 (nx10324), .A2 (nx11236)) ;
    dffr gen_8_cmp_mRegCmp_reg_Q_11 (.Q (gen_8_cmp_mReg_11), .QB (nx5901), .D (
         window_8__11), .CLK (start), .R (rst)) ;
    nor03_2x ix3361 (.Y (nx3360), .A0 (gen_8_cmp_mReg_11), .A1 (nx10780), .A2 (
             nx11244)) ;
    nand02 ix3397 (.Y (gen_8_cmp_BSCmp_op2_12), .A0 (nx5905), .A1 (nx5911)) ;
    nor02_2x ix5906 (.Y (nx5905), .A0 (nx3392), .A1 (nx3388)) ;
    nor03_2x ix3393 (.Y (nx3392), .A0 (gen_8_cmp_mReg_11), .A1 (nx10330), .A2 (
             nx11212)) ;
    nor03_2x ix3389 (.Y (nx3388), .A0 (nx5901), .A1 (nx11218), .A2 (nx11228)) ;
    nor02_2x ix5912 (.Y (nx5911), .A0 (nx3384), .A1 (nx3382)) ;
    nor03_2x ix3385 (.Y (nx3384), .A0 (nx5915), .A1 (nx10326), .A2 (nx11236)) ;
    dffr gen_8_cmp_mRegCmp_reg_Q_12 (.Q (gen_8_cmp_mReg_12), .QB (nx5915), .D (
         window_8__12), .CLK (start), .R (rst)) ;
    nor03_2x ix3383 (.Y (nx3382), .A0 (gen_8_cmp_mReg_12), .A1 (nx10780), .A2 (
             nx11244)) ;
    nand02 ix3419 (.Y (gen_8_cmp_BSCmp_op2_13), .A0 (nx5919), .A1 (nx5925)) ;
    nor02_2x ix5920 (.Y (nx5919), .A0 (nx3414), .A1 (nx3410)) ;
    nor03_2x ix3415 (.Y (nx3414), .A0 (gen_8_cmp_mReg_12), .A1 (nx10332), .A2 (
             nx11214)) ;
    nor03_2x ix3411 (.Y (nx3410), .A0 (nx5915), .A1 (nx11218), .A2 (nx11230)) ;
    nor02_2x ix5926 (.Y (nx5925), .A0 (nx3406), .A1 (nx3404)) ;
    nor03_2x ix3407 (.Y (nx3406), .A0 (nx5928), .A1 (nx10326), .A2 (nx11238)) ;
    dffr gen_8_cmp_mRegCmp_reg_Q_13 (.Q (gen_8_cmp_mReg_13), .QB (nx5928), .D (
         window_8__13), .CLK (start), .R (rst)) ;
    nor03_2x ix3405 (.Y (nx3404), .A0 (gen_8_cmp_mReg_13), .A1 (nx10780), .A2 (
             nx11246)) ;
    nand02 ix3441 (.Y (gen_8_cmp_BSCmp_op2_14), .A0 (nx5935), .A1 (nx5941)) ;
    nor02_2x ix5936 (.Y (nx5935), .A0 (nx3436), .A1 (nx3432)) ;
    nor03_2x ix3437 (.Y (nx3436), .A0 (gen_8_cmp_mReg_13), .A1 (nx10332), .A2 (
             nx11214)) ;
    nor03_2x ix3433 (.Y (nx3432), .A0 (nx5928), .A1 (nx11220), .A2 (nx11230)) ;
    nor02_2x ix5942 (.Y (nx5941), .A0 (nx3428), .A1 (nx3426)) ;
    nor03_2x ix3429 (.Y (nx3428), .A0 (nx5945), .A1 (nx10326), .A2 (nx11238)) ;
    dffr gen_8_cmp_mRegCmp_reg_Q_14 (.Q (gen_8_cmp_mReg_14), .QB (nx5945), .D (
         window_8__14), .CLK (start), .R (rst)) ;
    nor03_2x ix3427 (.Y (nx3426), .A0 (gen_8_cmp_mReg_14), .A1 (nx10780), .A2 (
             nx11246)) ;
    nand02 ix3463 (.Y (gen_8_cmp_BSCmp_op2_15), .A0 (nx5949), .A1 (nx5955)) ;
    nor02_2x ix5950 (.Y (nx5949), .A0 (nx3458), .A1 (nx3454)) ;
    nor03_2x ix3459 (.Y (nx3458), .A0 (gen_8_cmp_mReg_14), .A1 (nx10332), .A2 (
             nx11214)) ;
    nor03_2x ix3455 (.Y (nx3454), .A0 (nx5945), .A1 (nx11220), .A2 (nx11230)) ;
    nor02_2x ix5956 (.Y (nx5955), .A0 (nx3450), .A1 (nx3448)) ;
    nor03_2x ix3451 (.Y (nx3450), .A0 (nx5959), .A1 (nx10326), .A2 (nx11238)) ;
    dffr gen_8_cmp_mRegCmp_reg_Q_15 (.Q (gen_8_cmp_mReg_15), .QB (nx5959), .D (
         window_8__15), .CLK (start), .R (rst)) ;
    nor03_2x ix3449 (.Y (nx3448), .A0 (gen_8_cmp_mReg_15), .A1 (nx10782), .A2 (
             nx11246)) ;
    nand02 ix3473 (.Y (gen_8_cmp_BSCmp_op2_16), .A0 (nx5963), .A1 (nx5955)) ;
    nor02_2x ix5964 (.Y (nx5963), .A0 (nx3468), .A1 (nx3464)) ;
    nor03_2x ix3469 (.Y (nx3468), .A0 (gen_8_cmp_mReg_15), .A1 (nx10332), .A2 (
             nx11214)) ;
    nor03_2x ix3465 (.Y (nx3464), .A0 (nx5959), .A1 (nx11220), .A2 (nx11230)) ;
    nand02 ix3541 (.Y (gen_9_cmp_BSCmp_op2_1), .A0 (nx5970), .A1 (nx5989)) ;
    nor02_2x ix5971 (.Y (nx5970), .A0 (nx3536), .A1 (nx3532)) ;
    nor03_2x ix3537 (.Y (nx3536), .A0 (gen_9_cmp_mReg_0), .A1 (nx10316), .A2 (
             nx11250)) ;
    dffr gen_9_cmp_mRegCmp_reg_Q_0 (.Q (gen_9_cmp_mReg_0), .QB (nx5975), .D (
         window_9__0), .CLK (start), .R (rst)) ;
    inv01 ix5980 (.Y (nx5979), .A (gen_9_cmp_pMux_0)) ;
    nor03_2x ix3533 (.Y (nx3532), .A0 (nx5975), .A1 (nx11256), .A2 (nx11266)) ;
    inv02 ix5988 (.Y (nx5987), .A (gen_9_cmp_pMux_2)) ;
    nor02_2x ix5990 (.Y (nx5989), .A0 (nx3522), .A1 (nx3520)) ;
    nor03_2x ix3523 (.Y (nx3522), .A0 (nx5992), .A1 (nx10310), .A2 (nx11274)) ;
    dffr gen_9_cmp_mRegCmp_reg_Q_1 (.Q (gen_9_cmp_mReg_1), .QB (nx5992), .D (
         window_9__1), .CLK (start), .R (rst)) ;
    nor03_2x ix3521 (.Y (nx3520), .A0 (gen_9_cmp_mReg_1), .A1 (nx10784), .A2 (
             nx11282)) ;
    nor03_2x ix3481 (.Y (nx3480), .A0 (nx10316), .A1 (nx5987), .A2 (
             gen_9_cmp_pMux_0)) ;
    nand02 ix3563 (.Y (gen_9_cmp_BSCmp_op2_2), .A0 (nx6005), .A1 (nx6011)) ;
    nor02_2x ix6006 (.Y (nx6005), .A0 (nx3558), .A1 (nx3554)) ;
    nor03_2x ix3559 (.Y (nx3558), .A0 (gen_9_cmp_mReg_1), .A1 (nx10316), .A2 (
             nx11250)) ;
    nor03_2x ix3555 (.Y (nx3554), .A0 (nx5992), .A1 (nx11256), .A2 (nx11266)) ;
    nor02_2x ix6012 (.Y (nx6011), .A0 (nx3550), .A1 (nx3548)) ;
    nor03_2x ix3551 (.Y (nx3550), .A0 (nx6014), .A1 (nx10310), .A2 (nx11274)) ;
    dffr gen_9_cmp_mRegCmp_reg_Q_2 (.Q (gen_9_cmp_mReg_2), .QB (nx6014), .D (
         window_9__2), .CLK (start), .R (rst)) ;
    nor03_2x ix3549 (.Y (nx3548), .A0 (gen_9_cmp_mReg_2), .A1 (nx10784), .A2 (
             nx11282)) ;
    nand02 ix3585 (.Y (gen_9_cmp_BSCmp_op2_3), .A0 (nx6019), .A1 (nx6025)) ;
    nor02_2x ix6020 (.Y (nx6019), .A0 (nx3580), .A1 (nx3576)) ;
    nor03_2x ix3581 (.Y (nx3580), .A0 (gen_9_cmp_mReg_2), .A1 (nx10316), .A2 (
             nx11250)) ;
    nor03_2x ix3577 (.Y (nx3576), .A0 (nx6014), .A1 (nx11256), .A2 (nx11266)) ;
    nor02_2x ix6026 (.Y (nx6025), .A0 (nx3572), .A1 (nx3570)) ;
    nor03_2x ix3573 (.Y (nx3572), .A0 (nx6029), .A1 (nx10310), .A2 (nx11274)) ;
    dffr gen_9_cmp_mRegCmp_reg_Q_3 (.Q (gen_9_cmp_mReg_3), .QB (nx6029), .D (
         window_9__3), .CLK (start), .R (rst)) ;
    nor03_2x ix3571 (.Y (nx3570), .A0 (gen_9_cmp_mReg_3), .A1 (nx10784), .A2 (
             nx11282)) ;
    nand02 ix3607 (.Y (gen_9_cmp_BSCmp_op2_4), .A0 (nx6035), .A1 (nx6039)) ;
    nor02_2x ix6036 (.Y (nx6035), .A0 (nx3602), .A1 (nx3598)) ;
    nor03_2x ix3603 (.Y (nx3602), .A0 (gen_9_cmp_mReg_3), .A1 (nx10316), .A2 (
             nx11250)) ;
    nor03_2x ix3599 (.Y (nx3598), .A0 (nx6029), .A1 (nx11256), .A2 (nx11266)) ;
    nor02_2x ix6040 (.Y (nx6039), .A0 (nx3594), .A1 (nx3592)) ;
    nor03_2x ix3595 (.Y (nx3594), .A0 (nx6043), .A1 (nx10310), .A2 (nx11274)) ;
    dffr gen_9_cmp_mRegCmp_reg_Q_4 (.Q (gen_9_cmp_mReg_4), .QB (nx6043), .D (
         window_9__4), .CLK (start), .R (rst)) ;
    nor03_2x ix3593 (.Y (nx3592), .A0 (gen_9_cmp_mReg_4), .A1 (nx10784), .A2 (
             nx11282)) ;
    nand02 ix3629 (.Y (gen_9_cmp_BSCmp_op2_5), .A0 (nx6049), .A1 (nx6055)) ;
    nor02_2x ix6050 (.Y (nx6049), .A0 (nx3624), .A1 (nx3620)) ;
    nor03_2x ix3625 (.Y (nx3624), .A0 (gen_9_cmp_mReg_4), .A1 (nx10316), .A2 (
             nx11250)) ;
    nor03_2x ix3621 (.Y (nx3620), .A0 (nx6043), .A1 (nx11256), .A2 (nx11266)) ;
    nor02_2x ix6056 (.Y (nx6055), .A0 (nx3616), .A1 (nx3614)) ;
    nor03_2x ix3617 (.Y (nx3616), .A0 (nx6058), .A1 (nx10312), .A2 (nx11274)) ;
    dffr gen_9_cmp_mRegCmp_reg_Q_5 (.Q (gen_9_cmp_mReg_5), .QB (nx6058), .D (
         window_9__5), .CLK (start), .R (rst)) ;
    nor03_2x ix3615 (.Y (nx3614), .A0 (gen_9_cmp_mReg_5), .A1 (nx10784), .A2 (
             nx11282)) ;
    nand02 ix3651 (.Y (gen_9_cmp_BSCmp_op2_6), .A0 (nx6063), .A1 (nx6069)) ;
    nor02_2x ix6064 (.Y (nx6063), .A0 (nx3646), .A1 (nx3642)) ;
    nor03_2x ix3647 (.Y (nx3646), .A0 (gen_9_cmp_mReg_5), .A1 (nx10318), .A2 (
             nx11250)) ;
    nor03_2x ix3643 (.Y (nx3642), .A0 (nx6058), .A1 (nx11256), .A2 (nx11266)) ;
    nor02_2x ix6070 (.Y (nx6069), .A0 (nx3638), .A1 (nx3636)) ;
    nor03_2x ix3639 (.Y (nx3638), .A0 (nx6073), .A1 (nx10312), .A2 (nx11274)) ;
    dffr gen_9_cmp_mRegCmp_reg_Q_6 (.Q (gen_9_cmp_mReg_6), .QB (nx6073), .D (
         window_9__6), .CLK (start), .R (rst)) ;
    nor03_2x ix3637 (.Y (nx3636), .A0 (gen_9_cmp_mReg_6), .A1 (nx10784), .A2 (
             nx11282)) ;
    nand02 ix3673 (.Y (gen_9_cmp_BSCmp_op2_7), .A0 (nx6079), .A1 (nx6083)) ;
    nor02_2x ix6080 (.Y (nx6079), .A0 (nx3668), .A1 (nx3664)) ;
    nor03_2x ix3669 (.Y (nx3668), .A0 (gen_9_cmp_mReg_6), .A1 (nx10318), .A2 (
             nx11252)) ;
    nor03_2x ix3665 (.Y (nx3664), .A0 (nx6073), .A1 (nx11258), .A2 (nx11268)) ;
    nor02_2x ix6084 (.Y (nx6083), .A0 (nx3660), .A1 (nx3658)) ;
    nor03_2x ix3661 (.Y (nx3660), .A0 (nx6087), .A1 (nx10312), .A2 (nx11276)) ;
    dffr gen_9_cmp_mRegCmp_reg_Q_7 (.Q (gen_9_cmp_mReg_7), .QB (nx6087), .D (
         window_9__7), .CLK (start), .R (rst)) ;
    nor03_2x ix3659 (.Y (nx3658), .A0 (gen_9_cmp_mReg_7), .A1 (nx10784), .A2 (
             nx11284)) ;
    nand02 ix3695 (.Y (gen_9_cmp_BSCmp_op2_8), .A0 (nx6093), .A1 (nx6099)) ;
    nor02_2x ix6094 (.Y (nx6093), .A0 (nx3690), .A1 (nx3686)) ;
    nor03_2x ix3691 (.Y (nx3690), .A0 (gen_9_cmp_mReg_7), .A1 (nx10318), .A2 (
             nx11252)) ;
    nor03_2x ix3687 (.Y (nx3686), .A0 (nx6087), .A1 (nx11258), .A2 (nx11268)) ;
    nor02_2x ix6100 (.Y (nx6099), .A0 (nx3682), .A1 (nx3680)) ;
    nor03_2x ix3683 (.Y (nx3682), .A0 (nx6102), .A1 (nx10312), .A2 (nx11276)) ;
    dffr gen_9_cmp_mRegCmp_reg_Q_8 (.Q (gen_9_cmp_mReg_8), .QB (nx6102), .D (
         window_9__8), .CLK (start), .R (rst)) ;
    nor03_2x ix3681 (.Y (nx3680), .A0 (gen_9_cmp_mReg_8), .A1 (nx10786), .A2 (
             nx11284)) ;
    nand02 ix3717 (.Y (gen_9_cmp_BSCmp_op2_9), .A0 (nx6107), .A1 (nx6113)) ;
    nor02_2x ix6108 (.Y (nx6107), .A0 (nx3712), .A1 (nx3708)) ;
    nor03_2x ix3713 (.Y (nx3712), .A0 (gen_9_cmp_mReg_8), .A1 (nx10318), .A2 (
             nx11252)) ;
    nor03_2x ix3709 (.Y (nx3708), .A0 (nx6102), .A1 (nx11258), .A2 (nx11268)) ;
    nor02_2x ix6114 (.Y (nx6113), .A0 (nx3704), .A1 (nx3702)) ;
    nor03_2x ix3705 (.Y (nx3704), .A0 (nx6117), .A1 (nx10312), .A2 (nx11276)) ;
    dffr gen_9_cmp_mRegCmp_reg_Q_9 (.Q (gen_9_cmp_mReg_9), .QB (nx6117), .D (
         window_9__9), .CLK (start), .R (rst)) ;
    nor03_2x ix3703 (.Y (nx3702), .A0 (gen_9_cmp_mReg_9), .A1 (nx10786), .A2 (
             nx11284)) ;
    nand02 ix3739 (.Y (gen_9_cmp_BSCmp_op2_10), .A0 (nx6123), .A1 (nx6127)) ;
    nor02_2x ix6124 (.Y (nx6123), .A0 (nx3734), .A1 (nx3730)) ;
    nor03_2x ix3735 (.Y (nx3734), .A0 (gen_9_cmp_mReg_9), .A1 (nx10318), .A2 (
             nx11252)) ;
    nor03_2x ix3731 (.Y (nx3730), .A0 (nx6117), .A1 (nx11258), .A2 (nx11268)) ;
    nor02_2x ix6128 (.Y (nx6127), .A0 (nx3726), .A1 (nx3724)) ;
    nor03_2x ix3727 (.Y (nx3726), .A0 (nx6131), .A1 (nx10312), .A2 (nx11276)) ;
    dffr gen_9_cmp_mRegCmp_reg_Q_10 (.Q (gen_9_cmp_mReg_10), .QB (nx6131), .D (
         window_9__10), .CLK (start), .R (rst)) ;
    nor03_2x ix3725 (.Y (nx3724), .A0 (gen_9_cmp_mReg_10), .A1 (nx10786), .A2 (
             nx11284)) ;
    nand02 ix3761 (.Y (gen_9_cmp_BSCmp_op2_11), .A0 (nx6137), .A1 (nx6143)) ;
    nor02_2x ix6138 (.Y (nx6137), .A0 (nx3756), .A1 (nx3752)) ;
    nor03_2x ix3757 (.Y (nx3756), .A0 (gen_9_cmp_mReg_10), .A1 (nx10318), .A2 (
             nx11252)) ;
    nor03_2x ix3753 (.Y (nx3752), .A0 (nx6131), .A1 (nx11258), .A2 (nx11268)) ;
    nor02_2x ix6144 (.Y (nx6143), .A0 (nx3748), .A1 (nx3746)) ;
    nor03_2x ix3749 (.Y (nx3748), .A0 (nx6146), .A1 (nx10312), .A2 (nx11276)) ;
    dffr gen_9_cmp_mRegCmp_reg_Q_11 (.Q (gen_9_cmp_mReg_11), .QB (nx6146), .D (
         window_9__11), .CLK (start), .R (rst)) ;
    nor03_2x ix3747 (.Y (nx3746), .A0 (gen_9_cmp_mReg_11), .A1 (nx10786), .A2 (
             nx11284)) ;
    nand02 ix3783 (.Y (gen_9_cmp_BSCmp_op2_12), .A0 (nx6151), .A1 (nx6157)) ;
    nor02_2x ix6152 (.Y (nx6151), .A0 (nx3778), .A1 (nx3774)) ;
    nor03_2x ix3779 (.Y (nx3778), .A0 (gen_9_cmp_mReg_11), .A1 (nx10318), .A2 (
             nx11252)) ;
    nor03_2x ix3775 (.Y (nx3774), .A0 (nx6146), .A1 (nx11258), .A2 (nx11268)) ;
    nor02_2x ix6158 (.Y (nx6157), .A0 (nx3770), .A1 (nx3768)) ;
    nor03_2x ix3771 (.Y (nx3770), .A0 (nx6161), .A1 (nx10314), .A2 (nx11276)) ;
    dffr gen_9_cmp_mRegCmp_reg_Q_12 (.Q (gen_9_cmp_mReg_12), .QB (nx6161), .D (
         window_9__12), .CLK (start), .R (rst)) ;
    nor03_2x ix3769 (.Y (nx3768), .A0 (gen_9_cmp_mReg_12), .A1 (nx10786), .A2 (
             nx11284)) ;
    nand02 ix3805 (.Y (gen_9_cmp_BSCmp_op2_13), .A0 (nx6167), .A1 (nx6171)) ;
    nor02_2x ix6168 (.Y (nx6167), .A0 (nx3800), .A1 (nx3796)) ;
    nor03_2x ix3801 (.Y (nx3800), .A0 (gen_9_cmp_mReg_12), .A1 (nx10320), .A2 (
             nx11254)) ;
    nor03_2x ix3797 (.Y (nx3796), .A0 (nx6161), .A1 (nx11258), .A2 (nx11270)) ;
    nor02_2x ix6172 (.Y (nx6171), .A0 (nx3792), .A1 (nx3790)) ;
    nor03_2x ix3793 (.Y (nx3792), .A0 (nx6175), .A1 (nx10314), .A2 (nx11278)) ;
    dffr gen_9_cmp_mRegCmp_reg_Q_13 (.Q (gen_9_cmp_mReg_13), .QB (nx6175), .D (
         window_9__13), .CLK (start), .R (rst)) ;
    nor03_2x ix3791 (.Y (nx3790), .A0 (gen_9_cmp_mReg_13), .A1 (nx10786), .A2 (
             nx11286)) ;
    nand02 ix3827 (.Y (gen_9_cmp_BSCmp_op2_14), .A0 (nx6181), .A1 (nx6186)) ;
    nor02_2x ix6182 (.Y (nx6181), .A0 (nx3822), .A1 (nx3818)) ;
    nor03_2x ix3823 (.Y (nx3822), .A0 (gen_9_cmp_mReg_13), .A1 (nx10320), .A2 (
             nx11254)) ;
    nor03_2x ix3819 (.Y (nx3818), .A0 (nx6175), .A1 (nx11260), .A2 (nx11270)) ;
    nor02_2x ix6187 (.Y (nx6186), .A0 (nx3814), .A1 (nx3812)) ;
    nor03_2x ix3815 (.Y (nx3814), .A0 (nx6189), .A1 (nx10314), .A2 (nx11278)) ;
    dffr gen_9_cmp_mRegCmp_reg_Q_14 (.Q (gen_9_cmp_mReg_14), .QB (nx6189), .D (
         window_9__14), .CLK (start), .R (rst)) ;
    nor03_2x ix3813 (.Y (nx3812), .A0 (gen_9_cmp_mReg_14), .A1 (nx10786), .A2 (
             nx11286)) ;
    nand02 ix3849 (.Y (gen_9_cmp_BSCmp_op2_15), .A0 (nx6193), .A1 (nx6199)) ;
    nor02_2x ix6194 (.Y (nx6193), .A0 (nx3844), .A1 (nx3840)) ;
    nor03_2x ix3845 (.Y (nx3844), .A0 (gen_9_cmp_mReg_14), .A1 (nx10320), .A2 (
             nx11254)) ;
    nor03_2x ix3841 (.Y (nx3840), .A0 (nx6189), .A1 (nx11260), .A2 (nx11270)) ;
    nor02_2x ix6200 (.Y (nx6199), .A0 (nx3836), .A1 (nx3834)) ;
    nor03_2x ix3837 (.Y (nx3836), .A0 (nx6203), .A1 (nx10314), .A2 (nx11278)) ;
    dffr gen_9_cmp_mRegCmp_reg_Q_15 (.Q (gen_9_cmp_mReg_15), .QB (nx6203), .D (
         window_9__15), .CLK (start), .R (rst)) ;
    nor03_2x ix3835 (.Y (nx3834), .A0 (gen_9_cmp_mReg_15), .A1 (nx10788), .A2 (
             nx11286)) ;
    nand02 ix3859 (.Y (gen_9_cmp_BSCmp_op2_16), .A0 (nx6209), .A1 (nx6199)) ;
    nor02_2x ix6210 (.Y (nx6209), .A0 (nx3854), .A1 (nx3850)) ;
    nor03_2x ix3855 (.Y (nx3854), .A0 (gen_9_cmp_mReg_15), .A1 (nx10320), .A2 (
             nx11254)) ;
    nor03_2x ix3851 (.Y (nx3850), .A0 (nx6203), .A1 (nx11260), .A2 (nx11270)) ;
    nand02 ix3927 (.Y (gen_10_cmp_BSCmp_op2_1), .A0 (nx6217), .A1 (nx6235)) ;
    nor02_2x ix6218 (.Y (nx6217), .A0 (nx3922), .A1 (nx3918)) ;
    nor03_2x ix3923 (.Y (nx3922), .A0 (gen_10_cmp_mReg_0), .A1 (nx10304), .A2 (
             nx11290)) ;
    dffr gen_10_cmp_mRegCmp_reg_Q_0 (.Q (gen_10_cmp_mReg_0), .QB (nx6221), .D (
         window_10__0), .CLK (start), .R (rst)) ;
    inv01 ix6226 (.Y (nx6225), .A (gen_10_cmp_pMux_0)) ;
    nor03_2x ix3919 (.Y (nx3918), .A0 (nx6221), .A1 (nx11296), .A2 (nx11306)) ;
    inv02 ix6234 (.Y (nx6233), .A (gen_10_cmp_pMux_2)) ;
    nor02_2x ix6236 (.Y (nx6235), .A0 (nx3908), .A1 (nx3906)) ;
    nor03_2x ix3909 (.Y (nx3908), .A0 (nx6239), .A1 (nx10298), .A2 (nx11314)) ;
    dffr gen_10_cmp_mRegCmp_reg_Q_1 (.Q (gen_10_cmp_mReg_1), .QB (nx6239), .D (
         window_10__1), .CLK (start), .R (rst)) ;
    nor03_2x ix3907 (.Y (nx3906), .A0 (gen_10_cmp_mReg_1), .A1 (nx10790), .A2 (
             nx11322)) ;
    nor03_2x ix3867 (.Y (nx3866), .A0 (nx10304), .A1 (nx6233), .A2 (
             gen_10_cmp_pMux_0)) ;
    nand02 ix3949 (.Y (gen_10_cmp_BSCmp_op2_2), .A0 (nx6249), .A1 (nx6255)) ;
    nor02_2x ix6250 (.Y (nx6249), .A0 (nx3944), .A1 (nx3940)) ;
    nor03_2x ix3945 (.Y (nx3944), .A0 (gen_10_cmp_mReg_1), .A1 (nx10304), .A2 (
             nx11290)) ;
    nor03_2x ix3941 (.Y (nx3940), .A0 (nx6239), .A1 (nx11296), .A2 (nx11306)) ;
    nor02_2x ix6256 (.Y (nx6255), .A0 (nx3936), .A1 (nx3934)) ;
    nor03_2x ix3937 (.Y (nx3936), .A0 (nx6259), .A1 (nx10298), .A2 (nx11314)) ;
    dffr gen_10_cmp_mRegCmp_reg_Q_2 (.Q (gen_10_cmp_mReg_2), .QB (nx6259), .D (
         window_10__2), .CLK (start), .R (rst)) ;
    nor03_2x ix3935 (.Y (nx3934), .A0 (gen_10_cmp_mReg_2), .A1 (nx10790), .A2 (
             nx11322)) ;
    nand02 ix3971 (.Y (gen_10_cmp_BSCmp_op2_3), .A0 (nx6265), .A1 (nx6269)) ;
    nor02_2x ix6266 (.Y (nx6265), .A0 (nx3966), .A1 (nx3962)) ;
    nor03_2x ix3967 (.Y (nx3966), .A0 (gen_10_cmp_mReg_2), .A1 (nx10304), .A2 (
             nx11290)) ;
    nor03_2x ix3963 (.Y (nx3962), .A0 (nx6259), .A1 (nx11296), .A2 (nx11306)) ;
    nor02_2x ix6270 (.Y (nx6269), .A0 (nx3958), .A1 (nx3956)) ;
    nor03_2x ix3959 (.Y (nx3958), .A0 (nx6273), .A1 (nx10298), .A2 (nx11314)) ;
    dffr gen_10_cmp_mRegCmp_reg_Q_3 (.Q (gen_10_cmp_mReg_3), .QB (nx6273), .D (
         window_10__3), .CLK (start), .R (rst)) ;
    nor03_2x ix3957 (.Y (nx3956), .A0 (gen_10_cmp_mReg_3), .A1 (nx10790), .A2 (
             nx11322)) ;
    nand02 ix3993 (.Y (gen_10_cmp_BSCmp_op2_4), .A0 (nx6279), .A1 (nx6283)) ;
    nor02_2x ix6280 (.Y (nx6279), .A0 (nx3988), .A1 (nx3984)) ;
    nor03_2x ix3989 (.Y (nx3988), .A0 (gen_10_cmp_mReg_3), .A1 (nx10304), .A2 (
             nx11290)) ;
    nor03_2x ix3985 (.Y (nx3984), .A0 (nx6273), .A1 (nx11296), .A2 (nx11306)) ;
    nor02_2x ix6284 (.Y (nx6283), .A0 (nx3980), .A1 (nx3978)) ;
    nor03_2x ix3981 (.Y (nx3980), .A0 (nx6287), .A1 (nx10298), .A2 (nx11314)) ;
    dffr gen_10_cmp_mRegCmp_reg_Q_4 (.Q (gen_10_cmp_mReg_4), .QB (nx6287), .D (
         window_10__4), .CLK (start), .R (rst)) ;
    nor03_2x ix3979 (.Y (nx3978), .A0 (gen_10_cmp_mReg_4), .A1 (nx10790), .A2 (
             nx11322)) ;
    nand02 ix4015 (.Y (gen_10_cmp_BSCmp_op2_5), .A0 (nx6291), .A1 (nx6297)) ;
    nor02_2x ix6292 (.Y (nx6291), .A0 (nx4010), .A1 (nx4006)) ;
    nor03_2x ix4011 (.Y (nx4010), .A0 (gen_10_cmp_mReg_4), .A1 (nx10304), .A2 (
             nx11290)) ;
    nor03_2x ix4007 (.Y (nx4006), .A0 (nx6287), .A1 (nx11296), .A2 (nx11306)) ;
    nor02_2x ix6298 (.Y (nx6297), .A0 (nx4002), .A1 (nx4000)) ;
    nor03_2x ix4003 (.Y (nx4002), .A0 (nx6301), .A1 (nx10300), .A2 (nx11314)) ;
    dffr gen_10_cmp_mRegCmp_reg_Q_5 (.Q (gen_10_cmp_mReg_5), .QB (nx6301), .D (
         window_10__5), .CLK (start), .R (rst)) ;
    nor03_2x ix4001 (.Y (nx4000), .A0 (gen_10_cmp_mReg_5), .A1 (nx10790), .A2 (
             nx11322)) ;
    nand02 ix4037 (.Y (gen_10_cmp_BSCmp_op2_6), .A0 (nx6305), .A1 (nx6311)) ;
    nor02_2x ix6306 (.Y (nx6305), .A0 (nx4032), .A1 (nx4028)) ;
    nor03_2x ix4033 (.Y (nx4032), .A0 (gen_10_cmp_mReg_5), .A1 (nx10306), .A2 (
             nx11290)) ;
    nor03_2x ix4029 (.Y (nx4028), .A0 (nx6301), .A1 (nx11296), .A2 (nx11306)) ;
    nor02_2x ix6312 (.Y (nx6311), .A0 (nx4024), .A1 (nx4022)) ;
    nor03_2x ix4025 (.Y (nx4024), .A0 (nx6314), .A1 (nx10300), .A2 (nx11314)) ;
    dffr gen_10_cmp_mRegCmp_reg_Q_6 (.Q (gen_10_cmp_mReg_6), .QB (nx6314), .D (
         window_10__6), .CLK (start), .R (rst)) ;
    nor03_2x ix4023 (.Y (nx4022), .A0 (gen_10_cmp_mReg_6), .A1 (nx10790), .A2 (
             nx11322)) ;
    nand02 ix4059 (.Y (gen_10_cmp_BSCmp_op2_7), .A0 (nx6321), .A1 (nx6327)) ;
    nor02_2x ix6322 (.Y (nx6321), .A0 (nx4054), .A1 (nx4050)) ;
    nor03_2x ix4055 (.Y (nx4054), .A0 (gen_10_cmp_mReg_6), .A1 (nx10306), .A2 (
             nx11292)) ;
    nor03_2x ix4051 (.Y (nx4050), .A0 (nx6314), .A1 (nx11298), .A2 (nx11308)) ;
    nor02_2x ix6328 (.Y (nx6327), .A0 (nx4046), .A1 (nx4044)) ;
    nor03_2x ix4047 (.Y (nx4046), .A0 (nx6331), .A1 (nx10300), .A2 (nx11316)) ;
    dffr gen_10_cmp_mRegCmp_reg_Q_7 (.Q (gen_10_cmp_mReg_7), .QB (nx6331), .D (
         window_10__7), .CLK (start), .R (rst)) ;
    nor03_2x ix4045 (.Y (nx4044), .A0 (gen_10_cmp_mReg_7), .A1 (nx10790), .A2 (
             nx11324)) ;
    nand02 ix4081 (.Y (gen_10_cmp_BSCmp_op2_8), .A0 (nx6335), .A1 (nx6341)) ;
    nor02_2x ix6336 (.Y (nx6335), .A0 (nx4076), .A1 (nx4072)) ;
    nor03_2x ix4077 (.Y (nx4076), .A0 (gen_10_cmp_mReg_7), .A1 (nx10306), .A2 (
             nx11292)) ;
    nor03_2x ix4073 (.Y (nx4072), .A0 (nx6331), .A1 (nx11298), .A2 (nx11308)) ;
    nor02_2x ix6342 (.Y (nx6341), .A0 (nx4068), .A1 (nx4066)) ;
    nor03_2x ix4069 (.Y (nx4068), .A0 (nx6345), .A1 (nx10300), .A2 (nx11316)) ;
    dffr gen_10_cmp_mRegCmp_reg_Q_8 (.Q (gen_10_cmp_mReg_8), .QB (nx6345), .D (
         window_10__8), .CLK (start), .R (rst)) ;
    nor03_2x ix4067 (.Y (nx4066), .A0 (gen_10_cmp_mReg_8), .A1 (nx10792), .A2 (
             nx11324)) ;
    nand02 ix4103 (.Y (gen_10_cmp_BSCmp_op2_9), .A0 (nx6349), .A1 (nx6355)) ;
    nor02_2x ix6350 (.Y (nx6349), .A0 (nx4098), .A1 (nx4094)) ;
    nor03_2x ix4099 (.Y (nx4098), .A0 (gen_10_cmp_mReg_8), .A1 (nx10306), .A2 (
             nx11292)) ;
    nor03_2x ix4095 (.Y (nx4094), .A0 (nx6345), .A1 (nx11298), .A2 (nx11308)) ;
    nor02_2x ix6356 (.Y (nx6355), .A0 (nx4090), .A1 (nx4088)) ;
    nor03_2x ix4091 (.Y (nx4090), .A0 (nx6358), .A1 (nx10300), .A2 (nx11316)) ;
    dffr gen_10_cmp_mRegCmp_reg_Q_9 (.Q (gen_10_cmp_mReg_9), .QB (nx6358), .D (
         window_10__9), .CLK (start), .R (rst)) ;
    nor03_2x ix4089 (.Y (nx4088), .A0 (gen_10_cmp_mReg_9), .A1 (nx10792), .A2 (
             nx11324)) ;
    nand02 ix4125 (.Y (gen_10_cmp_BSCmp_op2_10), .A0 (nx6365), .A1 (nx6371)) ;
    nor02_2x ix6366 (.Y (nx6365), .A0 (nx4120), .A1 (nx4116)) ;
    nor03_2x ix4121 (.Y (nx4120), .A0 (gen_10_cmp_mReg_9), .A1 (nx10306), .A2 (
             nx11292)) ;
    nor03_2x ix4117 (.Y (nx4116), .A0 (nx6358), .A1 (nx11298), .A2 (nx11308)) ;
    nor02_2x ix6372 (.Y (nx6371), .A0 (nx4112), .A1 (nx4110)) ;
    nor03_2x ix4113 (.Y (nx4112), .A0 (nx6375), .A1 (nx10300), .A2 (nx11316)) ;
    dffr gen_10_cmp_mRegCmp_reg_Q_10 (.Q (gen_10_cmp_mReg_10), .QB (nx6375), .D (
         window_10__10), .CLK (start), .R (rst)) ;
    nor03_2x ix4111 (.Y (nx4110), .A0 (gen_10_cmp_mReg_10), .A1 (nx10792), .A2 (
             nx11324)) ;
    nand02 ix4147 (.Y (gen_10_cmp_BSCmp_op2_11), .A0 (nx6379), .A1 (nx6385)) ;
    nor02_2x ix6380 (.Y (nx6379), .A0 (nx4142), .A1 (nx4138)) ;
    nor03_2x ix4143 (.Y (nx4142), .A0 (gen_10_cmp_mReg_10), .A1 (nx10306), .A2 (
             nx11292)) ;
    nor03_2x ix4139 (.Y (nx4138), .A0 (nx6375), .A1 (nx11298), .A2 (nx11308)) ;
    nor02_2x ix6386 (.Y (nx6385), .A0 (nx4134), .A1 (nx4132)) ;
    nor03_2x ix4135 (.Y (nx4134), .A0 (nx6389), .A1 (nx10300), .A2 (nx11316)) ;
    dffr gen_10_cmp_mRegCmp_reg_Q_11 (.Q (gen_10_cmp_mReg_11), .QB (nx6389), .D (
         window_10__11), .CLK (start), .R (rst)) ;
    nor03_2x ix4133 (.Y (nx4132), .A0 (gen_10_cmp_mReg_11), .A1 (nx10792), .A2 (
             nx11324)) ;
    nand02 ix4169 (.Y (gen_10_cmp_BSCmp_op2_12), .A0 (nx6393), .A1 (nx6399)) ;
    nor02_2x ix6394 (.Y (nx6393), .A0 (nx4164), .A1 (nx4160)) ;
    nor03_2x ix4165 (.Y (nx4164), .A0 (gen_10_cmp_mReg_11), .A1 (nx10306), .A2 (
             nx11292)) ;
    nor03_2x ix4161 (.Y (nx4160), .A0 (nx6389), .A1 (nx11298), .A2 (nx11308)) ;
    nor02_2x ix6400 (.Y (nx6399), .A0 (nx4156), .A1 (nx4154)) ;
    nor03_2x ix4157 (.Y (nx4156), .A0 (nx6402), .A1 (nx10302), .A2 (nx11316)) ;
    dffr gen_10_cmp_mRegCmp_reg_Q_12 (.Q (gen_10_cmp_mReg_12), .QB (nx6402), .D (
         window_10__12), .CLK (start), .R (rst)) ;
    nor03_2x ix4155 (.Y (nx4154), .A0 (gen_10_cmp_mReg_12), .A1 (nx10792), .A2 (
             nx11324)) ;
    nand02 ix4191 (.Y (gen_10_cmp_BSCmp_op2_13), .A0 (nx6409), .A1 (nx6415)) ;
    nor02_2x ix6410 (.Y (nx6409), .A0 (nx4186), .A1 (nx4182)) ;
    nor03_2x ix4187 (.Y (nx4186), .A0 (gen_10_cmp_mReg_12), .A1 (nx10308), .A2 (
             nx11294)) ;
    nor03_2x ix4183 (.Y (nx4182), .A0 (nx6402), .A1 (nx11298), .A2 (nx11310)) ;
    nor02_2x ix6416 (.Y (nx6415), .A0 (nx4178), .A1 (nx4176)) ;
    nor03_2x ix4179 (.Y (nx4178), .A0 (nx6419), .A1 (nx10302), .A2 (nx11318)) ;
    dffr gen_10_cmp_mRegCmp_reg_Q_13 (.Q (gen_10_cmp_mReg_13), .QB (nx6419), .D (
         window_10__13), .CLK (start), .R (rst)) ;
    nor03_2x ix4177 (.Y (nx4176), .A0 (gen_10_cmp_mReg_13), .A1 (nx10792), .A2 (
             nx11326)) ;
    nand02 ix4213 (.Y (gen_10_cmp_BSCmp_op2_14), .A0 (nx6423), .A1 (nx6429)) ;
    nor02_2x ix6424 (.Y (nx6423), .A0 (nx4208), .A1 (nx4204)) ;
    nor03_2x ix4209 (.Y (nx4208), .A0 (gen_10_cmp_mReg_13), .A1 (nx10308), .A2 (
             nx11294)) ;
    nor03_2x ix4205 (.Y (nx4204), .A0 (nx6419), .A1 (nx11300), .A2 (nx11310)) ;
    nor02_2x ix6430 (.Y (nx6429), .A0 (nx4200), .A1 (nx4198)) ;
    nor03_2x ix4201 (.Y (nx4200), .A0 (nx6433), .A1 (nx10302), .A2 (nx11318)) ;
    dffr gen_10_cmp_mRegCmp_reg_Q_14 (.Q (gen_10_cmp_mReg_14), .QB (nx6433), .D (
         window_10__14), .CLK (start), .R (rst)) ;
    nor03_2x ix4199 (.Y (nx4198), .A0 (gen_10_cmp_mReg_14), .A1 (nx10792), .A2 (
             nx11326)) ;
    nand02 ix4235 (.Y (gen_10_cmp_BSCmp_op2_15), .A0 (nx6437), .A1 (nx6443)) ;
    nor02_2x ix6438 (.Y (nx6437), .A0 (nx4230), .A1 (nx4226)) ;
    nor03_2x ix4231 (.Y (nx4230), .A0 (gen_10_cmp_mReg_14), .A1 (nx10308), .A2 (
             nx11294)) ;
    nor03_2x ix4227 (.Y (nx4226), .A0 (nx6433), .A1 (nx11300), .A2 (nx11310)) ;
    nor02_2x ix6444 (.Y (nx6443), .A0 (nx4222), .A1 (nx4220)) ;
    nor03_2x ix4223 (.Y (nx4222), .A0 (nx6446), .A1 (nx10302), .A2 (nx11318)) ;
    dffr gen_10_cmp_mRegCmp_reg_Q_15 (.Q (gen_10_cmp_mReg_15), .QB (nx6446), .D (
         window_10__15), .CLK (start), .R (rst)) ;
    nor03_2x ix4221 (.Y (nx4220), .A0 (gen_10_cmp_mReg_15), .A1 (nx10794), .A2 (
             nx11326)) ;
    nand02 ix4245 (.Y (gen_10_cmp_BSCmp_op2_16), .A0 (nx6453), .A1 (nx6443)) ;
    nor02_2x ix6454 (.Y (nx6453), .A0 (nx4240), .A1 (nx4236)) ;
    nor03_2x ix4241 (.Y (nx4240), .A0 (gen_10_cmp_mReg_15), .A1 (nx10308), .A2 (
             nx11294)) ;
    nor03_2x ix4237 (.Y (nx4236), .A0 (nx6446), .A1 (nx11300), .A2 (nx11310)) ;
    nand02 ix4313 (.Y (gen_11_cmp_BSCmp_op2_1), .A0 (nx6459), .A1 (nx6479)) ;
    nor02_2x ix6460 (.Y (nx6459), .A0 (nx4308), .A1 (nx4304)) ;
    nor03_2x ix4309 (.Y (nx4308), .A0 (gen_11_cmp_mReg_0), .A1 (nx10292), .A2 (
             nx11330)) ;
    dffr gen_11_cmp_mRegCmp_reg_Q_0 (.Q (gen_11_cmp_mReg_0), .QB (nx6465), .D (
         window_11__0), .CLK (start), .R (rst)) ;
    inv01 ix6470 (.Y (nx6468), .A (gen_11_cmp_pMux_0)) ;
    nor03_2x ix4305 (.Y (nx4304), .A0 (nx6465), .A1 (nx11336), .A2 (nx11346)) ;
    inv02 ix6478 (.Y (nx6477), .A (gen_11_cmp_pMux_2)) ;
    nor02_2x ix6480 (.Y (nx6479), .A0 (nx4294), .A1 (nx4292)) ;
    nor03_2x ix4295 (.Y (nx4294), .A0 (nx6483), .A1 (nx10286), .A2 (nx11354)) ;
    dffr gen_11_cmp_mRegCmp_reg_Q_1 (.Q (gen_11_cmp_mReg_1), .QB (nx6483), .D (
         window_11__1), .CLK (start), .R (rst)) ;
    nor03_2x ix4293 (.Y (nx4292), .A0 (gen_11_cmp_mReg_1), .A1 (nx10796), .A2 (
             nx11362)) ;
    nor03_2x ix4253 (.Y (nx4252), .A0 (nx10292), .A1 (nx6477), .A2 (
             gen_11_cmp_pMux_0)) ;
    nand02 ix4335 (.Y (gen_11_cmp_BSCmp_op2_2), .A0 (nx6493), .A1 (nx6499)) ;
    nor02_2x ix6494 (.Y (nx6493), .A0 (nx4330), .A1 (nx4326)) ;
    nor03_2x ix4331 (.Y (nx4330), .A0 (gen_11_cmp_mReg_1), .A1 (nx10292), .A2 (
             nx11330)) ;
    nor03_2x ix4327 (.Y (nx4326), .A0 (nx6483), .A1 (nx11336), .A2 (nx11346)) ;
    nor02_2x ix6500 (.Y (nx6499), .A0 (nx4322), .A1 (nx4320)) ;
    nor03_2x ix4323 (.Y (nx4322), .A0 (nx6503), .A1 (nx10286), .A2 (nx11354)) ;
    dffr gen_11_cmp_mRegCmp_reg_Q_2 (.Q (gen_11_cmp_mReg_2), .QB (nx6503), .D (
         window_11__2), .CLK (start), .R (rst)) ;
    nor03_2x ix4321 (.Y (nx4320), .A0 (gen_11_cmp_mReg_2), .A1 (nx10796), .A2 (
             nx11362)) ;
    nand02 ix4357 (.Y (gen_11_cmp_BSCmp_op2_3), .A0 (nx6509), .A1 (nx6513)) ;
    nor02_2x ix6510 (.Y (nx6509), .A0 (nx4352), .A1 (nx4348)) ;
    nor03_2x ix4353 (.Y (nx4352), .A0 (gen_11_cmp_mReg_2), .A1 (nx10292), .A2 (
             nx11330)) ;
    nor03_2x ix4349 (.Y (nx4348), .A0 (nx6503), .A1 (nx11336), .A2 (nx11346)) ;
    nor02_2x ix6514 (.Y (nx6513), .A0 (nx4344), .A1 (nx4342)) ;
    nor03_2x ix4345 (.Y (nx4344), .A0 (nx6517), .A1 (nx10286), .A2 (nx11354)) ;
    dffr gen_11_cmp_mRegCmp_reg_Q_3 (.Q (gen_11_cmp_mReg_3), .QB (nx6517), .D (
         window_11__3), .CLK (start), .R (rst)) ;
    nor03_2x ix4343 (.Y (nx4342), .A0 (gen_11_cmp_mReg_3), .A1 (nx10796), .A2 (
             nx11362)) ;
    nand02 ix4379 (.Y (gen_11_cmp_BSCmp_op2_4), .A0 (nx6523), .A1 (nx6529)) ;
    nor02_2x ix6524 (.Y (nx6523), .A0 (nx4374), .A1 (nx4370)) ;
    nor03_2x ix4375 (.Y (nx4374), .A0 (gen_11_cmp_mReg_3), .A1 (nx10292), .A2 (
             nx11330)) ;
    nor03_2x ix4371 (.Y (nx4370), .A0 (nx6517), .A1 (nx11336), .A2 (nx11346)) ;
    nor02_2x ix6530 (.Y (nx6529), .A0 (nx4366), .A1 (nx4364)) ;
    nor03_2x ix4367 (.Y (nx4366), .A0 (nx6532), .A1 (nx10286), .A2 (nx11354)) ;
    dffr gen_11_cmp_mRegCmp_reg_Q_4 (.Q (gen_11_cmp_mReg_4), .QB (nx6532), .D (
         window_11__4), .CLK (start), .R (rst)) ;
    nor03_2x ix4365 (.Y (nx4364), .A0 (gen_11_cmp_mReg_4), .A1 (nx10796), .A2 (
             nx11362)) ;
    nand02 ix4401 (.Y (gen_11_cmp_BSCmp_op2_5), .A0 (nx6537), .A1 (nx6543)) ;
    nor02_2x ix6538 (.Y (nx6537), .A0 (nx4396), .A1 (nx4392)) ;
    nor03_2x ix4397 (.Y (nx4396), .A0 (gen_11_cmp_mReg_4), .A1 (nx10292), .A2 (
             nx11330)) ;
    nor03_2x ix4393 (.Y (nx4392), .A0 (nx6532), .A1 (nx11336), .A2 (nx11346)) ;
    nor02_2x ix6544 (.Y (nx6543), .A0 (nx4388), .A1 (nx4386)) ;
    nor03_2x ix4389 (.Y (nx4388), .A0 (nx6547), .A1 (nx10288), .A2 (nx11354)) ;
    dffr gen_11_cmp_mRegCmp_reg_Q_5 (.Q (gen_11_cmp_mReg_5), .QB (nx6547), .D (
         window_11__5), .CLK (start), .R (rst)) ;
    nor03_2x ix4387 (.Y (nx4386), .A0 (gen_11_cmp_mReg_5), .A1 (nx10796), .A2 (
             nx11362)) ;
    nand02 ix4423 (.Y (gen_11_cmp_BSCmp_op2_6), .A0 (nx6553), .A1 (nx6557)) ;
    nor02_2x ix6554 (.Y (nx6553), .A0 (nx4418), .A1 (nx4414)) ;
    nor03_2x ix4419 (.Y (nx4418), .A0 (gen_11_cmp_mReg_5), .A1 (nx10294), .A2 (
             nx11330)) ;
    nor03_2x ix4415 (.Y (nx4414), .A0 (nx6547), .A1 (nx11336), .A2 (nx11346)) ;
    nor02_2x ix6558 (.Y (nx6557), .A0 (nx4410), .A1 (nx4408)) ;
    nor03_2x ix4411 (.Y (nx4410), .A0 (nx6561), .A1 (nx10288), .A2 (nx11354)) ;
    dffr gen_11_cmp_mRegCmp_reg_Q_6 (.Q (gen_11_cmp_mReg_6), .QB (nx6561), .D (
         window_11__6), .CLK (start), .R (rst)) ;
    nor03_2x ix4409 (.Y (nx4408), .A0 (gen_11_cmp_mReg_6), .A1 (nx10796), .A2 (
             nx11362)) ;
    nand02 ix4445 (.Y (gen_11_cmp_BSCmp_op2_7), .A0 (nx6567), .A1 (nx6572)) ;
    nor02_2x ix6568 (.Y (nx6567), .A0 (nx4440), .A1 (nx4436)) ;
    nor03_2x ix4441 (.Y (nx4440), .A0 (gen_11_cmp_mReg_6), .A1 (nx10294), .A2 (
             nx11332)) ;
    nor03_2x ix4437 (.Y (nx4436), .A0 (nx6561), .A1 (nx11338), .A2 (nx11348)) ;
    nor02_2x ix6573 (.Y (nx6572), .A0 (nx4432), .A1 (nx4430)) ;
    nor03_2x ix4433 (.Y (nx4432), .A0 (nx6575), .A1 (nx10288), .A2 (nx11356)) ;
    dffr gen_11_cmp_mRegCmp_reg_Q_7 (.Q (gen_11_cmp_mReg_7), .QB (nx6575), .D (
         window_11__7), .CLK (start), .R (rst)) ;
    nor03_2x ix4431 (.Y (nx4430), .A0 (gen_11_cmp_mReg_7), .A1 (nx10796), .A2 (
             nx11364)) ;
    nand02 ix4467 (.Y (gen_11_cmp_BSCmp_op2_8), .A0 (nx6579), .A1 (nx6585)) ;
    nor02_2x ix6580 (.Y (nx6579), .A0 (nx4462), .A1 (nx4458)) ;
    nor03_2x ix4463 (.Y (nx4462), .A0 (gen_11_cmp_mReg_7), .A1 (nx10294), .A2 (
             nx11332)) ;
    nor03_2x ix4459 (.Y (nx4458), .A0 (nx6575), .A1 (nx11338), .A2 (nx11348)) ;
    nor02_2x ix6586 (.Y (nx6585), .A0 (nx4454), .A1 (nx4452)) ;
    nor03_2x ix4455 (.Y (nx4454), .A0 (nx6589), .A1 (nx10288), .A2 (nx11356)) ;
    dffr gen_11_cmp_mRegCmp_reg_Q_8 (.Q (gen_11_cmp_mReg_8), .QB (nx6589), .D (
         window_11__8), .CLK (start), .R (rst)) ;
    nor03_2x ix4453 (.Y (nx4452), .A0 (gen_11_cmp_mReg_8), .A1 (nx10798), .A2 (
             nx11364)) ;
    nand02 ix4489 (.Y (gen_11_cmp_BSCmp_op2_9), .A0 (nx6595), .A1 (nx6601)) ;
    nor02_2x ix6596 (.Y (nx6595), .A0 (nx4484), .A1 (nx4480)) ;
    nor03_2x ix4485 (.Y (nx4484), .A0 (gen_11_cmp_mReg_8), .A1 (nx10294), .A2 (
             nx11332)) ;
    nor03_2x ix4481 (.Y (nx4480), .A0 (nx6589), .A1 (nx11338), .A2 (nx11348)) ;
    nor02_2x ix6602 (.Y (nx6601), .A0 (nx4476), .A1 (nx4474)) ;
    nor03_2x ix4477 (.Y (nx4476), .A0 (nx6604), .A1 (nx10288), .A2 (nx11356)) ;
    dffr gen_11_cmp_mRegCmp_reg_Q_9 (.Q (gen_11_cmp_mReg_9), .QB (nx6604), .D (
         window_11__9), .CLK (start), .R (rst)) ;
    nor03_2x ix4475 (.Y (nx4474), .A0 (gen_11_cmp_mReg_9), .A1 (nx10798), .A2 (
             nx11364)) ;
    nand02 ix4511 (.Y (gen_11_cmp_BSCmp_op2_10), .A0 (nx6609), .A1 (nx6615)) ;
    nor02_2x ix6610 (.Y (nx6609), .A0 (nx4506), .A1 (nx4502)) ;
    nor03_2x ix4507 (.Y (nx4506), .A0 (gen_11_cmp_mReg_9), .A1 (nx10294), .A2 (
             nx11332)) ;
    nor03_2x ix4503 (.Y (nx4502), .A0 (nx6604), .A1 (nx11338), .A2 (nx11348)) ;
    nor02_2x ix6616 (.Y (nx6615), .A0 (nx4498), .A1 (nx4496)) ;
    nor03_2x ix4499 (.Y (nx4498), .A0 (nx6619), .A1 (nx10288), .A2 (nx11356)) ;
    dffr gen_11_cmp_mRegCmp_reg_Q_10 (.Q (gen_11_cmp_mReg_10), .QB (nx6619), .D (
         window_11__10), .CLK (start), .R (rst)) ;
    nor03_2x ix4497 (.Y (nx4496), .A0 (gen_11_cmp_mReg_10), .A1 (nx10798), .A2 (
             nx11364)) ;
    nand02 ix4533 (.Y (gen_11_cmp_BSCmp_op2_11), .A0 (nx6625), .A1 (nx6631)) ;
    nor02_2x ix6626 (.Y (nx6625), .A0 (nx4528), .A1 (nx4524)) ;
    nor03_2x ix4529 (.Y (nx4528), .A0 (gen_11_cmp_mReg_10), .A1 (nx10294), .A2 (
             nx11332)) ;
    nor03_2x ix4525 (.Y (nx4524), .A0 (nx6619), .A1 (nx11338), .A2 (nx11348)) ;
    nor02_2x ix6632 (.Y (nx6631), .A0 (nx4520), .A1 (nx4518)) ;
    nor03_2x ix4521 (.Y (nx4520), .A0 (nx6634), .A1 (nx10288), .A2 (nx11356)) ;
    dffr gen_11_cmp_mRegCmp_reg_Q_11 (.Q (gen_11_cmp_mReg_11), .QB (nx6634), .D (
         window_11__11), .CLK (start), .R (rst)) ;
    nor03_2x ix4519 (.Y (nx4518), .A0 (gen_11_cmp_mReg_11), .A1 (nx10798), .A2 (
             nx11364)) ;
    nand02 ix4555 (.Y (gen_11_cmp_BSCmp_op2_12), .A0 (nx6641), .A1 (nx6647)) ;
    nor02_2x ix6642 (.Y (nx6641), .A0 (nx4550), .A1 (nx4546)) ;
    nor03_2x ix4551 (.Y (nx4550), .A0 (gen_11_cmp_mReg_11), .A1 (nx10294), .A2 (
             nx11332)) ;
    nor03_2x ix4547 (.Y (nx4546), .A0 (nx6634), .A1 (nx11338), .A2 (nx11348)) ;
    nor02_2x ix6648 (.Y (nx6647), .A0 (nx4542), .A1 (nx4540)) ;
    nor03_2x ix4543 (.Y (nx4542), .A0 (nx6651), .A1 (nx10290), .A2 (nx11356)) ;
    dffr gen_11_cmp_mRegCmp_reg_Q_12 (.Q (gen_11_cmp_mReg_12), .QB (nx6651), .D (
         window_11__12), .CLK (start), .R (rst)) ;
    nor03_2x ix4541 (.Y (nx4540), .A0 (gen_11_cmp_mReg_12), .A1 (nx10798), .A2 (
             nx11364)) ;
    nand02 ix4577 (.Y (gen_11_cmp_BSCmp_op2_13), .A0 (nx6655), .A1 (nx6661)) ;
    nor02_2x ix6656 (.Y (nx6655), .A0 (nx4572), .A1 (nx4568)) ;
    nor03_2x ix4573 (.Y (nx4572), .A0 (gen_11_cmp_mReg_12), .A1 (nx10296), .A2 (
             nx11334)) ;
    nor03_2x ix4569 (.Y (nx4568), .A0 (nx6651), .A1 (nx11338), .A2 (nx11350)) ;
    nor02_2x ix6662 (.Y (nx6661), .A0 (nx4564), .A1 (nx4562)) ;
    nor03_2x ix4565 (.Y (nx4564), .A0 (nx6665), .A1 (nx10290), .A2 (nx11358)) ;
    dffr gen_11_cmp_mRegCmp_reg_Q_13 (.Q (gen_11_cmp_mReg_13), .QB (nx6665), .D (
         window_11__13), .CLK (start), .R (rst)) ;
    nor03_2x ix4563 (.Y (nx4562), .A0 (gen_11_cmp_mReg_13), .A1 (nx10798), .A2 (
             nx11366)) ;
    nand02 ix4599 (.Y (gen_11_cmp_BSCmp_op2_14), .A0 (nx6669), .A1 (nx6675)) ;
    nor02_2x ix6670 (.Y (nx6669), .A0 (nx4594), .A1 (nx4590)) ;
    nor03_2x ix4595 (.Y (nx4594), .A0 (gen_11_cmp_mReg_13), .A1 (nx10296), .A2 (
             nx11334)) ;
    nor03_2x ix4591 (.Y (nx4590), .A0 (nx6665), .A1 (nx11340), .A2 (nx11350)) ;
    nor02_2x ix6676 (.Y (nx6675), .A0 (nx4586), .A1 (nx4584)) ;
    nor03_2x ix4587 (.Y (nx4586), .A0 (nx6678), .A1 (nx10290), .A2 (nx11358)) ;
    dffr gen_11_cmp_mRegCmp_reg_Q_14 (.Q (gen_11_cmp_mReg_14), .QB (nx6678), .D (
         window_11__14), .CLK (start), .R (rst)) ;
    nor03_2x ix4585 (.Y (nx4584), .A0 (gen_11_cmp_mReg_14), .A1 (nx10798), .A2 (
             nx11366)) ;
    nand02 ix4621 (.Y (gen_11_cmp_BSCmp_op2_15), .A0 (nx6685), .A1 (nx6691)) ;
    nor02_2x ix6686 (.Y (nx6685), .A0 (nx4616), .A1 (nx4612)) ;
    nor03_2x ix4617 (.Y (nx4616), .A0 (gen_11_cmp_mReg_14), .A1 (nx10296), .A2 (
             nx11334)) ;
    nor03_2x ix4613 (.Y (nx4612), .A0 (nx6678), .A1 (nx11340), .A2 (nx11350)) ;
    nor02_2x ix6692 (.Y (nx6691), .A0 (nx4608), .A1 (nx4606)) ;
    nor03_2x ix4609 (.Y (nx4608), .A0 (nx6695), .A1 (nx10290), .A2 (nx11358)) ;
    dffr gen_11_cmp_mRegCmp_reg_Q_15 (.Q (gen_11_cmp_mReg_15), .QB (nx6695), .D (
         window_11__15), .CLK (start), .R (rst)) ;
    nor03_2x ix4607 (.Y (nx4606), .A0 (gen_11_cmp_mReg_15), .A1 (nx10800), .A2 (
             nx11366)) ;
    nand02 ix4631 (.Y (gen_11_cmp_BSCmp_op2_16), .A0 (nx6699), .A1 (nx6691)) ;
    nor02_2x ix6700 (.Y (nx6699), .A0 (nx4626), .A1 (nx4622)) ;
    nor03_2x ix4627 (.Y (nx4626), .A0 (gen_11_cmp_mReg_15), .A1 (nx10296), .A2 (
             nx11334)) ;
    nor03_2x ix4623 (.Y (nx4622), .A0 (nx6695), .A1 (nx11340), .A2 (nx11350)) ;
    nand02 ix4699 (.Y (gen_12_cmp_BSCmp_op2_1), .A0 (nx6707), .A1 (nx6727)) ;
    nor02_2x ix6708 (.Y (nx6707), .A0 (nx4694), .A1 (nx4690)) ;
    nor03_2x ix4695 (.Y (nx4694), .A0 (gen_12_cmp_mReg_0), .A1 (nx10280), .A2 (
             nx11370)) ;
    dffr gen_12_cmp_mRegCmp_reg_Q_0 (.Q (gen_12_cmp_mReg_0), .QB (nx6713), .D (
         window_12__0), .CLK (start), .R (rst)) ;
    inv01 ix6718 (.Y (nx6717), .A (gen_12_cmp_pMux_0)) ;
    nor03_2x ix4691 (.Y (nx4690), .A0 (nx6713), .A1 (nx11376), .A2 (nx11386)) ;
    inv02 ix6726 (.Y (nx6725), .A (gen_12_cmp_pMux_2)) ;
    nor02_2x ix6728 (.Y (nx6727), .A0 (nx4680), .A1 (nx4678)) ;
    nor03_2x ix4681 (.Y (nx4680), .A0 (nx6731), .A1 (nx10274), .A2 (nx11394)) ;
    dffr gen_12_cmp_mRegCmp_reg_Q_1 (.Q (gen_12_cmp_mReg_1), .QB (nx6731), .D (
         window_12__1), .CLK (start), .R (rst)) ;
    nor03_2x ix4679 (.Y (nx4678), .A0 (gen_12_cmp_mReg_1), .A1 (nx10802), .A2 (
             nx11402)) ;
    nor03_2x ix4639 (.Y (nx4638), .A0 (nx10280), .A1 (nx6725), .A2 (
             gen_12_cmp_pMux_0)) ;
    nand02 ix4721 (.Y (gen_12_cmp_BSCmp_op2_2), .A0 (nx6742), .A1 (nx6747)) ;
    nor02_2x ix6743 (.Y (nx6742), .A0 (nx4716), .A1 (nx4712)) ;
    nor03_2x ix4717 (.Y (nx4716), .A0 (gen_12_cmp_mReg_1), .A1 (nx10280), .A2 (
             nx11370)) ;
    nor03_2x ix4713 (.Y (nx4712), .A0 (nx6731), .A1 (nx11376), .A2 (nx11386)) ;
    nor02_2x ix6748 (.Y (nx6747), .A0 (nx4708), .A1 (nx4706)) ;
    nor03_2x ix4709 (.Y (nx4708), .A0 (nx6751), .A1 (nx10274), .A2 (nx11394)) ;
    dffr gen_12_cmp_mRegCmp_reg_Q_2 (.Q (gen_12_cmp_mReg_2), .QB (nx6751), .D (
         window_12__2), .CLK (start), .R (rst)) ;
    nor03_2x ix4707 (.Y (nx4706), .A0 (gen_12_cmp_mReg_2), .A1 (nx10802), .A2 (
             nx11402)) ;
    nand02 ix4743 (.Y (gen_12_cmp_BSCmp_op2_3), .A0 (nx6757), .A1 (nx6763)) ;
    nor02_2x ix6758 (.Y (nx6757), .A0 (nx4738), .A1 (nx4734)) ;
    nor03_2x ix4739 (.Y (nx4738), .A0 (gen_12_cmp_mReg_2), .A1 (nx10280), .A2 (
             nx11370)) ;
    nor03_2x ix4735 (.Y (nx4734), .A0 (nx6751), .A1 (nx11376), .A2 (nx11386)) ;
    nor02_2x ix6764 (.Y (nx6763), .A0 (nx4730), .A1 (nx4728)) ;
    nor03_2x ix4731 (.Y (nx4730), .A0 (nx6766), .A1 (nx10274), .A2 (nx11394)) ;
    dffr gen_12_cmp_mRegCmp_reg_Q_3 (.Q (gen_12_cmp_mReg_3), .QB (nx6766), .D (
         window_12__3), .CLK (start), .R (rst)) ;
    nor03_2x ix4729 (.Y (nx4728), .A0 (gen_12_cmp_mReg_3), .A1 (nx10802), .A2 (
             nx11402)) ;
    nand02 ix4765 (.Y (gen_12_cmp_BSCmp_op2_4), .A0 (nx6773), .A1 (nx6779)) ;
    nor02_2x ix6774 (.Y (nx6773), .A0 (nx4760), .A1 (nx4756)) ;
    nor03_2x ix4761 (.Y (nx4760), .A0 (gen_12_cmp_mReg_3), .A1 (nx10280), .A2 (
             nx11370)) ;
    nor03_2x ix4757 (.Y (nx4756), .A0 (nx6766), .A1 (nx11376), .A2 (nx11386)) ;
    nor02_2x ix6780 (.Y (nx6779), .A0 (nx4752), .A1 (nx4750)) ;
    nor03_2x ix4753 (.Y (nx4752), .A0 (nx6783), .A1 (nx10274), .A2 (nx11394)) ;
    dffr gen_12_cmp_mRegCmp_reg_Q_4 (.Q (gen_12_cmp_mReg_4), .QB (nx6783), .D (
         window_12__4), .CLK (start), .R (rst)) ;
    nor03_2x ix4751 (.Y (nx4750), .A0 (gen_12_cmp_mReg_4), .A1 (nx10802), .A2 (
             nx11402)) ;
    nand02 ix4787 (.Y (gen_12_cmp_BSCmp_op2_5), .A0 (nx6787), .A1 (nx6793)) ;
    nor02_2x ix6788 (.Y (nx6787), .A0 (nx4782), .A1 (nx4778)) ;
    nor03_2x ix4783 (.Y (nx4782), .A0 (gen_12_cmp_mReg_4), .A1 (nx10280), .A2 (
             nx11370)) ;
    nor03_2x ix4779 (.Y (nx4778), .A0 (nx6783), .A1 (nx11376), .A2 (nx11386)) ;
    nor02_2x ix6794 (.Y (nx6793), .A0 (nx4774), .A1 (nx4772)) ;
    nor03_2x ix4775 (.Y (nx4774), .A0 (nx6797), .A1 (nx10276), .A2 (nx11394)) ;
    dffr gen_12_cmp_mRegCmp_reg_Q_5 (.Q (gen_12_cmp_mReg_5), .QB (nx6797), .D (
         window_12__5), .CLK (start), .R (rst)) ;
    nor03_2x ix4773 (.Y (nx4772), .A0 (gen_12_cmp_mReg_5), .A1 (nx10802), .A2 (
             nx11402)) ;
    nand02 ix4809 (.Y (gen_12_cmp_BSCmp_op2_6), .A0 (nx6801), .A1 (nx6807)) ;
    nor02_2x ix6802 (.Y (nx6801), .A0 (nx4804), .A1 (nx4800)) ;
    nor03_2x ix4805 (.Y (nx4804), .A0 (gen_12_cmp_mReg_5), .A1 (nx10282), .A2 (
             nx11370)) ;
    nor03_2x ix4801 (.Y (nx4800), .A0 (nx6797), .A1 (nx11376), .A2 (nx11386)) ;
    nor02_2x ix6808 (.Y (nx6807), .A0 (nx4796), .A1 (nx4794)) ;
    nor03_2x ix4797 (.Y (nx4796), .A0 (nx6810), .A1 (nx10276), .A2 (nx11394)) ;
    dffr gen_12_cmp_mRegCmp_reg_Q_6 (.Q (gen_12_cmp_mReg_6), .QB (nx6810), .D (
         window_12__6), .CLK (start), .R (rst)) ;
    nor03_2x ix4795 (.Y (nx4794), .A0 (gen_12_cmp_mReg_6), .A1 (nx10802), .A2 (
             nx11402)) ;
    nand02 ix4831 (.Y (gen_12_cmp_BSCmp_op2_7), .A0 (nx6817), .A1 (nx6823)) ;
    nor02_2x ix6818 (.Y (nx6817), .A0 (nx4826), .A1 (nx4822)) ;
    nor03_2x ix4827 (.Y (nx4826), .A0 (gen_12_cmp_mReg_6), .A1 (nx10282), .A2 (
             nx11372)) ;
    nor03_2x ix4823 (.Y (nx4822), .A0 (nx6810), .A1 (nx11378), .A2 (nx11388)) ;
    nor02_2x ix6824 (.Y (nx6823), .A0 (nx4818), .A1 (nx4816)) ;
    nor03_2x ix4819 (.Y (nx4818), .A0 (nx6827), .A1 (nx10276), .A2 (nx11396)) ;
    dffr gen_12_cmp_mRegCmp_reg_Q_7 (.Q (gen_12_cmp_mReg_7), .QB (nx6827), .D (
         window_12__7), .CLK (start), .R (rst)) ;
    nor03_2x ix4817 (.Y (nx4816), .A0 (gen_12_cmp_mReg_7), .A1 (nx10802), .A2 (
             nx11404)) ;
    nand02 ix4853 (.Y (gen_12_cmp_BSCmp_op2_8), .A0 (nx6831), .A1 (nx6837)) ;
    nor02_2x ix6832 (.Y (nx6831), .A0 (nx4848), .A1 (nx4844)) ;
    nor03_2x ix4849 (.Y (nx4848), .A0 (gen_12_cmp_mReg_7), .A1 (nx10282), .A2 (
             nx11372)) ;
    nor03_2x ix4845 (.Y (nx4844), .A0 (nx6827), .A1 (nx11378), .A2 (nx11388)) ;
    nor02_2x ix6838 (.Y (nx6837), .A0 (nx4840), .A1 (nx4838)) ;
    nor03_2x ix4841 (.Y (nx4840), .A0 (nx6841), .A1 (nx10276), .A2 (nx11396)) ;
    dffr gen_12_cmp_mRegCmp_reg_Q_8 (.Q (gen_12_cmp_mReg_8), .QB (nx6841), .D (
         window_12__8), .CLK (start), .R (rst)) ;
    nor03_2x ix4839 (.Y (nx4838), .A0 (gen_12_cmp_mReg_8), .A1 (nx10804), .A2 (
             nx11404)) ;
    nand02 ix4875 (.Y (gen_12_cmp_BSCmp_op2_9), .A0 (nx6845), .A1 (nx6851)) ;
    nor02_2x ix6846 (.Y (nx6845), .A0 (nx4870), .A1 (nx4866)) ;
    nor03_2x ix4871 (.Y (nx4870), .A0 (gen_12_cmp_mReg_8), .A1 (nx10282), .A2 (
             nx11372)) ;
    nor03_2x ix4867 (.Y (nx4866), .A0 (nx6841), .A1 (nx11378), .A2 (nx11388)) ;
    nor02_2x ix6852 (.Y (nx6851), .A0 (nx4862), .A1 (nx4860)) ;
    nor03_2x ix4863 (.Y (nx4862), .A0 (nx6854), .A1 (nx10276), .A2 (nx11396)) ;
    dffr gen_12_cmp_mRegCmp_reg_Q_9 (.Q (gen_12_cmp_mReg_9), .QB (nx6854), .D (
         window_12__9), .CLK (start), .R (rst)) ;
    nor03_2x ix4861 (.Y (nx4860), .A0 (gen_12_cmp_mReg_9), .A1 (nx10804), .A2 (
             nx11404)) ;
    nand02 ix4897 (.Y (gen_12_cmp_BSCmp_op2_10), .A0 (nx6861), .A1 (nx6867)) ;
    nor02_2x ix6862 (.Y (nx6861), .A0 (nx4892), .A1 (nx4888)) ;
    nor03_2x ix4893 (.Y (nx4892), .A0 (gen_12_cmp_mReg_9), .A1 (nx10282), .A2 (
             nx11372)) ;
    nor03_2x ix4889 (.Y (nx4888), .A0 (nx6854), .A1 (nx11378), .A2 (nx11388)) ;
    nor02_2x ix6868 (.Y (nx6867), .A0 (nx4884), .A1 (nx4882)) ;
    nor03_2x ix4885 (.Y (nx4884), .A0 (nx6871), .A1 (nx10276), .A2 (nx11396)) ;
    dffr gen_12_cmp_mRegCmp_reg_Q_10 (.Q (gen_12_cmp_mReg_10), .QB (nx6871), .D (
         window_12__10), .CLK (start), .R (rst)) ;
    nor03_2x ix4883 (.Y (nx4882), .A0 (gen_12_cmp_mReg_10), .A1 (nx10804), .A2 (
             nx11404)) ;
    nand02 ix4919 (.Y (gen_12_cmp_BSCmp_op2_11), .A0 (nx6875), .A1 (nx6881)) ;
    nor02_2x ix6876 (.Y (nx6875), .A0 (nx4914), .A1 (nx4910)) ;
    nor03_2x ix4915 (.Y (nx4914), .A0 (gen_12_cmp_mReg_10), .A1 (nx10282), .A2 (
             nx11372)) ;
    nor03_2x ix4911 (.Y (nx4910), .A0 (nx6871), .A1 (nx11378), .A2 (nx11388)) ;
    nor02_2x ix6882 (.Y (nx6881), .A0 (nx4906), .A1 (nx4904)) ;
    nor03_2x ix4907 (.Y (nx4906), .A0 (nx6885), .A1 (nx10276), .A2 (nx11396)) ;
    dffr gen_12_cmp_mRegCmp_reg_Q_11 (.Q (gen_12_cmp_mReg_11), .QB (nx6885), .D (
         window_12__11), .CLK (start), .R (rst)) ;
    nor03_2x ix4905 (.Y (nx4904), .A0 (gen_12_cmp_mReg_11), .A1 (nx10804), .A2 (
             nx11404)) ;
    nand02 ix4941 (.Y (gen_12_cmp_BSCmp_op2_12), .A0 (nx6889), .A1 (nx6895)) ;
    nor02_2x ix6890 (.Y (nx6889), .A0 (nx4936), .A1 (nx4932)) ;
    nor03_2x ix4937 (.Y (nx4936), .A0 (gen_12_cmp_mReg_11), .A1 (nx10282), .A2 (
             nx11372)) ;
    nor03_2x ix4933 (.Y (nx4932), .A0 (nx6885), .A1 (nx11378), .A2 (nx11388)) ;
    nor02_2x ix6896 (.Y (nx6895), .A0 (nx4928), .A1 (nx4926)) ;
    nor03_2x ix4929 (.Y (nx4928), .A0 (nx6898), .A1 (nx10278), .A2 (nx11396)) ;
    dffr gen_12_cmp_mRegCmp_reg_Q_12 (.Q (gen_12_cmp_mReg_12), .QB (nx6898), .D (
         window_12__12), .CLK (start), .R (rst)) ;
    nor03_2x ix4927 (.Y (nx4926), .A0 (gen_12_cmp_mReg_12), .A1 (nx10804), .A2 (
             nx11404)) ;
    nand02 ix4963 (.Y (gen_12_cmp_BSCmp_op2_13), .A0 (nx6905), .A1 (nx6911)) ;
    nor02_2x ix6906 (.Y (nx6905), .A0 (nx4958), .A1 (nx4954)) ;
    nor03_2x ix4959 (.Y (nx4958), .A0 (gen_12_cmp_mReg_12), .A1 (nx10284), .A2 (
             nx11374)) ;
    nor03_2x ix4955 (.Y (nx4954), .A0 (nx6898), .A1 (nx11378), .A2 (nx11390)) ;
    nor02_2x ix6912 (.Y (nx6911), .A0 (nx4950), .A1 (nx4948)) ;
    nor03_2x ix4951 (.Y (nx4950), .A0 (nx6915), .A1 (nx10278), .A2 (nx11398)) ;
    dffr gen_12_cmp_mRegCmp_reg_Q_13 (.Q (gen_12_cmp_mReg_13), .QB (nx6915), .D (
         window_12__13), .CLK (start), .R (rst)) ;
    nor03_2x ix4949 (.Y (nx4948), .A0 (gen_12_cmp_mReg_13), .A1 (nx10804), .A2 (
             nx11406)) ;
    nand02 ix4985 (.Y (gen_12_cmp_BSCmp_op2_14), .A0 (nx6919), .A1 (nx6925)) ;
    nor02_2x ix6920 (.Y (nx6919), .A0 (nx4980), .A1 (nx4976)) ;
    nor03_2x ix4981 (.Y (nx4980), .A0 (gen_12_cmp_mReg_13), .A1 (nx10284), .A2 (
             nx11374)) ;
    nor03_2x ix4977 (.Y (nx4976), .A0 (nx6915), .A1 (nx11380), .A2 (nx11390)) ;
    nor02_2x ix6926 (.Y (nx6925), .A0 (nx4972), .A1 (nx4970)) ;
    nor03_2x ix4973 (.Y (nx4972), .A0 (nx6929), .A1 (nx10278), .A2 (nx11398)) ;
    dffr gen_12_cmp_mRegCmp_reg_Q_14 (.Q (gen_12_cmp_mReg_14), .QB (nx6929), .D (
         window_12__14), .CLK (start), .R (rst)) ;
    nor03_2x ix4971 (.Y (nx4970), .A0 (gen_12_cmp_mReg_14), .A1 (nx10804), .A2 (
             nx11406)) ;
    nand02 ix5007 (.Y (gen_12_cmp_BSCmp_op2_15), .A0 (nx6933), .A1 (nx6939)) ;
    nor02_2x ix6934 (.Y (nx6933), .A0 (nx5002), .A1 (nx4998)) ;
    nor03_2x ix5003 (.Y (nx5002), .A0 (gen_12_cmp_mReg_14), .A1 (nx10284), .A2 (
             nx11374)) ;
    nor03_2x ix4999 (.Y (nx4998), .A0 (nx6929), .A1 (nx11380), .A2 (nx11390)) ;
    nor02_2x ix6940 (.Y (nx6939), .A0 (nx4994), .A1 (nx4992)) ;
    nor03_2x ix4995 (.Y (nx4994), .A0 (nx6943), .A1 (nx10278), .A2 (nx11398)) ;
    dffr gen_12_cmp_mRegCmp_reg_Q_15 (.Q (gen_12_cmp_mReg_15), .QB (nx6943), .D (
         window_12__15), .CLK (start), .R (rst)) ;
    nor03_2x ix4993 (.Y (nx4992), .A0 (gen_12_cmp_mReg_15), .A1 (nx10806), .A2 (
             nx11406)) ;
    nand02 ix5017 (.Y (gen_12_cmp_BSCmp_op2_16), .A0 (nx6949), .A1 (nx6939)) ;
    nor02_2x ix6950 (.Y (nx6949), .A0 (nx5012), .A1 (nx5008)) ;
    nor03_2x ix5013 (.Y (nx5012), .A0 (gen_12_cmp_mReg_15), .A1 (nx10284), .A2 (
             nx11374)) ;
    nor03_2x ix5009 (.Y (nx5008), .A0 (nx6943), .A1 (nx11380), .A2 (nx11390)) ;
    nand02 ix5085 (.Y (gen_13_cmp_BSCmp_op2_1), .A0 (nx6957), .A1 (nx6975)) ;
    nor02_2x ix6958 (.Y (nx6957), .A0 (nx5080), .A1 (nx5076)) ;
    nor03_2x ix5081 (.Y (nx5080), .A0 (gen_13_cmp_mReg_0), .A1 (nx10268), .A2 (
             nx11410)) ;
    dffr gen_13_cmp_mRegCmp_reg_Q_0 (.Q (gen_13_cmp_mReg_0), .QB (nx6961), .D (
         window_13__0), .CLK (start), .R (rst)) ;
    inv01 ix6966 (.Y (nx6965), .A (gen_13_cmp_pMux_0)) ;
    nor03_2x ix5077 (.Y (nx5076), .A0 (nx6961), .A1 (nx11416), .A2 (nx11426)) ;
    inv02 ix6974 (.Y (nx6973), .A (gen_13_cmp_pMux_2)) ;
    nor02_2x ix6976 (.Y (nx6975), .A0 (nx5066), .A1 (nx5064)) ;
    nor03_2x ix5067 (.Y (nx5066), .A0 (nx6979), .A1 (nx10262), .A2 (nx11434)) ;
    dffr gen_13_cmp_mRegCmp_reg_Q_1 (.Q (gen_13_cmp_mReg_1), .QB (nx6979), .D (
         window_13__1), .CLK (start), .R (rst)) ;
    nor03_2x ix5065 (.Y (nx5064), .A0 (gen_13_cmp_mReg_1), .A1 (nx10808), .A2 (
             nx11442)) ;
    nor03_2x ix5025 (.Y (nx5024), .A0 (nx10268), .A1 (nx6973), .A2 (
             gen_13_cmp_pMux_0)) ;
    nand02 ix5107 (.Y (gen_13_cmp_BSCmp_op2_2), .A0 (nx6990), .A1 (nx6995)) ;
    nor02_2x ix6991 (.Y (nx6990), .A0 (nx5102), .A1 (nx5098)) ;
    nor03_2x ix5103 (.Y (nx5102), .A0 (gen_13_cmp_mReg_1), .A1 (nx10268), .A2 (
             nx11410)) ;
    nor03_2x ix5099 (.Y (nx5098), .A0 (nx6979), .A1 (nx11416), .A2 (nx11426)) ;
    nor02_2x ix6996 (.Y (nx6995), .A0 (nx5094), .A1 (nx5092)) ;
    nor03_2x ix5095 (.Y (nx5094), .A0 (nx6999), .A1 (nx10262), .A2 (nx11434)) ;
    dffr gen_13_cmp_mRegCmp_reg_Q_2 (.Q (gen_13_cmp_mReg_2), .QB (nx6999), .D (
         window_13__2), .CLK (start), .R (rst)) ;
    nor03_2x ix5093 (.Y (nx5092), .A0 (gen_13_cmp_mReg_2), .A1 (nx10808), .A2 (
             nx11442)) ;
    nand02 ix5129 (.Y (gen_13_cmp_BSCmp_op2_3), .A0 (nx7003), .A1 (nx7009)) ;
    nor02_2x ix7004 (.Y (nx7003), .A0 (nx5124), .A1 (nx5120)) ;
    nor03_2x ix5125 (.Y (nx5124), .A0 (gen_13_cmp_mReg_2), .A1 (nx10268), .A2 (
             nx11410)) ;
    nor03_2x ix5121 (.Y (nx5120), .A0 (nx6999), .A1 (nx11416), .A2 (nx11426)) ;
    nor02_2x ix7010 (.Y (nx7009), .A0 (nx5116), .A1 (nx5114)) ;
    nor03_2x ix5117 (.Y (nx5116), .A0 (nx7013), .A1 (nx10262), .A2 (nx11434)) ;
    dffr gen_13_cmp_mRegCmp_reg_Q_3 (.Q (gen_13_cmp_mReg_3), .QB (nx7013), .D (
         window_13__3), .CLK (start), .R (rst)) ;
    nor03_2x ix5115 (.Y (nx5114), .A0 (gen_13_cmp_mReg_3), .A1 (nx10808), .A2 (
             nx11442)) ;
    nand02 ix5151 (.Y (gen_13_cmp_BSCmp_op2_4), .A0 (nx7018), .A1 (nx7023)) ;
    nor02_2x ix7019 (.Y (nx7018), .A0 (nx5146), .A1 (nx5142)) ;
    nor03_2x ix5147 (.Y (nx5146), .A0 (gen_13_cmp_mReg_3), .A1 (nx10268), .A2 (
             nx11410)) ;
    nor03_2x ix5143 (.Y (nx5142), .A0 (nx7013), .A1 (nx11416), .A2 (nx11426)) ;
    nor02_2x ix7024 (.Y (nx7023), .A0 (nx5138), .A1 (nx5136)) ;
    nor03_2x ix5139 (.Y (nx5138), .A0 (nx7027), .A1 (nx10262), .A2 (nx11434)) ;
    dffr gen_13_cmp_mRegCmp_reg_Q_4 (.Q (gen_13_cmp_mReg_4), .QB (nx7027), .D (
         window_13__4), .CLK (start), .R (rst)) ;
    nor03_2x ix5137 (.Y (nx5136), .A0 (gen_13_cmp_mReg_4), .A1 (nx10808), .A2 (
             nx11442)) ;
    nand02 ix5173 (.Y (gen_13_cmp_BSCmp_op2_5), .A0 (nx7033), .A1 (nx7039)) ;
    nor02_2x ix7034 (.Y (nx7033), .A0 (nx5168), .A1 (nx5164)) ;
    nor03_2x ix5169 (.Y (nx5168), .A0 (gen_13_cmp_mReg_4), .A1 (nx10268), .A2 (
             nx11410)) ;
    nor03_2x ix5165 (.Y (nx5164), .A0 (nx7027), .A1 (nx11416), .A2 (nx11426)) ;
    nor02_2x ix7040 (.Y (nx7039), .A0 (nx5160), .A1 (nx5158)) ;
    nor03_2x ix5161 (.Y (nx5160), .A0 (nx7042), .A1 (nx10264), .A2 (nx11434)) ;
    dffr gen_13_cmp_mRegCmp_reg_Q_5 (.Q (gen_13_cmp_mReg_5), .QB (nx7042), .D (
         window_13__5), .CLK (start), .R (rst)) ;
    nor03_2x ix5159 (.Y (nx5158), .A0 (gen_13_cmp_mReg_5), .A1 (nx10808), .A2 (
             nx11442)) ;
    nand02 ix5195 (.Y (gen_13_cmp_BSCmp_op2_6), .A0 (nx7049), .A1 (nx7055)) ;
    nor02_2x ix7050 (.Y (nx7049), .A0 (nx5190), .A1 (nx5186)) ;
    nor03_2x ix5191 (.Y (nx5190), .A0 (gen_13_cmp_mReg_5), .A1 (nx10270), .A2 (
             nx11410)) ;
    nor03_2x ix5187 (.Y (nx5186), .A0 (nx7042), .A1 (nx11416), .A2 (nx11426)) ;
    nor02_2x ix7056 (.Y (nx7055), .A0 (nx5182), .A1 (nx5180)) ;
    nor03_2x ix5183 (.Y (nx5182), .A0 (nx7059), .A1 (nx10264), .A2 (nx11434)) ;
    dffr gen_13_cmp_mRegCmp_reg_Q_6 (.Q (gen_13_cmp_mReg_6), .QB (nx7059), .D (
         window_13__6), .CLK (start), .R (rst)) ;
    nor03_2x ix5181 (.Y (nx5180), .A0 (gen_13_cmp_mReg_6), .A1 (nx10808), .A2 (
             nx11442)) ;
    nand02 ix5217 (.Y (gen_13_cmp_BSCmp_op2_7), .A0 (nx7063), .A1 (nx7069)) ;
    nor02_2x ix7064 (.Y (nx7063), .A0 (nx5212), .A1 (nx5208)) ;
    nor03_2x ix5213 (.Y (nx5212), .A0 (gen_13_cmp_mReg_6), .A1 (nx10270), .A2 (
             nx11412)) ;
    nor03_2x ix5209 (.Y (nx5208), .A0 (nx7059), .A1 (nx11418), .A2 (nx11428)) ;
    nor02_2x ix7070 (.Y (nx7069), .A0 (nx5204), .A1 (nx5202)) ;
    nor03_2x ix5205 (.Y (nx5204), .A0 (nx7073), .A1 (nx10264), .A2 (nx11436)) ;
    dffr gen_13_cmp_mRegCmp_reg_Q_7 (.Q (gen_13_cmp_mReg_7), .QB (nx7073), .D (
         window_13__7), .CLK (start), .R (rst)) ;
    nor03_2x ix5203 (.Y (nx5202), .A0 (gen_13_cmp_mReg_7), .A1 (nx10808), .A2 (
             nx11444)) ;
    nand02 ix5239 (.Y (gen_13_cmp_BSCmp_op2_8), .A0 (nx7077), .A1 (nx7083)) ;
    nor02_2x ix7078 (.Y (nx7077), .A0 (nx5234), .A1 (nx5230)) ;
    nor03_2x ix5235 (.Y (nx5234), .A0 (gen_13_cmp_mReg_7), .A1 (nx10270), .A2 (
             nx11412)) ;
    nor03_2x ix5231 (.Y (nx5230), .A0 (nx7073), .A1 (nx11418), .A2 (nx11428)) ;
    nor02_2x ix7084 (.Y (nx7083), .A0 (nx5226), .A1 (nx5224)) ;
    nor03_2x ix5227 (.Y (nx5226), .A0 (nx7086), .A1 (nx10264), .A2 (nx11436)) ;
    dffr gen_13_cmp_mRegCmp_reg_Q_8 (.Q (gen_13_cmp_mReg_8), .QB (nx7086), .D (
         window_13__8), .CLK (start), .R (rst)) ;
    nor03_2x ix5225 (.Y (nx5224), .A0 (gen_13_cmp_mReg_8), .A1 (nx10810), .A2 (
             nx11444)) ;
    nand02 ix5261 (.Y (gen_13_cmp_BSCmp_op2_9), .A0 (nx7093), .A1 (nx7099)) ;
    nor02_2x ix7094 (.Y (nx7093), .A0 (nx5256), .A1 (nx5252)) ;
    nor03_2x ix5257 (.Y (nx5256), .A0 (gen_13_cmp_mReg_8), .A1 (nx10270), .A2 (
             nx11412)) ;
    nor03_2x ix5253 (.Y (nx5252), .A0 (nx7086), .A1 (nx11418), .A2 (nx11428)) ;
    nor02_2x ix7100 (.Y (nx7099), .A0 (nx5248), .A1 (nx5246)) ;
    nor03_2x ix5249 (.Y (nx5248), .A0 (nx7103), .A1 (nx10264), .A2 (nx11436)) ;
    dffr gen_13_cmp_mRegCmp_reg_Q_9 (.Q (gen_13_cmp_mReg_9), .QB (nx7103), .D (
         window_13__9), .CLK (start), .R (rst)) ;
    nor03_2x ix5247 (.Y (nx5246), .A0 (gen_13_cmp_mReg_9), .A1 (nx10810), .A2 (
             nx11444)) ;
    nand02 ix5283 (.Y (gen_13_cmp_BSCmp_op2_10), .A0 (nx7107), .A1 (nx7113)) ;
    nor02_2x ix7108 (.Y (nx7107), .A0 (nx5278), .A1 (nx5274)) ;
    nor03_2x ix5279 (.Y (nx5278), .A0 (gen_13_cmp_mReg_9), .A1 (nx10270), .A2 (
             nx11412)) ;
    nor03_2x ix5275 (.Y (nx5274), .A0 (nx7103), .A1 (nx11418), .A2 (nx11428)) ;
    nor02_2x ix7114 (.Y (nx7113), .A0 (nx5270), .A1 (nx5268)) ;
    nor03_2x ix5271 (.Y (nx5270), .A0 (nx7117), .A1 (nx10264), .A2 (nx11436)) ;
    dffr gen_13_cmp_mRegCmp_reg_Q_10 (.Q (gen_13_cmp_mReg_10), .QB (nx7117), .D (
         window_13__10), .CLK (start), .R (rst)) ;
    nor03_2x ix5269 (.Y (nx5268), .A0 (gen_13_cmp_mReg_10), .A1 (nx10810), .A2 (
             nx11444)) ;
    nand02 ix5305 (.Y (gen_13_cmp_BSCmp_op2_11), .A0 (nx7121), .A1 (nx7127)) ;
    nor02_2x ix7122 (.Y (nx7121), .A0 (nx5300), .A1 (nx5296)) ;
    nor03_2x ix5301 (.Y (nx5300), .A0 (gen_13_cmp_mReg_10), .A1 (nx10270), .A2 (
             nx11412)) ;
    nor03_2x ix5297 (.Y (nx5296), .A0 (nx7117), .A1 (nx11418), .A2 (nx11428)) ;
    nor02_2x ix7128 (.Y (nx7127), .A0 (nx5292), .A1 (nx5290)) ;
    nor03_2x ix5293 (.Y (nx5292), .A0 (nx7130), .A1 (nx10264), .A2 (nx11436)) ;
    dffr gen_13_cmp_mRegCmp_reg_Q_11 (.Q (gen_13_cmp_mReg_11), .QB (nx7130), .D (
         window_13__11), .CLK (start), .R (rst)) ;
    nor03_2x ix5291 (.Y (nx5290), .A0 (gen_13_cmp_mReg_11), .A1 (nx10810), .A2 (
             nx11444)) ;
    nand02 ix5327 (.Y (gen_13_cmp_BSCmp_op2_12), .A0 (nx7137), .A1 (nx7143)) ;
    nor02_2x ix7138 (.Y (nx7137), .A0 (nx5322), .A1 (nx5318)) ;
    nor03_2x ix5323 (.Y (nx5322), .A0 (gen_13_cmp_mReg_11), .A1 (nx10270), .A2 (
             nx11412)) ;
    nor03_2x ix5319 (.Y (nx5318), .A0 (nx7130), .A1 (nx11418), .A2 (nx11428)) ;
    nor02_2x ix7144 (.Y (nx7143), .A0 (nx5314), .A1 (nx5312)) ;
    nor03_2x ix5315 (.Y (nx5314), .A0 (nx7147), .A1 (nx10266), .A2 (nx11436)) ;
    dffr gen_13_cmp_mRegCmp_reg_Q_12 (.Q (gen_13_cmp_mReg_12), .QB (nx7147), .D (
         window_13__12), .CLK (start), .R (rst)) ;
    nor03_2x ix5313 (.Y (nx5312), .A0 (gen_13_cmp_mReg_12), .A1 (nx10810), .A2 (
             nx11444)) ;
    nand02 ix5349 (.Y (gen_13_cmp_BSCmp_op2_13), .A0 (nx7151), .A1 (nx7157)) ;
    nor02_2x ix7152 (.Y (nx7151), .A0 (nx5344), .A1 (nx5340)) ;
    nor03_2x ix5345 (.Y (nx5344), .A0 (gen_13_cmp_mReg_12), .A1 (nx10272), .A2 (
             nx11414)) ;
    nor03_2x ix5341 (.Y (nx5340), .A0 (nx7147), .A1 (nx11418), .A2 (nx11430)) ;
    nor02_2x ix7158 (.Y (nx7157), .A0 (nx5336), .A1 (nx5334)) ;
    nor03_2x ix5337 (.Y (nx5336), .A0 (nx7161), .A1 (nx10266), .A2 (nx11438)) ;
    dffr gen_13_cmp_mRegCmp_reg_Q_13 (.Q (gen_13_cmp_mReg_13), .QB (nx7161), .D (
         window_13__13), .CLK (start), .R (rst)) ;
    nor03_2x ix5335 (.Y (nx5334), .A0 (gen_13_cmp_mReg_13), .A1 (nx10810), .A2 (
             nx11446)) ;
    nand02 ix5371 (.Y (gen_13_cmp_BSCmp_op2_14), .A0 (nx7165), .A1 (nx7171)) ;
    nor02_2x ix7166 (.Y (nx7165), .A0 (nx5366), .A1 (nx5362)) ;
    nor03_2x ix5367 (.Y (nx5366), .A0 (gen_13_cmp_mReg_13), .A1 (nx10272), .A2 (
             nx11414)) ;
    nor03_2x ix5363 (.Y (nx5362), .A0 (nx7161), .A1 (nx11420), .A2 (nx11430)) ;
    nor02_2x ix7172 (.Y (nx7171), .A0 (nx5358), .A1 (nx5356)) ;
    nor03_2x ix5359 (.Y (nx5358), .A0 (nx7174), .A1 (nx10266), .A2 (nx11438)) ;
    dffr gen_13_cmp_mRegCmp_reg_Q_14 (.Q (gen_13_cmp_mReg_14), .QB (nx7174), .D (
         window_13__14), .CLK (start), .R (rst)) ;
    nor03_2x ix5357 (.Y (nx5356), .A0 (gen_13_cmp_mReg_14), .A1 (nx10810), .A2 (
             nx11446)) ;
    nand02 ix5393 (.Y (gen_13_cmp_BSCmp_op2_15), .A0 (nx7181), .A1 (nx7187)) ;
    nor02_2x ix7182 (.Y (nx7181), .A0 (nx5388), .A1 (nx5384)) ;
    nor03_2x ix5389 (.Y (nx5388), .A0 (gen_13_cmp_mReg_14), .A1 (nx10272), .A2 (
             nx11414)) ;
    nor03_2x ix5385 (.Y (nx5384), .A0 (nx7174), .A1 (nx11420), .A2 (nx11430)) ;
    nor02_2x ix7188 (.Y (nx7187), .A0 (nx5380), .A1 (nx5378)) ;
    nor03_2x ix5381 (.Y (nx5380), .A0 (nx7191), .A1 (nx10266), .A2 (nx11438)) ;
    dffr gen_13_cmp_mRegCmp_reg_Q_15 (.Q (gen_13_cmp_mReg_15), .QB (nx7191), .D (
         window_13__15), .CLK (start), .R (rst)) ;
    nor03_2x ix5379 (.Y (nx5378), .A0 (gen_13_cmp_mReg_15), .A1 (nx10812), .A2 (
             nx11446)) ;
    nand02 ix5403 (.Y (gen_13_cmp_BSCmp_op2_16), .A0 (nx7195), .A1 (nx7187)) ;
    nor02_2x ix7196 (.Y (nx7195), .A0 (nx5398), .A1 (nx5394)) ;
    nor03_2x ix5399 (.Y (nx5398), .A0 (gen_13_cmp_mReg_15), .A1 (nx10272), .A2 (
             nx11414)) ;
    nor03_2x ix5395 (.Y (nx5394), .A0 (nx7191), .A1 (nx11420), .A2 (nx11430)) ;
    nand02 ix5471 (.Y (gen_14_cmp_BSCmp_op2_1), .A0 (nx7203), .A1 (nx7223)) ;
    nor02_2x ix7204 (.Y (nx7203), .A0 (nx5466), .A1 (nx5462)) ;
    nor03_2x ix5467 (.Y (nx5466), .A0 (gen_14_cmp_mReg_0), .A1 (nx10256), .A2 (
             nx11450)) ;
    dffr gen_14_cmp_mRegCmp_reg_Q_0 (.Q (gen_14_cmp_mReg_0), .QB (nx7209), .D (
         window_14__0), .CLK (start), .R (rst)) ;
    inv01 ix7214 (.Y (nx7213), .A (gen_14_cmp_pMux_0)) ;
    nor03_2x ix5463 (.Y (nx5462), .A0 (nx7209), .A1 (nx11456), .A2 (nx11466)) ;
    inv02 ix7222 (.Y (nx7221), .A (gen_14_cmp_pMux_2)) ;
    nor02_2x ix7224 (.Y (nx7223), .A0 (nx5452), .A1 (nx5450)) ;
    nor03_2x ix5453 (.Y (nx5452), .A0 (nx7227), .A1 (nx10250), .A2 (nx11474)) ;
    dffr gen_14_cmp_mRegCmp_reg_Q_1 (.Q (gen_14_cmp_mReg_1), .QB (nx7227), .D (
         window_14__1), .CLK (start), .R (rst)) ;
    nor03_2x ix5451 (.Y (nx5450), .A0 (gen_14_cmp_mReg_1), .A1 (nx10814), .A2 (
             nx11482)) ;
    nor03_2x ix5411 (.Y (nx5410), .A0 (nx10256), .A1 (nx7221), .A2 (
             gen_14_cmp_pMux_0)) ;
    nand02 ix5493 (.Y (gen_14_cmp_BSCmp_op2_2), .A0 (nx7238), .A1 (nx7243)) ;
    nor02_2x ix7239 (.Y (nx7238), .A0 (nx5488), .A1 (nx5484)) ;
    nor03_2x ix5489 (.Y (nx5488), .A0 (gen_14_cmp_mReg_1), .A1 (nx10256), .A2 (
             nx11450)) ;
    nor03_2x ix5485 (.Y (nx5484), .A0 (nx7227), .A1 (nx11456), .A2 (nx11466)) ;
    nor02_2x ix7244 (.Y (nx7243), .A0 (nx5480), .A1 (nx5478)) ;
    nor03_2x ix5481 (.Y (nx5480), .A0 (nx7247), .A1 (nx10250), .A2 (nx11474)) ;
    dffr gen_14_cmp_mRegCmp_reg_Q_2 (.Q (gen_14_cmp_mReg_2), .QB (nx7247), .D (
         window_14__2), .CLK (start), .R (rst)) ;
    nor03_2x ix5479 (.Y (nx5478), .A0 (gen_14_cmp_mReg_2), .A1 (nx10814), .A2 (
             nx11482)) ;
    nand02 ix5515 (.Y (gen_14_cmp_BSCmp_op2_3), .A0 (nx7253), .A1 (nx7259)) ;
    nor02_2x ix7254 (.Y (nx7253), .A0 (nx5510), .A1 (nx5506)) ;
    nor03_2x ix5511 (.Y (nx5510), .A0 (gen_14_cmp_mReg_2), .A1 (nx10256), .A2 (
             nx11450)) ;
    nor03_2x ix5507 (.Y (nx5506), .A0 (nx7247), .A1 (nx11456), .A2 (nx11466)) ;
    nor02_2x ix7260 (.Y (nx7259), .A0 (nx5502), .A1 (nx5500)) ;
    nor03_2x ix5503 (.Y (nx5502), .A0 (nx7262), .A1 (nx10250), .A2 (nx11474)) ;
    dffr gen_14_cmp_mRegCmp_reg_Q_3 (.Q (gen_14_cmp_mReg_3), .QB (nx7262), .D (
         window_14__3), .CLK (start), .R (rst)) ;
    nor03_2x ix5501 (.Y (nx5500), .A0 (gen_14_cmp_mReg_3), .A1 (nx10814), .A2 (
             nx11482)) ;
    nand02 ix5537 (.Y (gen_14_cmp_BSCmp_op2_4), .A0 (nx7269), .A1 (nx7275)) ;
    nor02_2x ix7270 (.Y (nx7269), .A0 (nx5532), .A1 (nx5528)) ;
    nor03_2x ix5533 (.Y (nx5532), .A0 (gen_14_cmp_mReg_3), .A1 (nx10256), .A2 (
             nx11450)) ;
    nor03_2x ix5529 (.Y (nx5528), .A0 (nx7262), .A1 (nx11456), .A2 (nx11466)) ;
    nor02_2x ix7276 (.Y (nx7275), .A0 (nx5524), .A1 (nx5522)) ;
    nor03_2x ix5525 (.Y (nx5524), .A0 (nx7279), .A1 (nx10250), .A2 (nx11474)) ;
    dffr gen_14_cmp_mRegCmp_reg_Q_4 (.Q (gen_14_cmp_mReg_4), .QB (nx7279), .D (
         window_14__4), .CLK (start), .R (rst)) ;
    nor03_2x ix5523 (.Y (nx5522), .A0 (gen_14_cmp_mReg_4), .A1 (nx10814), .A2 (
             nx11482)) ;
    nand02 ix5559 (.Y (gen_14_cmp_BSCmp_op2_5), .A0 (nx7283), .A1 (nx7289)) ;
    nor02_2x ix7284 (.Y (nx7283), .A0 (nx5554), .A1 (nx5550)) ;
    nor03_2x ix5555 (.Y (nx5554), .A0 (gen_14_cmp_mReg_4), .A1 (nx10256), .A2 (
             nx11450)) ;
    nor03_2x ix5551 (.Y (nx5550), .A0 (nx7279), .A1 (nx11456), .A2 (nx11466)) ;
    nor02_2x ix7290 (.Y (nx7289), .A0 (nx5546), .A1 (nx5544)) ;
    nor03_2x ix5547 (.Y (nx5546), .A0 (nx7293), .A1 (nx10252), .A2 (nx11474)) ;
    dffr gen_14_cmp_mRegCmp_reg_Q_5 (.Q (gen_14_cmp_mReg_5), .QB (nx7293), .D (
         window_14__5), .CLK (start), .R (rst)) ;
    nor03_2x ix5545 (.Y (nx5544), .A0 (gen_14_cmp_mReg_5), .A1 (nx10814), .A2 (
             nx11482)) ;
    nand02 ix5581 (.Y (gen_14_cmp_BSCmp_op2_6), .A0 (nx7297), .A1 (nx7303)) ;
    nor02_2x ix7298 (.Y (nx7297), .A0 (nx5576), .A1 (nx5572)) ;
    nor03_2x ix5577 (.Y (nx5576), .A0 (gen_14_cmp_mReg_5), .A1 (nx10258), .A2 (
             nx11450)) ;
    nor03_2x ix5573 (.Y (nx5572), .A0 (nx7293), .A1 (nx11456), .A2 (nx11466)) ;
    nor02_2x ix7304 (.Y (nx7303), .A0 (nx5568), .A1 (nx5566)) ;
    nor03_2x ix5569 (.Y (nx5568), .A0 (nx7306), .A1 (nx10252), .A2 (nx11474)) ;
    dffr gen_14_cmp_mRegCmp_reg_Q_6 (.Q (gen_14_cmp_mReg_6), .QB (nx7306), .D (
         window_14__6), .CLK (start), .R (rst)) ;
    nor03_2x ix5567 (.Y (nx5566), .A0 (gen_14_cmp_mReg_6), .A1 (nx10814), .A2 (
             nx11482)) ;
    nand02 ix5603 (.Y (gen_14_cmp_BSCmp_op2_7), .A0 (nx7313), .A1 (nx7319)) ;
    nor02_2x ix7314 (.Y (nx7313), .A0 (nx5598), .A1 (nx5594)) ;
    nor03_2x ix5599 (.Y (nx5598), .A0 (gen_14_cmp_mReg_6), .A1 (nx10258), .A2 (
             nx11452)) ;
    nor03_2x ix5595 (.Y (nx5594), .A0 (nx7306), .A1 (nx11458), .A2 (nx11468)) ;
    nor02_2x ix7320 (.Y (nx7319), .A0 (nx5590), .A1 (nx5588)) ;
    nor03_2x ix5591 (.Y (nx5590), .A0 (nx7323), .A1 (nx10252), .A2 (nx11476)) ;
    dffr gen_14_cmp_mRegCmp_reg_Q_7 (.Q (gen_14_cmp_mReg_7), .QB (nx7323), .D (
         window_14__7), .CLK (start), .R (rst)) ;
    nor03_2x ix5589 (.Y (nx5588), .A0 (gen_14_cmp_mReg_7), .A1 (nx10814), .A2 (
             nx11484)) ;
    nand02 ix5625 (.Y (gen_14_cmp_BSCmp_op2_8), .A0 (nx7329), .A1 (nx7335)) ;
    nor02_2x ix7330 (.Y (nx7329), .A0 (nx5620), .A1 (nx5616)) ;
    nor03_2x ix5621 (.Y (nx5620), .A0 (gen_14_cmp_mReg_7), .A1 (nx10258), .A2 (
             nx11452)) ;
    nor03_2x ix5617 (.Y (nx5616), .A0 (nx7323), .A1 (nx11458), .A2 (nx11468)) ;
    nor02_2x ix7336 (.Y (nx7335), .A0 (nx5612), .A1 (nx5610)) ;
    nor03_2x ix5613 (.Y (nx5612), .A0 (nx7339), .A1 (nx10252), .A2 (nx11476)) ;
    dffr gen_14_cmp_mRegCmp_reg_Q_8 (.Q (gen_14_cmp_mReg_8), .QB (nx7339), .D (
         window_14__8), .CLK (start), .R (rst)) ;
    nor03_2x ix5611 (.Y (nx5610), .A0 (gen_14_cmp_mReg_8), .A1 (nx10816), .A2 (
             nx11484)) ;
    nand02 ix5647 (.Y (gen_14_cmp_BSCmp_op2_9), .A0 (nx7344), .A1 (nx7348)) ;
    nor02_2x ix7345 (.Y (nx7344), .A0 (nx5642), .A1 (nx5638)) ;
    nor03_2x ix5643 (.Y (nx5642), .A0 (gen_14_cmp_mReg_8), .A1 (nx10258), .A2 (
             nx11452)) ;
    nor03_2x ix5639 (.Y (nx5638), .A0 (nx7339), .A1 (nx11458), .A2 (nx11468)) ;
    nor02_2x ix7349 (.Y (nx7348), .A0 (nx5634), .A1 (nx5632)) ;
    nor03_2x ix5635 (.Y (nx5634), .A0 (nx7351), .A1 (nx10252), .A2 (nx11476)) ;
    dffr gen_14_cmp_mRegCmp_reg_Q_9 (.Q (gen_14_cmp_mReg_9), .QB (nx7351), .D (
         window_14__9), .CLK (start), .R (rst)) ;
    nor03_2x ix5633 (.Y (nx5632), .A0 (gen_14_cmp_mReg_9), .A1 (nx10816), .A2 (
             nx11484)) ;
    nand02 ix5669 (.Y (gen_14_cmp_BSCmp_op2_10), .A0 (nx7357), .A1 (nx7363)) ;
    nor02_2x ix7358 (.Y (nx7357), .A0 (nx5664), .A1 (nx5660)) ;
    nor03_2x ix5665 (.Y (nx5664), .A0 (gen_14_cmp_mReg_9), .A1 (nx10258), .A2 (
             nx11452)) ;
    nor03_2x ix5661 (.Y (nx5660), .A0 (nx7351), .A1 (nx11458), .A2 (nx11468)) ;
    nor02_2x ix7364 (.Y (nx7363), .A0 (nx5656), .A1 (nx5654)) ;
    nor03_2x ix5657 (.Y (nx5656), .A0 (nx7367), .A1 (nx10252), .A2 (nx11476)) ;
    dffr gen_14_cmp_mRegCmp_reg_Q_10 (.Q (gen_14_cmp_mReg_10), .QB (nx7367), .D (
         window_14__10), .CLK (start), .R (rst)) ;
    nor03_2x ix5655 (.Y (nx5654), .A0 (gen_14_cmp_mReg_10), .A1 (nx10816), .A2 (
             nx11484)) ;
    nand02 ix5691 (.Y (gen_14_cmp_BSCmp_op2_11), .A0 (nx7373), .A1 (nx7377)) ;
    nor02_2x ix7374 (.Y (nx7373), .A0 (nx5686), .A1 (nx5682)) ;
    nor03_2x ix5687 (.Y (nx5686), .A0 (gen_14_cmp_mReg_10), .A1 (nx10258), .A2 (
             nx11452)) ;
    nor03_2x ix5683 (.Y (nx5682), .A0 (nx7367), .A1 (nx11458), .A2 (nx11468)) ;
    nor02_2x ix7378 (.Y (nx7377), .A0 (nx5678), .A1 (nx5676)) ;
    nor03_2x ix5679 (.Y (nx5678), .A0 (nx7381), .A1 (nx10252), .A2 (nx11476)) ;
    dffr gen_14_cmp_mRegCmp_reg_Q_11 (.Q (gen_14_cmp_mReg_11), .QB (nx7381), .D (
         window_14__11), .CLK (start), .R (rst)) ;
    nor03_2x ix5677 (.Y (nx5676), .A0 (gen_14_cmp_mReg_11), .A1 (nx10816), .A2 (
             nx11484)) ;
    nand02 ix5713 (.Y (gen_14_cmp_BSCmp_op2_12), .A0 (nx7387), .A1 (nx7393)) ;
    nor02_2x ix7388 (.Y (nx7387), .A0 (nx5708), .A1 (nx5704)) ;
    nor03_2x ix5709 (.Y (nx5708), .A0 (gen_14_cmp_mReg_11), .A1 (nx10258), .A2 (
             nx11452)) ;
    nor03_2x ix5705 (.Y (nx5704), .A0 (nx7381), .A1 (nx11458), .A2 (nx11468)) ;
    nor02_2x ix7394 (.Y (nx7393), .A0 (nx5700), .A1 (nx5698)) ;
    nor03_2x ix5701 (.Y (nx5700), .A0 (nx7397), .A1 (nx10254), .A2 (nx11476)) ;
    dffr gen_14_cmp_mRegCmp_reg_Q_12 (.Q (gen_14_cmp_mReg_12), .QB (nx7397), .D (
         window_14__12), .CLK (start), .R (rst)) ;
    nor03_2x ix5699 (.Y (nx5698), .A0 (gen_14_cmp_mReg_12), .A1 (nx10816), .A2 (
             nx11484)) ;
    nand02 ix5735 (.Y (gen_14_cmp_BSCmp_op2_13), .A0 (nx7403), .A1 (nx7407)) ;
    nor02_2x ix7404 (.Y (nx7403), .A0 (nx5730), .A1 (nx5726)) ;
    nor03_2x ix5731 (.Y (nx5730), .A0 (gen_14_cmp_mReg_12), .A1 (nx10260), .A2 (
             nx11454)) ;
    nor03_2x ix5727 (.Y (nx5726), .A0 (nx7397), .A1 (nx11458), .A2 (nx11470)) ;
    nor02_2x ix7408 (.Y (nx7407), .A0 (nx5722), .A1 (nx5720)) ;
    nor03_2x ix5723 (.Y (nx5722), .A0 (nx7411), .A1 (nx10254), .A2 (nx11478)) ;
    dffr gen_14_cmp_mRegCmp_reg_Q_13 (.Q (gen_14_cmp_mReg_13), .QB (nx7411), .D (
         window_14__13), .CLK (start), .R (rst)) ;
    nor03_2x ix5721 (.Y (nx5720), .A0 (gen_14_cmp_mReg_13), .A1 (nx10816), .A2 (
             nx11486)) ;
    nand02 ix5757 (.Y (gen_14_cmp_BSCmp_op2_14), .A0 (nx7417), .A1 (nx7423)) ;
    nor02_2x ix7418 (.Y (nx7417), .A0 (nx5752), .A1 (nx5748)) ;
    nor03_2x ix5753 (.Y (nx5752), .A0 (gen_14_cmp_mReg_13), .A1 (nx10260), .A2 (
             nx11454)) ;
    nor03_2x ix5749 (.Y (nx5748), .A0 (nx7411), .A1 (nx11460), .A2 (nx11470)) ;
    nor02_2x ix7424 (.Y (nx7423), .A0 (nx5744), .A1 (nx5742)) ;
    nor03_2x ix5745 (.Y (nx5744), .A0 (nx7426), .A1 (nx10254), .A2 (nx11478)) ;
    dffr gen_14_cmp_mRegCmp_reg_Q_14 (.Q (gen_14_cmp_mReg_14), .QB (nx7426), .D (
         window_14__14), .CLK (start), .R (rst)) ;
    nor03_2x ix5743 (.Y (nx5742), .A0 (gen_14_cmp_mReg_14), .A1 (nx10816), .A2 (
             nx11486)) ;
    nand02 ix5779 (.Y (gen_14_cmp_BSCmp_op2_15), .A0 (nx7431), .A1 (nx7437)) ;
    nor02_2x ix7432 (.Y (nx7431), .A0 (nx5774), .A1 (nx5770)) ;
    nor03_2x ix5775 (.Y (nx5774), .A0 (gen_14_cmp_mReg_14), .A1 (nx10260), .A2 (
             nx11454)) ;
    nor03_2x ix5771 (.Y (nx5770), .A0 (nx7426), .A1 (nx11460), .A2 (nx11470)) ;
    nor02_2x ix7438 (.Y (nx7437), .A0 (nx5766), .A1 (nx5764)) ;
    nor03_2x ix5767 (.Y (nx5766), .A0 (nx7441), .A1 (nx10254), .A2 (nx11478)) ;
    dffr gen_14_cmp_mRegCmp_reg_Q_15 (.Q (gen_14_cmp_mReg_15), .QB (nx7441), .D (
         window_14__15), .CLK (start), .R (rst)) ;
    nor03_2x ix5765 (.Y (nx5764), .A0 (gen_14_cmp_mReg_15), .A1 (nx10818), .A2 (
             nx11486)) ;
    nand02 ix5789 (.Y (gen_14_cmp_BSCmp_op2_16), .A0 (nx7447), .A1 (nx7437)) ;
    nor02_2x ix7448 (.Y (nx7447), .A0 (nx5784), .A1 (nx5780)) ;
    nor03_2x ix5785 (.Y (nx5784), .A0 (gen_14_cmp_mReg_15), .A1 (nx10260), .A2 (
             nx11454)) ;
    nor03_2x ix5781 (.Y (nx5780), .A0 (nx7441), .A1 (nx11460), .A2 (nx11470)) ;
    nand02 ix5857 (.Y (gen_15_cmp_BSCmp_op2_1), .A0 (nx7453), .A1 (nx7473)) ;
    nor02_2x ix7454 (.Y (nx7453), .A0 (nx5852), .A1 (nx5848)) ;
    nor03_2x ix5853 (.Y (nx5852), .A0 (gen_15_cmp_mReg_0), .A1 (nx10244), .A2 (
             nx11490)) ;
    dffr gen_15_cmp_mRegCmp_reg_Q_0 (.Q (gen_15_cmp_mReg_0), .QB (nx7459), .D (
         window_15__0), .CLK (start), .R (rst)) ;
    inv01 ix7464 (.Y (nx7463), .A (gen_15_cmp_pMux_0)) ;
    nor03_2x ix5849 (.Y (nx5848), .A0 (nx7459), .A1 (nx11496), .A2 (nx11506)) ;
    inv02 ix7472 (.Y (nx7471), .A (gen_15_cmp_pMux_2)) ;
    nor02_2x ix7474 (.Y (nx7473), .A0 (nx5838), .A1 (nx5836)) ;
    nor03_2x ix5839 (.Y (nx5838), .A0 (nx7477), .A1 (nx10238), .A2 (nx11514)) ;
    dffr gen_15_cmp_mRegCmp_reg_Q_1 (.Q (gen_15_cmp_mReg_1), .QB (nx7477), .D (
         window_15__1), .CLK (start), .R (rst)) ;
    nor03_2x ix5837 (.Y (nx5836), .A0 (gen_15_cmp_mReg_1), .A1 (nx10820), .A2 (
             nx11522)) ;
    nor03_2x ix5797 (.Y (nx5796), .A0 (nx10244), .A1 (nx7471), .A2 (
             gen_15_cmp_pMux_0)) ;
    nand02 ix5879 (.Y (gen_15_cmp_BSCmp_op2_2), .A0 (nx7489), .A1 (nx7493)) ;
    nor02_2x ix7490 (.Y (nx7489), .A0 (nx5874), .A1 (nx5870)) ;
    nor03_2x ix5875 (.Y (nx5874), .A0 (gen_15_cmp_mReg_1), .A1 (nx10244), .A2 (
             nx11490)) ;
    nor03_2x ix5871 (.Y (nx5870), .A0 (nx7477), .A1 (nx11496), .A2 (nx11506)) ;
    nor02_2x ix7494 (.Y (nx7493), .A0 (nx5866), .A1 (nx5864)) ;
    nor03_2x ix5867 (.Y (nx5866), .A0 (nx7497), .A1 (nx10238), .A2 (nx11514)) ;
    dffr gen_15_cmp_mRegCmp_reg_Q_2 (.Q (gen_15_cmp_mReg_2), .QB (nx7497), .D (
         window_15__2), .CLK (start), .R (rst)) ;
    nor03_2x ix5865 (.Y (nx5864), .A0 (gen_15_cmp_mReg_2), .A1 (nx10820), .A2 (
             nx11522)) ;
    nand02 ix5901 (.Y (gen_15_cmp_BSCmp_op2_3), .A0 (nx7503), .A1 (nx7507)) ;
    nor02_2x ix7504 (.Y (nx7503), .A0 (nx5896), .A1 (nx5892)) ;
    nor03_2x ix5897 (.Y (nx5896), .A0 (gen_15_cmp_mReg_2), .A1 (nx10244), .A2 (
             nx11490)) ;
    nor03_2x ix5893 (.Y (nx5892), .A0 (nx7497), .A1 (nx11496), .A2 (nx11506)) ;
    nor02_2x ix7508 (.Y (nx7507), .A0 (nx5888), .A1 (nx5886)) ;
    nor03_2x ix5889 (.Y (nx5888), .A0 (nx7511), .A1 (nx10238), .A2 (nx11514)) ;
    dffr gen_15_cmp_mRegCmp_reg_Q_3 (.Q (gen_15_cmp_mReg_3), .QB (nx7511), .D (
         window_15__3), .CLK (start), .R (rst)) ;
    nor03_2x ix5887 (.Y (nx5886), .A0 (gen_15_cmp_mReg_3), .A1 (nx10820), .A2 (
             nx11522)) ;
    nand02 ix5923 (.Y (gen_15_cmp_BSCmp_op2_4), .A0 (nx7515), .A1 (nx7521)) ;
    nor02_2x ix7516 (.Y (nx7515), .A0 (nx5918), .A1 (nx5914)) ;
    nor03_2x ix5919 (.Y (nx5918), .A0 (gen_15_cmp_mReg_3), .A1 (nx10244), .A2 (
             nx11490)) ;
    nor03_2x ix5915 (.Y (nx5914), .A0 (nx7511), .A1 (nx11496), .A2 (nx11506)) ;
    nor02_2x ix7522 (.Y (nx7521), .A0 (nx5910), .A1 (nx5908)) ;
    nor03_2x ix5911 (.Y (nx5910), .A0 (nx7525), .A1 (nx10238), .A2 (nx11514)) ;
    dffr gen_15_cmp_mRegCmp_reg_Q_4 (.Q (gen_15_cmp_mReg_4), .QB (nx7525), .D (
         window_15__4), .CLK (start), .R (rst)) ;
    nor03_2x ix5909 (.Y (nx5908), .A0 (gen_15_cmp_mReg_4), .A1 (nx10820), .A2 (
             nx11522)) ;
    nand02 ix5945 (.Y (gen_15_cmp_BSCmp_op2_5), .A0 (nx7529), .A1 (nx7535)) ;
    nor02_2x ix7530 (.Y (nx7529), .A0 (nx5940), .A1 (nx5936)) ;
    nor03_2x ix5941 (.Y (nx5940), .A0 (gen_15_cmp_mReg_4), .A1 (nx10244), .A2 (
             nx11490)) ;
    nor03_2x ix5937 (.Y (nx5936), .A0 (nx7525), .A1 (nx11496), .A2 (nx11506)) ;
    nor02_2x ix7536 (.Y (nx7535), .A0 (nx5932), .A1 (nx5930)) ;
    nor03_2x ix5933 (.Y (nx5932), .A0 (nx7538), .A1 (nx10240), .A2 (nx11514)) ;
    dffr gen_15_cmp_mRegCmp_reg_Q_5 (.Q (gen_15_cmp_mReg_5), .QB (nx7538), .D (
         window_15__5), .CLK (start), .R (rst)) ;
    nor03_2x ix5931 (.Y (nx5930), .A0 (gen_15_cmp_mReg_5), .A1 (nx10820), .A2 (
             nx11522)) ;
    nand02 ix5967 (.Y (gen_15_cmp_BSCmp_op2_6), .A0 (nx7545), .A1 (nx7551)) ;
    nor02_2x ix7546 (.Y (nx7545), .A0 (nx5962), .A1 (nx5958)) ;
    nor03_2x ix5963 (.Y (nx5962), .A0 (gen_15_cmp_mReg_5), .A1 (nx10246), .A2 (
             nx11490)) ;
    nor03_2x ix5959 (.Y (nx5958), .A0 (nx7538), .A1 (nx11496), .A2 (nx11506)) ;
    nor02_2x ix7552 (.Y (nx7551), .A0 (nx5954), .A1 (nx5952)) ;
    nor03_2x ix5955 (.Y (nx5954), .A0 (nx7555), .A1 (nx10240), .A2 (nx11514)) ;
    dffr gen_15_cmp_mRegCmp_reg_Q_6 (.Q (gen_15_cmp_mReg_6), .QB (nx7555), .D (
         window_15__6), .CLK (start), .R (rst)) ;
    nor03_2x ix5953 (.Y (nx5952), .A0 (gen_15_cmp_mReg_6), .A1 (nx10820), .A2 (
             nx11522)) ;
    nand02 ix5989 (.Y (gen_15_cmp_BSCmp_op2_7), .A0 (nx7559), .A1 (nx7565)) ;
    nor02_2x ix7560 (.Y (nx7559), .A0 (nx5984), .A1 (nx5980)) ;
    nor03_2x ix5985 (.Y (nx5984), .A0 (gen_15_cmp_mReg_6), .A1 (nx10246), .A2 (
             nx11492)) ;
    nor03_2x ix5981 (.Y (nx5980), .A0 (nx7555), .A1 (nx11498), .A2 (nx11508)) ;
    nor02_2x ix7566 (.Y (nx7565), .A0 (nx5976), .A1 (nx5974)) ;
    nor03_2x ix5977 (.Y (nx5976), .A0 (nx7569), .A1 (nx10240), .A2 (nx11516)) ;
    dffr gen_15_cmp_mRegCmp_reg_Q_7 (.Q (gen_15_cmp_mReg_7), .QB (nx7569), .D (
         window_15__7), .CLK (start), .R (rst)) ;
    nor03_2x ix5975 (.Y (nx5974), .A0 (gen_15_cmp_mReg_7), .A1 (nx10820), .A2 (
             nx11524)) ;
    nand02 ix6011 (.Y (gen_15_cmp_BSCmp_op2_8), .A0 (nx7573), .A1 (nx7579)) ;
    nor02_2x ix7574 (.Y (nx7573), .A0 (nx6006), .A1 (nx6002)) ;
    nor03_2x ix6007 (.Y (nx6006), .A0 (gen_15_cmp_mReg_7), .A1 (nx10246), .A2 (
             nx11492)) ;
    nor03_2x ix6003 (.Y (nx6002), .A0 (nx7569), .A1 (nx11498), .A2 (nx11508)) ;
    nor02_2x ix7580 (.Y (nx7579), .A0 (nx5998), .A1 (nx5996)) ;
    nor03_2x ix5999 (.Y (nx5998), .A0 (nx7582), .A1 (nx10240), .A2 (nx11516)) ;
    dffr gen_15_cmp_mRegCmp_reg_Q_8 (.Q (gen_15_cmp_mReg_8), .QB (nx7582), .D (
         window_15__8), .CLK (start), .R (rst)) ;
    nor03_2x ix5997 (.Y (nx5996), .A0 (gen_15_cmp_mReg_8), .A1 (nx10822), .A2 (
             nx11524)) ;
    nand02 ix6033 (.Y (gen_15_cmp_BSCmp_op2_9), .A0 (nx7589), .A1 (nx7595)) ;
    nor02_2x ix7590 (.Y (nx7589), .A0 (nx6028), .A1 (nx6024)) ;
    nor03_2x ix6029 (.Y (nx6028), .A0 (gen_15_cmp_mReg_8), .A1 (nx10246), .A2 (
             nx11492)) ;
    nor03_2x ix6025 (.Y (nx6024), .A0 (nx7582), .A1 (nx11498), .A2 (nx11508)) ;
    nor02_2x ix7596 (.Y (nx7595), .A0 (nx6020), .A1 (nx6018)) ;
    nor03_2x ix6021 (.Y (nx6020), .A0 (nx7599), .A1 (nx10240), .A2 (nx11516)) ;
    dffr gen_15_cmp_mRegCmp_reg_Q_9 (.Q (gen_15_cmp_mReg_9), .QB (nx7599), .D (
         window_15__9), .CLK (start), .R (rst)) ;
    nor03_2x ix6019 (.Y (nx6018), .A0 (gen_15_cmp_mReg_9), .A1 (nx10822), .A2 (
             nx11524)) ;
    nand02 ix6055 (.Y (gen_15_cmp_BSCmp_op2_10), .A0 (nx7603), .A1 (nx7609)) ;
    nor02_2x ix7604 (.Y (nx7603), .A0 (nx6050), .A1 (nx6046)) ;
    nor03_2x ix6051 (.Y (nx6050), .A0 (gen_15_cmp_mReg_9), .A1 (nx10246), .A2 (
             nx11492)) ;
    nor03_2x ix6047 (.Y (nx6046), .A0 (nx7599), .A1 (nx11498), .A2 (nx11508)) ;
    nor02_2x ix7610 (.Y (nx7609), .A0 (nx6042), .A1 (nx6040)) ;
    nor03_2x ix6043 (.Y (nx6042), .A0 (nx7613), .A1 (nx10240), .A2 (nx11516)) ;
    dffr gen_15_cmp_mRegCmp_reg_Q_10 (.Q (gen_15_cmp_mReg_10), .QB (nx7613), .D (
         window_15__10), .CLK (start), .R (rst)) ;
    nor03_2x ix6041 (.Y (nx6040), .A0 (gen_15_cmp_mReg_10), .A1 (nx10822), .A2 (
             nx11524)) ;
    nand02 ix6077 (.Y (gen_15_cmp_BSCmp_op2_11), .A0 (nx7617), .A1 (nx7623)) ;
    nor02_2x ix7618 (.Y (nx7617), .A0 (nx6072), .A1 (nx6068)) ;
    nor03_2x ix6073 (.Y (nx6072), .A0 (gen_15_cmp_mReg_10), .A1 (nx10246), .A2 (
             nx11492)) ;
    nor03_2x ix6069 (.Y (nx6068), .A0 (nx7613), .A1 (nx11498), .A2 (nx11508)) ;
    nor02_2x ix7624 (.Y (nx7623), .A0 (nx6064), .A1 (nx6062)) ;
    nor03_2x ix6065 (.Y (nx6064), .A0 (nx7626), .A1 (nx10240), .A2 (nx11516)) ;
    dffr gen_15_cmp_mRegCmp_reg_Q_11 (.Q (gen_15_cmp_mReg_11), .QB (nx7626), .D (
         window_15__11), .CLK (start), .R (rst)) ;
    nor03_2x ix6063 (.Y (nx6062), .A0 (gen_15_cmp_mReg_11), .A1 (nx10822), .A2 (
             nx11524)) ;
    nand02 ix6099 (.Y (gen_15_cmp_BSCmp_op2_12), .A0 (nx7633), .A1 (nx7639)) ;
    nor02_2x ix7634 (.Y (nx7633), .A0 (nx6094), .A1 (nx6090)) ;
    nor03_2x ix6095 (.Y (nx6094), .A0 (gen_15_cmp_mReg_11), .A1 (nx10246), .A2 (
             nx11492)) ;
    nor03_2x ix6091 (.Y (nx6090), .A0 (nx7626), .A1 (nx11498), .A2 (nx11508)) ;
    nor02_2x ix7640 (.Y (nx7639), .A0 (nx6086), .A1 (nx6084)) ;
    nor03_2x ix6087 (.Y (nx6086), .A0 (nx7643), .A1 (nx10242), .A2 (nx11516)) ;
    dffr gen_15_cmp_mRegCmp_reg_Q_12 (.Q (gen_15_cmp_mReg_12), .QB (nx7643), .D (
         window_15__12), .CLK (start), .R (rst)) ;
    nor03_2x ix6085 (.Y (nx6084), .A0 (gen_15_cmp_mReg_12), .A1 (nx10822), .A2 (
             nx11524)) ;
    nand02 ix6121 (.Y (gen_15_cmp_BSCmp_op2_13), .A0 (nx7647), .A1 (nx7653)) ;
    nor02_2x ix7648 (.Y (nx7647), .A0 (nx6116), .A1 (nx6112)) ;
    nor03_2x ix6117 (.Y (nx6116), .A0 (gen_15_cmp_mReg_12), .A1 (nx10248), .A2 (
             nx11494)) ;
    nor03_2x ix6113 (.Y (nx6112), .A0 (nx7643), .A1 (nx11498), .A2 (nx11510)) ;
    nor02_2x ix7654 (.Y (nx7653), .A0 (nx6108), .A1 (nx6106)) ;
    nor03_2x ix6109 (.Y (nx6108), .A0 (nx7657), .A1 (nx10242), .A2 (nx11518)) ;
    dffr gen_15_cmp_mRegCmp_reg_Q_13 (.Q (gen_15_cmp_mReg_13), .QB (nx7657), .D (
         window_15__13), .CLK (start), .R (rst)) ;
    nor03_2x ix6107 (.Y (nx6106), .A0 (gen_15_cmp_mReg_13), .A1 (nx10822), .A2 (
             nx11526)) ;
    nand02 ix6143 (.Y (gen_15_cmp_BSCmp_op2_14), .A0 (nx7661), .A1 (nx7667)) ;
    nor02_2x ix7662 (.Y (nx7661), .A0 (nx6138), .A1 (nx6134)) ;
    nor03_2x ix6139 (.Y (nx6138), .A0 (gen_15_cmp_mReg_13), .A1 (nx10248), .A2 (
             nx11494)) ;
    nor03_2x ix6135 (.Y (nx6134), .A0 (nx7657), .A1 (nx11500), .A2 (nx11510)) ;
    nor02_2x ix7668 (.Y (nx7667), .A0 (nx6130), .A1 (nx6128)) ;
    nor03_2x ix6131 (.Y (nx6130), .A0 (nx7670), .A1 (nx10242), .A2 (nx11518)) ;
    dffr gen_15_cmp_mRegCmp_reg_Q_14 (.Q (gen_15_cmp_mReg_14), .QB (nx7670), .D (
         window_15__14), .CLK (start), .R (rst)) ;
    nor03_2x ix6129 (.Y (nx6128), .A0 (gen_15_cmp_mReg_14), .A1 (nx10822), .A2 (
             nx11526)) ;
    nand02 ix6165 (.Y (gen_15_cmp_BSCmp_op2_15), .A0 (nx7677), .A1 (nx7683)) ;
    nor02_2x ix7678 (.Y (nx7677), .A0 (nx6160), .A1 (nx6156)) ;
    nor03_2x ix6161 (.Y (nx6160), .A0 (gen_15_cmp_mReg_14), .A1 (nx10248), .A2 (
             nx11494)) ;
    nor03_2x ix6157 (.Y (nx6156), .A0 (nx7670), .A1 (nx11500), .A2 (nx11510)) ;
    nor02_2x ix7684 (.Y (nx7683), .A0 (nx6152), .A1 (nx6150)) ;
    nor03_2x ix6153 (.Y (nx6152), .A0 (nx7687), .A1 (nx10242), .A2 (nx11518)) ;
    dffr gen_15_cmp_mRegCmp_reg_Q_15 (.Q (gen_15_cmp_mReg_15), .QB (nx7687), .D (
         window_15__15), .CLK (start), .R (rst)) ;
    nor03_2x ix6151 (.Y (nx6150), .A0 (gen_15_cmp_mReg_15), .A1 (nx10824), .A2 (
             nx11526)) ;
    nand02 ix6175 (.Y (gen_15_cmp_BSCmp_op2_16), .A0 (nx7691), .A1 (nx7683)) ;
    nor02_2x ix7692 (.Y (nx7691), .A0 (nx6170), .A1 (nx6166)) ;
    nor03_2x ix6171 (.Y (nx6170), .A0 (gen_15_cmp_mReg_15), .A1 (nx10248), .A2 (
             nx11494)) ;
    nor03_2x ix6167 (.Y (nx6166), .A0 (nx7687), .A1 (nx11500), .A2 (nx11510)) ;
    nand02 ix6243 (.Y (gen_16_cmp_BSCmp_op2_1), .A0 (nx7699), .A1 (nx7719)) ;
    nor02_2x ix7700 (.Y (nx7699), .A0 (nx6238), .A1 (nx6234)) ;
    nor03_2x ix6239 (.Y (nx6238), .A0 (gen_16_cmp_mReg_0), .A1 (nx10232), .A2 (
             nx11530)) ;
    dffr gen_16_cmp_mRegCmp_reg_Q_0 (.Q (gen_16_cmp_mReg_0), .QB (nx7705), .D (
         window_16__0), .CLK (start), .R (rst)) ;
    inv01 ix7710 (.Y (nx7709), .A (gen_16_cmp_pMux_0)) ;
    nor03_2x ix6235 (.Y (nx6234), .A0 (nx7705), .A1 (nx11536), .A2 (nx11546)) ;
    inv02 ix7718 (.Y (nx7717), .A (gen_16_cmp_pMux_2)) ;
    nor02_2x ix7720 (.Y (nx7719), .A0 (nx6224), .A1 (nx6222)) ;
    nor03_2x ix6225 (.Y (nx6224), .A0 (nx7723), .A1 (nx10226), .A2 (nx11554)) ;
    dffr gen_16_cmp_mRegCmp_reg_Q_1 (.Q (gen_16_cmp_mReg_1), .QB (nx7723), .D (
         window_16__1), .CLK (start), .R (rst)) ;
    nor03_2x ix6223 (.Y (nx6222), .A0 (gen_16_cmp_mReg_1), .A1 (nx10826), .A2 (
             nx11562)) ;
    nor03_2x ix6183 (.Y (nx6182), .A0 (nx10232), .A1 (nx7717), .A2 (
             gen_16_cmp_pMux_0)) ;
    nand02 ix6265 (.Y (gen_16_cmp_BSCmp_op2_2), .A0 (nx7733), .A1 (nx7737)) ;
    nor02_2x ix7734 (.Y (nx7733), .A0 (nx6260), .A1 (nx6256)) ;
    nor03_2x ix6261 (.Y (nx6260), .A0 (gen_16_cmp_mReg_1), .A1 (nx10232), .A2 (
             nx11530)) ;
    nor03_2x ix6257 (.Y (nx6256), .A0 (nx7723), .A1 (nx11536), .A2 (nx11546)) ;
    nor02_2x ix7738 (.Y (nx7737), .A0 (nx6252), .A1 (nx6250)) ;
    nor03_2x ix6253 (.Y (nx6252), .A0 (nx7741), .A1 (nx10226), .A2 (nx11554)) ;
    dffr gen_16_cmp_mRegCmp_reg_Q_2 (.Q (gen_16_cmp_mReg_2), .QB (nx7741), .D (
         window_16__2), .CLK (start), .R (rst)) ;
    nor03_2x ix6251 (.Y (nx6250), .A0 (gen_16_cmp_mReg_2), .A1 (nx10826), .A2 (
             nx11562)) ;
    nand02 ix6287 (.Y (gen_16_cmp_BSCmp_op2_3), .A0 (nx7747), .A1 (nx7753)) ;
    nor02_2x ix7748 (.Y (nx7747), .A0 (nx6282), .A1 (nx6278)) ;
    nor03_2x ix6283 (.Y (nx6282), .A0 (gen_16_cmp_mReg_2), .A1 (nx10232), .A2 (
             nx11530)) ;
    nor03_2x ix6279 (.Y (nx6278), .A0 (nx7741), .A1 (nx11536), .A2 (nx11546)) ;
    nor02_2x ix7754 (.Y (nx7753), .A0 (nx6274), .A1 (nx6272)) ;
    nor03_2x ix6275 (.Y (nx6274), .A0 (nx7757), .A1 (nx10226), .A2 (nx11554)) ;
    dffr gen_16_cmp_mRegCmp_reg_Q_3 (.Q (gen_16_cmp_mReg_3), .QB (nx7757), .D (
         window_16__3), .CLK (start), .R (rst)) ;
    nor03_2x ix6273 (.Y (nx6272), .A0 (gen_16_cmp_mReg_3), .A1 (nx10826), .A2 (
             nx11562)) ;
    nand02 ix6309 (.Y (gen_16_cmp_BSCmp_op2_4), .A0 (nx7762), .A1 (nx7767)) ;
    nor02_2x ix7763 (.Y (nx7762), .A0 (nx6304), .A1 (nx6300)) ;
    nor03_2x ix6305 (.Y (nx6304), .A0 (gen_16_cmp_mReg_3), .A1 (nx10232), .A2 (
             nx11530)) ;
    nor03_2x ix6301 (.Y (nx6300), .A0 (nx7757), .A1 (nx11536), .A2 (nx11546)) ;
    nor02_2x ix7768 (.Y (nx7767), .A0 (nx6296), .A1 (nx6294)) ;
    nor03_2x ix6297 (.Y (nx6296), .A0 (nx7771), .A1 (nx10226), .A2 (nx11554)) ;
    dffr gen_16_cmp_mRegCmp_reg_Q_4 (.Q (gen_16_cmp_mReg_4), .QB (nx7771), .D (
         window_16__4), .CLK (start), .R (rst)) ;
    nor03_2x ix6295 (.Y (nx6294), .A0 (gen_16_cmp_mReg_4), .A1 (nx10826), .A2 (
             nx11562)) ;
    nand02 ix6331 (.Y (gen_16_cmp_BSCmp_op2_5), .A0 (nx7775), .A1 (nx7781)) ;
    nor02_2x ix7776 (.Y (nx7775), .A0 (nx6326), .A1 (nx6322)) ;
    nor03_2x ix6327 (.Y (nx6326), .A0 (gen_16_cmp_mReg_4), .A1 (nx10232), .A2 (
             nx11530)) ;
    nor03_2x ix6323 (.Y (nx6322), .A0 (nx7771), .A1 (nx11536), .A2 (nx11546)) ;
    nor02_2x ix7782 (.Y (nx7781), .A0 (nx6318), .A1 (nx6316)) ;
    nor03_2x ix6319 (.Y (nx6318), .A0 (nx7785), .A1 (nx10228), .A2 (nx11554)) ;
    dffr gen_16_cmp_mRegCmp_reg_Q_5 (.Q (gen_16_cmp_mReg_5), .QB (nx7785), .D (
         window_16__5), .CLK (start), .R (rst)) ;
    nor03_2x ix6317 (.Y (nx6316), .A0 (gen_16_cmp_mReg_5), .A1 (nx10826), .A2 (
             nx11562)) ;
    nand02 ix6353 (.Y (gen_16_cmp_BSCmp_op2_6), .A0 (nx7790), .A1 (nx7795)) ;
    nor02_2x ix7791 (.Y (nx7790), .A0 (nx6348), .A1 (nx6344)) ;
    nor03_2x ix6349 (.Y (nx6348), .A0 (gen_16_cmp_mReg_5), .A1 (nx10234), .A2 (
             nx11530)) ;
    nor03_2x ix6345 (.Y (nx6344), .A0 (nx7785), .A1 (nx11536), .A2 (nx11546)) ;
    nor02_2x ix7796 (.Y (nx7795), .A0 (nx6340), .A1 (nx6338)) ;
    nor03_2x ix6341 (.Y (nx6340), .A0 (nx7799), .A1 (nx10228), .A2 (nx11554)) ;
    dffr gen_16_cmp_mRegCmp_reg_Q_6 (.Q (gen_16_cmp_mReg_6), .QB (nx7799), .D (
         window_16__6), .CLK (start), .R (rst)) ;
    nor03_2x ix6339 (.Y (nx6338), .A0 (gen_16_cmp_mReg_6), .A1 (nx10826), .A2 (
             nx11562)) ;
    nand02 ix6375 (.Y (gen_16_cmp_BSCmp_op2_7), .A0 (nx7805), .A1 (nx7811)) ;
    nor02_2x ix7806 (.Y (nx7805), .A0 (nx6370), .A1 (nx6366)) ;
    nor03_2x ix6371 (.Y (nx6370), .A0 (gen_16_cmp_mReg_6), .A1 (nx10234), .A2 (
             nx11532)) ;
    nor03_2x ix6367 (.Y (nx6366), .A0 (nx7799), .A1 (nx11538), .A2 (nx11548)) ;
    nor02_2x ix7812 (.Y (nx7811), .A0 (nx6362), .A1 (nx6360)) ;
    nor03_2x ix6363 (.Y (nx6362), .A0 (nx7814), .A1 (nx10228), .A2 (nx11556)) ;
    dffr gen_16_cmp_mRegCmp_reg_Q_7 (.Q (gen_16_cmp_mReg_7), .QB (nx7814), .D (
         window_16__7), .CLK (start), .R (rst)) ;
    nor03_2x ix6361 (.Y (nx6360), .A0 (gen_16_cmp_mReg_7), .A1 (nx10826), .A2 (
             nx11564)) ;
    nand02 ix6397 (.Y (gen_16_cmp_BSCmp_op2_8), .A0 (nx7821), .A1 (nx7827)) ;
    nor02_2x ix7822 (.Y (nx7821), .A0 (nx6392), .A1 (nx6388)) ;
    nor03_2x ix6393 (.Y (nx6392), .A0 (gen_16_cmp_mReg_7), .A1 (nx10234), .A2 (
             nx11532)) ;
    nor03_2x ix6389 (.Y (nx6388), .A0 (nx7814), .A1 (nx11538), .A2 (nx11548)) ;
    nor02_2x ix7828 (.Y (nx7827), .A0 (nx6384), .A1 (nx6382)) ;
    nor03_2x ix6385 (.Y (nx6384), .A0 (nx7831), .A1 (nx10228), .A2 (nx11556)) ;
    dffr gen_16_cmp_mRegCmp_reg_Q_8 (.Q (gen_16_cmp_mReg_8), .QB (nx7831), .D (
         window_16__8), .CLK (start), .R (rst)) ;
    nor03_2x ix6383 (.Y (nx6382), .A0 (gen_16_cmp_mReg_8), .A1 (nx10828), .A2 (
             nx11564)) ;
    nand02 ix6419 (.Y (gen_16_cmp_BSCmp_op2_9), .A0 (nx7835), .A1 (nx7841)) ;
    nor02_2x ix7836 (.Y (nx7835), .A0 (nx6414), .A1 (nx6410)) ;
    nor03_2x ix6415 (.Y (nx6414), .A0 (gen_16_cmp_mReg_8), .A1 (nx10234), .A2 (
             nx11532)) ;
    nor03_2x ix6411 (.Y (nx6410), .A0 (nx7831), .A1 (nx11538), .A2 (nx11548)) ;
    nor02_2x ix7842 (.Y (nx7841), .A0 (nx6406), .A1 (nx6404)) ;
    nor03_2x ix6407 (.Y (nx6406), .A0 (nx7845), .A1 (nx10228), .A2 (nx11556)) ;
    dffr gen_16_cmp_mRegCmp_reg_Q_9 (.Q (gen_16_cmp_mReg_9), .QB (nx7845), .D (
         window_16__9), .CLK (start), .R (rst)) ;
    nor03_2x ix6405 (.Y (nx6404), .A0 (gen_16_cmp_mReg_9), .A1 (nx10828), .A2 (
             nx11564)) ;
    nand02 ix6441 (.Y (gen_16_cmp_BSCmp_op2_10), .A0 (nx7849), .A1 (nx7855)) ;
    nor02_2x ix7850 (.Y (nx7849), .A0 (nx6436), .A1 (nx6432)) ;
    nor03_2x ix6437 (.Y (nx6436), .A0 (gen_16_cmp_mReg_9), .A1 (nx10234), .A2 (
             nx11532)) ;
    nor03_2x ix6433 (.Y (nx6432), .A0 (nx7845), .A1 (nx11538), .A2 (nx11548)) ;
    nor02_2x ix7856 (.Y (nx7855), .A0 (nx6428), .A1 (nx6426)) ;
    nor03_2x ix6429 (.Y (nx6428), .A0 (nx7858), .A1 (nx10228), .A2 (nx11556)) ;
    dffr gen_16_cmp_mRegCmp_reg_Q_10 (.Q (gen_16_cmp_mReg_10), .QB (nx7858), .D (
         window_16__10), .CLK (start), .R (rst)) ;
    nor03_2x ix6427 (.Y (nx6426), .A0 (gen_16_cmp_mReg_10), .A1 (nx10828), .A2 (
             nx11564)) ;
    nand02 ix6463 (.Y (gen_16_cmp_BSCmp_op2_11), .A0 (nx7865), .A1 (nx7871)) ;
    nor02_2x ix7866 (.Y (nx7865), .A0 (nx6458), .A1 (nx6454)) ;
    nor03_2x ix6459 (.Y (nx6458), .A0 (gen_16_cmp_mReg_10), .A1 (nx10234), .A2 (
             nx11532)) ;
    nor03_2x ix6455 (.Y (nx6454), .A0 (nx7858), .A1 (nx11538), .A2 (nx11548)) ;
    nor02_2x ix7872 (.Y (nx7871), .A0 (nx6450), .A1 (nx6448)) ;
    nor03_2x ix6451 (.Y (nx6450), .A0 (nx7875), .A1 (nx10228), .A2 (nx11556)) ;
    dffr gen_16_cmp_mRegCmp_reg_Q_11 (.Q (gen_16_cmp_mReg_11), .QB (nx7875), .D (
         window_16__11), .CLK (start), .R (rst)) ;
    nor03_2x ix6449 (.Y (nx6448), .A0 (gen_16_cmp_mReg_11), .A1 (nx10828), .A2 (
             nx11564)) ;
    nand02 ix6485 (.Y (gen_16_cmp_BSCmp_op2_12), .A0 (nx7879), .A1 (nx7885)) ;
    nor02_2x ix7880 (.Y (nx7879), .A0 (nx6480), .A1 (nx6476)) ;
    nor03_2x ix6481 (.Y (nx6480), .A0 (gen_16_cmp_mReg_11), .A1 (nx10234), .A2 (
             nx11532)) ;
    nor03_2x ix6477 (.Y (nx6476), .A0 (nx7875), .A1 (nx11538), .A2 (nx11548)) ;
    nor02_2x ix7886 (.Y (nx7885), .A0 (nx6472), .A1 (nx6470)) ;
    nor03_2x ix6473 (.Y (nx6472), .A0 (nx7889), .A1 (nx10230), .A2 (nx11556)) ;
    dffr gen_16_cmp_mRegCmp_reg_Q_12 (.Q (gen_16_cmp_mReg_12), .QB (nx7889), .D (
         window_16__12), .CLK (start), .R (rst)) ;
    nor03_2x ix6471 (.Y (nx6470), .A0 (gen_16_cmp_mReg_12), .A1 (nx10828), .A2 (
             nx11564)) ;
    nand02 ix6507 (.Y (gen_16_cmp_BSCmp_op2_13), .A0 (nx7893), .A1 (nx7899)) ;
    nor02_2x ix7894 (.Y (nx7893), .A0 (nx6502), .A1 (nx6498)) ;
    nor03_2x ix6503 (.Y (nx6502), .A0 (gen_16_cmp_mReg_12), .A1 (nx10236), .A2 (
             nx11534)) ;
    nor03_2x ix6499 (.Y (nx6498), .A0 (nx7889), .A1 (nx11538), .A2 (nx11550)) ;
    nor02_2x ix7900 (.Y (nx7899), .A0 (nx6494), .A1 (nx6492)) ;
    nor03_2x ix6495 (.Y (nx6494), .A0 (nx7902), .A1 (nx10230), .A2 (nx11558)) ;
    dffr gen_16_cmp_mRegCmp_reg_Q_13 (.Q (gen_16_cmp_mReg_13), .QB (nx7902), .D (
         window_16__13), .CLK (start), .R (rst)) ;
    nor03_2x ix6493 (.Y (nx6492), .A0 (gen_16_cmp_mReg_13), .A1 (nx10828), .A2 (
             nx11566)) ;
    nand02 ix6529 (.Y (gen_16_cmp_BSCmp_op2_14), .A0 (nx7909), .A1 (nx7915)) ;
    nor02_2x ix7910 (.Y (nx7909), .A0 (nx6524), .A1 (nx6520)) ;
    nor03_2x ix6525 (.Y (nx6524), .A0 (gen_16_cmp_mReg_13), .A1 (nx10236), .A2 (
             nx11534)) ;
    nor03_2x ix6521 (.Y (nx6520), .A0 (nx7902), .A1 (nx11540), .A2 (nx11550)) ;
    nor02_2x ix7916 (.Y (nx7915), .A0 (nx6516), .A1 (nx6514)) ;
    nor03_2x ix6517 (.Y (nx6516), .A0 (nx7919), .A1 (nx10230), .A2 (nx11558)) ;
    dffr gen_16_cmp_mRegCmp_reg_Q_14 (.Q (gen_16_cmp_mReg_14), .QB (nx7919), .D (
         window_16__14), .CLK (start), .R (rst)) ;
    nor03_2x ix6515 (.Y (nx6514), .A0 (gen_16_cmp_mReg_14), .A1 (nx10828), .A2 (
             nx11566)) ;
    nand02 ix6551 (.Y (gen_16_cmp_BSCmp_op2_15), .A0 (nx7923), .A1 (nx7929)) ;
    nor02_2x ix7924 (.Y (nx7923), .A0 (nx6546), .A1 (nx6542)) ;
    nor03_2x ix6547 (.Y (nx6546), .A0 (gen_16_cmp_mReg_14), .A1 (nx10236), .A2 (
             nx11534)) ;
    nor03_2x ix6543 (.Y (nx6542), .A0 (nx7919), .A1 (nx11540), .A2 (nx11550)) ;
    nor02_2x ix7930 (.Y (nx7929), .A0 (nx6538), .A1 (nx6536)) ;
    nor03_2x ix6539 (.Y (nx6538), .A0 (nx7933), .A1 (nx10230), .A2 (nx11558)) ;
    dffr gen_16_cmp_mRegCmp_reg_Q_15 (.Q (gen_16_cmp_mReg_15), .QB (nx7933), .D (
         window_16__15), .CLK (start), .R (rst)) ;
    nor03_2x ix6537 (.Y (nx6536), .A0 (gen_16_cmp_mReg_15), .A1 (nx10830), .A2 (
             nx11566)) ;
    nand02 ix6561 (.Y (gen_16_cmp_BSCmp_op2_16), .A0 (nx7937), .A1 (nx7929)) ;
    nor02_2x ix7938 (.Y (nx7937), .A0 (nx6556), .A1 (nx6552)) ;
    nor03_2x ix6557 (.Y (nx6556), .A0 (gen_16_cmp_mReg_15), .A1 (nx10236), .A2 (
             nx11534)) ;
    nor03_2x ix6553 (.Y (nx6552), .A0 (nx7933), .A1 (nx11540), .A2 (nx11550)) ;
    nand02 ix6629 (.Y (gen_17_cmp_BSCmp_op2_1), .A0 (nx7944), .A1 (nx7963)) ;
    nor02_2x ix7945 (.Y (nx7944), .A0 (nx6624), .A1 (nx6620)) ;
    nor03_2x ix6625 (.Y (nx6624), .A0 (gen_17_cmp_mReg_0), .A1 (nx10220), .A2 (
             nx11570)) ;
    dffr gen_17_cmp_mRegCmp_reg_Q_0 (.Q (gen_17_cmp_mReg_0), .QB (nx7949), .D (
         window_17__0), .CLK (start), .R (rst)) ;
    inv01 ix7954 (.Y (nx7953), .A (gen_17_cmp_pMux_0)) ;
    nor03_2x ix6621 (.Y (nx6620), .A0 (nx7949), .A1 (nx11576), .A2 (nx11586)) ;
    inv02 ix7962 (.Y (nx7961), .A (gen_17_cmp_pMux_2)) ;
    nor02_2x ix7964 (.Y (nx7963), .A0 (nx6610), .A1 (nx6608)) ;
    nor03_2x ix6611 (.Y (nx6610), .A0 (nx7966), .A1 (nx10214), .A2 (nx11594)) ;
    dffr gen_17_cmp_mRegCmp_reg_Q_1 (.Q (gen_17_cmp_mReg_1), .QB (nx7966), .D (
         window_17__1), .CLK (start), .R (rst)) ;
    nor03_2x ix6609 (.Y (nx6608), .A0 (gen_17_cmp_mReg_1), .A1 (nx10832), .A2 (
             nx11602)) ;
    nor03_2x ix6569 (.Y (nx6568), .A0 (nx10220), .A1 (nx7961), .A2 (
             gen_17_cmp_pMux_0)) ;
    nand02 ix6651 (.Y (gen_17_cmp_BSCmp_op2_2), .A0 (nx7979), .A1 (nx7985)) ;
    nor02_2x ix7980 (.Y (nx7979), .A0 (nx6646), .A1 (nx6642)) ;
    nor03_2x ix6647 (.Y (nx6646), .A0 (gen_17_cmp_mReg_1), .A1 (nx10220), .A2 (
             nx11570)) ;
    nor03_2x ix6643 (.Y (nx6642), .A0 (nx7966), .A1 (nx11576), .A2 (nx11586)) ;
    nor02_2x ix7986 (.Y (nx7985), .A0 (nx6638), .A1 (nx6636)) ;
    nor03_2x ix6639 (.Y (nx6638), .A0 (nx7988), .A1 (nx10214), .A2 (nx11594)) ;
    dffr gen_17_cmp_mRegCmp_reg_Q_2 (.Q (gen_17_cmp_mReg_2), .QB (nx7988), .D (
         window_17__2), .CLK (start), .R (rst)) ;
    nor03_2x ix6637 (.Y (nx6636), .A0 (gen_17_cmp_mReg_2), .A1 (nx10832), .A2 (
             nx11602)) ;
    nand02 ix6673 (.Y (gen_17_cmp_BSCmp_op2_3), .A0 (nx7993), .A1 (nx7999)) ;
    nor02_2x ix7994 (.Y (nx7993), .A0 (nx6668), .A1 (nx6664)) ;
    nor03_2x ix6669 (.Y (nx6668), .A0 (gen_17_cmp_mReg_2), .A1 (nx10220), .A2 (
             nx11570)) ;
    nor03_2x ix6665 (.Y (nx6664), .A0 (nx7988), .A1 (nx11576), .A2 (nx11586)) ;
    nor02_2x ix8000 (.Y (nx7999), .A0 (nx6660), .A1 (nx6658)) ;
    nor03_2x ix6661 (.Y (nx6660), .A0 (nx8003), .A1 (nx10214), .A2 (nx11594)) ;
    dffr gen_17_cmp_mRegCmp_reg_Q_3 (.Q (gen_17_cmp_mReg_3), .QB (nx8003), .D (
         window_17__3), .CLK (start), .R (rst)) ;
    nor03_2x ix6659 (.Y (nx6658), .A0 (gen_17_cmp_mReg_3), .A1 (nx10832), .A2 (
             nx11602)) ;
    nand02 ix6695 (.Y (gen_17_cmp_BSCmp_op2_4), .A0 (nx8009), .A1 (nx8013)) ;
    nor02_2x ix8010 (.Y (nx8009), .A0 (nx6690), .A1 (nx6686)) ;
    nor03_2x ix6691 (.Y (nx6690), .A0 (gen_17_cmp_mReg_3), .A1 (nx10220), .A2 (
             nx11570)) ;
    nor03_2x ix6687 (.Y (nx6686), .A0 (nx8003), .A1 (nx11576), .A2 (nx11586)) ;
    nor02_2x ix8014 (.Y (nx8013), .A0 (nx6682), .A1 (nx6680)) ;
    nor03_2x ix6683 (.Y (nx6682), .A0 (nx8017), .A1 (nx10214), .A2 (nx11594)) ;
    dffr gen_17_cmp_mRegCmp_reg_Q_4 (.Q (gen_17_cmp_mReg_4), .QB (nx8017), .D (
         window_17__4), .CLK (start), .R (rst)) ;
    nor03_2x ix6681 (.Y (nx6680), .A0 (gen_17_cmp_mReg_4), .A1 (nx10832), .A2 (
             nx11602)) ;
    nand02 ix6717 (.Y (gen_17_cmp_BSCmp_op2_5), .A0 (nx8023), .A1 (nx8029)) ;
    nor02_2x ix8024 (.Y (nx8023), .A0 (nx6712), .A1 (nx6708)) ;
    nor03_2x ix6713 (.Y (nx6712), .A0 (gen_17_cmp_mReg_4), .A1 (nx10220), .A2 (
             nx11570)) ;
    nor03_2x ix6709 (.Y (nx6708), .A0 (nx8017), .A1 (nx11576), .A2 (nx11586)) ;
    nor02_2x ix8030 (.Y (nx8029), .A0 (nx6704), .A1 (nx6702)) ;
    nor03_2x ix6705 (.Y (nx6704), .A0 (nx8032), .A1 (nx10216), .A2 (nx11594)) ;
    dffr gen_17_cmp_mRegCmp_reg_Q_5 (.Q (gen_17_cmp_mReg_5), .QB (nx8032), .D (
         window_17__5), .CLK (start), .R (rst)) ;
    nor03_2x ix6703 (.Y (nx6702), .A0 (gen_17_cmp_mReg_5), .A1 (nx10832), .A2 (
             nx11602)) ;
    nand02 ix6739 (.Y (gen_17_cmp_BSCmp_op2_6), .A0 (nx8037), .A1 (nx8043)) ;
    nor02_2x ix8038 (.Y (nx8037), .A0 (nx6734), .A1 (nx6730)) ;
    nor03_2x ix6735 (.Y (nx6734), .A0 (gen_17_cmp_mReg_5), .A1 (nx10222), .A2 (
             nx11570)) ;
    nor03_2x ix6731 (.Y (nx6730), .A0 (nx8032), .A1 (nx11576), .A2 (nx11586)) ;
    nor02_2x ix8044 (.Y (nx8043), .A0 (nx6726), .A1 (nx6724)) ;
    nor03_2x ix6727 (.Y (nx6726), .A0 (nx8047), .A1 (nx10216), .A2 (nx11594)) ;
    dffr gen_17_cmp_mRegCmp_reg_Q_6 (.Q (gen_17_cmp_mReg_6), .QB (nx8047), .D (
         window_17__6), .CLK (start), .R (rst)) ;
    nor03_2x ix6725 (.Y (nx6724), .A0 (gen_17_cmp_mReg_6), .A1 (nx10832), .A2 (
             nx11602)) ;
    nand02 ix6761 (.Y (gen_17_cmp_BSCmp_op2_7), .A0 (nx8053), .A1 (nx8057)) ;
    nor02_2x ix8054 (.Y (nx8053), .A0 (nx6756), .A1 (nx6752)) ;
    nor03_2x ix6757 (.Y (nx6756), .A0 (gen_17_cmp_mReg_6), .A1 (nx10222), .A2 (
             nx11572)) ;
    nor03_2x ix6753 (.Y (nx6752), .A0 (nx8047), .A1 (nx11578), .A2 (nx11588)) ;
    nor02_2x ix8058 (.Y (nx8057), .A0 (nx6748), .A1 (nx6746)) ;
    nor03_2x ix6749 (.Y (nx6748), .A0 (nx8061), .A1 (nx10216), .A2 (nx11596)) ;
    dffr gen_17_cmp_mRegCmp_reg_Q_7 (.Q (gen_17_cmp_mReg_7), .QB (nx8061), .D (
         window_17__7), .CLK (start), .R (rst)) ;
    nor03_2x ix6747 (.Y (nx6746), .A0 (gen_17_cmp_mReg_7), .A1 (nx10832), .A2 (
             nx11604)) ;
    nand02 ix6783 (.Y (gen_17_cmp_BSCmp_op2_8), .A0 (nx8067), .A1 (nx8073)) ;
    nor02_2x ix8068 (.Y (nx8067), .A0 (nx6778), .A1 (nx6774)) ;
    nor03_2x ix6779 (.Y (nx6778), .A0 (gen_17_cmp_mReg_7), .A1 (nx10222), .A2 (
             nx11572)) ;
    nor03_2x ix6775 (.Y (nx6774), .A0 (nx8061), .A1 (nx11578), .A2 (nx11588)) ;
    nor02_2x ix8074 (.Y (nx8073), .A0 (nx6770), .A1 (nx6768)) ;
    nor03_2x ix6771 (.Y (nx6770), .A0 (nx8076), .A1 (nx10216), .A2 (nx11596)) ;
    dffr gen_17_cmp_mRegCmp_reg_Q_8 (.Q (gen_17_cmp_mReg_8), .QB (nx8076), .D (
         window_17__8), .CLK (start), .R (rst)) ;
    nor03_2x ix6769 (.Y (nx6768), .A0 (gen_17_cmp_mReg_8), .A1 (nx10834), .A2 (
             nx11604)) ;
    nand02 ix6805 (.Y (gen_17_cmp_BSCmp_op2_9), .A0 (nx8081), .A1 (nx8087)) ;
    nor02_2x ix8082 (.Y (nx8081), .A0 (nx6800), .A1 (nx6796)) ;
    nor03_2x ix6801 (.Y (nx6800), .A0 (gen_17_cmp_mReg_8), .A1 (nx10222), .A2 (
             nx11572)) ;
    nor03_2x ix6797 (.Y (nx6796), .A0 (nx8076), .A1 (nx11578), .A2 (nx11588)) ;
    nor02_2x ix8088 (.Y (nx8087), .A0 (nx6792), .A1 (nx6790)) ;
    nor03_2x ix6793 (.Y (nx6792), .A0 (nx8091), .A1 (nx10216), .A2 (nx11596)) ;
    dffr gen_17_cmp_mRegCmp_reg_Q_9 (.Q (gen_17_cmp_mReg_9), .QB (nx8091), .D (
         window_17__9), .CLK (start), .R (rst)) ;
    nor03_2x ix6791 (.Y (nx6790), .A0 (gen_17_cmp_mReg_9), .A1 (nx10834), .A2 (
             nx11604)) ;
    nand02 ix6827 (.Y (gen_17_cmp_BSCmp_op2_10), .A0 (nx8097), .A1 (nx8101)) ;
    nor02_2x ix8098 (.Y (nx8097), .A0 (nx6822), .A1 (nx6818)) ;
    nor03_2x ix6823 (.Y (nx6822), .A0 (gen_17_cmp_mReg_9), .A1 (nx10222), .A2 (
             nx11572)) ;
    nor03_2x ix6819 (.Y (nx6818), .A0 (nx8091), .A1 (nx11578), .A2 (nx11588)) ;
    nor02_2x ix8102 (.Y (nx8101), .A0 (nx6814), .A1 (nx6812)) ;
    nor03_2x ix6815 (.Y (nx6814), .A0 (nx8105), .A1 (nx10216), .A2 (nx11596)) ;
    dffr gen_17_cmp_mRegCmp_reg_Q_10 (.Q (gen_17_cmp_mReg_10), .QB (nx8105), .D (
         window_17__10), .CLK (start), .R (rst)) ;
    nor03_2x ix6813 (.Y (nx6812), .A0 (gen_17_cmp_mReg_10), .A1 (nx10834), .A2 (
             nx11604)) ;
    nand02 ix6849 (.Y (gen_17_cmp_BSCmp_op2_11), .A0 (nx8111), .A1 (nx8116)) ;
    nor02_2x ix8112 (.Y (nx8111), .A0 (nx6844), .A1 (nx6840)) ;
    nor03_2x ix6845 (.Y (nx6844), .A0 (gen_17_cmp_mReg_10), .A1 (nx10222), .A2 (
             nx11572)) ;
    nor03_2x ix6841 (.Y (nx6840), .A0 (nx8105), .A1 (nx11578), .A2 (nx11588)) ;
    nor02_2x ix8117 (.Y (nx8116), .A0 (nx6836), .A1 (nx6834)) ;
    nor03_2x ix6837 (.Y (nx6836), .A0 (nx8119), .A1 (nx10216), .A2 (nx11596)) ;
    dffr gen_17_cmp_mRegCmp_reg_Q_11 (.Q (gen_17_cmp_mReg_11), .QB (nx8119), .D (
         window_17__11), .CLK (start), .R (rst)) ;
    nor03_2x ix6835 (.Y (nx6834), .A0 (gen_17_cmp_mReg_11), .A1 (nx10834), .A2 (
             nx11604)) ;
    nand02 ix6871 (.Y (gen_17_cmp_BSCmp_op2_12), .A0 (nx8123), .A1 (nx8129)) ;
    nor02_2x ix8124 (.Y (nx8123), .A0 (nx6866), .A1 (nx6862)) ;
    nor03_2x ix6867 (.Y (nx6866), .A0 (gen_17_cmp_mReg_11), .A1 (nx10222), .A2 (
             nx11572)) ;
    nor03_2x ix6863 (.Y (nx6862), .A0 (nx8119), .A1 (nx11578), .A2 (nx11588)) ;
    nor02_2x ix8130 (.Y (nx8129), .A0 (nx6858), .A1 (nx6856)) ;
    nor03_2x ix6859 (.Y (nx6858), .A0 (nx8133), .A1 (nx10218), .A2 (nx11596)) ;
    dffr gen_17_cmp_mRegCmp_reg_Q_12 (.Q (gen_17_cmp_mReg_12), .QB (nx8133), .D (
         window_17__12), .CLK (start), .R (rst)) ;
    nor03_2x ix6857 (.Y (nx6856), .A0 (gen_17_cmp_mReg_12), .A1 (nx10834), .A2 (
             nx11604)) ;
    nand02 ix6893 (.Y (gen_17_cmp_BSCmp_op2_13), .A0 (nx8139), .A1 (nx8145)) ;
    nor02_2x ix8140 (.Y (nx8139), .A0 (nx6888), .A1 (nx6884)) ;
    nor03_2x ix6889 (.Y (nx6888), .A0 (gen_17_cmp_mReg_12), .A1 (nx10224), .A2 (
             nx11574)) ;
    nor03_2x ix6885 (.Y (nx6884), .A0 (nx8133), .A1 (nx11578), .A2 (nx11590)) ;
    nor02_2x ix8146 (.Y (nx8145), .A0 (nx6880), .A1 (nx6878)) ;
    nor03_2x ix6881 (.Y (nx6880), .A0 (nx8148), .A1 (nx10218), .A2 (nx11598)) ;
    dffr gen_17_cmp_mRegCmp_reg_Q_13 (.Q (gen_17_cmp_mReg_13), .QB (nx8148), .D (
         window_17__13), .CLK (start), .R (rst)) ;
    nor03_2x ix6879 (.Y (nx6878), .A0 (gen_17_cmp_mReg_13), .A1 (nx10834), .A2 (
             nx11606)) ;
    nand02 ix6915 (.Y (gen_17_cmp_BSCmp_op2_14), .A0 (nx8153), .A1 (nx8159)) ;
    nor02_2x ix8154 (.Y (nx8153), .A0 (nx6910), .A1 (nx6906)) ;
    nor03_2x ix6911 (.Y (nx6910), .A0 (gen_17_cmp_mReg_13), .A1 (nx10224), .A2 (
             nx11574)) ;
    nor03_2x ix6907 (.Y (nx6906), .A0 (nx8148), .A1 (nx11580), .A2 (nx11590)) ;
    nor02_2x ix8160 (.Y (nx8159), .A0 (nx6902), .A1 (nx6900)) ;
    nor03_2x ix6903 (.Y (nx6902), .A0 (nx8163), .A1 (nx10218), .A2 (nx11598)) ;
    dffr gen_17_cmp_mRegCmp_reg_Q_14 (.Q (gen_17_cmp_mReg_14), .QB (nx8163), .D (
         window_17__14), .CLK (start), .R (rst)) ;
    nor03_2x ix6901 (.Y (nx6900), .A0 (gen_17_cmp_mReg_14), .A1 (nx10834), .A2 (
             nx11606)) ;
    nand02 ix6937 (.Y (gen_17_cmp_BSCmp_op2_15), .A0 (nx8169), .A1 (nx8175)) ;
    nor02_2x ix8170 (.Y (nx8169), .A0 (nx6932), .A1 (nx6928)) ;
    nor03_2x ix6933 (.Y (nx6932), .A0 (gen_17_cmp_mReg_14), .A1 (nx10224), .A2 (
             nx11574)) ;
    nor03_2x ix6929 (.Y (nx6928), .A0 (nx8163), .A1 (nx11580), .A2 (nx11590)) ;
    nor02_2x ix8176 (.Y (nx8175), .A0 (nx6924), .A1 (nx6922)) ;
    nor03_2x ix6925 (.Y (nx6924), .A0 (nx8178), .A1 (nx10218), .A2 (nx11598)) ;
    dffr gen_17_cmp_mRegCmp_reg_Q_15 (.Q (gen_17_cmp_mReg_15), .QB (nx8178), .D (
         window_17__15), .CLK (start), .R (rst)) ;
    nor03_2x ix6923 (.Y (nx6922), .A0 (gen_17_cmp_mReg_15), .A1 (nx10836), .A2 (
             nx11606)) ;
    nand02 ix6947 (.Y (gen_17_cmp_BSCmp_op2_16), .A0 (nx8185), .A1 (nx8175)) ;
    nor02_2x ix8186 (.Y (nx8185), .A0 (nx6942), .A1 (nx6938)) ;
    nor03_2x ix6943 (.Y (nx6942), .A0 (gen_17_cmp_mReg_15), .A1 (nx10224), .A2 (
             nx11574)) ;
    nor03_2x ix6939 (.Y (nx6938), .A0 (nx8178), .A1 (nx11580), .A2 (nx11590)) ;
    nand02 ix7015 (.Y (gen_18_cmp_BSCmp_op2_1), .A0 (nx8191), .A1 (nx8211)) ;
    nor02_2x ix8192 (.Y (nx8191), .A0 (nx7010), .A1 (nx7006)) ;
    nor03_2x ix7011 (.Y (nx7010), .A0 (gen_18_cmp_mReg_0), .A1 (nx10208), .A2 (
             nx11610)) ;
    dffr gen_18_cmp_mRegCmp_reg_Q_0 (.Q (gen_18_cmp_mReg_0), .QB (nx8197), .D (
         window_18__0), .CLK (start), .R (rst)) ;
    inv01 ix8202 (.Y (nx8200), .A (gen_18_cmp_pMux_0)) ;
    nor03_2x ix7007 (.Y (nx7006), .A0 (nx8197), .A1 (nx11616), .A2 (nx11626)) ;
    inv02 ix8210 (.Y (nx8209), .A (gen_18_cmp_pMux_2)) ;
    nor02_2x ix8212 (.Y (nx8211), .A0 (nx6996), .A1 (nx6994)) ;
    nor03_2x ix6997 (.Y (nx6996), .A0 (nx8215), .A1 (nx10202), .A2 (nx11634)) ;
    dffr gen_18_cmp_mRegCmp_reg_Q_1 (.Q (gen_18_cmp_mReg_1), .QB (nx8215), .D (
         window_18__1), .CLK (start), .R (rst)) ;
    nor03_2x ix6995 (.Y (nx6994), .A0 (gen_18_cmp_mReg_1), .A1 (nx10838), .A2 (
             nx11642)) ;
    nor03_2x ix6955 (.Y (nx6954), .A0 (nx10208), .A1 (nx8209), .A2 (
             gen_18_cmp_pMux_0)) ;
    nand02 ix7037 (.Y (gen_18_cmp_BSCmp_op2_2), .A0 (nx8225), .A1 (nx8231)) ;
    nor02_2x ix8226 (.Y (nx8225), .A0 (nx7032), .A1 (nx7028)) ;
    nor03_2x ix7033 (.Y (nx7032), .A0 (gen_18_cmp_mReg_1), .A1 (nx10208), .A2 (
             nx11610)) ;
    nor03_2x ix7029 (.Y (nx7028), .A0 (nx8215), .A1 (nx11616), .A2 (nx11626)) ;
    nor02_2x ix8232 (.Y (nx8231), .A0 (nx7024), .A1 (nx7022)) ;
    nor03_2x ix7025 (.Y (nx7024), .A0 (nx8235), .A1 (nx10202), .A2 (nx11634)) ;
    dffr gen_18_cmp_mRegCmp_reg_Q_2 (.Q (gen_18_cmp_mReg_2), .QB (nx8235), .D (
         window_18__2), .CLK (start), .R (rst)) ;
    nor03_2x ix7023 (.Y (nx7022), .A0 (gen_18_cmp_mReg_2), .A1 (nx10838), .A2 (
             nx11642)) ;
    nand02 ix7059 (.Y (gen_18_cmp_BSCmp_op2_3), .A0 (nx8241), .A1 (nx8245)) ;
    nor02_2x ix8242 (.Y (nx8241), .A0 (nx7054), .A1 (nx7050)) ;
    nor03_2x ix7055 (.Y (nx7054), .A0 (gen_18_cmp_mReg_2), .A1 (nx10208), .A2 (
             nx11610)) ;
    nor03_2x ix7051 (.Y (nx7050), .A0 (nx8235), .A1 (nx11616), .A2 (nx11626)) ;
    nor02_2x ix8246 (.Y (nx8245), .A0 (nx7046), .A1 (nx7044)) ;
    nor03_2x ix7047 (.Y (nx7046), .A0 (nx8249), .A1 (nx10202), .A2 (nx11634)) ;
    dffr gen_18_cmp_mRegCmp_reg_Q_3 (.Q (gen_18_cmp_mReg_3), .QB (nx8249), .D (
         window_18__3), .CLK (start), .R (rst)) ;
    nor03_2x ix7045 (.Y (nx7044), .A0 (gen_18_cmp_mReg_3), .A1 (nx10838), .A2 (
             nx11642)) ;
    nand02 ix7081 (.Y (gen_18_cmp_BSCmp_op2_4), .A0 (nx8255), .A1 (nx8261)) ;
    nor02_2x ix8256 (.Y (nx8255), .A0 (nx7076), .A1 (nx7072)) ;
    nor03_2x ix7077 (.Y (nx7076), .A0 (gen_18_cmp_mReg_3), .A1 (nx10208), .A2 (
             nx11610)) ;
    nor03_2x ix7073 (.Y (nx7072), .A0 (nx8249), .A1 (nx11616), .A2 (nx11626)) ;
    nor02_2x ix8262 (.Y (nx8261), .A0 (nx7068), .A1 (nx7066)) ;
    nor03_2x ix7069 (.Y (nx7068), .A0 (nx8264), .A1 (nx10202), .A2 (nx11634)) ;
    dffr gen_18_cmp_mRegCmp_reg_Q_4 (.Q (gen_18_cmp_mReg_4), .QB (nx8264), .D (
         window_18__4), .CLK (start), .R (rst)) ;
    nor03_2x ix7067 (.Y (nx7066), .A0 (gen_18_cmp_mReg_4), .A1 (nx10838), .A2 (
             nx11642)) ;
    nand02 ix7103 (.Y (gen_18_cmp_BSCmp_op2_5), .A0 (nx8269), .A1 (nx8275)) ;
    nor02_2x ix8270 (.Y (nx8269), .A0 (nx7098), .A1 (nx7094)) ;
    nor03_2x ix7099 (.Y (nx7098), .A0 (gen_18_cmp_mReg_4), .A1 (nx10208), .A2 (
             nx11610)) ;
    nor03_2x ix7095 (.Y (nx7094), .A0 (nx8264), .A1 (nx11616), .A2 (nx11626)) ;
    nor02_2x ix8276 (.Y (nx8275), .A0 (nx7090), .A1 (nx7088)) ;
    nor03_2x ix7091 (.Y (nx7090), .A0 (nx8279), .A1 (nx10204), .A2 (nx11634)) ;
    dffr gen_18_cmp_mRegCmp_reg_Q_5 (.Q (gen_18_cmp_mReg_5), .QB (nx8279), .D (
         window_18__5), .CLK (start), .R (rst)) ;
    nor03_2x ix7089 (.Y (nx7088), .A0 (gen_18_cmp_mReg_5), .A1 (nx10838), .A2 (
             nx11642)) ;
    nand02 ix7125 (.Y (gen_18_cmp_BSCmp_op2_6), .A0 (nx8285), .A1 (nx8289)) ;
    nor02_2x ix8286 (.Y (nx8285), .A0 (nx7120), .A1 (nx7116)) ;
    nor03_2x ix7121 (.Y (nx7120), .A0 (gen_18_cmp_mReg_5), .A1 (nx10210), .A2 (
             nx11610)) ;
    nor03_2x ix7117 (.Y (nx7116), .A0 (nx8279), .A1 (nx11616), .A2 (nx11626)) ;
    nor02_2x ix8290 (.Y (nx8289), .A0 (nx7112), .A1 (nx7110)) ;
    nor03_2x ix7113 (.Y (nx7112), .A0 (nx8293), .A1 (nx10204), .A2 (nx11634)) ;
    dffr gen_18_cmp_mRegCmp_reg_Q_6 (.Q (gen_18_cmp_mReg_6), .QB (nx8293), .D (
         window_18__6), .CLK (start), .R (rst)) ;
    nor03_2x ix7111 (.Y (nx7110), .A0 (gen_18_cmp_mReg_6), .A1 (nx10838), .A2 (
             nx11642)) ;
    nand02 ix7147 (.Y (gen_18_cmp_BSCmp_op2_7), .A0 (nx8299), .A1 (nx8305)) ;
    nor02_2x ix8300 (.Y (nx8299), .A0 (nx7142), .A1 (nx7138)) ;
    nor03_2x ix7143 (.Y (nx7142), .A0 (gen_18_cmp_mReg_6), .A1 (nx10210), .A2 (
             nx11612)) ;
    nor03_2x ix7139 (.Y (nx7138), .A0 (nx8293), .A1 (nx11618), .A2 (nx11628)) ;
    nor02_2x ix8306 (.Y (nx8305), .A0 (nx7134), .A1 (nx7132)) ;
    nor03_2x ix7135 (.Y (nx7134), .A0 (nx8308), .A1 (nx10204), .A2 (nx11636)) ;
    dffr gen_18_cmp_mRegCmp_reg_Q_7 (.Q (gen_18_cmp_mReg_7), .QB (nx8308), .D (
         window_18__7), .CLK (start), .R (rst)) ;
    nor03_2x ix7133 (.Y (nx7132), .A0 (gen_18_cmp_mReg_7), .A1 (nx10838), .A2 (
             nx11644)) ;
    nand02 ix7169 (.Y (gen_18_cmp_BSCmp_op2_8), .A0 (nx8313), .A1 (nx8319)) ;
    nor02_2x ix8314 (.Y (nx8313), .A0 (nx7164), .A1 (nx7160)) ;
    nor03_2x ix7165 (.Y (nx7164), .A0 (gen_18_cmp_mReg_7), .A1 (nx10210), .A2 (
             nx11612)) ;
    nor03_2x ix7161 (.Y (nx7160), .A0 (nx8308), .A1 (nx11618), .A2 (nx11628)) ;
    nor02_2x ix8320 (.Y (nx8319), .A0 (nx7156), .A1 (nx7154)) ;
    nor03_2x ix7157 (.Y (nx7156), .A0 (nx8323), .A1 (nx10204), .A2 (nx11636)) ;
    dffr gen_18_cmp_mRegCmp_reg_Q_8 (.Q (gen_18_cmp_mReg_8), .QB (nx8323), .D (
         window_18__8), .CLK (start), .R (rst)) ;
    nor03_2x ix7155 (.Y (nx7154), .A0 (gen_18_cmp_mReg_8), .A1 (nx10840), .A2 (
             nx11644)) ;
    nand02 ix7191 (.Y (gen_18_cmp_BSCmp_op2_9), .A0 (nx8329), .A1 (nx8333)) ;
    nor02_2x ix8330 (.Y (nx8329), .A0 (nx7186), .A1 (nx7182)) ;
    nor03_2x ix7187 (.Y (nx7186), .A0 (gen_18_cmp_mReg_8), .A1 (nx10210), .A2 (
             nx11612)) ;
    nor03_2x ix7183 (.Y (nx7182), .A0 (nx8323), .A1 (nx11618), .A2 (nx11628)) ;
    nor02_2x ix8334 (.Y (nx8333), .A0 (nx7178), .A1 (nx7176)) ;
    nor03_2x ix7179 (.Y (nx7178), .A0 (nx8337), .A1 (nx10204), .A2 (nx11636)) ;
    dffr gen_18_cmp_mRegCmp_reg_Q_9 (.Q (gen_18_cmp_mReg_9), .QB (nx8337), .D (
         window_18__9), .CLK (start), .R (rst)) ;
    nor03_2x ix7177 (.Y (nx7176), .A0 (gen_18_cmp_mReg_9), .A1 (nx10840), .A2 (
             nx11644)) ;
    nand02 ix7213 (.Y (gen_18_cmp_BSCmp_op2_10), .A0 (nx8343), .A1 (nx8349)) ;
    nor02_2x ix8344 (.Y (nx8343), .A0 (nx7208), .A1 (nx7204)) ;
    nor03_2x ix7209 (.Y (nx7208), .A0 (gen_18_cmp_mReg_9), .A1 (nx10210), .A2 (
             nx11612)) ;
    nor03_2x ix7205 (.Y (nx7204), .A0 (nx8337), .A1 (nx11618), .A2 (nx11628)) ;
    nor02_2x ix8350 (.Y (nx8349), .A0 (nx7200), .A1 (nx7198)) ;
    nor03_2x ix7201 (.Y (nx7200), .A0 (nx8352), .A1 (nx10204), .A2 (nx11636)) ;
    dffr gen_18_cmp_mRegCmp_reg_Q_10 (.Q (gen_18_cmp_mReg_10), .QB (nx8352), .D (
         window_18__10), .CLK (start), .R (rst)) ;
    nor03_2x ix7199 (.Y (nx7198), .A0 (gen_18_cmp_mReg_10), .A1 (nx10840), .A2 (
             nx11644)) ;
    nand02 ix7235 (.Y (gen_18_cmp_BSCmp_op2_11), .A0 (nx8357), .A1 (nx8363)) ;
    nor02_2x ix8358 (.Y (nx8357), .A0 (nx7230), .A1 (nx7226)) ;
    nor03_2x ix7231 (.Y (nx7230), .A0 (gen_18_cmp_mReg_10), .A1 (nx10210), .A2 (
             nx11612)) ;
    nor03_2x ix7227 (.Y (nx7226), .A0 (nx8352), .A1 (nx11618), .A2 (nx11628)) ;
    nor02_2x ix8364 (.Y (nx8363), .A0 (nx7222), .A1 (nx7220)) ;
    nor03_2x ix7223 (.Y (nx7222), .A0 (nx8367), .A1 (nx10204), .A2 (nx11636)) ;
    dffr gen_18_cmp_mRegCmp_reg_Q_11 (.Q (gen_18_cmp_mReg_11), .QB (nx8367), .D (
         window_18__11), .CLK (start), .R (rst)) ;
    nor03_2x ix7221 (.Y (nx7220), .A0 (gen_18_cmp_mReg_11), .A1 (nx10840), .A2 (
             nx11644)) ;
    nand02 ix7257 (.Y (gen_18_cmp_BSCmp_op2_12), .A0 (nx8373), .A1 (nx8377)) ;
    nor02_2x ix8374 (.Y (nx8373), .A0 (nx7252), .A1 (nx7248)) ;
    nor03_2x ix7253 (.Y (nx7252), .A0 (gen_18_cmp_mReg_11), .A1 (nx10210), .A2 (
             nx11612)) ;
    nor03_2x ix7249 (.Y (nx7248), .A0 (nx8367), .A1 (nx11618), .A2 (nx11628)) ;
    nor02_2x ix8378 (.Y (nx8377), .A0 (nx7244), .A1 (nx7242)) ;
    nor03_2x ix7245 (.Y (nx7244), .A0 (nx8381), .A1 (nx10206), .A2 (nx11636)) ;
    dffr gen_18_cmp_mRegCmp_reg_Q_12 (.Q (gen_18_cmp_mReg_12), .QB (nx8381), .D (
         window_18__12), .CLK (start), .R (rst)) ;
    nor03_2x ix7243 (.Y (nx7242), .A0 (gen_18_cmp_mReg_12), .A1 (nx10840), .A2 (
             nx11644)) ;
    nand02 ix7279 (.Y (gen_18_cmp_BSCmp_op2_13), .A0 (nx8387), .A1 (nx8393)) ;
    nor02_2x ix8388 (.Y (nx8387), .A0 (nx7274), .A1 (nx7270)) ;
    nor03_2x ix7275 (.Y (nx7274), .A0 (gen_18_cmp_mReg_12), .A1 (nx10212), .A2 (
             nx11614)) ;
    nor03_2x ix7271 (.Y (nx7270), .A0 (nx8381), .A1 (nx11618), .A2 (nx11630)) ;
    nor02_2x ix8394 (.Y (nx8393), .A0 (nx7266), .A1 (nx7264)) ;
    nor03_2x ix7267 (.Y (nx7266), .A0 (nx8396), .A1 (nx10206), .A2 (nx11638)) ;
    dffr gen_18_cmp_mRegCmp_reg_Q_13 (.Q (gen_18_cmp_mReg_13), .QB (nx8396), .D (
         window_18__13), .CLK (start), .R (rst)) ;
    nor03_2x ix7265 (.Y (nx7264), .A0 (gen_18_cmp_mReg_13), .A1 (nx10840), .A2 (
             nx11646)) ;
    nand02 ix7301 (.Y (gen_18_cmp_BSCmp_op2_14), .A0 (nx8401), .A1 (nx8407)) ;
    nor02_2x ix8402 (.Y (nx8401), .A0 (nx7296), .A1 (nx7292)) ;
    nor03_2x ix7297 (.Y (nx7296), .A0 (gen_18_cmp_mReg_13), .A1 (nx10212), .A2 (
             nx11614)) ;
    nor03_2x ix7293 (.Y (nx7292), .A0 (nx8396), .A1 (nx11620), .A2 (nx11630)) ;
    nor02_2x ix8408 (.Y (nx8407), .A0 (nx7288), .A1 (nx7286)) ;
    nor03_2x ix7289 (.Y (nx7288), .A0 (nx8411), .A1 (nx10206), .A2 (nx11638)) ;
    dffr gen_18_cmp_mRegCmp_reg_Q_14 (.Q (gen_18_cmp_mReg_14), .QB (nx8411), .D (
         window_18__14), .CLK (start), .R (rst)) ;
    nor03_2x ix7287 (.Y (nx7286), .A0 (gen_18_cmp_mReg_14), .A1 (nx10840), .A2 (
             nx11646)) ;
    nand02 ix7323 (.Y (gen_18_cmp_BSCmp_op2_15), .A0 (nx8417), .A1 (nx8421)) ;
    nor02_2x ix8418 (.Y (nx8417), .A0 (nx7318), .A1 (nx7314)) ;
    nor03_2x ix7319 (.Y (nx7318), .A0 (gen_18_cmp_mReg_14), .A1 (nx10212), .A2 (
             nx11614)) ;
    nor03_2x ix7315 (.Y (nx7314), .A0 (nx8411), .A1 (nx11620), .A2 (nx11630)) ;
    nor02_2x ix8422 (.Y (nx8421), .A0 (nx7310), .A1 (nx7308)) ;
    nor03_2x ix7311 (.Y (nx7310), .A0 (nx8425), .A1 (nx10206), .A2 (nx11638)) ;
    dffr gen_18_cmp_mRegCmp_reg_Q_15 (.Q (gen_18_cmp_mReg_15), .QB (nx8425), .D (
         window_18__15), .CLK (start), .R (rst)) ;
    nor03_2x ix7309 (.Y (nx7308), .A0 (gen_18_cmp_mReg_15), .A1 (nx10842), .A2 (
             nx11646)) ;
    nand02 ix7333 (.Y (gen_18_cmp_BSCmp_op2_16), .A0 (nx8431), .A1 (nx8421)) ;
    nor02_2x ix8432 (.Y (nx8431), .A0 (nx7328), .A1 (nx7324)) ;
    nor03_2x ix7329 (.Y (nx7328), .A0 (gen_18_cmp_mReg_15), .A1 (nx10212), .A2 (
             nx11614)) ;
    nor03_2x ix7325 (.Y (nx7324), .A0 (nx8425), .A1 (nx11620), .A2 (nx11630)) ;
    nand02 ix7401 (.Y (gen_19_cmp_BSCmp_op2_1), .A0 (nx8439), .A1 (nx8457)) ;
    nor02_2x ix8440 (.Y (nx8439), .A0 (nx7396), .A1 (nx7392)) ;
    nor03_2x ix7397 (.Y (nx7396), .A0 (gen_19_cmp_mReg_0), .A1 (nx10196), .A2 (
             nx11650)) ;
    dffr gen_19_cmp_mRegCmp_reg_Q_0 (.Q (gen_19_cmp_mReg_0), .QB (nx8443), .D (
         window_19__0), .CLK (start), .R (rst)) ;
    inv01 ix8448 (.Y (nx8447), .A (gen_19_cmp_pMux_0)) ;
    nor03_2x ix7393 (.Y (nx7392), .A0 (nx8443), .A1 (nx11656), .A2 (nx11666)) ;
    inv02 ix8456 (.Y (nx8455), .A (gen_19_cmp_pMux_2)) ;
    nor02_2x ix8458 (.Y (nx8457), .A0 (nx7382), .A1 (nx7380)) ;
    nor03_2x ix7383 (.Y (nx7382), .A0 (nx8461), .A1 (nx10190), .A2 (nx11674)) ;
    dffr gen_19_cmp_mRegCmp_reg_Q_1 (.Q (gen_19_cmp_mReg_1), .QB (nx8461), .D (
         window_19__1), .CLK (start), .R (rst)) ;
    nor03_2x ix7381 (.Y (nx7380), .A0 (gen_19_cmp_mReg_1), .A1 (nx10844), .A2 (
             nx11682)) ;
    nor03_2x ix7341 (.Y (nx7340), .A0 (nx10196), .A1 (nx8455), .A2 (
             gen_19_cmp_pMux_0)) ;
    nand02 ix7423 (.Y (gen_19_cmp_BSCmp_op2_2), .A0 (nx8473), .A1 (nx8477)) ;
    nor02_2x ix8474 (.Y (nx8473), .A0 (nx7418), .A1 (nx7414)) ;
    nor03_2x ix7419 (.Y (nx7418), .A0 (gen_19_cmp_mReg_1), .A1 (nx10196), .A2 (
             nx11650)) ;
    nor03_2x ix7415 (.Y (nx7414), .A0 (nx8461), .A1 (nx11656), .A2 (nx11666)) ;
    nor02_2x ix8478 (.Y (nx8477), .A0 (nx7410), .A1 (nx7408)) ;
    nor03_2x ix7411 (.Y (nx7410), .A0 (nx8481), .A1 (nx10190), .A2 (nx11674)) ;
    dffr gen_19_cmp_mRegCmp_reg_Q_2 (.Q (gen_19_cmp_mReg_2), .QB (nx8481), .D (
         window_19__2), .CLK (start), .R (rst)) ;
    nor03_2x ix7409 (.Y (nx7408), .A0 (gen_19_cmp_mReg_2), .A1 (nx10844), .A2 (
             nx11682)) ;
    nand02 ix7445 (.Y (gen_19_cmp_BSCmp_op2_3), .A0 (nx8487), .A1 (nx8493)) ;
    nor02_2x ix8488 (.Y (nx8487), .A0 (nx7440), .A1 (nx7436)) ;
    nor03_2x ix7441 (.Y (nx7440), .A0 (gen_19_cmp_mReg_2), .A1 (nx10196), .A2 (
             nx11650)) ;
    nor03_2x ix7437 (.Y (nx7436), .A0 (nx8481), .A1 (nx11656), .A2 (nx11666)) ;
    nor02_2x ix8494 (.Y (nx8493), .A0 (nx7432), .A1 (nx7430)) ;
    nor03_2x ix7433 (.Y (nx7432), .A0 (nx8497), .A1 (nx10190), .A2 (nx11674)) ;
    dffr gen_19_cmp_mRegCmp_reg_Q_3 (.Q (gen_19_cmp_mReg_3), .QB (nx8497), .D (
         window_19__3), .CLK (start), .R (rst)) ;
    nor03_2x ix7431 (.Y (nx7430), .A0 (gen_19_cmp_mReg_3), .A1 (nx10844), .A2 (
             nx11682)) ;
    nand02 ix7467 (.Y (gen_19_cmp_BSCmp_op2_4), .A0 (nx8502), .A1 (nx8506)) ;
    nor02_2x ix8503 (.Y (nx8502), .A0 (nx7462), .A1 (nx7458)) ;
    nor03_2x ix7463 (.Y (nx7462), .A0 (gen_19_cmp_mReg_3), .A1 (nx10196), .A2 (
             nx11650)) ;
    nor03_2x ix7459 (.Y (nx7458), .A0 (nx8497), .A1 (nx11656), .A2 (nx11666)) ;
    nor02_2x ix8507 (.Y (nx8506), .A0 (nx7454), .A1 (nx7452)) ;
    nor03_2x ix7455 (.Y (nx7454), .A0 (nx8509), .A1 (nx10190), .A2 (nx11674)) ;
    dffr gen_19_cmp_mRegCmp_reg_Q_4 (.Q (gen_19_cmp_mReg_4), .QB (nx8509), .D (
         window_19__4), .CLK (start), .R (rst)) ;
    nor03_2x ix7453 (.Y (nx7452), .A0 (gen_19_cmp_mReg_4), .A1 (nx10844), .A2 (
             nx11682)) ;
    nand02 ix7489 (.Y (gen_19_cmp_BSCmp_op2_5), .A0 (nx8515), .A1 (nx8521)) ;
    nor02_2x ix8516 (.Y (nx8515), .A0 (nx7484), .A1 (nx7480)) ;
    nor03_2x ix7485 (.Y (nx7484), .A0 (gen_19_cmp_mReg_4), .A1 (nx10196), .A2 (
             nx11650)) ;
    nor03_2x ix7481 (.Y (nx7480), .A0 (nx8509), .A1 (nx11656), .A2 (nx11666)) ;
    nor02_2x ix8522 (.Y (nx8521), .A0 (nx7476), .A1 (nx7474)) ;
    nor03_2x ix7477 (.Y (nx7476), .A0 (nx8525), .A1 (nx10192), .A2 (nx11674)) ;
    dffr gen_19_cmp_mRegCmp_reg_Q_5 (.Q (gen_19_cmp_mReg_5), .QB (nx8525), .D (
         window_19__5), .CLK (start), .R (rst)) ;
    nor03_2x ix7475 (.Y (nx7474), .A0 (gen_19_cmp_mReg_5), .A1 (nx10844), .A2 (
             nx11682)) ;
    nand02 ix7511 (.Y (gen_19_cmp_BSCmp_op2_6), .A0 (nx8531), .A1 (nx8535)) ;
    nor02_2x ix8532 (.Y (nx8531), .A0 (nx7506), .A1 (nx7502)) ;
    nor03_2x ix7507 (.Y (nx7506), .A0 (gen_19_cmp_mReg_5), .A1 (nx10198), .A2 (
             nx11650)) ;
    nor03_2x ix7503 (.Y (nx7502), .A0 (nx8525), .A1 (nx11656), .A2 (nx11666)) ;
    nor02_2x ix8536 (.Y (nx8535), .A0 (nx7498), .A1 (nx7496)) ;
    nor03_2x ix7499 (.Y (nx7498), .A0 (nx8539), .A1 (nx10192), .A2 (nx11674)) ;
    dffr gen_19_cmp_mRegCmp_reg_Q_6 (.Q (gen_19_cmp_mReg_6), .QB (nx8539), .D (
         window_19__6), .CLK (start), .R (rst)) ;
    nor03_2x ix7497 (.Y (nx7496), .A0 (gen_19_cmp_mReg_6), .A1 (nx10844), .A2 (
             nx11682)) ;
    nand02 ix7533 (.Y (gen_19_cmp_BSCmp_op2_7), .A0 (nx8545), .A1 (nx8551)) ;
    nor02_2x ix8546 (.Y (nx8545), .A0 (nx7528), .A1 (nx7524)) ;
    nor03_2x ix7529 (.Y (nx7528), .A0 (gen_19_cmp_mReg_6), .A1 (nx10198), .A2 (
             nx11652)) ;
    nor03_2x ix7525 (.Y (nx7524), .A0 (nx8539), .A1 (nx11658), .A2 (nx11668)) ;
    nor02_2x ix8552 (.Y (nx8551), .A0 (nx7520), .A1 (nx7518)) ;
    nor03_2x ix7521 (.Y (nx7520), .A0 (nx8555), .A1 (nx10192), .A2 (nx11676)) ;
    dffr gen_19_cmp_mRegCmp_reg_Q_7 (.Q (gen_19_cmp_mReg_7), .QB (nx8555), .D (
         window_19__7), .CLK (start), .R (rst)) ;
    nor03_2x ix7519 (.Y (nx7518), .A0 (gen_19_cmp_mReg_7), .A1 (nx10844), .A2 (
             nx11684)) ;
    nand02 ix7555 (.Y (gen_19_cmp_BSCmp_op2_8), .A0 (nx8561), .A1 (nx8565)) ;
    nor02_2x ix8562 (.Y (nx8561), .A0 (nx7550), .A1 (nx7546)) ;
    nor03_2x ix7551 (.Y (nx7550), .A0 (gen_19_cmp_mReg_7), .A1 (nx10198), .A2 (
             nx11652)) ;
    nor03_2x ix7547 (.Y (nx7546), .A0 (nx8555), .A1 (nx11658), .A2 (nx11668)) ;
    nor02_2x ix8566 (.Y (nx8565), .A0 (nx7542), .A1 (nx7540)) ;
    nor03_2x ix7543 (.Y (nx7542), .A0 (nx8569), .A1 (nx10192), .A2 (nx11676)) ;
    dffr gen_19_cmp_mRegCmp_reg_Q_8 (.Q (gen_19_cmp_mReg_8), .QB (nx8569), .D (
         window_19__8), .CLK (start), .R (rst)) ;
    nor03_2x ix7541 (.Y (nx7540), .A0 (gen_19_cmp_mReg_8), .A1 (nx10846), .A2 (
             nx11684)) ;
    nand02 ix7577 (.Y (gen_19_cmp_BSCmp_op2_9), .A0 (nx8575), .A1 (nx8581)) ;
    nor02_2x ix8576 (.Y (nx8575), .A0 (nx7572), .A1 (nx7568)) ;
    nor03_2x ix7573 (.Y (nx7572), .A0 (gen_19_cmp_mReg_8), .A1 (nx10198), .A2 (
             nx11652)) ;
    nor03_2x ix7569 (.Y (nx7568), .A0 (nx8569), .A1 (nx11658), .A2 (nx11668)) ;
    nor02_2x ix8582 (.Y (nx8581), .A0 (nx7564), .A1 (nx7562)) ;
    nor03_2x ix7565 (.Y (nx7564), .A0 (nx8584), .A1 (nx10192), .A2 (nx11676)) ;
    dffr gen_19_cmp_mRegCmp_reg_Q_9 (.Q (gen_19_cmp_mReg_9), .QB (nx8584), .D (
         window_19__9), .CLK (start), .R (rst)) ;
    nor03_2x ix7563 (.Y (nx7562), .A0 (gen_19_cmp_mReg_9), .A1 (nx10846), .A2 (
             nx11684)) ;
    nand02 ix7599 (.Y (gen_19_cmp_BSCmp_op2_10), .A0 (nx8589), .A1 (nx8595)) ;
    nor02_2x ix8590 (.Y (nx8589), .A0 (nx7594), .A1 (nx7590)) ;
    nor03_2x ix7595 (.Y (nx7594), .A0 (gen_19_cmp_mReg_9), .A1 (nx10198), .A2 (
             nx11652)) ;
    nor03_2x ix7591 (.Y (nx7590), .A0 (nx8584), .A1 (nx11658), .A2 (nx11668)) ;
    nor02_2x ix8596 (.Y (nx8595), .A0 (nx7586), .A1 (nx7584)) ;
    nor03_2x ix7587 (.Y (nx7586), .A0 (nx8599), .A1 (nx10192), .A2 (nx11676)) ;
    dffr gen_19_cmp_mRegCmp_reg_Q_10 (.Q (gen_19_cmp_mReg_10), .QB (nx8599), .D (
         window_19__10), .CLK (start), .R (rst)) ;
    nor03_2x ix7585 (.Y (nx7584), .A0 (gen_19_cmp_mReg_10), .A1 (nx10846), .A2 (
             nx11684)) ;
    nand02 ix7621 (.Y (gen_19_cmp_BSCmp_op2_11), .A0 (nx8605), .A1 (nx8609)) ;
    nor02_2x ix8606 (.Y (nx8605), .A0 (nx7616), .A1 (nx7612)) ;
    nor03_2x ix7617 (.Y (nx7616), .A0 (gen_19_cmp_mReg_10), .A1 (nx10198), .A2 (
             nx11652)) ;
    nor03_2x ix7613 (.Y (nx7612), .A0 (nx8599), .A1 (nx11658), .A2 (nx11668)) ;
    nor02_2x ix8610 (.Y (nx8609), .A0 (nx7608), .A1 (nx7606)) ;
    nor03_2x ix7609 (.Y (nx7608), .A0 (nx8613), .A1 (nx10192), .A2 (nx11676)) ;
    dffr gen_19_cmp_mRegCmp_reg_Q_11 (.Q (gen_19_cmp_mReg_11), .QB (nx8613), .D (
         window_19__11), .CLK (start), .R (rst)) ;
    nor03_2x ix7607 (.Y (nx7606), .A0 (gen_19_cmp_mReg_11), .A1 (nx10846), .A2 (
             nx11684)) ;
    nand02 ix7643 (.Y (gen_19_cmp_BSCmp_op2_12), .A0 (nx8619), .A1 (nx8625)) ;
    nor02_2x ix8620 (.Y (nx8619), .A0 (nx7638), .A1 (nx7634)) ;
    nor03_2x ix7639 (.Y (nx7638), .A0 (gen_19_cmp_mReg_11), .A1 (nx10198), .A2 (
             nx11652)) ;
    nor03_2x ix7635 (.Y (nx7634), .A0 (nx8613), .A1 (nx11658), .A2 (nx11668)) ;
    nor02_2x ix8626 (.Y (nx8625), .A0 (nx7630), .A1 (nx7628)) ;
    nor03_2x ix7631 (.Y (nx7630), .A0 (nx8628), .A1 (nx10194), .A2 (nx11676)) ;
    dffr gen_19_cmp_mRegCmp_reg_Q_12 (.Q (gen_19_cmp_mReg_12), .QB (nx8628), .D (
         window_19__12), .CLK (start), .R (rst)) ;
    nor03_2x ix7629 (.Y (nx7628), .A0 (gen_19_cmp_mReg_12), .A1 (nx10846), .A2 (
             nx11684)) ;
    nand02 ix7665 (.Y (gen_19_cmp_BSCmp_op2_13), .A0 (nx8633), .A1 (nx8639)) ;
    nor02_2x ix8634 (.Y (nx8633), .A0 (nx7660), .A1 (nx7656)) ;
    nor03_2x ix7661 (.Y (nx7660), .A0 (gen_19_cmp_mReg_12), .A1 (nx10200), .A2 (
             nx11654)) ;
    nor03_2x ix7657 (.Y (nx7656), .A0 (nx8628), .A1 (nx11658), .A2 (nx11670)) ;
    nor02_2x ix8640 (.Y (nx8639), .A0 (nx7652), .A1 (nx7650)) ;
    nor03_2x ix7653 (.Y (nx7652), .A0 (nx8643), .A1 (nx10194), .A2 (nx11678)) ;
    dffr gen_19_cmp_mRegCmp_reg_Q_13 (.Q (gen_19_cmp_mReg_13), .QB (nx8643), .D (
         window_19__13), .CLK (start), .R (rst)) ;
    nor03_2x ix7651 (.Y (nx7650), .A0 (gen_19_cmp_mReg_13), .A1 (nx10846), .A2 (
             nx11686)) ;
    nand02 ix7687 (.Y (gen_19_cmp_BSCmp_op2_14), .A0 (nx8649), .A1 (nx8653)) ;
    nor02_2x ix8650 (.Y (nx8649), .A0 (nx7682), .A1 (nx7678)) ;
    nor03_2x ix7683 (.Y (nx7682), .A0 (gen_19_cmp_mReg_13), .A1 (nx10200), .A2 (
             nx11654)) ;
    nor03_2x ix7679 (.Y (nx7678), .A0 (nx8643), .A1 (nx11660), .A2 (nx11670)) ;
    nor02_2x ix8654 (.Y (nx8653), .A0 (nx7674), .A1 (nx7672)) ;
    nor03_2x ix7675 (.Y (nx7674), .A0 (nx8657), .A1 (nx10194), .A2 (nx11678)) ;
    dffr gen_19_cmp_mRegCmp_reg_Q_14 (.Q (gen_19_cmp_mReg_14), .QB (nx8657), .D (
         window_19__14), .CLK (start), .R (rst)) ;
    nor03_2x ix7673 (.Y (nx7672), .A0 (gen_19_cmp_mReg_14), .A1 (nx10846), .A2 (
             nx11686)) ;
    nand02 ix7709 (.Y (gen_19_cmp_BSCmp_op2_15), .A0 (nx8663), .A1 (nx8669)) ;
    nor02_2x ix8664 (.Y (nx8663), .A0 (nx7704), .A1 (nx7700)) ;
    nor03_2x ix7705 (.Y (nx7704), .A0 (gen_19_cmp_mReg_14), .A1 (nx10200), .A2 (
             nx11654)) ;
    nor03_2x ix7701 (.Y (nx7700), .A0 (nx8657), .A1 (nx11660), .A2 (nx11670)) ;
    nor02_2x ix8670 (.Y (nx8669), .A0 (nx7696), .A1 (nx7694)) ;
    nor03_2x ix7697 (.Y (nx7696), .A0 (nx8672), .A1 (nx10194), .A2 (nx11678)) ;
    dffr gen_19_cmp_mRegCmp_reg_Q_15 (.Q (gen_19_cmp_mReg_15), .QB (nx8672), .D (
         window_19__15), .CLK (start), .R (rst)) ;
    nor03_2x ix7695 (.Y (nx7694), .A0 (gen_19_cmp_mReg_15), .A1 (nx10848), .A2 (
             nx11686)) ;
    nand02 ix7719 (.Y (gen_19_cmp_BSCmp_op2_16), .A0 (nx8677), .A1 (nx8669)) ;
    nor02_2x ix8678 (.Y (nx8677), .A0 (nx7714), .A1 (nx7710)) ;
    nor03_2x ix7715 (.Y (nx7714), .A0 (gen_19_cmp_mReg_15), .A1 (nx10200), .A2 (
             nx11654)) ;
    nor03_2x ix7711 (.Y (nx7710), .A0 (nx8672), .A1 (nx11660), .A2 (nx11670)) ;
    nand02 ix7787 (.Y (gen_20_cmp_BSCmp_op2_1), .A0 (nx8685), .A1 (nx8703)) ;
    nor02_2x ix8686 (.Y (nx8685), .A0 (nx7782), .A1 (nx7778)) ;
    nor03_2x ix7783 (.Y (nx7782), .A0 (gen_20_cmp_mReg_0), .A1 (nx10184), .A2 (
             nx11690)) ;
    dffr gen_20_cmp_mRegCmp_reg_Q_0 (.Q (gen_20_cmp_mReg_0), .QB (nx8691), .D (
         window_20__0), .CLK (start), .R (rst)) ;
    inv01 ix8695 (.Y (nx8694), .A (gen_20_cmp_pMux_0)) ;
    nor03_2x ix7779 (.Y (nx7778), .A0 (nx8691), .A1 (nx11696), .A2 (nx11706)) ;
    inv02 ix8702 (.Y (nx8701), .A (gen_20_cmp_pMux_2)) ;
    nor02_2x ix8704 (.Y (nx8703), .A0 (nx7768), .A1 (nx7766)) ;
    nor03_2x ix7769 (.Y (nx7768), .A0 (nx8707), .A1 (nx10178), .A2 (nx11714)) ;
    dffr gen_20_cmp_mRegCmp_reg_Q_1 (.Q (gen_20_cmp_mReg_1), .QB (nx8707), .D (
         window_20__1), .CLK (start), .R (rst)) ;
    nor03_2x ix7767 (.Y (nx7766), .A0 (gen_20_cmp_mReg_1), .A1 (nx10850), .A2 (
             nx11722)) ;
    nor03_2x ix7727 (.Y (nx7726), .A0 (nx10184), .A1 (nx8701), .A2 (
             gen_20_cmp_pMux_0)) ;
    nand02 ix7809 (.Y (gen_20_cmp_BSCmp_op2_2), .A0 (nx8718), .A1 (nx8725)) ;
    nor02_2x ix8720 (.Y (nx8718), .A0 (nx7804), .A1 (nx7800)) ;
    nor03_2x ix7805 (.Y (nx7804), .A0 (gen_20_cmp_mReg_1), .A1 (nx10184), .A2 (
             nx11690)) ;
    nor03_2x ix7801 (.Y (nx7800), .A0 (nx8707), .A1 (nx11696), .A2 (nx11706)) ;
    nor02_2x ix8726 (.Y (nx8725), .A0 (nx7796), .A1 (nx7794)) ;
    nor03_2x ix7797 (.Y (nx7796), .A0 (nx8729), .A1 (nx10178), .A2 (nx11714)) ;
    dffr gen_20_cmp_mRegCmp_reg_Q_2 (.Q (gen_20_cmp_mReg_2), .QB (nx8729), .D (
         window_20__2), .CLK (start), .R (rst)) ;
    nor03_2x ix7795 (.Y (nx7794), .A0 (gen_20_cmp_mReg_2), .A1 (nx10850), .A2 (
             nx11722)) ;
    nand02 ix7831 (.Y (gen_20_cmp_BSCmp_op2_3), .A0 (nx8735), .A1 (nx8739)) ;
    nor02_2x ix8736 (.Y (nx8735), .A0 (nx7826), .A1 (nx7822)) ;
    nor03_2x ix7827 (.Y (nx7826), .A0 (gen_20_cmp_mReg_2), .A1 (nx10184), .A2 (
             nx11690)) ;
    nor03_2x ix7823 (.Y (nx7822), .A0 (nx8729), .A1 (nx11696), .A2 (nx11706)) ;
    nor02_2x ix8740 (.Y (nx8739), .A0 (nx7818), .A1 (nx7816)) ;
    nor03_2x ix7819 (.Y (nx7818), .A0 (nx8743), .A1 (nx10178), .A2 (nx11714)) ;
    dffr gen_20_cmp_mRegCmp_reg_Q_3 (.Q (gen_20_cmp_mReg_3), .QB (nx8743), .D (
         window_20__3), .CLK (start), .R (rst)) ;
    nor03_2x ix7817 (.Y (nx7816), .A0 (gen_20_cmp_mReg_3), .A1 (nx10850), .A2 (
             nx11722)) ;
    nand02 ix7853 (.Y (gen_20_cmp_BSCmp_op2_4), .A0 (nx8749), .A1 (nx8753)) ;
    nor02_2x ix8750 (.Y (nx8749), .A0 (nx7848), .A1 (nx7844)) ;
    nor03_2x ix7849 (.Y (nx7848), .A0 (gen_20_cmp_mReg_3), .A1 (nx10184), .A2 (
             nx11690)) ;
    nor03_2x ix7845 (.Y (nx7844), .A0 (nx8743), .A1 (nx11696), .A2 (nx11706)) ;
    nor02_2x ix8754 (.Y (nx8753), .A0 (nx7840), .A1 (nx7838)) ;
    nor03_2x ix7841 (.Y (nx7840), .A0 (nx8757), .A1 (nx10178), .A2 (nx11714)) ;
    dffr gen_20_cmp_mRegCmp_reg_Q_4 (.Q (gen_20_cmp_mReg_4), .QB (nx8757), .D (
         window_20__4), .CLK (start), .R (rst)) ;
    nor03_2x ix7839 (.Y (nx7838), .A0 (gen_20_cmp_mReg_4), .A1 (nx10850), .A2 (
             nx11722)) ;
    nand02 ix7875 (.Y (gen_20_cmp_BSCmp_op2_5), .A0 (nx8761), .A1 (nx8767)) ;
    nor02_2x ix8762 (.Y (nx8761), .A0 (nx7870), .A1 (nx7866)) ;
    nor03_2x ix7871 (.Y (nx7870), .A0 (gen_20_cmp_mReg_4), .A1 (nx10184), .A2 (
             nx11690)) ;
    nor03_2x ix7867 (.Y (nx7866), .A0 (nx8757), .A1 (nx11696), .A2 (nx11706)) ;
    nor02_2x ix8768 (.Y (nx8767), .A0 (nx7862), .A1 (nx7860)) ;
    nor03_2x ix7863 (.Y (nx7862), .A0 (nx8771), .A1 (nx10180), .A2 (nx11714)) ;
    dffr gen_20_cmp_mRegCmp_reg_Q_5 (.Q (gen_20_cmp_mReg_5), .QB (nx8771), .D (
         window_20__5), .CLK (start), .R (rst)) ;
    nor03_2x ix7861 (.Y (nx7860), .A0 (gen_20_cmp_mReg_5), .A1 (nx10850), .A2 (
             nx11722)) ;
    nand02 ix7897 (.Y (gen_20_cmp_BSCmp_op2_6), .A0 (nx8775), .A1 (nx8781)) ;
    nor02_2x ix8776 (.Y (nx8775), .A0 (nx7892), .A1 (nx7888)) ;
    nor03_2x ix7893 (.Y (nx7892), .A0 (gen_20_cmp_mReg_5), .A1 (nx10186), .A2 (
             nx11690)) ;
    nor03_2x ix7889 (.Y (nx7888), .A0 (nx8771), .A1 (nx11696), .A2 (nx11706)) ;
    nor02_2x ix8782 (.Y (nx8781), .A0 (nx7884), .A1 (nx7882)) ;
    nor03_2x ix7885 (.Y (nx7884), .A0 (nx8784), .A1 (nx10180), .A2 (nx11714)) ;
    dffr gen_20_cmp_mRegCmp_reg_Q_6 (.Q (gen_20_cmp_mReg_6), .QB (nx8784), .D (
         window_20__6), .CLK (start), .R (rst)) ;
    nor03_2x ix7883 (.Y (nx7882), .A0 (gen_20_cmp_mReg_6), .A1 (nx10850), .A2 (
             nx11722)) ;
    nand02 ix7919 (.Y (gen_20_cmp_BSCmp_op2_7), .A0 (nx8791), .A1 (nx8797)) ;
    nor02_2x ix8792 (.Y (nx8791), .A0 (nx7914), .A1 (nx7910)) ;
    nor03_2x ix7915 (.Y (nx7914), .A0 (gen_20_cmp_mReg_6), .A1 (nx10186), .A2 (
             nx11692)) ;
    nor03_2x ix7911 (.Y (nx7910), .A0 (nx8784), .A1 (nx11698), .A2 (nx11708)) ;
    nor02_2x ix8798 (.Y (nx8797), .A0 (nx7906), .A1 (nx7904)) ;
    nor03_2x ix7907 (.Y (nx7906), .A0 (nx8801), .A1 (nx10180), .A2 (nx11716)) ;
    dffr gen_20_cmp_mRegCmp_reg_Q_7 (.Q (gen_20_cmp_mReg_7), .QB (nx8801), .D (
         window_20__7), .CLK (start), .R (rst)) ;
    nor03_2x ix7905 (.Y (nx7904), .A0 (gen_20_cmp_mReg_7), .A1 (nx10850), .A2 (
             nx11724)) ;
    nand02 ix7941 (.Y (gen_20_cmp_BSCmp_op2_8), .A0 (nx8805), .A1 (nx8811)) ;
    nor02_2x ix8806 (.Y (nx8805), .A0 (nx7936), .A1 (nx7932)) ;
    nor03_2x ix7937 (.Y (nx7936), .A0 (gen_20_cmp_mReg_7), .A1 (nx10186), .A2 (
             nx11692)) ;
    nor03_2x ix7933 (.Y (nx7932), .A0 (nx8801), .A1 (nx11698), .A2 (nx11708)) ;
    nor02_2x ix8812 (.Y (nx8811), .A0 (nx7928), .A1 (nx7926)) ;
    nor03_2x ix7929 (.Y (nx7928), .A0 (nx8815), .A1 (nx10180), .A2 (nx11716)) ;
    dffr gen_20_cmp_mRegCmp_reg_Q_8 (.Q (gen_20_cmp_mReg_8), .QB (nx8815), .D (
         window_20__8), .CLK (start), .R (rst)) ;
    nor03_2x ix7927 (.Y (nx7926), .A0 (gen_20_cmp_mReg_8), .A1 (nx10852), .A2 (
             nx11724)) ;
    nand02 ix7963 (.Y (gen_20_cmp_BSCmp_op2_9), .A0 (nx8819), .A1 (nx8825)) ;
    nor02_2x ix8820 (.Y (nx8819), .A0 (nx7958), .A1 (nx7954)) ;
    nor03_2x ix7959 (.Y (nx7958), .A0 (gen_20_cmp_mReg_8), .A1 (nx10186), .A2 (
             nx11692)) ;
    nor03_2x ix7955 (.Y (nx7954), .A0 (nx8815), .A1 (nx11698), .A2 (nx11708)) ;
    nor02_2x ix8826 (.Y (nx8825), .A0 (nx7950), .A1 (nx7948)) ;
    nor03_2x ix7951 (.Y (nx7950), .A0 (nx8828), .A1 (nx10180), .A2 (nx11716)) ;
    dffr gen_20_cmp_mRegCmp_reg_Q_9 (.Q (gen_20_cmp_mReg_9), .QB (nx8828), .D (
         window_20__9), .CLK (start), .R (rst)) ;
    nor03_2x ix7949 (.Y (nx7948), .A0 (gen_20_cmp_mReg_9), .A1 (nx10852), .A2 (
             nx11724)) ;
    nand02 ix7985 (.Y (gen_20_cmp_BSCmp_op2_10), .A0 (nx8835), .A1 (nx8841)) ;
    nor02_2x ix8836 (.Y (nx8835), .A0 (nx7980), .A1 (nx7976)) ;
    nor03_2x ix7981 (.Y (nx7980), .A0 (gen_20_cmp_mReg_9), .A1 (nx10186), .A2 (
             nx11692)) ;
    nor03_2x ix7977 (.Y (nx7976), .A0 (nx8828), .A1 (nx11698), .A2 (nx11708)) ;
    nor02_2x ix8842 (.Y (nx8841), .A0 (nx7972), .A1 (nx7970)) ;
    nor03_2x ix7973 (.Y (nx7972), .A0 (nx8845), .A1 (nx10180), .A2 (nx11716)) ;
    dffr gen_20_cmp_mRegCmp_reg_Q_10 (.Q (gen_20_cmp_mReg_10), .QB (nx8845), .D (
         window_20__10), .CLK (start), .R (rst)) ;
    nor03_2x ix7971 (.Y (nx7970), .A0 (gen_20_cmp_mReg_10), .A1 (nx10852), .A2 (
             nx11724)) ;
    nand02 ix8007 (.Y (gen_20_cmp_BSCmp_op2_11), .A0 (nx8849), .A1 (nx8855)) ;
    nor02_2x ix8850 (.Y (nx8849), .A0 (nx8002), .A1 (nx7998)) ;
    nor03_2x ix8003 (.Y (nx8002), .A0 (gen_20_cmp_mReg_10), .A1 (nx10186), .A2 (
             nx11692)) ;
    nor03_2x ix7999 (.Y (nx7998), .A0 (nx8845), .A1 (nx11698), .A2 (nx11708)) ;
    nor02_2x ix8856 (.Y (nx8855), .A0 (nx7994), .A1 (nx7992)) ;
    nor03_2x ix7995 (.Y (nx7994), .A0 (nx8859), .A1 (nx10180), .A2 (nx11716)) ;
    dffr gen_20_cmp_mRegCmp_reg_Q_11 (.Q (gen_20_cmp_mReg_11), .QB (nx8859), .D (
         window_20__11), .CLK (start), .R (rst)) ;
    nor03_2x ix7993 (.Y (nx7992), .A0 (gen_20_cmp_mReg_11), .A1 (nx10852), .A2 (
             nx11724)) ;
    nand02 ix8029 (.Y (gen_20_cmp_BSCmp_op2_12), .A0 (nx8863), .A1 (nx8869)) ;
    nor02_2x ix8864 (.Y (nx8863), .A0 (nx8024), .A1 (nx8020)) ;
    nor03_2x ix8025 (.Y (nx8024), .A0 (gen_20_cmp_mReg_11), .A1 (nx10186), .A2 (
             nx11692)) ;
    nor03_2x ix8021 (.Y (nx8020), .A0 (nx8859), .A1 (nx11698), .A2 (nx11708)) ;
    nor02_2x ix8870 (.Y (nx8869), .A0 (nx8016), .A1 (nx8014)) ;
    nor03_2x ix8017 (.Y (nx8016), .A0 (nx8873), .A1 (nx10182), .A2 (nx11716)) ;
    dffr gen_20_cmp_mRegCmp_reg_Q_12 (.Q (gen_20_cmp_mReg_12), .QB (nx8873), .D (
         window_20__12), .CLK (start), .R (rst)) ;
    nor03_2x ix8015 (.Y (nx8014), .A0 (gen_20_cmp_mReg_12), .A1 (nx10852), .A2 (
             nx11724)) ;
    nand02 ix8051 (.Y (gen_20_cmp_BSCmp_op2_13), .A0 (nx8879), .A1 (nx8885)) ;
    nor02_2x ix8880 (.Y (nx8879), .A0 (nx8046), .A1 (nx8042)) ;
    nor03_2x ix8047 (.Y (nx8046), .A0 (gen_20_cmp_mReg_12), .A1 (nx10188), .A2 (
             nx11694)) ;
    nor03_2x ix8043 (.Y (nx8042), .A0 (nx8873), .A1 (nx11698), .A2 (nx11710)) ;
    nor02_2x ix8886 (.Y (nx8885), .A0 (nx8038), .A1 (nx8036)) ;
    nor03_2x ix8039 (.Y (nx8038), .A0 (nx8888), .A1 (nx10182), .A2 (nx11718)) ;
    dffr gen_20_cmp_mRegCmp_reg_Q_13 (.Q (gen_20_cmp_mReg_13), .QB (nx8888), .D (
         window_20__13), .CLK (start), .R (rst)) ;
    nor03_2x ix8037 (.Y (nx8036), .A0 (gen_20_cmp_mReg_13), .A1 (nx10852), .A2 (
             nx11726)) ;
    nand02 ix8073 (.Y (gen_20_cmp_BSCmp_op2_14), .A0 (nx8892), .A1 (nx8897)) ;
    nor02_2x ix8893 (.Y (nx8892), .A0 (nx8068), .A1 (nx8064)) ;
    nor03_2x ix8069 (.Y (nx8068), .A0 (gen_20_cmp_mReg_13), .A1 (nx10188), .A2 (
             nx11694)) ;
    nor03_2x ix8065 (.Y (nx8064), .A0 (nx8888), .A1 (nx11700), .A2 (nx11710)) ;
    nor02_2x ix8898 (.Y (nx8897), .A0 (nx8060), .A1 (nx8058)) ;
    nor03_2x ix8061 (.Y (nx8060), .A0 (nx8901), .A1 (nx10182), .A2 (nx11718)) ;
    dffr gen_20_cmp_mRegCmp_reg_Q_14 (.Q (gen_20_cmp_mReg_14), .QB (nx8901), .D (
         window_20__14), .CLK (start), .R (rst)) ;
    nor03_2x ix8059 (.Y (nx8058), .A0 (gen_20_cmp_mReg_14), .A1 (nx10852), .A2 (
             nx11726)) ;
    nand02 ix8095 (.Y (gen_20_cmp_BSCmp_op2_15), .A0 (nx8907), .A1 (nx8913)) ;
    nor02_2x ix8908 (.Y (nx8907), .A0 (nx8090), .A1 (nx8086)) ;
    nor03_2x ix8091 (.Y (nx8090), .A0 (gen_20_cmp_mReg_14), .A1 (nx10188), .A2 (
             nx11694)) ;
    nor03_2x ix8087 (.Y (nx8086), .A0 (nx8901), .A1 (nx11700), .A2 (nx11710)) ;
    nor02_2x ix8914 (.Y (nx8913), .A0 (nx8082), .A1 (nx8080)) ;
    nor03_2x ix8083 (.Y (nx8082), .A0 (nx8917), .A1 (nx10182), .A2 (nx11718)) ;
    dffr gen_20_cmp_mRegCmp_reg_Q_15 (.Q (gen_20_cmp_mReg_15), .QB (nx8917), .D (
         window_20__15), .CLK (start), .R (rst)) ;
    nor03_2x ix8081 (.Y (nx8080), .A0 (gen_20_cmp_mReg_15), .A1 (nx10854), .A2 (
             nx11726)) ;
    nand02 ix8105 (.Y (gen_20_cmp_BSCmp_op2_16), .A0 (nx8921), .A1 (nx8913)) ;
    nor02_2x ix8922 (.Y (nx8921), .A0 (nx8100), .A1 (nx8096)) ;
    nor03_2x ix8101 (.Y (nx8100), .A0 (gen_20_cmp_mReg_15), .A1 (nx10188), .A2 (
             nx11694)) ;
    nor03_2x ix8097 (.Y (nx8096), .A0 (nx8917), .A1 (nx11700), .A2 (nx11710)) ;
    nand02 ix8173 (.Y (gen_21_cmp_BSCmp_op2_1), .A0 (nx8929), .A1 (nx8947)) ;
    nor02_2x ix8930 (.Y (nx8929), .A0 (nx8168), .A1 (nx8164)) ;
    nor03_2x ix8169 (.Y (nx8168), .A0 (gen_21_cmp_mReg_0), .A1 (nx10172), .A2 (
             nx11730)) ;
    dffr gen_21_cmp_mRegCmp_reg_Q_0 (.Q (gen_21_cmp_mReg_0), .QB (nx8933), .D (
         window_21__0), .CLK (start), .R (rst)) ;
    inv01 ix8938 (.Y (nx8937), .A (gen_21_cmp_pMux_0)) ;
    nor03_2x ix8165 (.Y (nx8164), .A0 (nx8933), .A1 (nx11736), .A2 (nx11746)) ;
    inv02 ix8946 (.Y (nx8945), .A (gen_21_cmp_pMux_2)) ;
    nor02_2x ix8948 (.Y (nx8947), .A0 (nx8154), .A1 (nx8152)) ;
    nor03_2x ix8155 (.Y (nx8154), .A0 (nx8950), .A1 (nx10166), .A2 (nx11754)) ;
    dffr gen_21_cmp_mRegCmp_reg_Q_1 (.Q (gen_21_cmp_mReg_1), .QB (nx8950), .D (
         window_21__1), .CLK (start), .R (rst)) ;
    nor03_2x ix8153 (.Y (nx8152), .A0 (gen_21_cmp_mReg_1), .A1 (nx10856), .A2 (
             nx11762)) ;
    nor03_2x ix8113 (.Y (nx8112), .A0 (nx10172), .A1 (nx8945), .A2 (
             gen_21_cmp_pMux_0)) ;
    nand02 ix8195 (.Y (gen_21_cmp_BSCmp_op2_2), .A0 (nx8963), .A1 (nx8969)) ;
    nor02_2x ix8964 (.Y (nx8963), .A0 (nx8190), .A1 (nx8186)) ;
    nor03_2x ix8191 (.Y (nx8190), .A0 (gen_21_cmp_mReg_1), .A1 (nx10172), .A2 (
             nx11730)) ;
    nor03_2x ix8187 (.Y (nx8186), .A0 (nx8950), .A1 (nx11736), .A2 (nx11746)) ;
    nor02_2x ix8970 (.Y (nx8969), .A0 (nx8182), .A1 (nx8180)) ;
    nor03_2x ix8183 (.Y (nx8182), .A0 (nx8972), .A1 (nx10166), .A2 (nx11754)) ;
    dffr gen_21_cmp_mRegCmp_reg_Q_2 (.Q (gen_21_cmp_mReg_2), .QB (nx8972), .D (
         window_21__2), .CLK (start), .R (rst)) ;
    nor03_2x ix8181 (.Y (nx8180), .A0 (gen_21_cmp_mReg_2), .A1 (nx10856), .A2 (
             nx11762)) ;
    nand02 ix8217 (.Y (gen_21_cmp_BSCmp_op2_3), .A0 (nx8979), .A1 (nx8985)) ;
    nor02_2x ix8980 (.Y (nx8979), .A0 (nx8212), .A1 (nx8208)) ;
    nor03_2x ix8213 (.Y (nx8212), .A0 (gen_21_cmp_mReg_2), .A1 (nx10172), .A2 (
             nx11730)) ;
    nor03_2x ix8209 (.Y (nx8208), .A0 (nx8972), .A1 (nx11736), .A2 (nx11746)) ;
    nor02_2x ix8986 (.Y (nx8985), .A0 (nx8204), .A1 (nx8202)) ;
    nor03_2x ix8205 (.Y (nx8204), .A0 (nx8989), .A1 (nx10166), .A2 (nx11754)) ;
    dffr gen_21_cmp_mRegCmp_reg_Q_3 (.Q (gen_21_cmp_mReg_3), .QB (nx8989), .D (
         window_21__3), .CLK (start), .R (rst)) ;
    nor03_2x ix8203 (.Y (nx8202), .A0 (gen_21_cmp_mReg_3), .A1 (nx10856), .A2 (
             nx11762)) ;
    nand02 ix8239 (.Y (gen_21_cmp_BSCmp_op2_4), .A0 (nx8993), .A1 (nx8999)) ;
    nor02_2x ix8994 (.Y (nx8993), .A0 (nx8234), .A1 (nx8230)) ;
    nor03_2x ix8235 (.Y (nx8234), .A0 (gen_21_cmp_mReg_3), .A1 (nx10172), .A2 (
             nx11730)) ;
    nor03_2x ix8231 (.Y (nx8230), .A0 (nx8989), .A1 (nx11736), .A2 (nx11746)) ;
    nor02_2x ix9000 (.Y (nx8999), .A0 (nx8226), .A1 (nx8224)) ;
    nor03_2x ix8227 (.Y (nx8226), .A0 (nx9003), .A1 (nx10166), .A2 (nx11754)) ;
    dffr gen_21_cmp_mRegCmp_reg_Q_4 (.Q (gen_21_cmp_mReg_4), .QB (nx9003), .D (
         window_21__4), .CLK (start), .R (rst)) ;
    nor03_2x ix8225 (.Y (nx8224), .A0 (gen_21_cmp_mReg_4), .A1 (nx10856), .A2 (
             nx11762)) ;
    nand02 ix8261 (.Y (gen_21_cmp_BSCmp_op2_5), .A0 (nx9007), .A1 (nx9013)) ;
    nor02_2x ix9008 (.Y (nx9007), .A0 (nx8256), .A1 (nx8252)) ;
    nor03_2x ix8257 (.Y (nx8256), .A0 (gen_21_cmp_mReg_4), .A1 (nx10172), .A2 (
             nx11730)) ;
    nor03_2x ix8253 (.Y (nx8252), .A0 (nx9003), .A1 (nx11736), .A2 (nx11746)) ;
    nor02_2x ix9014 (.Y (nx9013), .A0 (nx8248), .A1 (nx8246)) ;
    nor03_2x ix8249 (.Y (nx8248), .A0 (nx9016), .A1 (nx10168), .A2 (nx11754)) ;
    dffr gen_21_cmp_mRegCmp_reg_Q_5 (.Q (gen_21_cmp_mReg_5), .QB (nx9016), .D (
         window_21__5), .CLK (start), .R (rst)) ;
    nor03_2x ix8247 (.Y (nx8246), .A0 (gen_21_cmp_mReg_5), .A1 (nx10856), .A2 (
             nx11762)) ;
    nand02 ix8283 (.Y (gen_21_cmp_BSCmp_op2_6), .A0 (nx9023), .A1 (nx9029)) ;
    nor02_2x ix9024 (.Y (nx9023), .A0 (nx8278), .A1 (nx8274)) ;
    nor03_2x ix8279 (.Y (nx8278), .A0 (gen_21_cmp_mReg_5), .A1 (nx10174), .A2 (
             nx11730)) ;
    nor03_2x ix8275 (.Y (nx8274), .A0 (nx9016), .A1 (nx11736), .A2 (nx11746)) ;
    nor02_2x ix9030 (.Y (nx9029), .A0 (nx8270), .A1 (nx8268)) ;
    nor03_2x ix8271 (.Y (nx8270), .A0 (nx9033), .A1 (nx10168), .A2 (nx11754)) ;
    dffr gen_21_cmp_mRegCmp_reg_Q_6 (.Q (gen_21_cmp_mReg_6), .QB (nx9033), .D (
         window_21__6), .CLK (start), .R (rst)) ;
    nor03_2x ix8269 (.Y (nx8268), .A0 (gen_21_cmp_mReg_6), .A1 (nx10856), .A2 (
             nx11762)) ;
    nand02 ix8305 (.Y (gen_21_cmp_BSCmp_op2_7), .A0 (nx9037), .A1 (nx9043)) ;
    nor02_2x ix9038 (.Y (nx9037), .A0 (nx8300), .A1 (nx8296)) ;
    nor03_2x ix8301 (.Y (nx8300), .A0 (gen_21_cmp_mReg_6), .A1 (nx10174), .A2 (
             nx11732)) ;
    nor03_2x ix8297 (.Y (nx8296), .A0 (nx9033), .A1 (nx11738), .A2 (nx11748)) ;
    nor02_2x ix9044 (.Y (nx9043), .A0 (nx8292), .A1 (nx8290)) ;
    nor03_2x ix8293 (.Y (nx8292), .A0 (nx9047), .A1 (nx10168), .A2 (nx11756)) ;
    dffr gen_21_cmp_mRegCmp_reg_Q_7 (.Q (gen_21_cmp_mReg_7), .QB (nx9047), .D (
         window_21__7), .CLK (start), .R (rst)) ;
    nor03_2x ix8291 (.Y (nx8290), .A0 (gen_21_cmp_mReg_7), .A1 (nx10856), .A2 (
             nx11764)) ;
    nand02 ix8327 (.Y (gen_21_cmp_BSCmp_op2_8), .A0 (nx9051), .A1 (nx9057)) ;
    nor02_2x ix9052 (.Y (nx9051), .A0 (nx8322), .A1 (nx8318)) ;
    nor03_2x ix8323 (.Y (nx8322), .A0 (gen_21_cmp_mReg_7), .A1 (nx10174), .A2 (
             nx11732)) ;
    nor03_2x ix8319 (.Y (nx8318), .A0 (nx9047), .A1 (nx11738), .A2 (nx11748)) ;
    nor02_2x ix9058 (.Y (nx9057), .A0 (nx8314), .A1 (nx8312)) ;
    nor03_2x ix8315 (.Y (nx8314), .A0 (nx9060), .A1 (nx10168), .A2 (nx11756)) ;
    dffr gen_21_cmp_mRegCmp_reg_Q_8 (.Q (gen_21_cmp_mReg_8), .QB (nx9060), .D (
         window_21__8), .CLK (start), .R (rst)) ;
    nor03_2x ix8313 (.Y (nx8312), .A0 (gen_21_cmp_mReg_8), .A1 (nx10858), .A2 (
             nx11764)) ;
    nand02 ix8349 (.Y (gen_21_cmp_BSCmp_op2_9), .A0 (nx9067), .A1 (nx9073)) ;
    nor02_2x ix9068 (.Y (nx9067), .A0 (nx8344), .A1 (nx8340)) ;
    nor03_2x ix8345 (.Y (nx8344), .A0 (gen_21_cmp_mReg_8), .A1 (nx10174), .A2 (
             nx11732)) ;
    nor03_2x ix8341 (.Y (nx8340), .A0 (nx9060), .A1 (nx11738), .A2 (nx11748)) ;
    nor02_2x ix9074 (.Y (nx9073), .A0 (nx8336), .A1 (nx8334)) ;
    nor03_2x ix8337 (.Y (nx8336), .A0 (nx9077), .A1 (nx10168), .A2 (nx11756)) ;
    dffr gen_21_cmp_mRegCmp_reg_Q_9 (.Q (gen_21_cmp_mReg_9), .QB (nx9077), .D (
         window_21__9), .CLK (start), .R (rst)) ;
    nor03_2x ix8335 (.Y (nx8334), .A0 (gen_21_cmp_mReg_9), .A1 (nx10858), .A2 (
             nx11764)) ;
    nand02 ix8371 (.Y (gen_21_cmp_BSCmp_op2_10), .A0 (nx9081), .A1 (nx9087)) ;
    nor02_2x ix9082 (.Y (nx9081), .A0 (nx8366), .A1 (nx8362)) ;
    nor03_2x ix8367 (.Y (nx8366), .A0 (gen_21_cmp_mReg_9), .A1 (nx10174), .A2 (
             nx11732)) ;
    nor03_2x ix8363 (.Y (nx8362), .A0 (nx9077), .A1 (nx11738), .A2 (nx11748)) ;
    nor02_2x ix9088 (.Y (nx9087), .A0 (nx8358), .A1 (nx8356)) ;
    nor03_2x ix8359 (.Y (nx8358), .A0 (nx9091), .A1 (nx10168), .A2 (nx11756)) ;
    dffr gen_21_cmp_mRegCmp_reg_Q_10 (.Q (gen_21_cmp_mReg_10), .QB (nx9091), .D (
         window_21__10), .CLK (start), .R (rst)) ;
    nor03_2x ix8357 (.Y (nx8356), .A0 (gen_21_cmp_mReg_10), .A1 (nx10858), .A2 (
             nx11764)) ;
    nand02 ix8393 (.Y (gen_21_cmp_BSCmp_op2_11), .A0 (nx9095), .A1 (nx9101)) ;
    nor02_2x ix9096 (.Y (nx9095), .A0 (nx8388), .A1 (nx8384)) ;
    nor03_2x ix8389 (.Y (nx8388), .A0 (gen_21_cmp_mReg_10), .A1 (nx10174), .A2 (
             nx11732)) ;
    nor03_2x ix8385 (.Y (nx8384), .A0 (nx9091), .A1 (nx11738), .A2 (nx11748)) ;
    nor02_2x ix9102 (.Y (nx9101), .A0 (nx8380), .A1 (nx8378)) ;
    nor03_2x ix8381 (.Y (nx8380), .A0 (nx9104), .A1 (nx10168), .A2 (nx11756)) ;
    dffr gen_21_cmp_mRegCmp_reg_Q_11 (.Q (gen_21_cmp_mReg_11), .QB (nx9104), .D (
         window_21__11), .CLK (start), .R (rst)) ;
    nor03_2x ix8379 (.Y (nx8378), .A0 (gen_21_cmp_mReg_11), .A1 (nx10858), .A2 (
             nx11764)) ;
    nand02 ix8415 (.Y (gen_21_cmp_BSCmp_op2_12), .A0 (nx9111), .A1 (nx9117)) ;
    nor02_2x ix9112 (.Y (nx9111), .A0 (nx8410), .A1 (nx8406)) ;
    nor03_2x ix8411 (.Y (nx8410), .A0 (gen_21_cmp_mReg_11), .A1 (nx10174), .A2 (
             nx11732)) ;
    nor03_2x ix8407 (.Y (nx8406), .A0 (nx9104), .A1 (nx11738), .A2 (nx11748)) ;
    nor02_2x ix9118 (.Y (nx9117), .A0 (nx8402), .A1 (nx8400)) ;
    nor03_2x ix8403 (.Y (nx8402), .A0 (nx9121), .A1 (nx10170), .A2 (nx11756)) ;
    dffr gen_21_cmp_mRegCmp_reg_Q_12 (.Q (gen_21_cmp_mReg_12), .QB (nx9121), .D (
         window_21__12), .CLK (start), .R (rst)) ;
    nor03_2x ix8401 (.Y (nx8400), .A0 (gen_21_cmp_mReg_12), .A1 (nx10858), .A2 (
             nx11764)) ;
    nand02 ix8437 (.Y (gen_21_cmp_BSCmp_op2_13), .A0 (nx9125), .A1 (nx9131)) ;
    nor02_2x ix9126 (.Y (nx9125), .A0 (nx8432), .A1 (nx8428)) ;
    nor03_2x ix8433 (.Y (nx8432), .A0 (gen_21_cmp_mReg_12), .A1 (nx10176), .A2 (
             nx11734)) ;
    nor03_2x ix8429 (.Y (nx8428), .A0 (nx9121), .A1 (nx11738), .A2 (nx11750)) ;
    nor02_2x ix9132 (.Y (nx9131), .A0 (nx8424), .A1 (nx8422)) ;
    nor03_2x ix8425 (.Y (nx8424), .A0 (nx9135), .A1 (nx10170), .A2 (nx11758)) ;
    dffr gen_21_cmp_mRegCmp_reg_Q_13 (.Q (gen_21_cmp_mReg_13), .QB (nx9135), .D (
         window_21__13), .CLK (start), .R (rst)) ;
    nor03_2x ix8423 (.Y (nx8422), .A0 (gen_21_cmp_mReg_13), .A1 (nx10858), .A2 (
             nx11766)) ;
    nand02 ix8459 (.Y (gen_21_cmp_BSCmp_op2_14), .A0 (nx9139), .A1 (nx9145)) ;
    nor02_2x ix9140 (.Y (nx9139), .A0 (nx8454), .A1 (nx8450)) ;
    nor03_2x ix8455 (.Y (nx8454), .A0 (gen_21_cmp_mReg_13), .A1 (nx10176), .A2 (
             nx11734)) ;
    nor03_2x ix8451 (.Y (nx8450), .A0 (nx9135), .A1 (nx11740), .A2 (nx11750)) ;
    nor02_2x ix9146 (.Y (nx9145), .A0 (nx8446), .A1 (nx8444)) ;
    nor03_2x ix8447 (.Y (nx8446), .A0 (nx9148), .A1 (nx10170), .A2 (nx11758)) ;
    dffr gen_21_cmp_mRegCmp_reg_Q_14 (.Q (gen_21_cmp_mReg_14), .QB (nx9148), .D (
         window_21__14), .CLK (start), .R (rst)) ;
    nor03_2x ix8445 (.Y (nx8444), .A0 (gen_21_cmp_mReg_14), .A1 (nx10858), .A2 (
             nx11766)) ;
    nand02 ix8481 (.Y (gen_21_cmp_BSCmp_op2_15), .A0 (nx9155), .A1 (nx9161)) ;
    nor02_2x ix9156 (.Y (nx9155), .A0 (nx8476), .A1 (nx8472)) ;
    nor03_2x ix8477 (.Y (nx8476), .A0 (gen_21_cmp_mReg_14), .A1 (nx10176), .A2 (
             nx11734)) ;
    nor03_2x ix8473 (.Y (nx8472), .A0 (nx9148), .A1 (nx11740), .A2 (nx11750)) ;
    nor02_2x ix9162 (.Y (nx9161), .A0 (nx8468), .A1 (nx8466)) ;
    nor03_2x ix8469 (.Y (nx8468), .A0 (nx9165), .A1 (nx10170), .A2 (nx11758)) ;
    dffr gen_21_cmp_mRegCmp_reg_Q_15 (.Q (gen_21_cmp_mReg_15), .QB (nx9165), .D (
         window_21__15), .CLK (start), .R (rst)) ;
    nor03_2x ix8467 (.Y (nx8466), .A0 (gen_21_cmp_mReg_15), .A1 (nx10860), .A2 (
             nx11766)) ;
    nand02 ix8491 (.Y (gen_21_cmp_BSCmp_op2_16), .A0 (nx9169), .A1 (nx9161)) ;
    nor02_2x ix9170 (.Y (nx9169), .A0 (nx8486), .A1 (nx8482)) ;
    nor03_2x ix8487 (.Y (nx8486), .A0 (gen_21_cmp_mReg_15), .A1 (nx10176), .A2 (
             nx11734)) ;
    nor03_2x ix8483 (.Y (nx8482), .A0 (nx9165), .A1 (nx11740), .A2 (nx11750)) ;
    nand02 ix8559 (.Y (gen_22_cmp_BSCmp_op2_1), .A0 (nx9177), .A1 (nx9197)) ;
    nor02_2x ix9178 (.Y (nx9177), .A0 (nx8554), .A1 (nx8550)) ;
    nor03_2x ix8555 (.Y (nx8554), .A0 (gen_22_cmp_mReg_0), .A1 (nx10160), .A2 (
             nx11770)) ;
    dffr gen_22_cmp_mRegCmp_reg_Q_0 (.Q (gen_22_cmp_mReg_0), .QB (nx9183), .D (
         window_22__0), .CLK (start), .R (rst)) ;
    inv01 ix9188 (.Y (nx9187), .A (gen_22_cmp_pMux_0)) ;
    nor03_2x ix8551 (.Y (nx8550), .A0 (nx9183), .A1 (nx11776), .A2 (nx11786)) ;
    inv02 ix9196 (.Y (nx9195), .A (gen_22_cmp_pMux_2)) ;
    nor02_2x ix9198 (.Y (nx9197), .A0 (nx8540), .A1 (nx8538)) ;
    nor03_2x ix8541 (.Y (nx8540), .A0 (nx9201), .A1 (nx10154), .A2 (nx11794)) ;
    dffr gen_22_cmp_mRegCmp_reg_Q_1 (.Q (gen_22_cmp_mReg_1), .QB (nx9201), .D (
         window_22__1), .CLK (start), .R (rst)) ;
    nor03_2x ix8539 (.Y (nx8538), .A0 (gen_22_cmp_mReg_1), .A1 (nx10862), .A2 (
             nx11802)) ;
    nor03_2x ix8499 (.Y (nx8498), .A0 (nx10160), .A1 (nx9195), .A2 (
             gen_22_cmp_pMux_0)) ;
    nand02 ix8581 (.Y (gen_22_cmp_BSCmp_op2_2), .A0 (nx9212), .A1 (nx9217)) ;
    nor02_2x ix9213 (.Y (nx9212), .A0 (nx8576), .A1 (nx8572)) ;
    nor03_2x ix8577 (.Y (nx8576), .A0 (gen_22_cmp_mReg_1), .A1 (nx10160), .A2 (
             nx11770)) ;
    nor03_2x ix8573 (.Y (nx8572), .A0 (nx9201), .A1 (nx11776), .A2 (nx11786)) ;
    nor02_2x ix9218 (.Y (nx9217), .A0 (nx8568), .A1 (nx8566)) ;
    nor03_2x ix8569 (.Y (nx8568), .A0 (nx9221), .A1 (nx10154), .A2 (nx11794)) ;
    dffr gen_22_cmp_mRegCmp_reg_Q_2 (.Q (gen_22_cmp_mReg_2), .QB (nx9221), .D (
         window_22__2), .CLK (start), .R (rst)) ;
    nor03_2x ix8567 (.Y (nx8566), .A0 (gen_22_cmp_mReg_2), .A1 (nx10862), .A2 (
             nx11802)) ;
    nand02 ix8603 (.Y (gen_22_cmp_BSCmp_op2_3), .A0 (nx9227), .A1 (nx9233)) ;
    nor02_2x ix9228 (.Y (nx9227), .A0 (nx8598), .A1 (nx8594)) ;
    nor03_2x ix8599 (.Y (nx8598), .A0 (gen_22_cmp_mReg_2), .A1 (nx10160), .A2 (
             nx11770)) ;
    nor03_2x ix8595 (.Y (nx8594), .A0 (nx9221), .A1 (nx11776), .A2 (nx11786)) ;
    nor02_2x ix9234 (.Y (nx9233), .A0 (nx8590), .A1 (nx8588)) ;
    nor03_2x ix8591 (.Y (nx8590), .A0 (nx9236), .A1 (nx10154), .A2 (nx11794)) ;
    dffr gen_22_cmp_mRegCmp_reg_Q_3 (.Q (gen_22_cmp_mReg_3), .QB (nx9236), .D (
         window_22__3), .CLK (start), .R (rst)) ;
    nor03_2x ix8589 (.Y (nx8588), .A0 (gen_22_cmp_mReg_3), .A1 (nx10862), .A2 (
             nx11802)) ;
    nand02 ix8625 (.Y (gen_22_cmp_BSCmp_op2_4), .A0 (nx9243), .A1 (nx9249)) ;
    nor02_2x ix9244 (.Y (nx9243), .A0 (nx8620), .A1 (nx8616)) ;
    nor03_2x ix8621 (.Y (nx8620), .A0 (gen_22_cmp_mReg_3), .A1 (nx10160), .A2 (
             nx11770)) ;
    nor03_2x ix8617 (.Y (nx8616), .A0 (nx9236), .A1 (nx11776), .A2 (nx11786)) ;
    nor02_2x ix9250 (.Y (nx9249), .A0 (nx8612), .A1 (nx8610)) ;
    nor03_2x ix8613 (.Y (nx8612), .A0 (nx9253), .A1 (nx10154), .A2 (nx11794)) ;
    dffr gen_22_cmp_mRegCmp_reg_Q_4 (.Q (gen_22_cmp_mReg_4), .QB (nx9253), .D (
         window_22__4), .CLK (start), .R (rst)) ;
    nor03_2x ix8611 (.Y (nx8610), .A0 (gen_22_cmp_mReg_4), .A1 (nx10862), .A2 (
             nx11802)) ;
    nand02 ix8647 (.Y (gen_22_cmp_BSCmp_op2_5), .A0 (nx9259), .A1 (nx9265)) ;
    nor02_2x ix9260 (.Y (nx9259), .A0 (nx8642), .A1 (nx8638)) ;
    nor03_2x ix8643 (.Y (nx8642), .A0 (gen_22_cmp_mReg_4), .A1 (nx10160), .A2 (
             nx11770)) ;
    nor03_2x ix8639 (.Y (nx8638), .A0 (nx9253), .A1 (nx11776), .A2 (nx11786)) ;
    nor02_2x ix9266 (.Y (nx9265), .A0 (nx8634), .A1 (nx8632)) ;
    nor03_2x ix8635 (.Y (nx8634), .A0 (nx9269), .A1 (nx10156), .A2 (nx11794)) ;
    dffr gen_22_cmp_mRegCmp_reg_Q_5 (.Q (gen_22_cmp_mReg_5), .QB (nx9269), .D (
         window_22__5), .CLK (start), .R (rst)) ;
    nor03_2x ix8633 (.Y (nx8632), .A0 (gen_22_cmp_mReg_5), .A1 (nx10862), .A2 (
             nx11802)) ;
    nand02 ix8669 (.Y (gen_22_cmp_BSCmp_op2_6), .A0 (nx9274), .A1 (nx9278)) ;
    nor02_2x ix9275 (.Y (nx9274), .A0 (nx8664), .A1 (nx8660)) ;
    nor03_2x ix8665 (.Y (nx8664), .A0 (gen_22_cmp_mReg_5), .A1 (nx10162), .A2 (
             nx11770)) ;
    nor03_2x ix8661 (.Y (nx8660), .A0 (nx9269), .A1 (nx11776), .A2 (nx11786)) ;
    nor02_2x ix9279 (.Y (nx9278), .A0 (nx8656), .A1 (nx8654)) ;
    nor03_2x ix8657 (.Y (nx8656), .A0 (nx9281), .A1 (nx10156), .A2 (nx11794)) ;
    dffr gen_22_cmp_mRegCmp_reg_Q_6 (.Q (gen_22_cmp_mReg_6), .QB (nx9281), .D (
         window_22__6), .CLK (start), .R (rst)) ;
    nor03_2x ix8655 (.Y (nx8654), .A0 (gen_22_cmp_mReg_6), .A1 (nx10862), .A2 (
             nx11802)) ;
    nand02 ix8691 (.Y (gen_22_cmp_BSCmp_op2_7), .A0 (nx9287), .A1 (nx9293)) ;
    nor02_2x ix9288 (.Y (nx9287), .A0 (nx8686), .A1 (nx8682)) ;
    nor03_2x ix8687 (.Y (nx8686), .A0 (gen_22_cmp_mReg_6), .A1 (nx10162), .A2 (
             nx11772)) ;
    nor03_2x ix8683 (.Y (nx8682), .A0 (nx9281), .A1 (nx11778), .A2 (nx11788)) ;
    nor02_2x ix9294 (.Y (nx9293), .A0 (nx8678), .A1 (nx8676)) ;
    nor03_2x ix8679 (.Y (nx8678), .A0 (nx9297), .A1 (nx10156), .A2 (nx11796)) ;
    dffr gen_22_cmp_mRegCmp_reg_Q_7 (.Q (gen_22_cmp_mReg_7), .QB (nx9297), .D (
         window_22__7), .CLK (start), .R (rst)) ;
    nor03_2x ix8677 (.Y (nx8676), .A0 (gen_22_cmp_mReg_7), .A1 (nx10862), .A2 (
             nx11804)) ;
    nand02 ix8713 (.Y (gen_22_cmp_BSCmp_op2_8), .A0 (nx9303), .A1 (nx9307)) ;
    nor02_2x ix9304 (.Y (nx9303), .A0 (nx8708), .A1 (nx8704)) ;
    nor03_2x ix8709 (.Y (nx8708), .A0 (gen_22_cmp_mReg_7), .A1 (nx10162), .A2 (
             nx11772)) ;
    nor03_2x ix8705 (.Y (nx8704), .A0 (nx9297), .A1 (nx11778), .A2 (nx11788)) ;
    nor02_2x ix9308 (.Y (nx9307), .A0 (nx8700), .A1 (nx8698)) ;
    nor03_2x ix8701 (.Y (nx8700), .A0 (nx9311), .A1 (nx10156), .A2 (nx11796)) ;
    dffr gen_22_cmp_mRegCmp_reg_Q_8 (.Q (gen_22_cmp_mReg_8), .QB (nx9311), .D (
         window_22__8), .CLK (start), .R (rst)) ;
    nor03_2x ix8699 (.Y (nx8698), .A0 (gen_22_cmp_mReg_8), .A1 (nx10864), .A2 (
             nx11804)) ;
    nand02 ix8735 (.Y (gen_22_cmp_BSCmp_op2_9), .A0 (nx9317), .A1 (nx9323)) ;
    nor02_2x ix9318 (.Y (nx9317), .A0 (nx8730), .A1 (nx8726)) ;
    nor03_2x ix8731 (.Y (nx8730), .A0 (gen_22_cmp_mReg_8), .A1 (nx10162), .A2 (
             nx11772)) ;
    nor03_2x ix8727 (.Y (nx8726), .A0 (nx9311), .A1 (nx11778), .A2 (nx11788)) ;
    nor02_2x ix9324 (.Y (nx9323), .A0 (nx8722), .A1 (nx8720)) ;
    nor03_2x ix8723 (.Y (nx8722), .A0 (nx9327), .A1 (nx10156), .A2 (nx11796)) ;
    dffr gen_22_cmp_mRegCmp_reg_Q_9 (.Q (gen_22_cmp_mReg_9), .QB (nx9327), .D (
         window_22__9), .CLK (start), .R (rst)) ;
    nor03_2x ix8721 (.Y (nx8720), .A0 (gen_22_cmp_mReg_9), .A1 (nx10864), .A2 (
             nx11804)) ;
    nand02 ix8757 (.Y (gen_22_cmp_BSCmp_op2_10), .A0 (nx9333), .A1 (nx9337)) ;
    nor02_2x ix9334 (.Y (nx9333), .A0 (nx8752), .A1 (nx8748)) ;
    nor03_2x ix8753 (.Y (nx8752), .A0 (gen_22_cmp_mReg_9), .A1 (nx10162), .A2 (
             nx11772)) ;
    nor03_2x ix8749 (.Y (nx8748), .A0 (nx9327), .A1 (nx11778), .A2 (nx11788)) ;
    nor02_2x ix9338 (.Y (nx9337), .A0 (nx8744), .A1 (nx8742)) ;
    nor03_2x ix8745 (.Y (nx8744), .A0 (nx9341), .A1 (nx10156), .A2 (nx11796)) ;
    dffr gen_22_cmp_mRegCmp_reg_Q_10 (.Q (gen_22_cmp_mReg_10), .QB (nx9341), .D (
         window_22__10), .CLK (start), .R (rst)) ;
    nor03_2x ix8743 (.Y (nx8742), .A0 (gen_22_cmp_mReg_10), .A1 (nx10864), .A2 (
             nx11804)) ;
    nand02 ix8779 (.Y (gen_22_cmp_BSCmp_op2_11), .A0 (nx9347), .A1 (nx9353)) ;
    nor02_2x ix9348 (.Y (nx9347), .A0 (nx8774), .A1 (nx8770)) ;
    nor03_2x ix8775 (.Y (nx8774), .A0 (gen_22_cmp_mReg_10), .A1 (nx10162), .A2 (
             nx11772)) ;
    nor03_2x ix8771 (.Y (nx8770), .A0 (nx9341), .A1 (nx11778), .A2 (nx11788)) ;
    nor02_2x ix9354 (.Y (nx9353), .A0 (nx8766), .A1 (nx8764)) ;
    nor03_2x ix8767 (.Y (nx8766), .A0 (nx9356), .A1 (nx10156), .A2 (nx11796)) ;
    dffr gen_22_cmp_mRegCmp_reg_Q_11 (.Q (gen_22_cmp_mReg_11), .QB (nx9356), .D (
         window_22__11), .CLK (start), .R (rst)) ;
    nor03_2x ix8765 (.Y (nx8764), .A0 (gen_22_cmp_mReg_11), .A1 (nx10864), .A2 (
             nx11804)) ;
    nand02 ix8801 (.Y (gen_22_cmp_BSCmp_op2_12), .A0 (nx9361), .A1 (nx9367)) ;
    nor02_2x ix9362 (.Y (nx9361), .A0 (nx8796), .A1 (nx8792)) ;
    nor03_2x ix8797 (.Y (nx8796), .A0 (gen_22_cmp_mReg_11), .A1 (nx10162), .A2 (
             nx11772)) ;
    nor03_2x ix8793 (.Y (nx8792), .A0 (nx9356), .A1 (nx11778), .A2 (nx11788)) ;
    nor02_2x ix9368 (.Y (nx9367), .A0 (nx8788), .A1 (nx8786)) ;
    nor03_2x ix8789 (.Y (nx8788), .A0 (nx9371), .A1 (nx10158), .A2 (nx11796)) ;
    dffr gen_22_cmp_mRegCmp_reg_Q_12 (.Q (gen_22_cmp_mReg_12), .QB (nx9371), .D (
         window_22__12), .CLK (start), .R (rst)) ;
    nor03_2x ix8787 (.Y (nx8786), .A0 (gen_22_cmp_mReg_12), .A1 (nx10864), .A2 (
             nx11804)) ;
    nand02 ix8823 (.Y (gen_22_cmp_BSCmp_op2_13), .A0 (nx9377), .A1 (nx9381)) ;
    nor02_2x ix9378 (.Y (nx9377), .A0 (nx8818), .A1 (nx8814)) ;
    nor03_2x ix8819 (.Y (nx8818), .A0 (gen_22_cmp_mReg_12), .A1 (nx10164), .A2 (
             nx11774)) ;
    nor03_2x ix8815 (.Y (nx8814), .A0 (nx9371), .A1 (nx11778), .A2 (nx11790)) ;
    nor02_2x ix9382 (.Y (nx9381), .A0 (nx8810), .A1 (nx8808)) ;
    nor03_2x ix8811 (.Y (nx8810), .A0 (nx9385), .A1 (nx10158), .A2 (nx11798)) ;
    dffr gen_22_cmp_mRegCmp_reg_Q_13 (.Q (gen_22_cmp_mReg_13), .QB (nx9385), .D (
         window_22__13), .CLK (start), .R (rst)) ;
    nor03_2x ix8809 (.Y (nx8808), .A0 (gen_22_cmp_mReg_13), .A1 (nx10864), .A2 (
             nx11806)) ;
    nand02 ix8845 (.Y (gen_22_cmp_BSCmp_op2_14), .A0 (nx9391), .A1 (nx9397)) ;
    nor02_2x ix9392 (.Y (nx9391), .A0 (nx8840), .A1 (nx8836)) ;
    nor03_2x ix8841 (.Y (nx8840), .A0 (gen_22_cmp_mReg_13), .A1 (nx10164), .A2 (
             nx11774)) ;
    nor03_2x ix8837 (.Y (nx8836), .A0 (nx9385), .A1 (nx11780), .A2 (nx11790)) ;
    nor02_2x ix9398 (.Y (nx9397), .A0 (nx8832), .A1 (nx8830)) ;
    nor03_2x ix8833 (.Y (nx8832), .A0 (nx9400), .A1 (nx10158), .A2 (nx11798)) ;
    dffr gen_22_cmp_mRegCmp_reg_Q_14 (.Q (gen_22_cmp_mReg_14), .QB (nx9400), .D (
         window_22__14), .CLK (start), .R (rst)) ;
    nor03_2x ix8831 (.Y (nx8830), .A0 (gen_22_cmp_mReg_14), .A1 (nx10864), .A2 (
             nx11806)) ;
    nand02 ix8867 (.Y (gen_22_cmp_BSCmp_op2_15), .A0 (nx9405), .A1 (nx9411)) ;
    nor02_2x ix9406 (.Y (nx9405), .A0 (nx8862), .A1 (nx8858)) ;
    nor03_2x ix8863 (.Y (nx8862), .A0 (gen_22_cmp_mReg_14), .A1 (nx10164), .A2 (
             nx11774)) ;
    nor03_2x ix8859 (.Y (nx8858), .A0 (nx9400), .A1 (nx11780), .A2 (nx11790)) ;
    nor02_2x ix9412 (.Y (nx9411), .A0 (nx8854), .A1 (nx8852)) ;
    nor03_2x ix8855 (.Y (nx8854), .A0 (nx9415), .A1 (nx10158), .A2 (nx11798)) ;
    dffr gen_22_cmp_mRegCmp_reg_Q_15 (.Q (gen_22_cmp_mReg_15), .QB (nx9415), .D (
         window_22__15), .CLK (start), .R (rst)) ;
    nor03_2x ix8853 (.Y (nx8852), .A0 (gen_22_cmp_mReg_15), .A1 (nx10866), .A2 (
             nx11806)) ;
    nand02 ix8877 (.Y (gen_22_cmp_BSCmp_op2_16), .A0 (nx9421), .A1 (nx9411)) ;
    nor02_2x ix9422 (.Y (nx9421), .A0 (nx8872), .A1 (nx8868)) ;
    nor03_2x ix8873 (.Y (nx8872), .A0 (gen_22_cmp_mReg_15), .A1 (nx10164), .A2 (
             nx11774)) ;
    nor03_2x ix8869 (.Y (nx8868), .A0 (nx9415), .A1 (nx11780), .A2 (nx11790)) ;
    nand02 ix8945 (.Y (gen_23_cmp_BSCmp_op2_1), .A0 (nx9427), .A1 (nx9447)) ;
    nor02_2x ix9428 (.Y (nx9427), .A0 (nx8940), .A1 (nx8936)) ;
    nor03_2x ix8941 (.Y (nx8940), .A0 (gen_23_cmp_mReg_0), .A1 (nx10148), .A2 (
             nx11810)) ;
    dffr gen_23_cmp_mRegCmp_reg_Q_0 (.Q (gen_23_cmp_mReg_0), .QB (nx9433), .D (
         window_23__0), .CLK (start), .R (rst)) ;
    inv01 ix9438 (.Y (nx9437), .A (gen_23_cmp_pMux_0)) ;
    nor03_2x ix8937 (.Y (nx8936), .A0 (nx9433), .A1 (nx11816), .A2 (nx11826)) ;
    inv02 ix9446 (.Y (nx9445), .A (gen_23_cmp_pMux_2)) ;
    nor02_2x ix9448 (.Y (nx9447), .A0 (nx8926), .A1 (nx8924)) ;
    nor03_2x ix8927 (.Y (nx8926), .A0 (nx9451), .A1 (nx10142), .A2 (nx11834)) ;
    dffr gen_23_cmp_mRegCmp_reg_Q_1 (.Q (gen_23_cmp_mReg_1), .QB (nx9451), .D (
         window_23__1), .CLK (start), .R (rst)) ;
    nor03_2x ix8925 (.Y (nx8924), .A0 (gen_23_cmp_mReg_1), .A1 (nx10868), .A2 (
             nx11842)) ;
    nor03_2x ix8885 (.Y (nx8884), .A0 (nx10148), .A1 (nx9445), .A2 (
             gen_23_cmp_pMux_0)) ;
    nand02 ix8967 (.Y (gen_23_cmp_BSCmp_op2_2), .A0 (nx9463), .A1 (nx9467)) ;
    nor02_2x ix9464 (.Y (nx9463), .A0 (nx8962), .A1 (nx8958)) ;
    nor03_2x ix8963 (.Y (nx8962), .A0 (gen_23_cmp_mReg_1), .A1 (nx10148), .A2 (
             nx11810)) ;
    nor03_2x ix8959 (.Y (nx8958), .A0 (nx9451), .A1 (nx11816), .A2 (nx11826)) ;
    nor02_2x ix9468 (.Y (nx9467), .A0 (nx8954), .A1 (nx8952)) ;
    nor03_2x ix8955 (.Y (nx8954), .A0 (nx9471), .A1 (nx10142), .A2 (nx11834)) ;
    dffr gen_23_cmp_mRegCmp_reg_Q_2 (.Q (gen_23_cmp_mReg_2), .QB (nx9471), .D (
         window_23__2), .CLK (start), .R (rst)) ;
    nor03_2x ix8953 (.Y (nx8952), .A0 (gen_23_cmp_mReg_2), .A1 (nx10868), .A2 (
             nx11842)) ;
    nand02 ix8989 (.Y (gen_23_cmp_BSCmp_op2_3), .A0 (nx9477), .A1 (nx9481)) ;
    nor02_2x ix9478 (.Y (nx9477), .A0 (nx8984), .A1 (nx8980)) ;
    nor03_2x ix8985 (.Y (nx8984), .A0 (gen_23_cmp_mReg_2), .A1 (nx10148), .A2 (
             nx11810)) ;
    nor03_2x ix8981 (.Y (nx8980), .A0 (nx9471), .A1 (nx11816), .A2 (nx11826)) ;
    nor02_2x ix9482 (.Y (nx9481), .A0 (nx8976), .A1 (nx8974)) ;
    nor03_2x ix8977 (.Y (nx8976), .A0 (nx9485), .A1 (nx10142), .A2 (nx11834)) ;
    dffr gen_23_cmp_mRegCmp_reg_Q_3 (.Q (gen_23_cmp_mReg_3), .QB (nx9485), .D (
         window_23__3), .CLK (start), .R (rst)) ;
    nor03_2x ix8975 (.Y (nx8974), .A0 (gen_23_cmp_mReg_3), .A1 (nx10868), .A2 (
             nx11842)) ;
    nand02 ix9011 (.Y (gen_23_cmp_BSCmp_op2_4), .A0 (nx9489), .A1 (nx9495)) ;
    nor02_2x ix9490 (.Y (nx9489), .A0 (nx9006), .A1 (nx9002)) ;
    nor03_2x ix9007 (.Y (nx9006), .A0 (gen_23_cmp_mReg_3), .A1 (nx10148), .A2 (
             nx11810)) ;
    nor03_2x ix9003 (.Y (nx9002), .A0 (nx9485), .A1 (nx11816), .A2 (nx11826)) ;
    nor02_2x ix9496 (.Y (nx9495), .A0 (nx8998), .A1 (nx8996)) ;
    nor03_2x ix8999 (.Y (nx8998), .A0 (nx9499), .A1 (nx10142), .A2 (nx11834)) ;
    dffr gen_23_cmp_mRegCmp_reg_Q_4 (.Q (gen_23_cmp_mReg_4), .QB (nx9499), .D (
         window_23__4), .CLK (start), .R (rst)) ;
    nor03_2x ix8997 (.Y (nx8996), .A0 (gen_23_cmp_mReg_4), .A1 (nx10868), .A2 (
             nx11842)) ;
    nand02 ix9033 (.Y (gen_23_cmp_BSCmp_op2_5), .A0 (nx9503), .A1 (nx9509)) ;
    nor02_2x ix9504 (.Y (nx9503), .A0 (nx9028), .A1 (nx9024)) ;
    nor03_2x ix9029 (.Y (nx9028), .A0 (gen_23_cmp_mReg_4), .A1 (nx10148), .A2 (
             nx11810)) ;
    nor03_2x ix9025 (.Y (nx9024), .A0 (nx9499), .A1 (nx11816), .A2 (nx11826)) ;
    nor02_2x ix9510 (.Y (nx9509), .A0 (nx9020), .A1 (nx9018)) ;
    nor03_2x ix9021 (.Y (nx9020), .A0 (nx9512), .A1 (nx10144), .A2 (nx11834)) ;
    dffr gen_23_cmp_mRegCmp_reg_Q_5 (.Q (gen_23_cmp_mReg_5), .QB (nx9512), .D (
         window_23__5), .CLK (start), .R (rst)) ;
    nor03_2x ix9019 (.Y (nx9018), .A0 (gen_23_cmp_mReg_5), .A1 (nx10868), .A2 (
             nx11842)) ;
    nand02 ix9055 (.Y (gen_23_cmp_BSCmp_op2_6), .A0 (nx9519), .A1 (nx9525)) ;
    nor02_2x ix9520 (.Y (nx9519), .A0 (nx9050), .A1 (nx9046)) ;
    nor03_2x ix9051 (.Y (nx9050), .A0 (gen_23_cmp_mReg_5), .A1 (nx10150), .A2 (
             nx11810)) ;
    nor03_2x ix9047 (.Y (nx9046), .A0 (nx9512), .A1 (nx11816), .A2 (nx11826)) ;
    nor02_2x ix9526 (.Y (nx9525), .A0 (nx9042), .A1 (nx9040)) ;
    nor03_2x ix9043 (.Y (nx9042), .A0 (nx9529), .A1 (nx10144), .A2 (nx11834)) ;
    dffr gen_23_cmp_mRegCmp_reg_Q_6 (.Q (gen_23_cmp_mReg_6), .QB (nx9529), .D (
         window_23__6), .CLK (start), .R (rst)) ;
    nor03_2x ix9041 (.Y (nx9040), .A0 (gen_23_cmp_mReg_6), .A1 (nx10868), .A2 (
             nx11842)) ;
    nand02 ix9077 (.Y (gen_23_cmp_BSCmp_op2_7), .A0 (nx9533), .A1 (nx9539)) ;
    nor02_2x ix9534 (.Y (nx9533), .A0 (nx9072), .A1 (nx9068)) ;
    nor03_2x ix9073 (.Y (nx9072), .A0 (gen_23_cmp_mReg_6), .A1 (nx10150), .A2 (
             nx11812)) ;
    nor03_2x ix9069 (.Y (nx9068), .A0 (nx9529), .A1 (nx11818), .A2 (nx11828)) ;
    nor02_2x ix9540 (.Y (nx9539), .A0 (nx9064), .A1 (nx9062)) ;
    nor03_2x ix9065 (.Y (nx9064), .A0 (nx9543), .A1 (nx10144), .A2 (nx11836)) ;
    dffr gen_23_cmp_mRegCmp_reg_Q_7 (.Q (gen_23_cmp_mReg_7), .QB (nx9543), .D (
         window_23__7), .CLK (start), .R (rst)) ;
    nor03_2x ix9063 (.Y (nx9062), .A0 (gen_23_cmp_mReg_7), .A1 (nx10868), .A2 (
             nx11844)) ;
    nand02 ix9099 (.Y (gen_23_cmp_BSCmp_op2_8), .A0 (nx9547), .A1 (nx9553)) ;
    nor02_2x ix9548 (.Y (nx9547), .A0 (nx9094), .A1 (nx9090)) ;
    nor03_2x ix9095 (.Y (nx9094), .A0 (gen_23_cmp_mReg_7), .A1 (nx10150), .A2 (
             nx11812)) ;
    nor03_2x ix9091 (.Y (nx9090), .A0 (nx9543), .A1 (nx11818), .A2 (nx11828)) ;
    nor02_2x ix9554 (.Y (nx9553), .A0 (nx9086), .A1 (nx9084)) ;
    nor03_2x ix9087 (.Y (nx9086), .A0 (nx9556), .A1 (nx10144), .A2 (nx11836)) ;
    dffr gen_23_cmp_mRegCmp_reg_Q_8 (.Q (gen_23_cmp_mReg_8), .QB (nx9556), .D (
         window_23__8), .CLK (start), .R (rst)) ;
    nor03_2x ix9085 (.Y (nx9084), .A0 (gen_23_cmp_mReg_8), .A1 (nx10870), .A2 (
             nx11844)) ;
    nand02 ix9121 (.Y (gen_23_cmp_BSCmp_op2_9), .A0 (nx9563), .A1 (nx9569)) ;
    nor02_2x ix9564 (.Y (nx9563), .A0 (nx9116), .A1 (nx9112)) ;
    nor03_2x ix9117 (.Y (nx9116), .A0 (gen_23_cmp_mReg_8), .A1 (nx10150), .A2 (
             nx11812)) ;
    nor03_2x ix9113 (.Y (nx9112), .A0 (nx9556), .A1 (nx11818), .A2 (nx11828)) ;
    nor02_2x ix9570 (.Y (nx9569), .A0 (nx9108), .A1 (nx9106)) ;
    nor03_2x ix9109 (.Y (nx9108), .A0 (nx9573), .A1 (nx10144), .A2 (nx11836)) ;
    dffr gen_23_cmp_mRegCmp_reg_Q_9 (.Q (gen_23_cmp_mReg_9), .QB (nx9573), .D (
         window_23__9), .CLK (start), .R (rst)) ;
    nor03_2x ix9107 (.Y (nx9106), .A0 (gen_23_cmp_mReg_9), .A1 (nx10870), .A2 (
             nx11844)) ;
    nand02 ix9143 (.Y (gen_23_cmp_BSCmp_op2_10), .A0 (nx9577), .A1 (nx9583)) ;
    nor02_2x ix9578 (.Y (nx9577), .A0 (nx9138), .A1 (nx9134)) ;
    nor03_2x ix9139 (.Y (nx9138), .A0 (gen_23_cmp_mReg_9), .A1 (nx10150), .A2 (
             nx11812)) ;
    nor03_2x ix9135 (.Y (nx9134), .A0 (nx9573), .A1 (nx11818), .A2 (nx11828)) ;
    nor02_2x ix9584 (.Y (nx9583), .A0 (nx9130), .A1 (nx9128)) ;
    nor03_2x ix9131 (.Y (nx9130), .A0 (nx9587), .A1 (nx10144), .A2 (nx11836)) ;
    dffr gen_23_cmp_mRegCmp_reg_Q_10 (.Q (gen_23_cmp_mReg_10), .QB (nx9587), .D (
         window_23__10), .CLK (start), .R (rst)) ;
    nor03_2x ix9129 (.Y (nx9128), .A0 (gen_23_cmp_mReg_10), .A1 (nx10870), .A2 (
             nx11844)) ;
    nand02 ix9165 (.Y (gen_23_cmp_BSCmp_op2_11), .A0 (nx9591), .A1 (nx9597)) ;
    nor02_2x ix9592 (.Y (nx9591), .A0 (nx9160), .A1 (nx9156)) ;
    nor03_2x ix9161 (.Y (nx9160), .A0 (gen_23_cmp_mReg_10), .A1 (nx10150), .A2 (
             nx11812)) ;
    nor03_2x ix9157 (.Y (nx9156), .A0 (nx9587), .A1 (nx11818), .A2 (nx11828)) ;
    nor02_2x ix9598 (.Y (nx9597), .A0 (nx9152), .A1 (nx9150)) ;
    nor03_2x ix9153 (.Y (nx9152), .A0 (nx9600), .A1 (nx10144), .A2 (nx11836)) ;
    dffr gen_23_cmp_mRegCmp_reg_Q_11 (.Q (gen_23_cmp_mReg_11), .QB (nx9600), .D (
         window_23__11), .CLK (start), .R (rst)) ;
    nor03_2x ix9151 (.Y (nx9150), .A0 (gen_23_cmp_mReg_11), .A1 (nx10870), .A2 (
             nx11844)) ;
    nand02 ix9187 (.Y (gen_23_cmp_BSCmp_op2_12), .A0 (nx9607), .A1 (nx9613)) ;
    nor02_2x ix9608 (.Y (nx9607), .A0 (nx9182), .A1 (nx9178)) ;
    nor03_2x ix9183 (.Y (nx9182), .A0 (gen_23_cmp_mReg_11), .A1 (nx10150), .A2 (
             nx11812)) ;
    nor03_2x ix9179 (.Y (nx9178), .A0 (nx9600), .A1 (nx11818), .A2 (nx11828)) ;
    nor02_2x ix9614 (.Y (nx9613), .A0 (nx9174), .A1 (nx9172)) ;
    nor03_2x ix9175 (.Y (nx9174), .A0 (nx9617), .A1 (nx10146), .A2 (nx11836)) ;
    dffr gen_23_cmp_mRegCmp_reg_Q_12 (.Q (gen_23_cmp_mReg_12), .QB (nx9617), .D (
         window_23__12), .CLK (start), .R (rst)) ;
    nor03_2x ix9173 (.Y (nx9172), .A0 (gen_23_cmp_mReg_12), .A1 (nx10870), .A2 (
             nx11844)) ;
    nand02 ix9209 (.Y (gen_23_cmp_BSCmp_op2_13), .A0 (nx9621), .A1 (nx9627)) ;
    nor02_2x ix9622 (.Y (nx9621), .A0 (nx9204), .A1 (nx9200)) ;
    nor03_2x ix9205 (.Y (nx9204), .A0 (gen_23_cmp_mReg_12), .A1 (nx10152), .A2 (
             nx11814)) ;
    nor03_2x ix9201 (.Y (nx9200), .A0 (nx9617), .A1 (nx11818), .A2 (nx11830)) ;
    nor02_2x ix9628 (.Y (nx9627), .A0 (nx9196), .A1 (nx9194)) ;
    nor03_2x ix9197 (.Y (nx9196), .A0 (nx9631), .A1 (nx10146), .A2 (nx11838)) ;
    dffr gen_23_cmp_mRegCmp_reg_Q_13 (.Q (gen_23_cmp_mReg_13), .QB (nx9631), .D (
         window_23__13), .CLK (start), .R (rst)) ;
    nor03_2x ix9195 (.Y (nx9194), .A0 (gen_23_cmp_mReg_13), .A1 (nx10870), .A2 (
             nx11846)) ;
    nand02 ix9231 (.Y (gen_23_cmp_BSCmp_op2_14), .A0 (nx9635), .A1 (nx9641)) ;
    nor02_2x ix9636 (.Y (nx9635), .A0 (nx9226), .A1 (nx9222)) ;
    nor03_2x ix9227 (.Y (nx9226), .A0 (gen_23_cmp_mReg_13), .A1 (nx10152), .A2 (
             nx11814)) ;
    nor03_2x ix9223 (.Y (nx9222), .A0 (nx9631), .A1 (nx11820), .A2 (nx11830)) ;
    nor02_2x ix9642 (.Y (nx9641), .A0 (nx9218), .A1 (nx9216)) ;
    nor03_2x ix9219 (.Y (nx9218), .A0 (nx9645), .A1 (nx10146), .A2 (nx11838)) ;
    dffr gen_23_cmp_mRegCmp_reg_Q_14 (.Q (gen_23_cmp_mReg_14), .QB (nx9645), .D (
         window_23__14), .CLK (start), .R (rst)) ;
    nor03_2x ix9217 (.Y (nx9216), .A0 (gen_23_cmp_mReg_14), .A1 (nx10870), .A2 (
             nx11846)) ;
    nand02 ix9253 (.Y (gen_23_cmp_BSCmp_op2_15), .A0 (nx9651), .A1 (nx9655)) ;
    nor02_2x ix9652 (.Y (nx9651), .A0 (nx9248), .A1 (nx9244)) ;
    nor03_2x ix9249 (.Y (nx9248), .A0 (gen_23_cmp_mReg_14), .A1 (nx10152), .A2 (
             nx11814)) ;
    nor03_2x ix9245 (.Y (nx9244), .A0 (nx9645), .A1 (nx11820), .A2 (nx11830)) ;
    nor02_2x ix9656 (.Y (nx9655), .A0 (nx9240), .A1 (nx9238)) ;
    nor03_2x ix9241 (.Y (nx9240), .A0 (nx9658), .A1 (nx10146), .A2 (nx11838)) ;
    dffr gen_23_cmp_mRegCmp_reg_Q_15 (.Q (gen_23_cmp_mReg_15), .QB (nx9658), .D (
         window_23__15), .CLK (start), .R (rst)) ;
    nor03_2x ix9239 (.Y (nx9238), .A0 (gen_23_cmp_mReg_15), .A1 (nx10872), .A2 (
             nx11846)) ;
    nand02 ix9263 (.Y (gen_23_cmp_BSCmp_op2_16), .A0 (nx9663), .A1 (nx9655)) ;
    nor02_2x ix9664 (.Y (nx9663), .A0 (nx9258), .A1 (nx9254)) ;
    nor03_2x ix9259 (.Y (nx9258), .A0 (gen_23_cmp_mReg_15), .A1 (nx10152), .A2 (
             nx11814)) ;
    nor03_2x ix9255 (.Y (nx9254), .A0 (nx9658), .A1 (nx11820), .A2 (nx11830)) ;
    nand02 ix9331 (.Y (gen_24_cmp_BSCmp_op2_1), .A0 (nx9669), .A1 (nx9685)) ;
    nor02_2x ix9670 (.Y (nx9669), .A0 (nx9326), .A1 (nx9322)) ;
    nor03_2x ix9327 (.Y (nx9326), .A0 (gen_24_cmp_mReg_0), .A1 (nx10136), .A2 (
             nx11850)) ;
    dffr gen_24_cmp_mRegCmp_reg_Q_0 (.Q (gen_24_cmp_mReg_0), .QB (nx9673), .D (
         window_24__0), .CLK (start), .R (rst)) ;
    inv01 ix9677 (.Y (nx9676), .A (gen_24_cmp_pMux_0)) ;
    nor03_2x ix9323 (.Y (nx9322), .A0 (nx9673), .A1 (nx11856), .A2 (nx11866)) ;
    inv02 ix9684 (.Y (nx9683), .A (gen_24_cmp_pMux_2)) ;
    nor02_2x ix9686 (.Y (nx9685), .A0 (nx9312), .A1 (nx9310)) ;
    nor03_2x ix9313 (.Y (nx9312), .A0 (nx9688), .A1 (nx10130), .A2 (nx11874)) ;
    dffr gen_24_cmp_mRegCmp_reg_Q_1 (.Q (gen_24_cmp_mReg_1), .QB (nx9688), .D (
         window_24__1), .CLK (start), .R (rst)) ;
    nor03_2x ix9311 (.Y (nx9310), .A0 (gen_24_cmp_mReg_1), .A1 (nx10874), .A2 (
             nx11882)) ;
    nor03_2x ix9271 (.Y (nx9270), .A0 (nx10136), .A1 (nx9683), .A2 (
             gen_24_cmp_pMux_0)) ;
    nand02 ix9353 (.Y (gen_24_cmp_BSCmp_op2_2), .A0 (nx9698), .A1 (nx9702)) ;
    nor02_2x ix9699 (.Y (nx9698), .A0 (nx9348), .A1 (nx9344)) ;
    nor03_2x ix9349 (.Y (nx9348), .A0 (gen_24_cmp_mReg_1), .A1 (nx10136), .A2 (
             nx11850)) ;
    nor03_2x ix9345 (.Y (nx9344), .A0 (nx9688), .A1 (nx11856), .A2 (nx11866)) ;
    nor02_2x ix9703 (.Y (nx9702), .A0 (nx9340), .A1 (nx9338)) ;
    nor03_2x ix9341 (.Y (nx9340), .A0 (nx9705), .A1 (nx10130), .A2 (nx11874)) ;
    dffr gen_24_cmp_mRegCmp_reg_Q_2 (.Q (gen_24_cmp_mReg_2), .QB (nx9705), .D (
         window_24__2), .CLK (start), .R (rst)) ;
    nor03_2x ix9339 (.Y (nx9338), .A0 (gen_24_cmp_mReg_2), .A1 (nx10874), .A2 (
             nx11882)) ;
    nand02 ix9375 (.Y (gen_24_cmp_BSCmp_op2_3), .A0 (nx9709), .A1 (nx9713)) ;
    nor02_2x ix9710 (.Y (nx9709), .A0 (nx9370), .A1 (nx9366)) ;
    nor03_2x ix9371 (.Y (nx9370), .A0 (gen_24_cmp_mReg_2), .A1 (nx10136), .A2 (
             nx11850)) ;
    nor03_2x ix9367 (.Y (nx9366), .A0 (nx9705), .A1 (nx11856), .A2 (nx11866)) ;
    nor02_2x ix9714 (.Y (nx9713), .A0 (nx9362), .A1 (nx9360)) ;
    nor03_2x ix9363 (.Y (nx9362), .A0 (nx9716), .A1 (nx10130), .A2 (nx11874)) ;
    dffr gen_24_cmp_mRegCmp_reg_Q_3 (.Q (gen_24_cmp_mReg_3), .QB (nx9716), .D (
         window_24__3), .CLK (start), .R (rst)) ;
    nor03_2x ix9361 (.Y (nx9360), .A0 (gen_24_cmp_mReg_3), .A1 (nx10874), .A2 (
             nx11882)) ;
    nand02 ix9397 (.Y (gen_24_cmp_BSCmp_op2_4), .A0 (nx9720), .A1 (nx9724)) ;
    nor02_2x ix9721 (.Y (nx9720), .A0 (nx9392), .A1 (nx9388)) ;
    nor03_2x ix9393 (.Y (nx9392), .A0 (gen_24_cmp_mReg_3), .A1 (nx10136), .A2 (
             nx11850)) ;
    nor03_2x ix9389 (.Y (nx9388), .A0 (nx9716), .A1 (nx11856), .A2 (nx11866)) ;
    nor02_2x ix9725 (.Y (nx9724), .A0 (nx9384), .A1 (nx9382)) ;
    nor03_2x ix9385 (.Y (nx9384), .A0 (nx9727), .A1 (nx10130), .A2 (nx11874)) ;
    dffr gen_24_cmp_mRegCmp_reg_Q_4 (.Q (gen_24_cmp_mReg_4), .QB (nx9727), .D (
         window_24__4), .CLK (start), .R (rst)) ;
    nor03_2x ix9383 (.Y (nx9382), .A0 (gen_24_cmp_mReg_4), .A1 (nx10874), .A2 (
             nx11882)) ;
    nand02 ix9419 (.Y (gen_24_cmp_BSCmp_op2_5), .A0 (nx9731), .A1 (nx9735)) ;
    nor02_2x ix9732 (.Y (nx9731), .A0 (nx9414), .A1 (nx9410)) ;
    nor03_2x ix9415 (.Y (nx9414), .A0 (gen_24_cmp_mReg_4), .A1 (nx10136), .A2 (
             nx11850)) ;
    nor03_2x ix9411 (.Y (nx9410), .A0 (nx9727), .A1 (nx11856), .A2 (nx11866)) ;
    nor02_2x ix9736 (.Y (nx9735), .A0 (nx9406), .A1 (nx9404)) ;
    nor03_2x ix9407 (.Y (nx9406), .A0 (nx9738), .A1 (nx10132), .A2 (nx11874)) ;
    dffr gen_24_cmp_mRegCmp_reg_Q_5 (.Q (gen_24_cmp_mReg_5), .QB (nx9738), .D (
         window_24__5), .CLK (start), .R (rst)) ;
    nor03_2x ix9405 (.Y (nx9404), .A0 (gen_24_cmp_mReg_5), .A1 (nx10874), .A2 (
             nx11882)) ;
    nand02 ix9441 (.Y (gen_24_cmp_BSCmp_op2_6), .A0 (nx9742), .A1 (nx9746)) ;
    nor02_2x ix9743 (.Y (nx9742), .A0 (nx9436), .A1 (nx9432)) ;
    nor03_2x ix9437 (.Y (nx9436), .A0 (gen_24_cmp_mReg_5), .A1 (nx10138), .A2 (
             nx11850)) ;
    nor03_2x ix9433 (.Y (nx9432), .A0 (nx9738), .A1 (nx11856), .A2 (nx11866)) ;
    nor02_2x ix9747 (.Y (nx9746), .A0 (nx9428), .A1 (nx9426)) ;
    nor03_2x ix9429 (.Y (nx9428), .A0 (nx9749), .A1 (nx10132), .A2 (nx11874)) ;
    dffr gen_24_cmp_mRegCmp_reg_Q_6 (.Q (gen_24_cmp_mReg_6), .QB (nx9749), .D (
         window_24__6), .CLK (start), .R (rst)) ;
    nor03_2x ix9427 (.Y (nx9426), .A0 (gen_24_cmp_mReg_6), .A1 (nx10874), .A2 (
             nx11882)) ;
    nand02 ix9463 (.Y (gen_24_cmp_BSCmp_op2_7), .A0 (nx9753), .A1 (nx9757)) ;
    nor02_2x ix9754 (.Y (nx9753), .A0 (nx9458), .A1 (nx9454)) ;
    nor03_2x ix9459 (.Y (nx9458), .A0 (gen_24_cmp_mReg_6), .A1 (nx10138), .A2 (
             nx11852)) ;
    nor03_2x ix9455 (.Y (nx9454), .A0 (nx9749), .A1 (nx11858), .A2 (nx11868)) ;
    nor02_2x ix9758 (.Y (nx9757), .A0 (nx9450), .A1 (nx9448)) ;
    nor03_2x ix9451 (.Y (nx9450), .A0 (nx9760), .A1 (nx10132), .A2 (nx11876)) ;
    dffr gen_24_cmp_mRegCmp_reg_Q_7 (.Q (gen_24_cmp_mReg_7), .QB (nx9760), .D (
         window_24__7), .CLK (start), .R (rst)) ;
    nor03_2x ix9449 (.Y (nx9448), .A0 (gen_24_cmp_mReg_7), .A1 (nx10874), .A2 (
             nx11884)) ;
    nand02 ix9485 (.Y (gen_24_cmp_BSCmp_op2_8), .A0 (nx9764), .A1 (nx9768)) ;
    nor02_2x ix9765 (.Y (nx9764), .A0 (nx9480), .A1 (nx9476)) ;
    nor03_2x ix9481 (.Y (nx9480), .A0 (gen_24_cmp_mReg_7), .A1 (nx10138), .A2 (
             nx11852)) ;
    nor03_2x ix9477 (.Y (nx9476), .A0 (nx9760), .A1 (nx11858), .A2 (nx11868)) ;
    nor02_2x ix9769 (.Y (nx9768), .A0 (nx9472), .A1 (nx9470)) ;
    nor03_2x ix9473 (.Y (nx9472), .A0 (nx9771), .A1 (nx10132), .A2 (nx11876)) ;
    dffr gen_24_cmp_mRegCmp_reg_Q_8 (.Q (gen_24_cmp_mReg_8), .QB (nx9771), .D (
         window_24__8), .CLK (start), .R (rst)) ;
    nor03_2x ix9471 (.Y (nx9470), .A0 (gen_24_cmp_mReg_8), .A1 (nx10876), .A2 (
             nx11884)) ;
    nand02 ix9507 (.Y (gen_24_cmp_BSCmp_op2_9), .A0 (nx9775), .A1 (nx9779)) ;
    nor02_2x ix9776 (.Y (nx9775), .A0 (nx9502), .A1 (nx9498)) ;
    nor03_2x ix9503 (.Y (nx9502), .A0 (gen_24_cmp_mReg_8), .A1 (nx10138), .A2 (
             nx11852)) ;
    nor03_2x ix9499 (.Y (nx9498), .A0 (nx9771), .A1 (nx11858), .A2 (nx11868)) ;
    nor02_2x ix9780 (.Y (nx9779), .A0 (nx9494), .A1 (nx9492)) ;
    nor03_2x ix9495 (.Y (nx9494), .A0 (nx9782), .A1 (nx10132), .A2 (nx11876)) ;
    dffr gen_24_cmp_mRegCmp_reg_Q_9 (.Q (gen_24_cmp_mReg_9), .QB (nx9782), .D (
         window_24__9), .CLK (start), .R (rst)) ;
    nor03_2x ix9493 (.Y (nx9492), .A0 (gen_24_cmp_mReg_9), .A1 (nx10876), .A2 (
             nx11884)) ;
    nand02 ix9529 (.Y (gen_24_cmp_BSCmp_op2_10), .A0 (nx9786), .A1 (nx9790)) ;
    nor02_2x ix9787 (.Y (nx9786), .A0 (nx9524), .A1 (nx9520)) ;
    nor03_2x ix9525 (.Y (nx9524), .A0 (gen_24_cmp_mReg_9), .A1 (nx10138), .A2 (
             nx11852)) ;
    nor03_2x ix9521 (.Y (nx9520), .A0 (nx9782), .A1 (nx11858), .A2 (nx11868)) ;
    nor02_2x ix9791 (.Y (nx9790), .A0 (nx9516), .A1 (nx9514)) ;
    nor03_2x ix9517 (.Y (nx9516), .A0 (nx9793), .A1 (nx10132), .A2 (nx11876)) ;
    dffr gen_24_cmp_mRegCmp_reg_Q_10 (.Q (gen_24_cmp_mReg_10), .QB (nx9793), .D (
         window_24__10), .CLK (start), .R (rst)) ;
    nor03_2x ix9515 (.Y (nx9514), .A0 (gen_24_cmp_mReg_10), .A1 (nx10876), .A2 (
             nx11884)) ;
    nand02 ix9551 (.Y (gen_24_cmp_BSCmp_op2_11), .A0 (nx9797), .A1 (nx9801)) ;
    nor02_2x ix9798 (.Y (nx9797), .A0 (nx9546), .A1 (nx9542)) ;
    nor03_2x ix9547 (.Y (nx9546), .A0 (gen_24_cmp_mReg_10), .A1 (nx10138), .A2 (
             nx11852)) ;
    nor03_2x ix9543 (.Y (nx9542), .A0 (nx9793), .A1 (nx11858), .A2 (nx11868)) ;
    nor02_2x ix9802 (.Y (nx9801), .A0 (nx9538), .A1 (nx9536)) ;
    nor03_2x ix9539 (.Y (nx9538), .A0 (nx9804), .A1 (nx10132), .A2 (nx11876)) ;
    dffr gen_24_cmp_mRegCmp_reg_Q_11 (.Q (gen_24_cmp_mReg_11), .QB (nx9804), .D (
         window_24__11), .CLK (start), .R (rst)) ;
    nor03_2x ix9537 (.Y (nx9536), .A0 (gen_24_cmp_mReg_11), .A1 (nx10876), .A2 (
             nx11884)) ;
    nand02 ix9573 (.Y (gen_24_cmp_BSCmp_op2_12), .A0 (nx9808), .A1 (nx9812)) ;
    nor02_2x ix9809 (.Y (nx9808), .A0 (nx9568), .A1 (nx9564)) ;
    nor03_2x ix9569 (.Y (nx9568), .A0 (gen_24_cmp_mReg_11), .A1 (nx10138), .A2 (
             nx11852)) ;
    nor03_2x ix9565 (.Y (nx9564), .A0 (nx9804), .A1 (nx11858), .A2 (nx11868)) ;
    nor02_2x ix9813 (.Y (nx9812), .A0 (nx9560), .A1 (nx9558)) ;
    nor03_2x ix9561 (.Y (nx9560), .A0 (nx9815), .A1 (nx10134), .A2 (nx11876)) ;
    dffr gen_24_cmp_mRegCmp_reg_Q_12 (.Q (gen_24_cmp_mReg_12), .QB (nx9815), .D (
         window_24__12), .CLK (start), .R (rst)) ;
    nor03_2x ix9559 (.Y (nx9558), .A0 (gen_24_cmp_mReg_12), .A1 (nx10876), .A2 (
             nx11884)) ;
    nand02 ix9595 (.Y (gen_24_cmp_BSCmp_op2_13), .A0 (nx9819), .A1 (nx9823)) ;
    nor02_2x ix9820 (.Y (nx9819), .A0 (nx9590), .A1 (nx9586)) ;
    nor03_2x ix9591 (.Y (nx9590), .A0 (gen_24_cmp_mReg_12), .A1 (nx10140), .A2 (
             nx11854)) ;
    nor03_2x ix9587 (.Y (nx9586), .A0 (nx9815), .A1 (nx11858), .A2 (nx11870)) ;
    nor02_2x ix9824 (.Y (nx9823), .A0 (nx9582), .A1 (nx9580)) ;
    nor03_2x ix9583 (.Y (nx9582), .A0 (nx9826), .A1 (nx10134), .A2 (nx11878)) ;
    dffr gen_24_cmp_mRegCmp_reg_Q_13 (.Q (gen_24_cmp_mReg_13), .QB (nx9826), .D (
         window_24__13), .CLK (start), .R (rst)) ;
    nor03_2x ix9581 (.Y (nx9580), .A0 (gen_24_cmp_mReg_13), .A1 (nx10876), .A2 (
             nx11886)) ;
    nand02 ix9617 (.Y (gen_24_cmp_BSCmp_op2_14), .A0 (nx9830), .A1 (nx9834)) ;
    nor02_2x ix9831 (.Y (nx9830), .A0 (nx9612), .A1 (nx9608)) ;
    nor03_2x ix9613 (.Y (nx9612), .A0 (gen_24_cmp_mReg_13), .A1 (nx10140), .A2 (
             nx11854)) ;
    nor03_2x ix9609 (.Y (nx9608), .A0 (nx9826), .A1 (nx11860), .A2 (nx11870)) ;
    nor02_2x ix9835 (.Y (nx9834), .A0 (nx9604), .A1 (nx9602)) ;
    nor03_2x ix9605 (.Y (nx9604), .A0 (nx9837), .A1 (nx10134), .A2 (nx11878)) ;
    dffr gen_24_cmp_mRegCmp_reg_Q_14 (.Q (gen_24_cmp_mReg_14), .QB (nx9837), .D (
         window_24__14), .CLK (start), .R (rst)) ;
    nor03_2x ix9603 (.Y (nx9602), .A0 (gen_24_cmp_mReg_14), .A1 (nx10876), .A2 (
             nx11886)) ;
    nand02 ix9639 (.Y (gen_24_cmp_BSCmp_op2_15), .A0 (nx9841), .A1 (nx9845)) ;
    nor02_2x ix9842 (.Y (nx9841), .A0 (nx9634), .A1 (nx9630)) ;
    nor03_2x ix9635 (.Y (nx9634), .A0 (gen_24_cmp_mReg_14), .A1 (nx10140), .A2 (
             nx11854)) ;
    nor03_2x ix9631 (.Y (nx9630), .A0 (nx9837), .A1 (nx11860), .A2 (nx11870)) ;
    nor02_2x ix9846 (.Y (nx9845), .A0 (nx9626), .A1 (nx9624)) ;
    nor03_2x ix9627 (.Y (nx9626), .A0 (nx9848), .A1 (nx10134), .A2 (nx11878)) ;
    dffr gen_24_cmp_mRegCmp_reg_Q_15 (.Q (gen_24_cmp_mReg_15), .QB (nx9848), .D (
         window_24__15), .CLK (start), .R (rst)) ;
    nor03_2x ix9625 (.Y (nx9624), .A0 (gen_24_cmp_mReg_15), .A1 (nx10878), .A2 (
             nx11886)) ;
    nand02 ix9649 (.Y (gen_24_cmp_BSCmp_op2_16), .A0 (nx9852), .A1 (nx9845)) ;
    nor02_2x ix9853 (.Y (nx9852), .A0 (nx9644), .A1 (nx9640)) ;
    nor03_2x ix9645 (.Y (nx9644), .A0 (gen_24_cmp_mReg_15), .A1 (nx10140), .A2 (
             nx11854)) ;
    nor03_2x ix9641 (.Y (nx9640), .A0 (nx9848), .A1 (nx11860), .A2 (nx11870)) ;
    nor02_2x ix19 (.Y (gen_0_cmp_BSCmp_carryIn), .A0 (nx3769), .A1 (nx9857)) ;
    nor02_2x ix9858 (.Y (nx9857), .A0 (nx10900), .A1 (nx3761)) ;
    nand02 ix39 (.Y (gen_0_cmp_BSCmp_op2_0), .A0 (nx9860), .A1 (nx9864)) ;
    nor02_2x ix9861 (.Y (nx9860), .A0 (nx34), .A1 (nx26)) ;
    nor03_2x ix35 (.Y (nx34), .A0 (nx3757), .A1 (nx10422), .A2 (nx10918)) ;
    nor03_2x ix27 (.Y (nx26), .A0 (gen_0_cmp_mReg_0), .A1 (nx10734), .A2 (
             nx10926)) ;
    nand03 ix9865 (.Y (nx9864), .A0 (nx10900), .A1 (nx10422), .A2 (nx3761)) ;
    nor02_2x ix405 (.Y (gen_1_cmp_BSCmp_carryIn), .A0 (nx4013), .A1 (nx9867)) ;
    nor02_2x ix9868 (.Y (nx9867), .A0 (nx10940), .A1 (nx4005)) ;
    nand02 ix425 (.Y (gen_1_cmp_BSCmp_op2_0), .A0 (nx9870), .A1 (nx9874)) ;
    nor02_2x ix9871 (.Y (nx9870), .A0 (nx420), .A1 (nx412)) ;
    nor03_2x ix421 (.Y (nx420), .A0 (nx4001), .A1 (nx10410), .A2 (nx10958)) ;
    nor03_2x ix413 (.Y (nx412), .A0 (gen_1_cmp_mReg_0), .A1 (nx10740), .A2 (
             nx10966)) ;
    nand03 ix9875 (.Y (nx9874), .A0 (nx10940), .A1 (nx10410), .A2 (nx4005)) ;
    nor02_2x ix791 (.Y (gen_2_cmp_BSCmp_carryIn), .A0 (nx4260), .A1 (nx9877)) ;
    nor02_2x ix9878 (.Y (nx9877), .A0 (nx10980), .A1 (nx4253)) ;
    nand02 ix811 (.Y (gen_2_cmp_BSCmp_op2_0), .A0 (nx9880), .A1 (nx9884)) ;
    nor02_2x ix9881 (.Y (nx9880), .A0 (nx806), .A1 (nx798)) ;
    nor03_2x ix807 (.Y (nx806), .A0 (nx4249), .A1 (nx10398), .A2 (nx10998)) ;
    nor03_2x ix799 (.Y (nx798), .A0 (gen_2_cmp_mReg_0), .A1 (nx10746), .A2 (
             nx11006)) ;
    nand03 ix9885 (.Y (nx9884), .A0 (nx10980), .A1 (nx10398), .A2 (nx4253)) ;
    nor02_2x ix1177 (.Y (gen_3_cmp_BSCmp_carryIn), .A0 (nx4509), .A1 (nx9887)) ;
    nor02_2x ix9888 (.Y (nx9887), .A0 (nx11020), .A1 (nx4501)) ;
    nand02 ix1197 (.Y (gen_3_cmp_BSCmp_op2_0), .A0 (nx9890), .A1 (nx9894)) ;
    nor02_2x ix9891 (.Y (nx9890), .A0 (nx1192), .A1 (nx1184)) ;
    nor03_2x ix1193 (.Y (nx1192), .A0 (nx4497), .A1 (nx10386), .A2 (nx11038)) ;
    nor03_2x ix1185 (.Y (nx1184), .A0 (gen_3_cmp_mReg_0), .A1 (nx10752), .A2 (
             nx11046)) ;
    nand03 ix9895 (.Y (nx9894), .A0 (nx11020), .A1 (nx10386), .A2 (nx4501)) ;
    nor02_2x ix1563 (.Y (gen_4_cmp_BSCmp_carryIn), .A0 (nx4757), .A1 (nx9897)) ;
    nor02_2x ix9898 (.Y (nx9897), .A0 (nx11060), .A1 (nx4748)) ;
    nand02 ix1583 (.Y (gen_4_cmp_BSCmp_op2_0), .A0 (nx9900), .A1 (nx9904)) ;
    nor02_2x ix9901 (.Y (nx9900), .A0 (nx1578), .A1 (nx1570)) ;
    nor03_2x ix1579 (.Y (nx1578), .A0 (nx4745), .A1 (nx10374), .A2 (nx11078)) ;
    nor03_2x ix1571 (.Y (nx1570), .A0 (gen_4_cmp_mReg_0), .A1 (nx10758), .A2 (
             nx11086)) ;
    nand03 ix9905 (.Y (nx9904), .A0 (nx11060), .A1 (nx10374), .A2 (nx4748)) ;
    nor02_2x ix1949 (.Y (gen_5_cmp_BSCmp_carryIn), .A0 (nx5003), .A1 (nx9907)) ;
    nor02_2x ix9908 (.Y (nx9907), .A0 (nx11100), .A1 (nx4995)) ;
    nand02 ix1969 (.Y (gen_5_cmp_BSCmp_op2_0), .A0 (nx9910), .A1 (nx9914)) ;
    nor02_2x ix9911 (.Y (nx9910), .A0 (nx1964), .A1 (nx1956)) ;
    nor03_2x ix1965 (.Y (nx1964), .A0 (nx4991), .A1 (nx10362), .A2 (nx11118)) ;
    nor03_2x ix1957 (.Y (nx1956), .A0 (gen_5_cmp_mReg_0), .A1 (nx10764), .A2 (
             nx11126)) ;
    nand03 ix9915 (.Y (nx9914), .A0 (nx11100), .A1 (nx10362), .A2 (nx4995)) ;
    nor02_2x ix2335 (.Y (gen_6_cmp_BSCmp_carryIn), .A0 (nx5253), .A1 (nx9917)) ;
    nor02_2x ix9918 (.Y (nx9917), .A0 (nx11140), .A1 (nx5244)) ;
    nand02 ix2355 (.Y (gen_6_cmp_BSCmp_op2_0), .A0 (nx9920), .A1 (nx9924)) ;
    nor02_2x ix9921 (.Y (nx9920), .A0 (nx2350), .A1 (nx2342)) ;
    nor03_2x ix2351 (.Y (nx2350), .A0 (nx5241), .A1 (nx10350), .A2 (nx11158)) ;
    nor03_2x ix2343 (.Y (nx2342), .A0 (gen_6_cmp_mReg_0), .A1 (nx10770), .A2 (
             nx11166)) ;
    nand03 ix9925 (.Y (nx9924), .A0 (nx11140), .A1 (nx10350), .A2 (nx5244)) ;
    nor02_2x ix2721 (.Y (gen_7_cmp_BSCmp_carryIn), .A0 (nx5499), .A1 (nx9927)) ;
    nor02_2x ix9928 (.Y (nx9927), .A0 (nx11180), .A1 (nx5491)) ;
    nand02 ix2741 (.Y (gen_7_cmp_BSCmp_op2_0), .A0 (nx9930), .A1 (nx9934)) ;
    nor02_2x ix9931 (.Y (nx9930), .A0 (nx2736), .A1 (nx2728)) ;
    nor03_2x ix2737 (.Y (nx2736), .A0 (nx5487), .A1 (nx10338), .A2 (nx11198)) ;
    nor03_2x ix2729 (.Y (nx2728), .A0 (gen_7_cmp_mReg_0), .A1 (nx10776), .A2 (
             nx11206)) ;
    nand03 ix9935 (.Y (nx9934), .A0 (nx11180), .A1 (nx10338), .A2 (nx5491)) ;
    nor02_2x ix3107 (.Y (gen_8_cmp_BSCmp_carryIn), .A0 (nx5743), .A1 (nx9937)) ;
    nor02_2x ix9938 (.Y (nx9937), .A0 (nx11220), .A1 (nx5735)) ;
    nand02 ix3127 (.Y (gen_8_cmp_BSCmp_op2_0), .A0 (nx9940), .A1 (nx9944)) ;
    nor02_2x ix9941 (.Y (nx9940), .A0 (nx3122), .A1 (nx3114)) ;
    nor03_2x ix3123 (.Y (nx3122), .A0 (nx5731), .A1 (nx10326), .A2 (nx11238)) ;
    nor03_2x ix3115 (.Y (nx3114), .A0 (gen_8_cmp_mReg_0), .A1 (nx10782), .A2 (
             nx11246)) ;
    nand03 ix9945 (.Y (nx9944), .A0 (nx11220), .A1 (nx10326), .A2 (nx5735)) ;
    nor02_2x ix3493 (.Y (gen_9_cmp_BSCmp_carryIn), .A0 (nx5987), .A1 (nx9947)) ;
    nor02_2x ix9948 (.Y (nx9947), .A0 (nx11260), .A1 (nx5979)) ;
    nand02 ix3513 (.Y (gen_9_cmp_BSCmp_op2_0), .A0 (nx9950), .A1 (nx9954)) ;
    nor02_2x ix9951 (.Y (nx9950), .A0 (nx3508), .A1 (nx3500)) ;
    nor03_2x ix3509 (.Y (nx3508), .A0 (nx5975), .A1 (nx10314), .A2 (nx11278)) ;
    nor03_2x ix3501 (.Y (nx3500), .A0 (gen_9_cmp_mReg_0), .A1 (nx10788), .A2 (
             nx11286)) ;
    nand03 ix9955 (.Y (nx9954), .A0 (nx11260), .A1 (nx10314), .A2 (nx5979)) ;
    nor02_2x ix3879 (.Y (gen_10_cmp_BSCmp_carryIn), .A0 (nx6233), .A1 (nx9957)
             ) ;
    nor02_2x ix9958 (.Y (nx9957), .A0 (nx11300), .A1 (nx6225)) ;
    nand02 ix3899 (.Y (gen_10_cmp_BSCmp_op2_0), .A0 (nx9960), .A1 (nx9964)) ;
    nor02_2x ix9961 (.Y (nx9960), .A0 (nx3894), .A1 (nx3886)) ;
    nor03_2x ix3895 (.Y (nx3894), .A0 (nx6221), .A1 (nx10302), .A2 (nx11318)) ;
    nor03_2x ix3887 (.Y (nx3886), .A0 (gen_10_cmp_mReg_0), .A1 (nx10794), .A2 (
             nx11326)) ;
    nand03 ix9965 (.Y (nx9964), .A0 (nx11300), .A1 (nx10302), .A2 (nx6225)) ;
    nor02_2x ix4265 (.Y (gen_11_cmp_BSCmp_carryIn), .A0 (nx6477), .A1 (nx9967)
             ) ;
    nor02_2x ix9968 (.Y (nx9967), .A0 (nx11340), .A1 (nx6468)) ;
    nand02 ix4285 (.Y (gen_11_cmp_BSCmp_op2_0), .A0 (nx9970), .A1 (nx9974)) ;
    nor02_2x ix9971 (.Y (nx9970), .A0 (nx4280), .A1 (nx4272)) ;
    nor03_2x ix4281 (.Y (nx4280), .A0 (nx6465), .A1 (nx10290), .A2 (nx11358)) ;
    nor03_2x ix4273 (.Y (nx4272), .A0 (gen_11_cmp_mReg_0), .A1 (nx10800), .A2 (
             nx11366)) ;
    nand03 ix9975 (.Y (nx9974), .A0 (nx11340), .A1 (nx10290), .A2 (nx6468)) ;
    nor02_2x ix4651 (.Y (gen_12_cmp_BSCmp_carryIn), .A0 (nx6725), .A1 (nx9977)
             ) ;
    nor02_2x ix9978 (.Y (nx9977), .A0 (nx11380), .A1 (nx6717)) ;
    nand02 ix4671 (.Y (gen_12_cmp_BSCmp_op2_0), .A0 (nx9980), .A1 (nx9984)) ;
    nor02_2x ix9981 (.Y (nx9980), .A0 (nx4666), .A1 (nx4658)) ;
    nor03_2x ix4667 (.Y (nx4666), .A0 (nx6713), .A1 (nx10278), .A2 (nx11398)) ;
    nor03_2x ix4659 (.Y (nx4658), .A0 (gen_12_cmp_mReg_0), .A1 (nx10806), .A2 (
             nx11406)) ;
    nand03 ix9985 (.Y (nx9984), .A0 (nx11380), .A1 (nx10278), .A2 (nx6717)) ;
    nor02_2x ix5037 (.Y (gen_13_cmp_BSCmp_carryIn), .A0 (nx6973), .A1 (nx9987)
             ) ;
    nor02_2x ix9988 (.Y (nx9987), .A0 (nx11420), .A1 (nx6965)) ;
    nand02 ix5057 (.Y (gen_13_cmp_BSCmp_op2_0), .A0 (nx9990), .A1 (nx9994)) ;
    nor02_2x ix9991 (.Y (nx9990), .A0 (nx5052), .A1 (nx5044)) ;
    nor03_2x ix5053 (.Y (nx5052), .A0 (nx6961), .A1 (nx10266), .A2 (nx11438)) ;
    nor03_2x ix5045 (.Y (nx5044), .A0 (gen_13_cmp_mReg_0), .A1 (nx10812), .A2 (
             nx11446)) ;
    nand03 ix9995 (.Y (nx9994), .A0 (nx11420), .A1 (nx10266), .A2 (nx6965)) ;
    nor02_2x ix5423 (.Y (gen_14_cmp_BSCmp_carryIn), .A0 (nx7221), .A1 (nx9997)
             ) ;
    nor02_2x ix9998 (.Y (nx9997), .A0 (nx11460), .A1 (nx7213)) ;
    nand02 ix5443 (.Y (gen_14_cmp_BSCmp_op2_0), .A0 (nx10000), .A1 (nx10004)) ;
    nor02_2x ix10001 (.Y (nx10000), .A0 (nx5438), .A1 (nx5430)) ;
    nor03_2x ix5439 (.Y (nx5438), .A0 (nx7209), .A1 (nx10254), .A2 (nx11478)) ;
    nor03_2x ix5431 (.Y (nx5430), .A0 (gen_14_cmp_mReg_0), .A1 (nx10818), .A2 (
             nx11486)) ;
    nand03 ix10005 (.Y (nx10004), .A0 (nx11460), .A1 (nx10254), .A2 (nx7213)) ;
    nor02_2x ix5809 (.Y (gen_15_cmp_BSCmp_carryIn), .A0 (nx7471), .A1 (nx10007)
             ) ;
    nor02_2x ix10008 (.Y (nx10007), .A0 (nx11500), .A1 (nx7463)) ;
    nand02 ix5829 (.Y (gen_15_cmp_BSCmp_op2_0), .A0 (nx10010), .A1 (nx10014)) ;
    nor02_2x ix10011 (.Y (nx10010), .A0 (nx5824), .A1 (nx5816)) ;
    nor03_2x ix5825 (.Y (nx5824), .A0 (nx7459), .A1 (nx10242), .A2 (nx11518)) ;
    nor03_2x ix5817 (.Y (nx5816), .A0 (gen_15_cmp_mReg_0), .A1 (nx10824), .A2 (
             nx11526)) ;
    nand03 ix10015 (.Y (nx10014), .A0 (nx11500), .A1 (nx10242), .A2 (nx7463)) ;
    nor02_2x ix6195 (.Y (gen_16_cmp_BSCmp_carryIn), .A0 (nx7717), .A1 (nx10017)
             ) ;
    nor02_2x ix10018 (.Y (nx10017), .A0 (nx11540), .A1 (nx7709)) ;
    nand02 ix6215 (.Y (gen_16_cmp_BSCmp_op2_0), .A0 (nx10020), .A1 (nx10024)) ;
    nor02_2x ix10021 (.Y (nx10020), .A0 (nx6210), .A1 (nx6202)) ;
    nor03_2x ix6211 (.Y (nx6210), .A0 (nx7705), .A1 (nx10230), .A2 (nx11558)) ;
    nor03_2x ix6203 (.Y (nx6202), .A0 (gen_16_cmp_mReg_0), .A1 (nx10830), .A2 (
             nx11566)) ;
    nand03 ix10025 (.Y (nx10024), .A0 (nx11540), .A1 (nx10230), .A2 (nx7709)) ;
    nor02_2x ix6581 (.Y (gen_17_cmp_BSCmp_carryIn), .A0 (nx7961), .A1 (nx10027)
             ) ;
    nor02_2x ix10028 (.Y (nx10027), .A0 (nx11580), .A1 (nx7953)) ;
    nand02 ix6601 (.Y (gen_17_cmp_BSCmp_op2_0), .A0 (nx10030), .A1 (nx10034)) ;
    nor02_2x ix10031 (.Y (nx10030), .A0 (nx6596), .A1 (nx6588)) ;
    nor03_2x ix6597 (.Y (nx6596), .A0 (nx7949), .A1 (nx10218), .A2 (nx11598)) ;
    nor03_2x ix6589 (.Y (nx6588), .A0 (gen_17_cmp_mReg_0), .A1 (nx10836), .A2 (
             nx11606)) ;
    nand03 ix10035 (.Y (nx10034), .A0 (nx11580), .A1 (nx10218), .A2 (nx7953)) ;
    nor02_2x ix6967 (.Y (gen_18_cmp_BSCmp_carryIn), .A0 (nx8209), .A1 (nx10037)
             ) ;
    nor02_2x ix10038 (.Y (nx10037), .A0 (nx11620), .A1 (nx8200)) ;
    nand02 ix6987 (.Y (gen_18_cmp_BSCmp_op2_0), .A0 (nx10040), .A1 (nx10044)) ;
    nor02_2x ix10041 (.Y (nx10040), .A0 (nx6982), .A1 (nx6974)) ;
    nor03_2x ix6983 (.Y (nx6982), .A0 (nx8197), .A1 (nx10206), .A2 (nx11638)) ;
    nor03_2x ix6975 (.Y (nx6974), .A0 (gen_18_cmp_mReg_0), .A1 (nx10842), .A2 (
             nx11646)) ;
    nand03 ix10045 (.Y (nx10044), .A0 (nx11620), .A1 (nx10206), .A2 (nx8200)) ;
    nor02_2x ix7353 (.Y (gen_19_cmp_BSCmp_carryIn), .A0 (nx8455), .A1 (nx10047)
             ) ;
    nor02_2x ix10048 (.Y (nx10047), .A0 (nx11660), .A1 (nx8447)) ;
    nand02 ix7373 (.Y (gen_19_cmp_BSCmp_op2_0), .A0 (nx10050), .A1 (nx10054)) ;
    nor02_2x ix10051 (.Y (nx10050), .A0 (nx7368), .A1 (nx7360)) ;
    nor03_2x ix7369 (.Y (nx7368), .A0 (nx8443), .A1 (nx10194), .A2 (nx11678)) ;
    nor03_2x ix7361 (.Y (nx7360), .A0 (gen_19_cmp_mReg_0), .A1 (nx10848), .A2 (
             nx11686)) ;
    nand03 ix10055 (.Y (nx10054), .A0 (nx11660), .A1 (nx10194), .A2 (nx8447)) ;
    nor02_2x ix7739 (.Y (gen_20_cmp_BSCmp_carryIn), .A0 (nx8701), .A1 (nx10057)
             ) ;
    nor02_2x ix10058 (.Y (nx10057), .A0 (nx11700), .A1 (nx8694)) ;
    nand02 ix7759 (.Y (gen_20_cmp_BSCmp_op2_0), .A0 (nx10060), .A1 (nx10064)) ;
    nor02_2x ix10061 (.Y (nx10060), .A0 (nx7754), .A1 (nx7746)) ;
    nor03_2x ix7755 (.Y (nx7754), .A0 (nx8691), .A1 (nx10182), .A2 (nx11718)) ;
    nor03_2x ix7747 (.Y (nx7746), .A0 (gen_20_cmp_mReg_0), .A1 (nx10854), .A2 (
             nx11726)) ;
    nand03 ix10065 (.Y (nx10064), .A0 (nx11700), .A1 (nx10182), .A2 (nx8694)) ;
    nor02_2x ix8125 (.Y (gen_21_cmp_BSCmp_carryIn), .A0 (nx8945), .A1 (nx10067)
             ) ;
    nor02_2x ix10068 (.Y (nx10067), .A0 (nx11740), .A1 (nx8937)) ;
    nand02 ix8145 (.Y (gen_21_cmp_BSCmp_op2_0), .A0 (nx10070), .A1 (nx10074)) ;
    nor02_2x ix10071 (.Y (nx10070), .A0 (nx8140), .A1 (nx8132)) ;
    nor03_2x ix8141 (.Y (nx8140), .A0 (nx8933), .A1 (nx10170), .A2 (nx11758)) ;
    nor03_2x ix8133 (.Y (nx8132), .A0 (gen_21_cmp_mReg_0), .A1 (nx10860), .A2 (
             nx11766)) ;
    nand03 ix10075 (.Y (nx10074), .A0 (nx11740), .A1 (nx10170), .A2 (nx8937)) ;
    nor02_2x ix8511 (.Y (gen_22_cmp_BSCmp_carryIn), .A0 (nx9195), .A1 (nx10077)
             ) ;
    nor02_2x ix10078 (.Y (nx10077), .A0 (nx11780), .A1 (nx9187)) ;
    nand02 ix8531 (.Y (gen_22_cmp_BSCmp_op2_0), .A0 (nx10080), .A1 (nx10084)) ;
    nor02_2x ix10081 (.Y (nx10080), .A0 (nx8526), .A1 (nx8518)) ;
    nor03_2x ix8527 (.Y (nx8526), .A0 (nx9183), .A1 (nx10158), .A2 (nx11798)) ;
    nor03_2x ix8519 (.Y (nx8518), .A0 (gen_22_cmp_mReg_0), .A1 (nx10866), .A2 (
             nx11806)) ;
    nand03 ix10085 (.Y (nx10084), .A0 (nx11780), .A1 (nx10158), .A2 (nx9187)) ;
    nor02_2x ix8897 (.Y (gen_23_cmp_BSCmp_carryIn), .A0 (nx9445), .A1 (nx10087)
             ) ;
    nor02_2x ix10088 (.Y (nx10087), .A0 (nx11820), .A1 (nx9437)) ;
    nand02 ix8917 (.Y (gen_23_cmp_BSCmp_op2_0), .A0 (nx10090), .A1 (nx10094)) ;
    nor02_2x ix10091 (.Y (nx10090), .A0 (nx8912), .A1 (nx8904)) ;
    nor03_2x ix8913 (.Y (nx8912), .A0 (nx9433), .A1 (nx10146), .A2 (nx11838)) ;
    nor03_2x ix8905 (.Y (nx8904), .A0 (gen_23_cmp_mReg_0), .A1 (nx10872), .A2 (
             nx11846)) ;
    nand03 ix10095 (.Y (nx10094), .A0 (nx11820), .A1 (nx10146), .A2 (nx9437)) ;
    nor02_2x ix9283 (.Y (gen_24_cmp_BSCmp_carryIn), .A0 (nx9683), .A1 (nx10097)
             ) ;
    nor02_2x ix10098 (.Y (nx10097), .A0 (nx11860), .A1 (nx9676)) ;
    nand02 ix9303 (.Y (gen_24_cmp_BSCmp_op2_0), .A0 (nx10100), .A1 (nx10104)) ;
    nor02_2x ix10101 (.Y (nx10100), .A0 (nx9298), .A1 (nx9290)) ;
    nor03_2x ix9299 (.Y (nx9298), .A0 (nx9673), .A1 (nx10134), .A2 (nx11878)) ;
    nor03_2x ix9291 (.Y (nx9290), .A0 (gen_24_cmp_mReg_0), .A1 (nx10878), .A2 (
             nx11886)) ;
    nand03 ix10105 (.Y (nx10104), .A0 (nx11860), .A1 (nx10134), .A2 (nx9676)) ;
    nor02_2x ix9695 (.Y (working), .A0 (nx10107), .A1 (nx11934)) ;
    dffr firtStartLachCmp_reg_Q_0 (.Q (\$dummy [130]), .QB (nx10107), .D (nx9650
         ), .CLK (start), .R (rst)) ;
    inv01 ix10119 (.Y (nx10120), .A (nx3745)) ;
    inv01 ix10121 (.Y (nx10122), .A (clk)) ;
    inv01 ix10123 (.Y (nx10124), .A (clk)) ;
    inv01 ix10125 (.Y (nx10126), .A (clk)) ;
    inv01 ix10127 (.Y (nx10128), .A (clk)) ;
    inv04 ix10129 (.Y (nx10130), .A (nx9683)) ;
    inv04 ix10131 (.Y (nx10132), .A (nx9683)) ;
    inv04 ix10133 (.Y (nx10134), .A (nx9683)) ;
    inv04 ix10135 (.Y (nx10136), .A (nx11860)) ;
    inv04 ix10137 (.Y (nx10138), .A (nx11860)) ;
    inv04 ix10139 (.Y (nx10140), .A (nx11862)) ;
    inv04 ix10141 (.Y (nx10142), .A (nx9445)) ;
    inv04 ix10143 (.Y (nx10144), .A (nx9445)) ;
    inv04 ix10145 (.Y (nx10146), .A (nx9445)) ;
    inv04 ix10147 (.Y (nx10148), .A (nx11820)) ;
    inv04 ix10149 (.Y (nx10150), .A (nx11820)) ;
    inv04 ix10151 (.Y (nx10152), .A (nx11822)) ;
    inv04 ix10153 (.Y (nx10154), .A (nx9195)) ;
    inv04 ix10155 (.Y (nx10156), .A (nx9195)) ;
    inv04 ix10157 (.Y (nx10158), .A (nx9195)) ;
    inv04 ix10159 (.Y (nx10160), .A (nx11780)) ;
    inv04 ix10161 (.Y (nx10162), .A (nx11780)) ;
    inv04 ix10163 (.Y (nx10164), .A (nx11782)) ;
    inv04 ix10165 (.Y (nx10166), .A (nx8945)) ;
    inv04 ix10167 (.Y (nx10168), .A (nx8945)) ;
    inv04 ix10169 (.Y (nx10170), .A (nx8945)) ;
    inv04 ix10171 (.Y (nx10172), .A (nx11740)) ;
    inv04 ix10173 (.Y (nx10174), .A (nx11740)) ;
    inv04 ix10175 (.Y (nx10176), .A (nx11742)) ;
    inv04 ix10177 (.Y (nx10178), .A (nx8701)) ;
    inv04 ix10179 (.Y (nx10180), .A (nx8701)) ;
    inv04 ix10181 (.Y (nx10182), .A (nx8701)) ;
    inv04 ix10183 (.Y (nx10184), .A (nx11700)) ;
    inv04 ix10185 (.Y (nx10186), .A (nx11700)) ;
    inv04 ix10187 (.Y (nx10188), .A (nx11702)) ;
    inv04 ix10189 (.Y (nx10190), .A (nx8455)) ;
    inv04 ix10191 (.Y (nx10192), .A (nx8455)) ;
    inv04 ix10193 (.Y (nx10194), .A (nx8455)) ;
    inv04 ix10195 (.Y (nx10196), .A (nx11660)) ;
    inv04 ix10197 (.Y (nx10198), .A (nx11660)) ;
    inv04 ix10199 (.Y (nx10200), .A (nx11662)) ;
    inv04 ix10201 (.Y (nx10202), .A (nx8209)) ;
    inv04 ix10203 (.Y (nx10204), .A (nx8209)) ;
    inv04 ix10205 (.Y (nx10206), .A (nx8209)) ;
    inv04 ix10207 (.Y (nx10208), .A (nx11620)) ;
    inv04 ix10209 (.Y (nx10210), .A (nx11620)) ;
    inv04 ix10211 (.Y (nx10212), .A (nx11622)) ;
    inv04 ix10213 (.Y (nx10214), .A (nx7961)) ;
    inv04 ix10215 (.Y (nx10216), .A (nx7961)) ;
    inv04 ix10217 (.Y (nx10218), .A (nx7961)) ;
    inv04 ix10219 (.Y (nx10220), .A (nx11580)) ;
    inv04 ix10221 (.Y (nx10222), .A (nx11580)) ;
    inv04 ix10223 (.Y (nx10224), .A (nx11582)) ;
    inv04 ix10225 (.Y (nx10226), .A (nx7717)) ;
    inv04 ix10227 (.Y (nx10228), .A (nx7717)) ;
    inv04 ix10229 (.Y (nx10230), .A (nx7717)) ;
    inv04 ix10231 (.Y (nx10232), .A (nx11540)) ;
    inv04 ix10233 (.Y (nx10234), .A (nx11540)) ;
    inv04 ix10235 (.Y (nx10236), .A (nx11542)) ;
    inv04 ix10237 (.Y (nx10238), .A (nx7471)) ;
    inv04 ix10239 (.Y (nx10240), .A (nx7471)) ;
    inv04 ix10241 (.Y (nx10242), .A (nx7471)) ;
    inv04 ix10243 (.Y (nx10244), .A (nx11500)) ;
    inv04 ix10245 (.Y (nx10246), .A (nx11500)) ;
    inv04 ix10247 (.Y (nx10248), .A (nx11502)) ;
    inv04 ix10249 (.Y (nx10250), .A (nx7221)) ;
    inv04 ix10251 (.Y (nx10252), .A (nx7221)) ;
    inv04 ix10253 (.Y (nx10254), .A (nx7221)) ;
    inv04 ix10255 (.Y (nx10256), .A (nx11460)) ;
    inv04 ix10257 (.Y (nx10258), .A (nx11460)) ;
    inv04 ix10259 (.Y (nx10260), .A (nx11462)) ;
    inv04 ix10261 (.Y (nx10262), .A (nx6973)) ;
    inv04 ix10263 (.Y (nx10264), .A (nx6973)) ;
    inv04 ix10265 (.Y (nx10266), .A (nx6973)) ;
    inv04 ix10267 (.Y (nx10268), .A (nx11420)) ;
    inv04 ix10269 (.Y (nx10270), .A (nx11420)) ;
    inv04 ix10271 (.Y (nx10272), .A (nx11422)) ;
    inv04 ix10273 (.Y (nx10274), .A (nx6725)) ;
    inv04 ix10275 (.Y (nx10276), .A (nx6725)) ;
    inv04 ix10277 (.Y (nx10278), .A (nx6725)) ;
    inv04 ix10279 (.Y (nx10280), .A (nx11380)) ;
    inv04 ix10281 (.Y (nx10282), .A (nx11380)) ;
    inv04 ix10283 (.Y (nx10284), .A (nx11382)) ;
    inv04 ix10285 (.Y (nx10286), .A (nx6477)) ;
    inv04 ix10287 (.Y (nx10288), .A (nx6477)) ;
    inv04 ix10289 (.Y (nx10290), .A (nx6477)) ;
    inv04 ix10291 (.Y (nx10292), .A (nx11340)) ;
    inv04 ix10293 (.Y (nx10294), .A (nx11340)) ;
    inv04 ix10295 (.Y (nx10296), .A (nx11342)) ;
    inv04 ix10297 (.Y (nx10298), .A (nx6233)) ;
    inv04 ix10299 (.Y (nx10300), .A (nx6233)) ;
    inv04 ix10301 (.Y (nx10302), .A (nx6233)) ;
    inv04 ix10303 (.Y (nx10304), .A (nx11300)) ;
    inv04 ix10305 (.Y (nx10306), .A (nx11300)) ;
    inv04 ix10307 (.Y (nx10308), .A (nx11302)) ;
    inv04 ix10309 (.Y (nx10310), .A (nx5987)) ;
    inv04 ix10311 (.Y (nx10312), .A (nx5987)) ;
    inv04 ix10313 (.Y (nx10314), .A (nx5987)) ;
    inv04 ix10315 (.Y (nx10316), .A (nx11260)) ;
    inv04 ix10317 (.Y (nx10318), .A (nx11260)) ;
    inv04 ix10319 (.Y (nx10320), .A (nx11262)) ;
    inv04 ix10321 (.Y (nx10322), .A (nx5743)) ;
    inv04 ix10323 (.Y (nx10324), .A (nx5743)) ;
    inv04 ix10325 (.Y (nx10326), .A (nx5743)) ;
    inv04 ix10327 (.Y (nx10328), .A (nx11220)) ;
    inv04 ix10329 (.Y (nx10330), .A (nx11220)) ;
    inv04 ix10331 (.Y (nx10332), .A (nx11222)) ;
    inv04 ix10333 (.Y (nx10334), .A (nx5499)) ;
    inv04 ix10335 (.Y (nx10336), .A (nx5499)) ;
    inv04 ix10337 (.Y (nx10338), .A (nx5499)) ;
    inv04 ix10339 (.Y (nx10340), .A (nx11180)) ;
    inv04 ix10341 (.Y (nx10342), .A (nx11180)) ;
    inv04 ix10343 (.Y (nx10344), .A (nx11182)) ;
    inv04 ix10345 (.Y (nx10346), .A (nx5253)) ;
    inv04 ix10347 (.Y (nx10348), .A (nx5253)) ;
    inv04 ix10349 (.Y (nx10350), .A (nx5253)) ;
    inv04 ix10351 (.Y (nx10352), .A (nx11140)) ;
    inv04 ix10353 (.Y (nx10354), .A (nx11140)) ;
    inv04 ix10355 (.Y (nx10356), .A (nx11142)) ;
    inv04 ix10357 (.Y (nx10358), .A (nx5003)) ;
    inv04 ix10359 (.Y (nx10360), .A (nx5003)) ;
    inv04 ix10361 (.Y (nx10362), .A (nx5003)) ;
    inv04 ix10363 (.Y (nx10364), .A (nx11100)) ;
    inv04 ix10365 (.Y (nx10366), .A (nx11100)) ;
    inv04 ix10367 (.Y (nx10368), .A (nx11102)) ;
    inv04 ix10369 (.Y (nx10370), .A (nx4757)) ;
    inv04 ix10371 (.Y (nx10372), .A (nx4757)) ;
    inv04 ix10373 (.Y (nx10374), .A (nx4757)) ;
    inv04 ix10375 (.Y (nx10376), .A (nx11060)) ;
    inv04 ix10377 (.Y (nx10378), .A (nx11060)) ;
    inv04 ix10379 (.Y (nx10380), .A (nx11062)) ;
    inv04 ix10381 (.Y (nx10382), .A (nx4509)) ;
    inv04 ix10383 (.Y (nx10384), .A (nx4509)) ;
    inv04 ix10385 (.Y (nx10386), .A (nx4509)) ;
    inv04 ix10387 (.Y (nx10388), .A (nx11020)) ;
    inv04 ix10389 (.Y (nx10390), .A (nx11020)) ;
    inv04 ix10391 (.Y (nx10392), .A (nx11022)) ;
    inv04 ix10393 (.Y (nx10394), .A (nx4260)) ;
    inv04 ix10395 (.Y (nx10396), .A (nx4260)) ;
    inv04 ix10397 (.Y (nx10398), .A (nx4260)) ;
    inv04 ix10399 (.Y (nx10400), .A (nx10980)) ;
    inv04 ix10401 (.Y (nx10402), .A (nx10980)) ;
    inv04 ix10403 (.Y (nx10404), .A (nx10982)) ;
    inv04 ix10405 (.Y (nx10406), .A (nx4013)) ;
    inv04 ix10407 (.Y (nx10408), .A (nx4013)) ;
    inv04 ix10409 (.Y (nx10410), .A (nx4013)) ;
    inv04 ix10411 (.Y (nx10412), .A (nx10940)) ;
    inv04 ix10413 (.Y (nx10414), .A (nx10940)) ;
    inv04 ix10415 (.Y (nx10416), .A (nx10942)) ;
    inv04 ix10417 (.Y (nx10418), .A (nx3769)) ;
    inv04 ix10419 (.Y (nx10420), .A (nx3769)) ;
    inv04 ix10421 (.Y (nx10422), .A (nx3769)) ;
    inv04 ix10423 (.Y (nx10424), .A (nx10900)) ;
    inv04 ix10425 (.Y (nx10426), .A (nx10900)) ;
    inv04 ix10427 (.Y (nx10428), .A (nx10902)) ;
    inv01 ix10429 (.Y (nx10430), .A (gen_24_cmp_BSCmp_op2_16)) ;
    inv02 ix10431 (.Y (nx10432), .A (nx10430)) ;
    inv02 ix10433 (.Y (nx10434), .A (nx10430)) ;
    inv02 ix10435 (.Y (nx10436), .A (nx10430)) ;
    inv02 ix10437 (.Y (nx10438), .A (nx10430)) ;
    inv02 ix10439 (.Y (nx10440), .A (nx10430)) ;
    inv01 ix10441 (.Y (nx10442), .A (gen_23_cmp_BSCmp_op2_16)) ;
    inv02 ix10443 (.Y (nx10444), .A (nx10442)) ;
    inv02 ix10445 (.Y (nx10446), .A (nx10442)) ;
    inv02 ix10447 (.Y (nx10448), .A (nx10442)) ;
    inv02 ix10449 (.Y (nx10450), .A (nx10442)) ;
    inv02 ix10451 (.Y (nx10452), .A (nx10442)) ;
    inv01 ix10453 (.Y (nx10454), .A (gen_22_cmp_BSCmp_op2_16)) ;
    inv02 ix10455 (.Y (nx10456), .A (nx10454)) ;
    inv02 ix10457 (.Y (nx10458), .A (nx10454)) ;
    inv02 ix10459 (.Y (nx10460), .A (nx10454)) ;
    inv02 ix10461 (.Y (nx10462), .A (nx10454)) ;
    inv02 ix10463 (.Y (nx10464), .A (nx10454)) ;
    inv01 ix10465 (.Y (nx10466), .A (gen_21_cmp_BSCmp_op2_16)) ;
    inv02 ix10467 (.Y (nx10468), .A (nx10466)) ;
    inv02 ix10469 (.Y (nx10470), .A (nx10466)) ;
    inv02 ix10471 (.Y (nx10472), .A (nx10466)) ;
    inv02 ix10473 (.Y (nx10474), .A (nx10466)) ;
    inv02 ix10475 (.Y (nx10476), .A (nx10466)) ;
    inv01 ix10477 (.Y (nx10478), .A (gen_20_cmp_BSCmp_op2_16)) ;
    inv02 ix10479 (.Y (nx10480), .A (nx10478)) ;
    inv02 ix10481 (.Y (nx10482), .A (nx10478)) ;
    inv02 ix10483 (.Y (nx10484), .A (nx10478)) ;
    inv02 ix10485 (.Y (nx10486), .A (nx10478)) ;
    inv02 ix10487 (.Y (nx10488), .A (nx10478)) ;
    inv01 ix10489 (.Y (nx10490), .A (gen_19_cmp_BSCmp_op2_16)) ;
    inv02 ix10491 (.Y (nx10492), .A (nx10490)) ;
    inv02 ix10493 (.Y (nx10494), .A (nx10490)) ;
    inv02 ix10495 (.Y (nx10496), .A (nx10490)) ;
    inv02 ix10497 (.Y (nx10498), .A (nx10490)) ;
    inv02 ix10499 (.Y (nx10500), .A (nx10490)) ;
    inv01 ix10501 (.Y (nx10502), .A (gen_18_cmp_BSCmp_op2_16)) ;
    inv02 ix10503 (.Y (nx10504), .A (nx10502)) ;
    inv02 ix10505 (.Y (nx10506), .A (nx10502)) ;
    inv02 ix10507 (.Y (nx10508), .A (nx10502)) ;
    inv02 ix10509 (.Y (nx10510), .A (nx10502)) ;
    inv02 ix10511 (.Y (nx10512), .A (nx10502)) ;
    inv01 ix10513 (.Y (nx10514), .A (gen_17_cmp_BSCmp_op2_16)) ;
    inv02 ix10515 (.Y (nx10516), .A (nx10514)) ;
    inv02 ix10517 (.Y (nx10518), .A (nx10514)) ;
    inv02 ix10519 (.Y (nx10520), .A (nx10514)) ;
    inv02 ix10521 (.Y (nx10522), .A (nx10514)) ;
    inv02 ix10523 (.Y (nx10524), .A (nx10514)) ;
    inv01 ix10525 (.Y (nx10526), .A (gen_16_cmp_BSCmp_op2_16)) ;
    inv02 ix10527 (.Y (nx10528), .A (nx10526)) ;
    inv02 ix10529 (.Y (nx10530), .A (nx10526)) ;
    inv02 ix10531 (.Y (nx10532), .A (nx10526)) ;
    inv02 ix10533 (.Y (nx10534), .A (nx10526)) ;
    inv02 ix10535 (.Y (nx10536), .A (nx10526)) ;
    inv01 ix10537 (.Y (nx10538), .A (gen_15_cmp_BSCmp_op2_16)) ;
    inv02 ix10539 (.Y (nx10540), .A (nx10538)) ;
    inv02 ix10541 (.Y (nx10542), .A (nx10538)) ;
    inv02 ix10543 (.Y (nx10544), .A (nx10538)) ;
    inv02 ix10545 (.Y (nx10546), .A (nx10538)) ;
    inv02 ix10547 (.Y (nx10548), .A (nx10538)) ;
    inv01 ix10549 (.Y (nx10550), .A (gen_14_cmp_BSCmp_op2_16)) ;
    inv02 ix10551 (.Y (nx10552), .A (nx10550)) ;
    inv02 ix10553 (.Y (nx10554), .A (nx10550)) ;
    inv02 ix10555 (.Y (nx10556), .A (nx10550)) ;
    inv02 ix10557 (.Y (nx10558), .A (nx10550)) ;
    inv02 ix10559 (.Y (nx10560), .A (nx10550)) ;
    inv01 ix10561 (.Y (nx10562), .A (gen_13_cmp_BSCmp_op2_16)) ;
    inv02 ix10563 (.Y (nx10564), .A (nx10562)) ;
    inv02 ix10565 (.Y (nx10566), .A (nx10562)) ;
    inv02 ix10567 (.Y (nx10568), .A (nx10562)) ;
    inv02 ix10569 (.Y (nx10570), .A (nx10562)) ;
    inv02 ix10571 (.Y (nx10572), .A (nx10562)) ;
    inv01 ix10573 (.Y (nx10574), .A (gen_12_cmp_BSCmp_op2_16)) ;
    inv02 ix10575 (.Y (nx10576), .A (nx10574)) ;
    inv02 ix10577 (.Y (nx10578), .A (nx10574)) ;
    inv02 ix10579 (.Y (nx10580), .A (nx10574)) ;
    inv02 ix10581 (.Y (nx10582), .A (nx10574)) ;
    inv02 ix10583 (.Y (nx10584), .A (nx10574)) ;
    inv01 ix10585 (.Y (nx10586), .A (gen_11_cmp_BSCmp_op2_16)) ;
    inv02 ix10587 (.Y (nx10588), .A (nx10586)) ;
    inv02 ix10589 (.Y (nx10590), .A (nx10586)) ;
    inv02 ix10591 (.Y (nx10592), .A (nx10586)) ;
    inv02 ix10593 (.Y (nx10594), .A (nx10586)) ;
    inv02 ix10595 (.Y (nx10596), .A (nx10586)) ;
    inv01 ix10597 (.Y (nx10598), .A (gen_10_cmp_BSCmp_op2_16)) ;
    inv02 ix10599 (.Y (nx10600), .A (nx10598)) ;
    inv02 ix10601 (.Y (nx10602), .A (nx10598)) ;
    inv02 ix10603 (.Y (nx10604), .A (nx10598)) ;
    inv02 ix10605 (.Y (nx10606), .A (nx10598)) ;
    inv02 ix10607 (.Y (nx10608), .A (nx10598)) ;
    inv01 ix10609 (.Y (nx10610), .A (gen_9_cmp_BSCmp_op2_16)) ;
    inv02 ix10611 (.Y (nx10612), .A (nx10610)) ;
    inv02 ix10613 (.Y (nx10614), .A (nx10610)) ;
    inv02 ix10615 (.Y (nx10616), .A (nx10610)) ;
    inv02 ix10617 (.Y (nx10618), .A (nx10610)) ;
    inv02 ix10619 (.Y (nx10620), .A (nx10610)) ;
    inv01 ix10621 (.Y (nx10622), .A (gen_8_cmp_BSCmp_op2_16)) ;
    inv02 ix10623 (.Y (nx10624), .A (nx10622)) ;
    inv02 ix10625 (.Y (nx10626), .A (nx10622)) ;
    inv02 ix10627 (.Y (nx10628), .A (nx10622)) ;
    inv02 ix10629 (.Y (nx10630), .A (nx10622)) ;
    inv02 ix10631 (.Y (nx10632), .A (nx10622)) ;
    inv01 ix10633 (.Y (nx10634), .A (gen_7_cmp_BSCmp_op2_16)) ;
    inv02 ix10635 (.Y (nx10636), .A (nx10634)) ;
    inv02 ix10637 (.Y (nx10638), .A (nx10634)) ;
    inv02 ix10639 (.Y (nx10640), .A (nx10634)) ;
    inv02 ix10641 (.Y (nx10642), .A (nx10634)) ;
    inv02 ix10643 (.Y (nx10644), .A (nx10634)) ;
    inv01 ix10645 (.Y (nx10646), .A (gen_6_cmp_BSCmp_op2_16)) ;
    inv02 ix10647 (.Y (nx10648), .A (nx10646)) ;
    inv02 ix10649 (.Y (nx10650), .A (nx10646)) ;
    inv02 ix10651 (.Y (nx10652), .A (nx10646)) ;
    inv02 ix10653 (.Y (nx10654), .A (nx10646)) ;
    inv02 ix10655 (.Y (nx10656), .A (nx10646)) ;
    inv01 ix10657 (.Y (nx10658), .A (gen_5_cmp_BSCmp_op2_16)) ;
    inv02 ix10659 (.Y (nx10660), .A (nx10658)) ;
    inv02 ix10661 (.Y (nx10662), .A (nx10658)) ;
    inv02 ix10663 (.Y (nx10664), .A (nx10658)) ;
    inv02 ix10665 (.Y (nx10666), .A (nx10658)) ;
    inv02 ix10667 (.Y (nx10668), .A (nx10658)) ;
    inv01 ix10669 (.Y (nx10670), .A (gen_4_cmp_BSCmp_op2_16)) ;
    inv02 ix10671 (.Y (nx10672), .A (nx10670)) ;
    inv02 ix10673 (.Y (nx10674), .A (nx10670)) ;
    inv02 ix10675 (.Y (nx10676), .A (nx10670)) ;
    inv02 ix10677 (.Y (nx10678), .A (nx10670)) ;
    inv02 ix10679 (.Y (nx10680), .A (nx10670)) ;
    inv01 ix10681 (.Y (nx10682), .A (gen_3_cmp_BSCmp_op2_16)) ;
    inv02 ix10683 (.Y (nx10684), .A (nx10682)) ;
    inv02 ix10685 (.Y (nx10686), .A (nx10682)) ;
    inv02 ix10687 (.Y (nx10688), .A (nx10682)) ;
    inv02 ix10689 (.Y (nx10690), .A (nx10682)) ;
    inv02 ix10691 (.Y (nx10692), .A (nx10682)) ;
    inv01 ix10693 (.Y (nx10694), .A (gen_2_cmp_BSCmp_op2_16)) ;
    inv02 ix10695 (.Y (nx10696), .A (nx10694)) ;
    inv02 ix10697 (.Y (nx10698), .A (nx10694)) ;
    inv02 ix10699 (.Y (nx10700), .A (nx10694)) ;
    inv02 ix10701 (.Y (nx10702), .A (nx10694)) ;
    inv02 ix10703 (.Y (nx10704), .A (nx10694)) ;
    inv01 ix10705 (.Y (nx10706), .A (gen_1_cmp_BSCmp_op2_16)) ;
    inv02 ix10707 (.Y (nx10708), .A (nx10706)) ;
    inv02 ix10709 (.Y (nx10710), .A (nx10706)) ;
    inv02 ix10711 (.Y (nx10712), .A (nx10706)) ;
    inv02 ix10713 (.Y (nx10714), .A (nx10706)) ;
    inv02 ix10715 (.Y (nx10716), .A (nx10706)) ;
    inv01 ix10717 (.Y (nx10718), .A (gen_0_cmp_BSCmp_op2_16)) ;
    inv02 ix10719 (.Y (nx10720), .A (nx10718)) ;
    inv02 ix10721 (.Y (nx10722), .A (nx10718)) ;
    inv02 ix10723 (.Y (nx10724), .A (nx10718)) ;
    inv02 ix10725 (.Y (nx10726), .A (nx10718)) ;
    inv02 ix10727 (.Y (nx10728), .A (nx10718)) ;
    buf02 ix10729 (.Y (nx10730), .A (nx6)) ;
    buf02 ix10731 (.Y (nx10732), .A (nx6)) ;
    buf02 ix10733 (.Y (nx10734), .A (nx6)) ;
    buf02 ix10735 (.Y (nx10736), .A (nx392)) ;
    buf02 ix10737 (.Y (nx10738), .A (nx392)) ;
    buf02 ix10739 (.Y (nx10740), .A (nx392)) ;
    buf02 ix10741 (.Y (nx10742), .A (nx778)) ;
    buf02 ix10743 (.Y (nx10744), .A (nx778)) ;
    buf02 ix10745 (.Y (nx10746), .A (nx778)) ;
    buf02 ix10747 (.Y (nx10748), .A (nx1164)) ;
    buf02 ix10749 (.Y (nx10750), .A (nx1164)) ;
    buf02 ix10751 (.Y (nx10752), .A (nx1164)) ;
    buf02 ix10753 (.Y (nx10754), .A (nx1550)) ;
    buf02 ix10755 (.Y (nx10756), .A (nx1550)) ;
    buf02 ix10757 (.Y (nx10758), .A (nx1550)) ;
    buf02 ix10759 (.Y (nx10760), .A (nx1936)) ;
    buf02 ix10761 (.Y (nx10762), .A (nx1936)) ;
    buf02 ix10763 (.Y (nx10764), .A (nx1936)) ;
    buf02 ix10765 (.Y (nx10766), .A (nx2322)) ;
    buf02 ix10767 (.Y (nx10768), .A (nx2322)) ;
    buf02 ix10769 (.Y (nx10770), .A (nx2322)) ;
    buf02 ix10771 (.Y (nx10772), .A (nx2708)) ;
    buf02 ix10773 (.Y (nx10774), .A (nx2708)) ;
    buf02 ix10775 (.Y (nx10776), .A (nx2708)) ;
    buf02 ix10777 (.Y (nx10778), .A (nx3094)) ;
    buf02 ix10779 (.Y (nx10780), .A (nx3094)) ;
    buf02 ix10781 (.Y (nx10782), .A (nx3094)) ;
    buf02 ix10783 (.Y (nx10784), .A (nx3480)) ;
    buf02 ix10785 (.Y (nx10786), .A (nx3480)) ;
    buf02 ix10787 (.Y (nx10788), .A (nx3480)) ;
    buf02 ix10789 (.Y (nx10790), .A (nx3866)) ;
    buf02 ix10791 (.Y (nx10792), .A (nx3866)) ;
    buf02 ix10793 (.Y (nx10794), .A (nx3866)) ;
    buf02 ix10795 (.Y (nx10796), .A (nx4252)) ;
    buf02 ix10797 (.Y (nx10798), .A (nx4252)) ;
    buf02 ix10799 (.Y (nx10800), .A (nx4252)) ;
    buf02 ix10801 (.Y (nx10802), .A (nx4638)) ;
    buf02 ix10803 (.Y (nx10804), .A (nx4638)) ;
    buf02 ix10805 (.Y (nx10806), .A (nx4638)) ;
    buf02 ix10807 (.Y (nx10808), .A (nx5024)) ;
    buf02 ix10809 (.Y (nx10810), .A (nx5024)) ;
    buf02 ix10811 (.Y (nx10812), .A (nx5024)) ;
    buf02 ix10813 (.Y (nx10814), .A (nx5410)) ;
    buf02 ix10815 (.Y (nx10816), .A (nx5410)) ;
    buf02 ix10817 (.Y (nx10818), .A (nx5410)) ;
    buf02 ix10819 (.Y (nx10820), .A (nx5796)) ;
    buf02 ix10821 (.Y (nx10822), .A (nx5796)) ;
    buf02 ix10823 (.Y (nx10824), .A (nx5796)) ;
    buf02 ix10825 (.Y (nx10826), .A (nx6182)) ;
    buf02 ix10827 (.Y (nx10828), .A (nx6182)) ;
    buf02 ix10829 (.Y (nx10830), .A (nx6182)) ;
    buf02 ix10831 (.Y (nx10832), .A (nx6568)) ;
    buf02 ix10833 (.Y (nx10834), .A (nx6568)) ;
    buf02 ix10835 (.Y (nx10836), .A (nx6568)) ;
    buf02 ix10837 (.Y (nx10838), .A (nx6954)) ;
    buf02 ix10839 (.Y (nx10840), .A (nx6954)) ;
    buf02 ix10841 (.Y (nx10842), .A (nx6954)) ;
    buf02 ix10843 (.Y (nx10844), .A (nx7340)) ;
    buf02 ix10845 (.Y (nx10846), .A (nx7340)) ;
    buf02 ix10847 (.Y (nx10848), .A (nx7340)) ;
    buf02 ix10849 (.Y (nx10850), .A (nx7726)) ;
    buf02 ix10851 (.Y (nx10852), .A (nx7726)) ;
    buf02 ix10853 (.Y (nx10854), .A (nx7726)) ;
    buf02 ix10855 (.Y (nx10856), .A (nx8112)) ;
    buf02 ix10857 (.Y (nx10858), .A (nx8112)) ;
    buf02 ix10859 (.Y (nx10860), .A (nx8112)) ;
    buf02 ix10861 (.Y (nx10862), .A (nx8498)) ;
    buf02 ix10863 (.Y (nx10864), .A (nx8498)) ;
    buf02 ix10865 (.Y (nx10866), .A (nx8498)) ;
    buf02 ix10867 (.Y (nx10868), .A (nx8884)) ;
    buf02 ix10869 (.Y (nx10870), .A (nx8884)) ;
    buf02 ix10871 (.Y (nx10872), .A (nx8884)) ;
    buf02 ix10873 (.Y (nx10874), .A (nx9270)) ;
    buf02 ix10875 (.Y (nx10876), .A (nx9270)) ;
    buf02 ix10877 (.Y (nx10878), .A (nx9270)) ;
    inv02 ix10879 (.Y (nx10880), .A (done)) ;
    inv02 ix10881 (.Y (nx10882), .A (nx11934)) ;
    inv02 ix10883 (.Y (nx10884), .A (nx11934)) ;
    inv02 ix10885 (.Y (nx10886), .A (nx11934)) ;
    inv02 ix10889 (.Y (nx10890), .A (nx10888)) ;
    inv02 ix10891 (.Y (nx10892), .A (nx10888)) ;
    inv02 ix10893 (.Y (nx10894), .A (nx10888)) ;
    inv04 ix10895 (.Y (nx10896), .A (gen_0_cmp_pMux_1)) ;
    inv04 ix10897 (.Y (nx10898), .A (gen_0_cmp_pMux_1)) ;
    inv04 ix10899 (.Y (nx10900), .A (gen_0_cmp_pMux_1)) ;
    inv04 ix10901 (.Y (nx10902), .A (gen_0_cmp_pMux_1)) ;
    inv02 ix10905 (.Y (nx10906), .A (nx10904)) ;
    inv02 ix10907 (.Y (nx10908), .A (nx10904)) ;
    inv02 ix10909 (.Y (nx10910), .A (nx10904)) ;
    inv02 ix10913 (.Y (nx10914), .A (nx10912)) ;
    inv02 ix10915 (.Y (nx10916), .A (nx10912)) ;
    inv02 ix10917 (.Y (nx10918), .A (nx10912)) ;
    inv02 ix10921 (.Y (nx10922), .A (nx10920)) ;
    inv02 ix10923 (.Y (nx10924), .A (nx10920)) ;
    inv02 ix10925 (.Y (nx10926), .A (nx10920)) ;
    inv02 ix10929 (.Y (nx10930), .A (nx10928)) ;
    inv02 ix10931 (.Y (nx10932), .A (nx10928)) ;
    inv02 ix10933 (.Y (nx10934), .A (nx10928)) ;
    inv04 ix10935 (.Y (nx10936), .A (gen_1_cmp_pMux_1)) ;
    inv04 ix10937 (.Y (nx10938), .A (gen_1_cmp_pMux_1)) ;
    inv04 ix10939 (.Y (nx10940), .A (gen_1_cmp_pMux_1)) ;
    inv04 ix10941 (.Y (nx10942), .A (gen_1_cmp_pMux_1)) ;
    inv02 ix10945 (.Y (nx10946), .A (nx10944)) ;
    inv02 ix10947 (.Y (nx10948), .A (nx10944)) ;
    inv02 ix10949 (.Y (nx10950), .A (nx10944)) ;
    inv02 ix10953 (.Y (nx10954), .A (nx10952)) ;
    inv02 ix10955 (.Y (nx10956), .A (nx10952)) ;
    inv02 ix10957 (.Y (nx10958), .A (nx10952)) ;
    inv02 ix10961 (.Y (nx10962), .A (nx10960)) ;
    inv02 ix10963 (.Y (nx10964), .A (nx10960)) ;
    inv02 ix10965 (.Y (nx10966), .A (nx10960)) ;
    inv02 ix10969 (.Y (nx10970), .A (nx10968)) ;
    inv02 ix10971 (.Y (nx10972), .A (nx10968)) ;
    inv02 ix10973 (.Y (nx10974), .A (nx10968)) ;
    inv04 ix10975 (.Y (nx10976), .A (gen_2_cmp_pMux_1)) ;
    inv04 ix10977 (.Y (nx10978), .A (gen_2_cmp_pMux_1)) ;
    inv04 ix10979 (.Y (nx10980), .A (gen_2_cmp_pMux_1)) ;
    inv04 ix10981 (.Y (nx10982), .A (gen_2_cmp_pMux_1)) ;
    inv02 ix10985 (.Y (nx10986), .A (nx10984)) ;
    inv02 ix10987 (.Y (nx10988), .A (nx10984)) ;
    inv02 ix10989 (.Y (nx10990), .A (nx10984)) ;
    inv02 ix10993 (.Y (nx10994), .A (nx10992)) ;
    inv02 ix10995 (.Y (nx10996), .A (nx10992)) ;
    inv02 ix10997 (.Y (nx10998), .A (nx10992)) ;
    inv02 ix11001 (.Y (nx11002), .A (nx11000)) ;
    inv02 ix11003 (.Y (nx11004), .A (nx11000)) ;
    inv02 ix11005 (.Y (nx11006), .A (nx11000)) ;
    inv02 ix11009 (.Y (nx11010), .A (nx11008)) ;
    inv02 ix11011 (.Y (nx11012), .A (nx11008)) ;
    inv02 ix11013 (.Y (nx11014), .A (nx11008)) ;
    inv04 ix11015 (.Y (nx11016), .A (gen_3_cmp_pMux_1)) ;
    inv04 ix11017 (.Y (nx11018), .A (gen_3_cmp_pMux_1)) ;
    inv04 ix11019 (.Y (nx11020), .A (gen_3_cmp_pMux_1)) ;
    inv04 ix11021 (.Y (nx11022), .A (gen_3_cmp_pMux_1)) ;
    inv02 ix11025 (.Y (nx11026), .A (nx11024)) ;
    inv02 ix11027 (.Y (nx11028), .A (nx11024)) ;
    inv02 ix11029 (.Y (nx11030), .A (nx11024)) ;
    inv02 ix11033 (.Y (nx11034), .A (nx11032)) ;
    inv02 ix11035 (.Y (nx11036), .A (nx11032)) ;
    inv02 ix11037 (.Y (nx11038), .A (nx11032)) ;
    inv02 ix11041 (.Y (nx11042), .A (nx11040)) ;
    inv02 ix11043 (.Y (nx11044), .A (nx11040)) ;
    inv02 ix11045 (.Y (nx11046), .A (nx11040)) ;
    inv02 ix11049 (.Y (nx11050), .A (nx11048)) ;
    inv02 ix11051 (.Y (nx11052), .A (nx11048)) ;
    inv02 ix11053 (.Y (nx11054), .A (nx11048)) ;
    inv04 ix11055 (.Y (nx11056), .A (gen_4_cmp_pMux_1)) ;
    inv04 ix11057 (.Y (nx11058), .A (gen_4_cmp_pMux_1)) ;
    inv04 ix11059 (.Y (nx11060), .A (gen_4_cmp_pMux_1)) ;
    inv04 ix11061 (.Y (nx11062), .A (gen_4_cmp_pMux_1)) ;
    inv02 ix11065 (.Y (nx11066), .A (nx11064)) ;
    inv02 ix11067 (.Y (nx11068), .A (nx11064)) ;
    inv02 ix11069 (.Y (nx11070), .A (nx11064)) ;
    inv02 ix11073 (.Y (nx11074), .A (nx11072)) ;
    inv02 ix11075 (.Y (nx11076), .A (nx11072)) ;
    inv02 ix11077 (.Y (nx11078), .A (nx11072)) ;
    inv02 ix11081 (.Y (nx11082), .A (nx11080)) ;
    inv02 ix11083 (.Y (nx11084), .A (nx11080)) ;
    inv02 ix11085 (.Y (nx11086), .A (nx11080)) ;
    inv02 ix11089 (.Y (nx11090), .A (nx11088)) ;
    inv02 ix11091 (.Y (nx11092), .A (nx11088)) ;
    inv02 ix11093 (.Y (nx11094), .A (nx11088)) ;
    inv04 ix11095 (.Y (nx11096), .A (gen_5_cmp_pMux_1)) ;
    inv04 ix11097 (.Y (nx11098), .A (gen_5_cmp_pMux_1)) ;
    inv04 ix11099 (.Y (nx11100), .A (gen_5_cmp_pMux_1)) ;
    inv04 ix11101 (.Y (nx11102), .A (gen_5_cmp_pMux_1)) ;
    inv02 ix11105 (.Y (nx11106), .A (nx11104)) ;
    inv02 ix11107 (.Y (nx11108), .A (nx11104)) ;
    inv02 ix11109 (.Y (nx11110), .A (nx11104)) ;
    inv02 ix11113 (.Y (nx11114), .A (nx11112)) ;
    inv02 ix11115 (.Y (nx11116), .A (nx11112)) ;
    inv02 ix11117 (.Y (nx11118), .A (nx11112)) ;
    inv02 ix11121 (.Y (nx11122), .A (nx11120)) ;
    inv02 ix11123 (.Y (nx11124), .A (nx11120)) ;
    inv02 ix11125 (.Y (nx11126), .A (nx11120)) ;
    inv02 ix11129 (.Y (nx11130), .A (nx11128)) ;
    inv02 ix11131 (.Y (nx11132), .A (nx11128)) ;
    inv02 ix11133 (.Y (nx11134), .A (nx11128)) ;
    inv04 ix11135 (.Y (nx11136), .A (gen_6_cmp_pMux_1)) ;
    inv04 ix11137 (.Y (nx11138), .A (gen_6_cmp_pMux_1)) ;
    inv04 ix11139 (.Y (nx11140), .A (gen_6_cmp_pMux_1)) ;
    inv04 ix11141 (.Y (nx11142), .A (gen_6_cmp_pMux_1)) ;
    inv02 ix11145 (.Y (nx11146), .A (nx11144)) ;
    inv02 ix11147 (.Y (nx11148), .A (nx11144)) ;
    inv02 ix11149 (.Y (nx11150), .A (nx11144)) ;
    inv02 ix11153 (.Y (nx11154), .A (nx11152)) ;
    inv02 ix11155 (.Y (nx11156), .A (nx11152)) ;
    inv02 ix11157 (.Y (nx11158), .A (nx11152)) ;
    inv02 ix11161 (.Y (nx11162), .A (nx11160)) ;
    inv02 ix11163 (.Y (nx11164), .A (nx11160)) ;
    inv02 ix11165 (.Y (nx11166), .A (nx11160)) ;
    inv02 ix11169 (.Y (nx11170), .A (nx11168)) ;
    inv02 ix11171 (.Y (nx11172), .A (nx11168)) ;
    inv02 ix11173 (.Y (nx11174), .A (nx11168)) ;
    inv04 ix11175 (.Y (nx11176), .A (gen_7_cmp_pMux_1)) ;
    inv04 ix11177 (.Y (nx11178), .A (gen_7_cmp_pMux_1)) ;
    inv04 ix11179 (.Y (nx11180), .A (gen_7_cmp_pMux_1)) ;
    inv04 ix11181 (.Y (nx11182), .A (gen_7_cmp_pMux_1)) ;
    inv02 ix11185 (.Y (nx11186), .A (nx11184)) ;
    inv02 ix11187 (.Y (nx11188), .A (nx11184)) ;
    inv02 ix11189 (.Y (nx11190), .A (nx11184)) ;
    inv02 ix11193 (.Y (nx11194), .A (nx11192)) ;
    inv02 ix11195 (.Y (nx11196), .A (nx11192)) ;
    inv02 ix11197 (.Y (nx11198), .A (nx11192)) ;
    inv02 ix11201 (.Y (nx11202), .A (nx11200)) ;
    inv02 ix11203 (.Y (nx11204), .A (nx11200)) ;
    inv02 ix11205 (.Y (nx11206), .A (nx11200)) ;
    inv02 ix11209 (.Y (nx11210), .A (nx11208)) ;
    inv02 ix11211 (.Y (nx11212), .A (nx11208)) ;
    inv02 ix11213 (.Y (nx11214), .A (nx11208)) ;
    inv04 ix11215 (.Y (nx11216), .A (gen_8_cmp_pMux_1)) ;
    inv04 ix11217 (.Y (nx11218), .A (gen_8_cmp_pMux_1)) ;
    inv04 ix11219 (.Y (nx11220), .A (gen_8_cmp_pMux_1)) ;
    inv04 ix11221 (.Y (nx11222), .A (gen_8_cmp_pMux_1)) ;
    inv02 ix11225 (.Y (nx11226), .A (nx11224)) ;
    inv02 ix11227 (.Y (nx11228), .A (nx11224)) ;
    inv02 ix11229 (.Y (nx11230), .A (nx11224)) ;
    inv02 ix11233 (.Y (nx11234), .A (nx11232)) ;
    inv02 ix11235 (.Y (nx11236), .A (nx11232)) ;
    inv02 ix11237 (.Y (nx11238), .A (nx11232)) ;
    inv02 ix11241 (.Y (nx11242), .A (nx11240)) ;
    inv02 ix11243 (.Y (nx11244), .A (nx11240)) ;
    inv02 ix11245 (.Y (nx11246), .A (nx11240)) ;
    inv02 ix11249 (.Y (nx11250), .A (nx11248)) ;
    inv02 ix11251 (.Y (nx11252), .A (nx11248)) ;
    inv02 ix11253 (.Y (nx11254), .A (nx11248)) ;
    inv04 ix11255 (.Y (nx11256), .A (gen_9_cmp_pMux_1)) ;
    inv04 ix11257 (.Y (nx11258), .A (gen_9_cmp_pMux_1)) ;
    inv04 ix11259 (.Y (nx11260), .A (gen_9_cmp_pMux_1)) ;
    inv04 ix11261 (.Y (nx11262), .A (gen_9_cmp_pMux_1)) ;
    inv02 ix11265 (.Y (nx11266), .A (nx11264)) ;
    inv02 ix11267 (.Y (nx11268), .A (nx11264)) ;
    inv02 ix11269 (.Y (nx11270), .A (nx11264)) ;
    inv02 ix11273 (.Y (nx11274), .A (nx11272)) ;
    inv02 ix11275 (.Y (nx11276), .A (nx11272)) ;
    inv02 ix11277 (.Y (nx11278), .A (nx11272)) ;
    inv02 ix11281 (.Y (nx11282), .A (nx11280)) ;
    inv02 ix11283 (.Y (nx11284), .A (nx11280)) ;
    inv02 ix11285 (.Y (nx11286), .A (nx11280)) ;
    inv02 ix11289 (.Y (nx11290), .A (nx11288)) ;
    inv02 ix11291 (.Y (nx11292), .A (nx11288)) ;
    inv02 ix11293 (.Y (nx11294), .A (nx11288)) ;
    inv04 ix11295 (.Y (nx11296), .A (gen_10_cmp_pMux_1)) ;
    inv04 ix11297 (.Y (nx11298), .A (gen_10_cmp_pMux_1)) ;
    inv04 ix11299 (.Y (nx11300), .A (gen_10_cmp_pMux_1)) ;
    inv04 ix11301 (.Y (nx11302), .A (gen_10_cmp_pMux_1)) ;
    inv02 ix11305 (.Y (nx11306), .A (nx11304)) ;
    inv02 ix11307 (.Y (nx11308), .A (nx11304)) ;
    inv02 ix11309 (.Y (nx11310), .A (nx11304)) ;
    inv02 ix11313 (.Y (nx11314), .A (nx11312)) ;
    inv02 ix11315 (.Y (nx11316), .A (nx11312)) ;
    inv02 ix11317 (.Y (nx11318), .A (nx11312)) ;
    inv02 ix11321 (.Y (nx11322), .A (nx11320)) ;
    inv02 ix11323 (.Y (nx11324), .A (nx11320)) ;
    inv02 ix11325 (.Y (nx11326), .A (nx11320)) ;
    inv02 ix11329 (.Y (nx11330), .A (nx11328)) ;
    inv02 ix11331 (.Y (nx11332), .A (nx11328)) ;
    inv02 ix11333 (.Y (nx11334), .A (nx11328)) ;
    inv04 ix11335 (.Y (nx11336), .A (gen_11_cmp_pMux_1)) ;
    inv04 ix11337 (.Y (nx11338), .A (gen_11_cmp_pMux_1)) ;
    inv04 ix11339 (.Y (nx11340), .A (gen_11_cmp_pMux_1)) ;
    inv04 ix11341 (.Y (nx11342), .A (gen_11_cmp_pMux_1)) ;
    inv02 ix11345 (.Y (nx11346), .A (nx11344)) ;
    inv02 ix11347 (.Y (nx11348), .A (nx11344)) ;
    inv02 ix11349 (.Y (nx11350), .A (nx11344)) ;
    inv02 ix11353 (.Y (nx11354), .A (nx11352)) ;
    inv02 ix11355 (.Y (nx11356), .A (nx11352)) ;
    inv02 ix11357 (.Y (nx11358), .A (nx11352)) ;
    inv02 ix11361 (.Y (nx11362), .A (nx11360)) ;
    inv02 ix11363 (.Y (nx11364), .A (nx11360)) ;
    inv02 ix11365 (.Y (nx11366), .A (nx11360)) ;
    inv02 ix11369 (.Y (nx11370), .A (nx11368)) ;
    inv02 ix11371 (.Y (nx11372), .A (nx11368)) ;
    inv02 ix11373 (.Y (nx11374), .A (nx11368)) ;
    inv04 ix11375 (.Y (nx11376), .A (gen_12_cmp_pMux_1)) ;
    inv04 ix11377 (.Y (nx11378), .A (gen_12_cmp_pMux_1)) ;
    inv04 ix11379 (.Y (nx11380), .A (gen_12_cmp_pMux_1)) ;
    inv04 ix11381 (.Y (nx11382), .A (gen_12_cmp_pMux_1)) ;
    inv02 ix11385 (.Y (nx11386), .A (nx11384)) ;
    inv02 ix11387 (.Y (nx11388), .A (nx11384)) ;
    inv02 ix11389 (.Y (nx11390), .A (nx11384)) ;
    inv02 ix11393 (.Y (nx11394), .A (nx11392)) ;
    inv02 ix11395 (.Y (nx11396), .A (nx11392)) ;
    inv02 ix11397 (.Y (nx11398), .A (nx11392)) ;
    inv02 ix11401 (.Y (nx11402), .A (nx11400)) ;
    inv02 ix11403 (.Y (nx11404), .A (nx11400)) ;
    inv02 ix11405 (.Y (nx11406), .A (nx11400)) ;
    inv02 ix11409 (.Y (nx11410), .A (nx11408)) ;
    inv02 ix11411 (.Y (nx11412), .A (nx11408)) ;
    inv02 ix11413 (.Y (nx11414), .A (nx11408)) ;
    inv04 ix11415 (.Y (nx11416), .A (gen_13_cmp_pMux_1)) ;
    inv04 ix11417 (.Y (nx11418), .A (gen_13_cmp_pMux_1)) ;
    inv04 ix11419 (.Y (nx11420), .A (gen_13_cmp_pMux_1)) ;
    inv04 ix11421 (.Y (nx11422), .A (gen_13_cmp_pMux_1)) ;
    inv02 ix11425 (.Y (nx11426), .A (nx11424)) ;
    inv02 ix11427 (.Y (nx11428), .A (nx11424)) ;
    inv02 ix11429 (.Y (nx11430), .A (nx11424)) ;
    inv02 ix11433 (.Y (nx11434), .A (nx11432)) ;
    inv02 ix11435 (.Y (nx11436), .A (nx11432)) ;
    inv02 ix11437 (.Y (nx11438), .A (nx11432)) ;
    inv02 ix11441 (.Y (nx11442), .A (nx11440)) ;
    inv02 ix11443 (.Y (nx11444), .A (nx11440)) ;
    inv02 ix11445 (.Y (nx11446), .A (nx11440)) ;
    inv02 ix11449 (.Y (nx11450), .A (nx11448)) ;
    inv02 ix11451 (.Y (nx11452), .A (nx11448)) ;
    inv02 ix11453 (.Y (nx11454), .A (nx11448)) ;
    inv04 ix11455 (.Y (nx11456), .A (gen_14_cmp_pMux_1)) ;
    inv04 ix11457 (.Y (nx11458), .A (gen_14_cmp_pMux_1)) ;
    inv04 ix11459 (.Y (nx11460), .A (gen_14_cmp_pMux_1)) ;
    inv04 ix11461 (.Y (nx11462), .A (gen_14_cmp_pMux_1)) ;
    inv02 ix11465 (.Y (nx11466), .A (nx11464)) ;
    inv02 ix11467 (.Y (nx11468), .A (nx11464)) ;
    inv02 ix11469 (.Y (nx11470), .A (nx11464)) ;
    inv02 ix11473 (.Y (nx11474), .A (nx11472)) ;
    inv02 ix11475 (.Y (nx11476), .A (nx11472)) ;
    inv02 ix11477 (.Y (nx11478), .A (nx11472)) ;
    inv02 ix11481 (.Y (nx11482), .A (nx11480)) ;
    inv02 ix11483 (.Y (nx11484), .A (nx11480)) ;
    inv02 ix11485 (.Y (nx11486), .A (nx11480)) ;
    inv02 ix11489 (.Y (nx11490), .A (nx11488)) ;
    inv02 ix11491 (.Y (nx11492), .A (nx11488)) ;
    inv02 ix11493 (.Y (nx11494), .A (nx11488)) ;
    inv04 ix11495 (.Y (nx11496), .A (gen_15_cmp_pMux_1)) ;
    inv04 ix11497 (.Y (nx11498), .A (gen_15_cmp_pMux_1)) ;
    inv04 ix11499 (.Y (nx11500), .A (gen_15_cmp_pMux_1)) ;
    inv04 ix11501 (.Y (nx11502), .A (gen_15_cmp_pMux_1)) ;
    inv02 ix11505 (.Y (nx11506), .A (nx11504)) ;
    inv02 ix11507 (.Y (nx11508), .A (nx11504)) ;
    inv02 ix11509 (.Y (nx11510), .A (nx11504)) ;
    inv02 ix11513 (.Y (nx11514), .A (nx11512)) ;
    inv02 ix11515 (.Y (nx11516), .A (nx11512)) ;
    inv02 ix11517 (.Y (nx11518), .A (nx11512)) ;
    inv02 ix11521 (.Y (nx11522), .A (nx11520)) ;
    inv02 ix11523 (.Y (nx11524), .A (nx11520)) ;
    inv02 ix11525 (.Y (nx11526), .A (nx11520)) ;
    inv02 ix11529 (.Y (nx11530), .A (nx11528)) ;
    inv02 ix11531 (.Y (nx11532), .A (nx11528)) ;
    inv02 ix11533 (.Y (nx11534), .A (nx11528)) ;
    inv04 ix11535 (.Y (nx11536), .A (gen_16_cmp_pMux_1)) ;
    inv04 ix11537 (.Y (nx11538), .A (gen_16_cmp_pMux_1)) ;
    inv04 ix11539 (.Y (nx11540), .A (gen_16_cmp_pMux_1)) ;
    inv04 ix11541 (.Y (nx11542), .A (gen_16_cmp_pMux_1)) ;
    inv02 ix11545 (.Y (nx11546), .A (nx11544)) ;
    inv02 ix11547 (.Y (nx11548), .A (nx11544)) ;
    inv02 ix11549 (.Y (nx11550), .A (nx11544)) ;
    inv02 ix11553 (.Y (nx11554), .A (nx11552)) ;
    inv02 ix11555 (.Y (nx11556), .A (nx11552)) ;
    inv02 ix11557 (.Y (nx11558), .A (nx11552)) ;
    inv02 ix11561 (.Y (nx11562), .A (nx11560)) ;
    inv02 ix11563 (.Y (nx11564), .A (nx11560)) ;
    inv02 ix11565 (.Y (nx11566), .A (nx11560)) ;
    inv02 ix11569 (.Y (nx11570), .A (nx11568)) ;
    inv02 ix11571 (.Y (nx11572), .A (nx11568)) ;
    inv02 ix11573 (.Y (nx11574), .A (nx11568)) ;
    inv04 ix11575 (.Y (nx11576), .A (gen_17_cmp_pMux_1)) ;
    inv04 ix11577 (.Y (nx11578), .A (gen_17_cmp_pMux_1)) ;
    inv04 ix11579 (.Y (nx11580), .A (gen_17_cmp_pMux_1)) ;
    inv04 ix11581 (.Y (nx11582), .A (gen_17_cmp_pMux_1)) ;
    inv02 ix11585 (.Y (nx11586), .A (nx11584)) ;
    inv02 ix11587 (.Y (nx11588), .A (nx11584)) ;
    inv02 ix11589 (.Y (nx11590), .A (nx11584)) ;
    inv02 ix11593 (.Y (nx11594), .A (nx11592)) ;
    inv02 ix11595 (.Y (nx11596), .A (nx11592)) ;
    inv02 ix11597 (.Y (nx11598), .A (nx11592)) ;
    inv02 ix11601 (.Y (nx11602), .A (nx11600)) ;
    inv02 ix11603 (.Y (nx11604), .A (nx11600)) ;
    inv02 ix11605 (.Y (nx11606), .A (nx11600)) ;
    inv02 ix11609 (.Y (nx11610), .A (nx11608)) ;
    inv02 ix11611 (.Y (nx11612), .A (nx11608)) ;
    inv02 ix11613 (.Y (nx11614), .A (nx11608)) ;
    inv04 ix11615 (.Y (nx11616), .A (gen_18_cmp_pMux_1)) ;
    inv04 ix11617 (.Y (nx11618), .A (gen_18_cmp_pMux_1)) ;
    inv04 ix11619 (.Y (nx11620), .A (gen_18_cmp_pMux_1)) ;
    inv04 ix11621 (.Y (nx11622), .A (gen_18_cmp_pMux_1)) ;
    inv02 ix11625 (.Y (nx11626), .A (nx11624)) ;
    inv02 ix11627 (.Y (nx11628), .A (nx11624)) ;
    inv02 ix11629 (.Y (nx11630), .A (nx11624)) ;
    inv02 ix11633 (.Y (nx11634), .A (nx11632)) ;
    inv02 ix11635 (.Y (nx11636), .A (nx11632)) ;
    inv02 ix11637 (.Y (nx11638), .A (nx11632)) ;
    inv02 ix11641 (.Y (nx11642), .A (nx11640)) ;
    inv02 ix11643 (.Y (nx11644), .A (nx11640)) ;
    inv02 ix11645 (.Y (nx11646), .A (nx11640)) ;
    inv02 ix11649 (.Y (nx11650), .A (nx11648)) ;
    inv02 ix11651 (.Y (nx11652), .A (nx11648)) ;
    inv02 ix11653 (.Y (nx11654), .A (nx11648)) ;
    inv04 ix11655 (.Y (nx11656), .A (gen_19_cmp_pMux_1)) ;
    inv04 ix11657 (.Y (nx11658), .A (gen_19_cmp_pMux_1)) ;
    inv04 ix11659 (.Y (nx11660), .A (gen_19_cmp_pMux_1)) ;
    inv04 ix11661 (.Y (nx11662), .A (gen_19_cmp_pMux_1)) ;
    inv02 ix11665 (.Y (nx11666), .A (nx11664)) ;
    inv02 ix11667 (.Y (nx11668), .A (nx11664)) ;
    inv02 ix11669 (.Y (nx11670), .A (nx11664)) ;
    inv02 ix11673 (.Y (nx11674), .A (nx11672)) ;
    inv02 ix11675 (.Y (nx11676), .A (nx11672)) ;
    inv02 ix11677 (.Y (nx11678), .A (nx11672)) ;
    inv02 ix11681 (.Y (nx11682), .A (nx11680)) ;
    inv02 ix11683 (.Y (nx11684), .A (nx11680)) ;
    inv02 ix11685 (.Y (nx11686), .A (nx11680)) ;
    inv02 ix11689 (.Y (nx11690), .A (nx11688)) ;
    inv02 ix11691 (.Y (nx11692), .A (nx11688)) ;
    inv02 ix11693 (.Y (nx11694), .A (nx11688)) ;
    inv04 ix11695 (.Y (nx11696), .A (gen_20_cmp_pMux_1)) ;
    inv04 ix11697 (.Y (nx11698), .A (gen_20_cmp_pMux_1)) ;
    inv04 ix11699 (.Y (nx11700), .A (gen_20_cmp_pMux_1)) ;
    inv04 ix11701 (.Y (nx11702), .A (gen_20_cmp_pMux_1)) ;
    inv02 ix11705 (.Y (nx11706), .A (nx11704)) ;
    inv02 ix11707 (.Y (nx11708), .A (nx11704)) ;
    inv02 ix11709 (.Y (nx11710), .A (nx11704)) ;
    inv02 ix11713 (.Y (nx11714), .A (nx11712)) ;
    inv02 ix11715 (.Y (nx11716), .A (nx11712)) ;
    inv02 ix11717 (.Y (nx11718), .A (nx11712)) ;
    inv02 ix11721 (.Y (nx11722), .A (nx11720)) ;
    inv02 ix11723 (.Y (nx11724), .A (nx11720)) ;
    inv02 ix11725 (.Y (nx11726), .A (nx11720)) ;
    inv02 ix11729 (.Y (nx11730), .A (nx11728)) ;
    inv02 ix11731 (.Y (nx11732), .A (nx11728)) ;
    inv02 ix11733 (.Y (nx11734), .A (nx11728)) ;
    inv04 ix11735 (.Y (nx11736), .A (gen_21_cmp_pMux_1)) ;
    inv04 ix11737 (.Y (nx11738), .A (gen_21_cmp_pMux_1)) ;
    inv04 ix11739 (.Y (nx11740), .A (gen_21_cmp_pMux_1)) ;
    inv04 ix11741 (.Y (nx11742), .A (gen_21_cmp_pMux_1)) ;
    inv02 ix11745 (.Y (nx11746), .A (nx11744)) ;
    inv02 ix11747 (.Y (nx11748), .A (nx11744)) ;
    inv02 ix11749 (.Y (nx11750), .A (nx11744)) ;
    inv02 ix11753 (.Y (nx11754), .A (nx11752)) ;
    inv02 ix11755 (.Y (nx11756), .A (nx11752)) ;
    inv02 ix11757 (.Y (nx11758), .A (nx11752)) ;
    inv02 ix11761 (.Y (nx11762), .A (nx11760)) ;
    inv02 ix11763 (.Y (nx11764), .A (nx11760)) ;
    inv02 ix11765 (.Y (nx11766), .A (nx11760)) ;
    inv02 ix11769 (.Y (nx11770), .A (nx11768)) ;
    inv02 ix11771 (.Y (nx11772), .A (nx11768)) ;
    inv02 ix11773 (.Y (nx11774), .A (nx11768)) ;
    inv04 ix11775 (.Y (nx11776), .A (gen_22_cmp_pMux_1)) ;
    inv04 ix11777 (.Y (nx11778), .A (gen_22_cmp_pMux_1)) ;
    inv04 ix11779 (.Y (nx11780), .A (gen_22_cmp_pMux_1)) ;
    inv04 ix11781 (.Y (nx11782), .A (gen_22_cmp_pMux_1)) ;
    inv02 ix11785 (.Y (nx11786), .A (nx11784)) ;
    inv02 ix11787 (.Y (nx11788), .A (nx11784)) ;
    inv02 ix11789 (.Y (nx11790), .A (nx11784)) ;
    inv02 ix11793 (.Y (nx11794), .A (nx11792)) ;
    inv02 ix11795 (.Y (nx11796), .A (nx11792)) ;
    inv02 ix11797 (.Y (nx11798), .A (nx11792)) ;
    inv02 ix11801 (.Y (nx11802), .A (nx11800)) ;
    inv02 ix11803 (.Y (nx11804), .A (nx11800)) ;
    inv02 ix11805 (.Y (nx11806), .A (nx11800)) ;
    inv02 ix11809 (.Y (nx11810), .A (nx11808)) ;
    inv02 ix11811 (.Y (nx11812), .A (nx11808)) ;
    inv02 ix11813 (.Y (nx11814), .A (nx11808)) ;
    inv04 ix11815 (.Y (nx11816), .A (gen_23_cmp_pMux_1)) ;
    inv04 ix11817 (.Y (nx11818), .A (gen_23_cmp_pMux_1)) ;
    inv04 ix11819 (.Y (nx11820), .A (gen_23_cmp_pMux_1)) ;
    inv04 ix11821 (.Y (nx11822), .A (gen_23_cmp_pMux_1)) ;
    inv02 ix11825 (.Y (nx11826), .A (nx11824)) ;
    inv02 ix11827 (.Y (nx11828), .A (nx11824)) ;
    inv02 ix11829 (.Y (nx11830), .A (nx11824)) ;
    inv02 ix11833 (.Y (nx11834), .A (nx11832)) ;
    inv02 ix11835 (.Y (nx11836), .A (nx11832)) ;
    inv02 ix11837 (.Y (nx11838), .A (nx11832)) ;
    inv02 ix11841 (.Y (nx11842), .A (nx11840)) ;
    inv02 ix11843 (.Y (nx11844), .A (nx11840)) ;
    inv02 ix11845 (.Y (nx11846), .A (nx11840)) ;
    inv02 ix11849 (.Y (nx11850), .A (nx11848)) ;
    inv02 ix11851 (.Y (nx11852), .A (nx11848)) ;
    inv02 ix11853 (.Y (nx11854), .A (nx11848)) ;
    inv04 ix11855 (.Y (nx11856), .A (gen_24_cmp_pMux_1)) ;
    inv04 ix11857 (.Y (nx11858), .A (gen_24_cmp_pMux_1)) ;
    inv04 ix11859 (.Y (nx11860), .A (gen_24_cmp_pMux_1)) ;
    inv04 ix11861 (.Y (nx11862), .A (gen_24_cmp_pMux_1)) ;
    inv02 ix11865 (.Y (nx11866), .A (nx11864)) ;
    inv02 ix11867 (.Y (nx11868), .A (nx11864)) ;
    inv02 ix11869 (.Y (nx11870), .A (nx11864)) ;
    inv02 ix11873 (.Y (nx11874), .A (nx11872)) ;
    inv02 ix11875 (.Y (nx11876), .A (nx11872)) ;
    inv02 ix11877 (.Y (nx11878), .A (nx11872)) ;
    inv02 ix11881 (.Y (nx11882), .A (nx11880)) ;
    inv02 ix11883 (.Y (nx11884), .A (nx11880)) ;
    inv02 ix11885 (.Y (nx11886), .A (nx11880)) ;
    nor02_2x ix3760 (.Y (nx10888), .A0 (nx3769), .A1 (gen_0_cmp_pMux_0)) ;
    nor02_2x ix3768 (.Y (nx10904), .A0 (gen_0_cmp_pMux_2), .A1 (nx3761)) ;
    xnor2 ix3778 (.Y (nx10912), .A0 (gen_0_cmp_pMux_0), .A1 (nx10900)) ;
    aoi21 ix3784 (.Y (nx10920), .A0 (gen_0_cmp_pMux_1), .A1 (gen_0_cmp_pMux_0), 
          .B0 (nx3769)) ;
    nor02_2x ix4004 (.Y (nx10928), .A0 (nx4013), .A1 (gen_1_cmp_pMux_0)) ;
    nor02_2x ix4012 (.Y (nx10944), .A0 (gen_1_cmp_pMux_2), .A1 (nx4005)) ;
    xnor2 ix4022 (.Y (nx10952), .A0 (gen_1_cmp_pMux_0), .A1 (nx10940)) ;
    aoi21 ix4028 (.Y (nx10960), .A0 (gen_1_cmp_pMux_1), .A1 (gen_1_cmp_pMux_0), 
          .B0 (nx4013)) ;
    nor02_2x ix4252 (.Y (nx10968), .A0 (nx4260), .A1 (gen_2_cmp_pMux_0)) ;
    nor02_2x ix4259 (.Y (nx10984), .A0 (gen_2_cmp_pMux_2), .A1 (nx4253)) ;
    xnor2 ix4270 (.Y (nx10992), .A0 (gen_2_cmp_pMux_0), .A1 (nx10980)) ;
    aoi21 ix4276 (.Y (nx11000), .A0 (gen_2_cmp_pMux_1), .A1 (gen_2_cmp_pMux_0), 
          .B0 (nx4260)) ;
    nor02_2x ix4500 (.Y (nx11008), .A0 (nx4509), .A1 (gen_3_cmp_pMux_0)) ;
    nor02_2x ix4508 (.Y (nx11024), .A0 (gen_3_cmp_pMux_2), .A1 (nx4501)) ;
    xnor2 ix4518 (.Y (nx11032), .A0 (gen_3_cmp_pMux_0), .A1 (nx11020)) ;
    aoi21 ix4524 (.Y (nx11040), .A0 (gen_3_cmp_pMux_1), .A1 (gen_3_cmp_pMux_0), 
          .B0 (nx4509)) ;
    nor02_2x ix4747 (.Y (nx11048), .A0 (nx4757), .A1 (gen_4_cmp_pMux_0)) ;
    nor02_2x ix4756 (.Y (nx11064), .A0 (gen_4_cmp_pMux_2), .A1 (nx4748)) ;
    xnor2 ix4766 (.Y (nx11072), .A0 (gen_4_cmp_pMux_0), .A1 (nx11060)) ;
    aoi21 ix4770 (.Y (nx11080), .A0 (gen_4_cmp_pMux_1), .A1 (gen_4_cmp_pMux_0), 
          .B0 (nx4757)) ;
    nor02_2x ix4994 (.Y (nx11088), .A0 (nx5003), .A1 (gen_5_cmp_pMux_0)) ;
    nor02_2x ix5002 (.Y (nx11104), .A0 (gen_5_cmp_pMux_2), .A1 (nx4995)) ;
    xnor2 ix5012 (.Y (nx11112), .A0 (gen_5_cmp_pMux_0), .A1 (nx11100)) ;
    aoi21 ix5018 (.Y (nx11120), .A0 (gen_5_cmp_pMux_1), .A1 (gen_5_cmp_pMux_0), 
          .B0 (nx5003)) ;
    nor02_2x ix5243 (.Y (nx11128), .A0 (nx5253), .A1 (gen_6_cmp_pMux_0)) ;
    nor02_2x ix5252 (.Y (nx11144), .A0 (gen_6_cmp_pMux_2), .A1 (nx5244)) ;
    xnor2 ix5262 (.Y (nx11152), .A0 (gen_6_cmp_pMux_0), .A1 (nx11140)) ;
    aoi21 ix5266 (.Y (nx11160), .A0 (gen_6_cmp_pMux_1), .A1 (gen_6_cmp_pMux_0), 
          .B0 (nx5253)) ;
    nor02_2x ix5490 (.Y (nx11168), .A0 (nx5499), .A1 (gen_7_cmp_pMux_0)) ;
    nor02_2x ix5498 (.Y (nx11184), .A0 (gen_7_cmp_pMux_2), .A1 (nx5491)) ;
    xnor2 ix5508 (.Y (nx11192), .A0 (gen_7_cmp_pMux_0), .A1 (nx11180)) ;
    aoi21 ix5512 (.Y (nx11200), .A0 (gen_7_cmp_pMux_1), .A1 (gen_7_cmp_pMux_0), 
          .B0 (nx5499)) ;
    nor02_2x ix5734 (.Y (nx11208), .A0 (nx5743), .A1 (gen_8_cmp_pMux_0)) ;
    nor02_2x ix5742 (.Y (nx11224), .A0 (gen_8_cmp_pMux_2), .A1 (nx5735)) ;
    xnor2 ix5752 (.Y (nx11232), .A0 (gen_8_cmp_pMux_0), .A1 (nx11220)) ;
    aoi21 ix5758 (.Y (nx11240), .A0 (gen_8_cmp_pMux_1), .A1 (gen_8_cmp_pMux_0), 
          .B0 (nx5743)) ;
    nor02_2x ix5978 (.Y (nx11248), .A0 (nx5987), .A1 (gen_9_cmp_pMux_0)) ;
    nor02_2x ix5986 (.Y (nx11264), .A0 (gen_9_cmp_pMux_2), .A1 (nx5979)) ;
    xnor2 ix5996 (.Y (nx11272), .A0 (gen_9_cmp_pMux_0), .A1 (nx11260)) ;
    aoi21 ix6002 (.Y (nx11280), .A0 (gen_9_cmp_pMux_1), .A1 (gen_9_cmp_pMux_0), 
          .B0 (nx5987)) ;
    nor02_2x ix6224 (.Y (nx11288), .A0 (nx6233), .A1 (gen_10_cmp_pMux_0)) ;
    nor02_2x ix6232 (.Y (nx11304), .A0 (gen_10_cmp_pMux_2), .A1 (nx6225)) ;
    xnor2 ix6242 (.Y (nx11312), .A0 (gen_10_cmp_pMux_0), .A1 (nx11300)) ;
    aoi21 ix6247 (.Y (nx11320), .A0 (gen_10_cmp_pMux_1), .A1 (gen_10_cmp_pMux_0)
          , .B0 (nx6233)) ;
    nor02_2x ix6467 (.Y (nx11328), .A0 (nx6477), .A1 (gen_11_cmp_pMux_0)) ;
    nor02_2x ix6476 (.Y (nx11344), .A0 (gen_11_cmp_pMux_2), .A1 (nx6468)) ;
    xnor2 ix6486 (.Y (nx11352), .A0 (gen_11_cmp_pMux_0), .A1 (nx11340)) ;
    aoi21 ix6490 (.Y (nx11360), .A0 (gen_11_cmp_pMux_1), .A1 (gen_11_cmp_pMux_0)
          , .B0 (nx6477)) ;
    nor02_2x ix6716 (.Y (nx11368), .A0 (nx6725), .A1 (gen_12_cmp_pMux_0)) ;
    nor02_2x ix6724 (.Y (nx11384), .A0 (gen_12_cmp_pMux_2), .A1 (nx6717)) ;
    xnor2 ix6734 (.Y (nx11392), .A0 (gen_12_cmp_pMux_0), .A1 (nx11380)) ;
    aoi21 ix6740 (.Y (nx11400), .A0 (gen_12_cmp_pMux_1), .A1 (gen_12_cmp_pMux_0)
          , .B0 (nx6725)) ;
    nor02_2x ix6963 (.Y (nx11408), .A0 (nx6973), .A1 (gen_13_cmp_pMux_0)) ;
    nor02_2x ix6972 (.Y (nx11424), .A0 (gen_13_cmp_pMux_2), .A1 (nx6965)) ;
    xnor2 ix6982 (.Y (nx11432), .A0 (gen_13_cmp_pMux_0), .A1 (nx11420)) ;
    aoi21 ix6988 (.Y (nx11440), .A0 (gen_13_cmp_pMux_1), .A1 (gen_13_cmp_pMux_0)
          , .B0 (nx6973)) ;
    nor02_2x ix7212 (.Y (nx11448), .A0 (nx7221), .A1 (gen_14_cmp_pMux_0)) ;
    nor02_2x ix7220 (.Y (nx11464), .A0 (gen_14_cmp_pMux_2), .A1 (nx7213)) ;
    xnor2 ix7230 (.Y (nx11472), .A0 (gen_14_cmp_pMux_0), .A1 (nx11460)) ;
    aoi21 ix7236 (.Y (nx11480), .A0 (gen_14_cmp_pMux_1), .A1 (gen_14_cmp_pMux_0)
          , .B0 (nx7221)) ;
    nor02_2x ix7461 (.Y (nx11488), .A0 (nx7471), .A1 (gen_15_cmp_pMux_0)) ;
    nor02_2x ix7470 (.Y (nx11504), .A0 (gen_15_cmp_pMux_2), .A1 (nx7463)) ;
    xnor2 ix7480 (.Y (nx11512), .A0 (gen_15_cmp_pMux_0), .A1 (nx11500)) ;
    aoi21 ix7486 (.Y (nx11520), .A0 (gen_15_cmp_pMux_1), .A1 (gen_15_cmp_pMux_0)
          , .B0 (nx7471)) ;
    nor02_2x ix7708 (.Y (nx11528), .A0 (nx7717), .A1 (gen_16_cmp_pMux_0)) ;
    nor02_2x ix7716 (.Y (nx11544), .A0 (gen_16_cmp_pMux_2), .A1 (nx7709)) ;
    xnor2 ix7726 (.Y (nx11552), .A0 (gen_16_cmp_pMux_0), .A1 (nx11540)) ;
    aoi21 ix7731 (.Y (nx11560), .A0 (gen_16_cmp_pMux_1), .A1 (gen_16_cmp_pMux_0)
          , .B0 (nx7717)) ;
    nor02_2x ix7952 (.Y (nx11568), .A0 (nx7961), .A1 (gen_17_cmp_pMux_0)) ;
    nor02_2x ix7960 (.Y (nx11584), .A0 (gen_17_cmp_pMux_2), .A1 (nx7953)) ;
    xnor2 ix7970 (.Y (nx11592), .A0 (gen_17_cmp_pMux_0), .A1 (nx11580)) ;
    aoi21 ix7976 (.Y (nx11600), .A0 (gen_17_cmp_pMux_1), .A1 (gen_17_cmp_pMux_0)
          , .B0 (nx7961)) ;
    nor02_2x ix8199 (.Y (nx11608), .A0 (nx8209), .A1 (gen_18_cmp_pMux_0)) ;
    nor02_2x ix8208 (.Y (nx11624), .A0 (gen_18_cmp_pMux_2), .A1 (nx8200)) ;
    xnor2 ix8218 (.Y (nx11632), .A0 (gen_18_cmp_pMux_0), .A1 (nx11620)) ;
    aoi21 ix8222 (.Y (nx11640), .A0 (gen_18_cmp_pMux_1), .A1 (gen_18_cmp_pMux_0)
          , .B0 (nx8209)) ;
    nor02_2x ix8446 (.Y (nx11648), .A0 (nx8455), .A1 (gen_19_cmp_pMux_0)) ;
    nor02_2x ix8454 (.Y (nx11664), .A0 (gen_19_cmp_pMux_2), .A1 (nx8447)) ;
    xnor2 ix8464 (.Y (nx11672), .A0 (gen_19_cmp_pMux_0), .A1 (nx11660)) ;
    aoi21 ix8470 (.Y (nx11680), .A0 (gen_19_cmp_pMux_1), .A1 (gen_19_cmp_pMux_0)
          , .B0 (nx8455)) ;
    nor02_2x ix8693 (.Y (nx11688), .A0 (nx8701), .A1 (gen_20_cmp_pMux_0)) ;
    nor02_2x ix8700 (.Y (nx11704), .A0 (gen_20_cmp_pMux_2), .A1 (nx8694)) ;
    xnor2 ix8710 (.Y (nx11712), .A0 (gen_20_cmp_pMux_0), .A1 (nx11700)) ;
    aoi21 ix8716 (.Y (nx11720), .A0 (gen_20_cmp_pMux_1), .A1 (gen_20_cmp_pMux_0)
          , .B0 (nx8701)) ;
    nor02_2x ix8936 (.Y (nx11728), .A0 (nx8945), .A1 (gen_21_cmp_pMux_0)) ;
    nor02_2x ix8944 (.Y (nx11744), .A0 (gen_21_cmp_pMux_2), .A1 (nx8937)) ;
    xnor2 ix8954 (.Y (nx11752), .A0 (gen_21_cmp_pMux_0), .A1 (nx11740)) ;
    aoi21 ix8960 (.Y (nx11760), .A0 (gen_21_cmp_pMux_1), .A1 (gen_21_cmp_pMux_0)
          , .B0 (nx8945)) ;
    nor02_2x ix9186 (.Y (nx11768), .A0 (nx9195), .A1 (gen_22_cmp_pMux_0)) ;
    nor02_2x ix9194 (.Y (nx11784), .A0 (gen_22_cmp_pMux_2), .A1 (nx9187)) ;
    xnor2 ix9204 (.Y (nx11792), .A0 (gen_22_cmp_pMux_0), .A1 (nx11780)) ;
    aoi21 ix9210 (.Y (nx11800), .A0 (gen_22_cmp_pMux_1), .A1 (gen_22_cmp_pMux_0)
          , .B0 (nx9195)) ;
    nor02_2x ix9435 (.Y (nx11808), .A0 (nx9445), .A1 (gen_23_cmp_pMux_0)) ;
    nor02_2x ix9444 (.Y (nx11824), .A0 (gen_23_cmp_pMux_2), .A1 (nx9437)) ;
    xnor2 ix9454 (.Y (nx11832), .A0 (gen_23_cmp_pMux_0), .A1 (nx11820)) ;
    aoi21 ix9460 (.Y (nx11840), .A0 (gen_23_cmp_pMux_1), .A1 (gen_23_cmp_pMux_0)
          , .B0 (nx9445)) ;
    nor02_2x ix9675 (.Y (nx11848), .A0 (nx9683), .A1 (gen_24_cmp_pMux_0)) ;
    nor02_2x ix9682 (.Y (nx11864), .A0 (gen_24_cmp_pMux_2), .A1 (nx9676)) ;
    xnor2 ix9691 (.Y (nx11872), .A0 (gen_24_cmp_pMux_0), .A1 (nx11860)) ;
    aoi21 ix9696 (.Y (nx11880), .A0 (gen_24_cmp_pMux_1), .A1 (gen_24_cmp_pMux_0)
          , .B0 (nx9683)) ;
    inv02 ix11895 (.Y (nx11896), .A (nx11938)) ;
    inv02 ix11897 (.Y (nx11898), .A (nx11938)) ;
    inv02 ix11899 (.Y (nx11900), .A (nx11938)) ;
    inv02 ix11901 (.Y (nx11902), .A (nx11938)) ;
    inv02 ix11903 (.Y (nx11904), .A (nx11938)) ;
    inv02 ix11905 (.Y (nx11906), .A (nx11938)) ;
    inv02 ix11907 (.Y (nx11908), .A (nx11940)) ;
    inv02 ix11909 (.Y (nx11910), .A (nx11940)) ;
    inv02 ix11911 (.Y (nx11912), .A (nx11940)) ;
    inv01 ix11913 (.Y (nx11914), .A (nx11940)) ;
    inv02 ix11915 (.Y (nx11916), .A (nx11934)) ;
    inv02 ix11917 (.Y (nx11918), .A (nx11936)) ;
    inv02 ix11919 (.Y (nx11920), .A (nx11936)) ;
    inv02 ix11921 (.Y (nx11922), .A (nx11936)) ;
    inv02 ix11923 (.Y (nx11924), .A (nx11936)) ;
    inv02 ix11925 (.Y (nx11926), .A (nx11936)) ;
    inv02 ix11927 (.Y (nx11928), .A (nx11936)) ;
    inv02 ix11933 (.Y (nx11934), .A (nx10880)) ;
    inv02 ix11935 (.Y (nx11936), .A (nx10880)) ;
    inv02 ix11937 (.Y (nx11938), .A (nx10120)) ;
    inv02 ix11939 (.Y (nx11940), .A (nx10120)) ;
endmodule


module NBitAdder_24 ( a, b, carryIn, sum, carryOut ) ;

    input [23:0]a ;
    input [23:0]b ;
    input carryIn ;
    output [23:0]sum ;
    output carryOut ;

    wire nx6, nx8, nx16, nx18, nx22, nx24, nx30, nx32, nx38, nx40, nx46, nx48, 
         nx54, nx56, nx62, nx64, nx70, nx72, nx78, nx80, nx86, nx88, nx94, nx96, 
         nx102, nx104, nx110, nx112, nx118, nx120, nx126, nx128, nx134, nx136, 
         nx142, nx144, nx150, nx152, nx158, nx160, nx166, nx168, nx170, nx172, 
         nx103, nx109, nx111, nx113, nx115, nx119, nx123, nx127, nx133, nx135, 
         nx137, nx141, nx145, nx149, nx155, nx157, nx159, nx163, nx167, nx171, 
         nx177, nx179, nx181, nx185, nx189, nx193, nx199, nx201, nx203, nx207, 
         nx211, nx215, nx221, nx223, nx225, nx229, nx232, nx235, nx239, nx241, 
         nx243, nx246, nx249, nx252, nx256, nx258, nx260, nx263, nx266, nx269, 
         nx273, nx275, nx277, nx280, nx283, nx286, nx290, nx292, nx294, nx297, 
         nx300, nx303, nx307, nx309, nx311, nx314, nx317, nx320, nx323, nx326, 
         nx329, nx332, nx335, nx338, nx341, nx344, nx347, nx350, nx353, nx356, 
         nx358, nx360, nx362, nx364, nx366, nx368, nx370, nx372;



    fake_gnd ix44 (.Y (carryOut)) ;
    xnor2 ix229 (.Y (sum[0]), .A0 (carryIn), .A1 (nx103)) ;
    xnor2 ix104 (.Y (nx103), .A0 (a[0]), .A1 (b[0])) ;
    xnor2 ix227 (.Y (sum[1]), .A0 (nx6), .A1 (nx115)) ;
    oai22 ix7 (.Y (nx6), .A0 (nx109), .A1 (nx103), .B0 (nx111), .B1 (nx113)) ;
    inv01 ix110 (.Y (nx109), .A (carryIn)) ;
    inv01 ix112 (.Y (nx111), .A (b[0])) ;
    inv01 ix114 (.Y (nx113), .A (a[0])) ;
    xnor2 ix116 (.Y (nx115), .A0 (a[1]), .A1 (b[1])) ;
    xnor2 ix225 (.Y (sum[2]), .A0 (nx119), .A1 (nx16)) ;
    aoi22 ix120 (.Y (nx119), .A0 (b[1]), .A1 (a[1]), .B0 (nx6), .B1 (nx8)) ;
    xnor2 ix9 (.Y (nx8), .A0 (a[1]), .A1 (nx123)) ;
    inv01 ix124 (.Y (nx123), .A (b[1])) ;
    xnor2 ix17 (.Y (nx16), .A0 (a[2]), .A1 (nx127)) ;
    inv01 ix128 (.Y (nx127), .A (b[2])) ;
    xnor2 ix223 (.Y (sum[3]), .A0 (nx22), .A1 (nx137)) ;
    oai21 ix23 (.Y (nx22), .A0 (nx119), .A1 (nx133), .B0 (nx135)) ;
    xnor2 ix134 (.Y (nx133), .A0 (a[2]), .A1 (b[2])) ;
    nand02 ix136 (.Y (nx135), .A0 (b[2]), .A1 (a[2])) ;
    xnor2 ix138 (.Y (nx137), .A0 (a[3]), .A1 (b[3])) ;
    xnor2 ix221 (.Y (sum[4]), .A0 (nx141), .A1 (nx32)) ;
    aoi22 ix142 (.Y (nx141), .A0 (b[3]), .A1 (a[3]), .B0 (nx22), .B1 (nx24)) ;
    xnor2 ix25 (.Y (nx24), .A0 (a[3]), .A1 (nx145)) ;
    inv01 ix146 (.Y (nx145), .A (b[3])) ;
    xnor2 ix33 (.Y (nx32), .A0 (a[4]), .A1 (nx149)) ;
    inv01 ix150 (.Y (nx149), .A (b[4])) ;
    xnor2 ix219 (.Y (sum[5]), .A0 (nx38), .A1 (nx159)) ;
    oai21 ix39 (.Y (nx38), .A0 (nx141), .A1 (nx155), .B0 (nx157)) ;
    xnor2 ix156 (.Y (nx155), .A0 (a[4]), .A1 (b[4])) ;
    nand02 ix158 (.Y (nx157), .A0 (b[4]), .A1 (a[4])) ;
    xnor2 ix160 (.Y (nx159), .A0 (a[5]), .A1 (b[5])) ;
    xnor2 ix217 (.Y (sum[6]), .A0 (nx163), .A1 (nx48)) ;
    aoi22 ix164 (.Y (nx163), .A0 (b[5]), .A1 (a[5]), .B0 (nx38), .B1 (nx40)) ;
    xnor2 ix41 (.Y (nx40), .A0 (a[5]), .A1 (nx167)) ;
    inv01 ix168 (.Y (nx167), .A (b[5])) ;
    xnor2 ix49 (.Y (nx48), .A0 (a[6]), .A1 (nx171)) ;
    inv01 ix172 (.Y (nx171), .A (b[6])) ;
    xnor2 ix215 (.Y (sum[7]), .A0 (nx54), .A1 (nx181)) ;
    oai21 ix55 (.Y (nx54), .A0 (nx163), .A1 (nx177), .B0 (nx179)) ;
    xnor2 ix178 (.Y (nx177), .A0 (a[6]), .A1 (b[6])) ;
    nand02 ix180 (.Y (nx179), .A0 (b[6]), .A1 (a[6])) ;
    xnor2 ix182 (.Y (nx181), .A0 (a[7]), .A1 (b[7])) ;
    xnor2 ix213 (.Y (sum[8]), .A0 (nx185), .A1 (nx64)) ;
    aoi22 ix186 (.Y (nx185), .A0 (b[7]), .A1 (a[7]), .B0 (nx54), .B1 (nx56)) ;
    xnor2 ix57 (.Y (nx56), .A0 (a[7]), .A1 (nx189)) ;
    inv01 ix190 (.Y (nx189), .A (b[7])) ;
    xnor2 ix65 (.Y (nx64), .A0 (a[8]), .A1 (nx193)) ;
    inv01 ix194 (.Y (nx193), .A (b[8])) ;
    xnor2 ix211 (.Y (sum[9]), .A0 (nx70), .A1 (nx203)) ;
    oai21 ix71 (.Y (nx70), .A0 (nx185), .A1 (nx199), .B0 (nx201)) ;
    xnor2 ix200 (.Y (nx199), .A0 (a[8]), .A1 (b[8])) ;
    nand02 ix202 (.Y (nx201), .A0 (b[8]), .A1 (a[8])) ;
    xnor2 ix204 (.Y (nx203), .A0 (a[9]), .A1 (b[9])) ;
    xnor2 ix209 (.Y (sum[10]), .A0 (nx207), .A1 (nx80)) ;
    aoi22 ix208 (.Y (nx207), .A0 (b[9]), .A1 (a[9]), .B0 (nx70), .B1 (nx72)) ;
    xnor2 ix73 (.Y (nx72), .A0 (a[9]), .A1 (nx211)) ;
    inv01 ix212 (.Y (nx211), .A (b[9])) ;
    xnor2 ix81 (.Y (nx80), .A0 (a[10]), .A1 (nx215)) ;
    inv01 ix216 (.Y (nx215), .A (b[10])) ;
    xnor2 ix207 (.Y (sum[11]), .A0 (nx86), .A1 (nx225)) ;
    oai21 ix87 (.Y (nx86), .A0 (nx207), .A1 (nx221), .B0 (nx223)) ;
    xnor2 ix222 (.Y (nx221), .A0 (a[10]), .A1 (b[10])) ;
    nand02 ix224 (.Y (nx223), .A0 (b[10]), .A1 (a[10])) ;
    xnor2 ix226 (.Y (nx225), .A0 (a[11]), .A1 (b[11])) ;
    xnor2 ix205 (.Y (sum[12]), .A0 (nx229), .A1 (nx96)) ;
    aoi22 ix230 (.Y (nx229), .A0 (b[11]), .A1 (a[11]), .B0 (nx86), .B1 (nx88)) ;
    xnor2 ix89 (.Y (nx88), .A0 (a[11]), .A1 (nx232)) ;
    inv01 ix233 (.Y (nx232), .A (b[11])) ;
    xnor2 ix97 (.Y (nx96), .A0 (a[12]), .A1 (nx235)) ;
    inv01 ix236 (.Y (nx235), .A (b[12])) ;
    xnor2 ix203 (.Y (sum[13]), .A0 (nx102), .A1 (nx243)) ;
    oai21 ix103 (.Y (nx102), .A0 (nx229), .A1 (nx239), .B0 (nx241)) ;
    xnor2 ix240 (.Y (nx239), .A0 (a[12]), .A1 (b[12])) ;
    nand02 ix242 (.Y (nx241), .A0 (b[12]), .A1 (a[12])) ;
    xnor2 ix244 (.Y (nx243), .A0 (a[13]), .A1 (b[13])) ;
    xnor2 ix201 (.Y (sum[14]), .A0 (nx246), .A1 (nx112)) ;
    aoi22 ix247 (.Y (nx246), .A0 (b[13]), .A1 (a[13]), .B0 (nx102), .B1 (nx104)
          ) ;
    xnor2 ix105 (.Y (nx104), .A0 (a[13]), .A1 (nx249)) ;
    inv01 ix250 (.Y (nx249), .A (b[13])) ;
    xnor2 ix113 (.Y (nx112), .A0 (a[14]), .A1 (nx252)) ;
    inv01 ix253 (.Y (nx252), .A (b[14])) ;
    xnor2 ix199 (.Y (sum[15]), .A0 (nx118), .A1 (nx260)) ;
    oai21 ix119 (.Y (nx118), .A0 (nx246), .A1 (nx256), .B0 (nx258)) ;
    xnor2 ix257 (.Y (nx256), .A0 (a[14]), .A1 (b[14])) ;
    nand02 ix259 (.Y (nx258), .A0 (b[14]), .A1 (a[14])) ;
    xnor2 ix261 (.Y (nx260), .A0 (a[15]), .A1 (b[15])) ;
    xnor2 ix197 (.Y (sum[16]), .A0 (nx263), .A1 (nx128)) ;
    aoi22 ix264 (.Y (nx263), .A0 (b[15]), .A1 (a[15]), .B0 (nx118), .B1 (nx120)
          ) ;
    xnor2 ix121 (.Y (nx120), .A0 (a[15]), .A1 (nx266)) ;
    inv01 ix267 (.Y (nx266), .A (b[15])) ;
    xnor2 ix129 (.Y (nx128), .A0 (a[16]), .A1 (nx269)) ;
    inv01 ix270 (.Y (nx269), .A (b[16])) ;
    xnor2 ix195 (.Y (sum[17]), .A0 (nx134), .A1 (nx277)) ;
    oai21 ix135 (.Y (nx134), .A0 (nx263), .A1 (nx273), .B0 (nx275)) ;
    xnor2 ix274 (.Y (nx273), .A0 (a[16]), .A1 (b[16])) ;
    nand02 ix276 (.Y (nx275), .A0 (b[16]), .A1 (a[16])) ;
    xnor2 ix278 (.Y (nx277), .A0 (a[17]), .A1 (b[17])) ;
    xnor2 ix193 (.Y (sum[18]), .A0 (nx280), .A1 (nx144)) ;
    aoi22 ix281 (.Y (nx280), .A0 (b[17]), .A1 (a[17]), .B0 (nx134), .B1 (nx136)
          ) ;
    xnor2 ix137 (.Y (nx136), .A0 (a[17]), .A1 (nx283)) ;
    inv01 ix284 (.Y (nx283), .A (b[17])) ;
    xnor2 ix145 (.Y (nx144), .A0 (a[18]), .A1 (nx286)) ;
    inv01 ix287 (.Y (nx286), .A (b[18])) ;
    xnor2 ix191 (.Y (sum[19]), .A0 (nx150), .A1 (nx294)) ;
    oai21 ix151 (.Y (nx150), .A0 (nx280), .A1 (nx290), .B0 (nx292)) ;
    xnor2 ix291 (.Y (nx290), .A0 (a[18]), .A1 (b[18])) ;
    nand02 ix293 (.Y (nx292), .A0 (b[18]), .A1 (a[18])) ;
    xnor2 ix295 (.Y (nx294), .A0 (a[19]), .A1 (b[19])) ;
    xnor2 ix189 (.Y (sum[20]), .A0 (nx297), .A1 (nx160)) ;
    aoi22 ix298 (.Y (nx297), .A0 (b[19]), .A1 (a[19]), .B0 (nx150), .B1 (nx152)
          ) ;
    xnor2 ix153 (.Y (nx152), .A0 (a[19]), .A1 (nx300)) ;
    inv01 ix301 (.Y (nx300), .A (b[19])) ;
    xnor2 ix161 (.Y (nx160), .A0 (a[20]), .A1 (nx303)) ;
    inv01 ix304 (.Y (nx303), .A (b[20])) ;
    xnor2 ix187 (.Y (sum[21]), .A0 (nx166), .A1 (nx311)) ;
    oai21 ix167 (.Y (nx166), .A0 (nx297), .A1 (nx307), .B0 (nx309)) ;
    xnor2 ix308 (.Y (nx307), .A0 (a[20]), .A1 (b[20])) ;
    nand02 ix310 (.Y (nx309), .A0 (b[20]), .A1 (a[20])) ;
    xnor2 ix312 (.Y (nx311), .A0 (a[21]), .A1 (b[21])) ;
    xnor2 ix185 (.Y (sum[22]), .A0 (b[22]), .A1 (nx314)) ;
    aoi22 ix315 (.Y (nx314), .A0 (b[21]), .A1 (a[21]), .B0 (nx166), .B1 (nx168)
          ) ;
    xnor2 ix169 (.Y (nx168), .A0 (a[21]), .A1 (nx317)) ;
    inv01 ix318 (.Y (nx317), .A (b[21])) ;
    xnor2 ix179 (.Y (sum[23]), .A0 (b[23]), .A1 (nx320)) ;
    oai21 ix321 (.Y (nx320), .A0 (nx172), .A1 (nx170), .B0 (b[22])) ;
    nor02_2x ix173 (.Y (nx172), .A0 (nx317), .A1 (nx323)) ;
    inv01 ix324 (.Y (nx323), .A (a[21])) ;
    nor02ii ix171 (.Y (nx170), .A0 (nx326), .A1 (nx168)) ;
    aoi22 ix327 (.Y (nx326), .A0 (b[20]), .A1 (a[20]), .B0 (nx158), .B1 (nx160)
          ) ;
    oai21 ix159 (.Y (nx158), .A0 (nx329), .A1 (nx294), .B0 (nx372)) ;
    aoi22 ix330 (.Y (nx329), .A0 (b[18]), .A1 (a[18]), .B0 (nx142), .B1 (nx144)
          ) ;
    oai21 ix143 (.Y (nx142), .A0 (nx332), .A1 (nx277), .B0 (nx370)) ;
    aoi22 ix333 (.Y (nx332), .A0 (b[16]), .A1 (a[16]), .B0 (nx126), .B1 (nx128)
          ) ;
    oai21 ix127 (.Y (nx126), .A0 (nx335), .A1 (nx260), .B0 (nx368)) ;
    aoi22 ix336 (.Y (nx335), .A0 (b[14]), .A1 (a[14]), .B0 (nx110), .B1 (nx112)
          ) ;
    oai21 ix111 (.Y (nx110), .A0 (nx338), .A1 (nx243), .B0 (nx366)) ;
    aoi22 ix339 (.Y (nx338), .A0 (b[12]), .A1 (a[12]), .B0 (nx94), .B1 (nx96)) ;
    oai21 ix95 (.Y (nx94), .A0 (nx341), .A1 (nx225), .B0 (nx364)) ;
    aoi22 ix342 (.Y (nx341), .A0 (b[10]), .A1 (a[10]), .B0 (nx78), .B1 (nx80)) ;
    oai21 ix79 (.Y (nx78), .A0 (nx344), .A1 (nx203), .B0 (nx362)) ;
    aoi22 ix345 (.Y (nx344), .A0 (b[8]), .A1 (a[8]), .B0 (nx62), .B1 (nx64)) ;
    oai21 ix63 (.Y (nx62), .A0 (nx347), .A1 (nx181), .B0 (nx360)) ;
    aoi22 ix348 (.Y (nx347), .A0 (b[6]), .A1 (a[6]), .B0 (nx46), .B1 (nx48)) ;
    oai21 ix47 (.Y (nx46), .A0 (nx350), .A1 (nx159), .B0 (nx358)) ;
    aoi22 ix351 (.Y (nx350), .A0 (b[4]), .A1 (a[4]), .B0 (nx30), .B1 (nx32)) ;
    oai21 ix31 (.Y (nx30), .A0 (nx353), .A1 (nx137), .B0 (nx356)) ;
    aoi21 ix354 (.Y (nx353), .A0 (b[2]), .A1 (a[2]), .B0 (nx18)) ;
    nor02ii ix19 (.Y (nx18), .A0 (nx119), .A1 (nx16)) ;
    nand02 ix357 (.Y (nx356), .A0 (b[3]), .A1 (a[3])) ;
    nand02 ix359 (.Y (nx358), .A0 (b[5]), .A1 (a[5])) ;
    nand02 ix361 (.Y (nx360), .A0 (b[7]), .A1 (a[7])) ;
    nand02 ix363 (.Y (nx362), .A0 (b[9]), .A1 (a[9])) ;
    nand02 ix365 (.Y (nx364), .A0 (b[11]), .A1 (a[11])) ;
    nand02 ix367 (.Y (nx366), .A0 (b[13]), .A1 (a[13])) ;
    nand02 ix369 (.Y (nx368), .A0 (b[15]), .A1 (a[15])) ;
    nand02 ix371 (.Y (nx370), .A0 (b[17]), .A1 (a[17])) ;
    nand02 ix373 (.Y (nx372), .A0 (b[19]), .A1 (a[19])) ;
endmodule


module BinaryMux_33 ( a, b, sel, f ) ;

    input [32:0]a ;
    input [32:0]b ;
    input sel ;
    output [32:0]f ;

    wire nx93, nx97, nx99, nx105, nx107, nx111, nx113, nx117, nx119, nx123, 
         nx125, nx129, nx131, nx135, nx137, nx141, nx143, nx147, nx151, nx155, 
         nx158, nx161, nx164, nx167, nx170, nx173, nx176, nx179, nx182, nx185, 
         nx188, nx191, nx194, nx197, nx200, nx203, nx206, nx209, nx212, nx219, 
         nx221, nx223, nx225, nx227, nx229, nx231;



    assign f[31] = f[32] ;
    fake_gnd ix44 (.Y (f[32])) ;
    nor02_2x ix3 (.Y (f[0]), .A0 (nx93), .A1 (nx219)) ;
    inv01 ix94 (.Y (nx93), .A (a[0])) ;
    nand02_2x ix99 (.Y (f[1]), .A0 (nx97), .A1 (nx99)) ;
    nand02 ix98 (.Y (nx97), .A0 (b[1]), .A1 (nx219)) ;
    nand02 ix100 (.Y (nx99), .A0 (a[1]), .A1 (nx229)) ;
    nand02 ix107 (.Y (f[2]), .A0 (nx105), .A1 (nx107)) ;
    nand02 ix106 (.Y (nx105), .A0 (b[2]), .A1 (nx219)) ;
    nand02 ix108 (.Y (nx107), .A0 (a[2]), .A1 (nx229)) ;
    nand02 ix115 (.Y (f[3]), .A0 (nx111), .A1 (nx113)) ;
    nand02 ix112 (.Y (nx111), .A0 (b[3]), .A1 (nx219)) ;
    nand02 ix114 (.Y (nx113), .A0 (a[3]), .A1 (nx229)) ;
    nand02 ix123 (.Y (f[4]), .A0 (nx117), .A1 (nx119)) ;
    nand02 ix118 (.Y (nx117), .A0 (b[4]), .A1 (nx219)) ;
    nand02 ix120 (.Y (nx119), .A0 (a[4]), .A1 (nx229)) ;
    nand02 ix131 (.Y (f[5]), .A0 (nx123), .A1 (nx125)) ;
    nand02 ix124 (.Y (nx123), .A0 (b[5]), .A1 (nx219)) ;
    nand02 ix126 (.Y (nx125), .A0 (a[5]), .A1 (nx229)) ;
    nand02 ix139 (.Y (f[6]), .A0 (nx129), .A1 (nx131)) ;
    nand02 ix130 (.Y (nx129), .A0 (b[6]), .A1 (nx219)) ;
    nand02 ix132 (.Y (nx131), .A0 (a[6]), .A1 (nx229)) ;
    nand02 ix147 (.Y (f[7]), .A0 (nx135), .A1 (nx137)) ;
    nand02 ix136 (.Y (nx135), .A0 (b[7]), .A1 (nx221)) ;
    nand02 ix138 (.Y (nx137), .A0 (a[7]), .A1 (nx229)) ;
    nand02 ix155 (.Y (f[8]), .A0 (nx141), .A1 (nx143)) ;
    nand02 ix142 (.Y (nx141), .A0 (nx221), .A1 (b[8])) ;
    nand02 ix144 (.Y (nx143), .A0 (nx231), .A1 (a[8])) ;
    nor02_2x ix7 (.Y (f[9]), .A0 (nx147), .A1 (nx221)) ;
    inv01 ix148 (.Y (nx147), .A (a[9])) ;
    nor02_2x ix11 (.Y (f[10]), .A0 (nx151), .A1 (nx221)) ;
    inv01 ix152 (.Y (nx151), .A (a[10])) ;
    nor02_2x ix15 (.Y (f[11]), .A0 (nx155), .A1 (nx221)) ;
    inv01 ix156 (.Y (nx155), .A (a[11])) ;
    nor02_2x ix19 (.Y (f[12]), .A0 (nx158), .A1 (nx221)) ;
    inv01 ix159 (.Y (nx158), .A (a[12])) ;
    nor02_2x ix23 (.Y (f[13]), .A0 (nx161), .A1 (nx221)) ;
    inv01 ix162 (.Y (nx161), .A (a[13])) ;
    nor02_2x ix27 (.Y (f[14]), .A0 (nx164), .A1 (nx223)) ;
    inv01 ix165 (.Y (nx164), .A (a[14])) ;
    nor02_2x ix31 (.Y (f[15]), .A0 (nx167), .A1 (nx223)) ;
    inv01 ix168 (.Y (nx167), .A (a[15])) ;
    nor02_2x ix35 (.Y (f[16]), .A0 (nx170), .A1 (nx223)) ;
    inv01 ix171 (.Y (nx170), .A (a[16])) ;
    nor02_2x ix39 (.Y (f[17]), .A0 (nx173), .A1 (nx223)) ;
    inv01 ix174 (.Y (nx173), .A (a[17])) ;
    nor02_2x ix43 (.Y (f[18]), .A0 (nx176), .A1 (nx223)) ;
    inv01 ix177 (.Y (nx176), .A (a[18])) ;
    nor02_2x ix47 (.Y (f[19]), .A0 (nx179), .A1 (nx223)) ;
    inv01 ix180 (.Y (nx179), .A (a[19])) ;
    nor02_2x ix51 (.Y (f[20]), .A0 (nx182), .A1 (nx223)) ;
    inv01 ix183 (.Y (nx182), .A (a[20])) ;
    nor02_2x ix55 (.Y (f[21]), .A0 (nx185), .A1 (nx225)) ;
    inv01 ix186 (.Y (nx185), .A (a[21])) ;
    nor02_2x ix59 (.Y (f[22]), .A0 (nx188), .A1 (nx225)) ;
    inv01 ix189 (.Y (nx188), .A (a[22])) ;
    nor02_2x ix63 (.Y (f[23]), .A0 (nx191), .A1 (nx225)) ;
    inv01 ix192 (.Y (nx191), .A (a[23])) ;
    nor02_2x ix67 (.Y (f[24]), .A0 (nx194), .A1 (nx225)) ;
    inv01 ix195 (.Y (nx194), .A (a[24])) ;
    nor02_2x ix71 (.Y (f[25]), .A0 (nx197), .A1 (nx225)) ;
    inv01 ix198 (.Y (nx197), .A (a[25])) ;
    nor02_2x ix75 (.Y (f[26]), .A0 (nx200), .A1 (nx225)) ;
    inv01 ix201 (.Y (nx200), .A (a[26])) ;
    nor02_2x ix79 (.Y (f[27]), .A0 (nx203), .A1 (nx225)) ;
    inv01 ix204 (.Y (nx203), .A (a[27])) ;
    nor02_2x ix83 (.Y (f[28]), .A0 (nx206), .A1 (nx227)) ;
    inv01 ix207 (.Y (nx206), .A (a[28])) ;
    nor02_2x ix87 (.Y (f[29]), .A0 (nx209), .A1 (nx227)) ;
    inv01 ix210 (.Y (nx209), .A (a[29])) ;
    nor02_2x ix91 (.Y (f[30]), .A0 (nx212), .A1 (nx227)) ;
    inv01 ix213 (.Y (nx212), .A (a[30])) ;
    inv02 ix218 (.Y (nx219), .A (nx231)) ;
    inv02 ix220 (.Y (nx221), .A (nx231)) ;
    inv02 ix222 (.Y (nx223), .A (nx231)) ;
    inv02 ix224 (.Y (nx225), .A (nx231)) ;
    inv02 ix226 (.Y (nx227), .A (nx231)) ;
    inv02 ix228 (.Y (nx229), .A (sel)) ;
    inv02 ix230 (.Y (nx231), .A (sel)) ;
endmodule


module Reg_33 ( D, en, clk, rst, Q ) ;

    input [32:0]D ;
    input en ;
    input clk ;
    input rst ;
    output [32:0]Q ;

    wire nx115, nx125, nx135, nx145, nx155, nx165, nx175, nx185, nx195, nx205, 
         nx215, nx225, nx235, nx245, nx255, nx265, nx275, nx285, nx295, nx305, 
         nx315, nx325, nx335, nx345, nx355, nx365, nx375, nx385, nx395, nx405, 
         nx415, nx427, nx431, nx436, nx438, nx443, nx445, nx450, nx452, nx457, 
         nx459, nx464, nx466, nx471, nx473, nx478, nx480, nx485, nx487, nx492, 
         nx494, nx499, nx501, nx506, nx508, nx513, nx515, nx520, nx522, nx527, 
         nx529, nx534, nx536, nx541, nx543, nx548, nx550, nx555, nx557, nx562, 
         nx564, nx569, nx571, nx576, nx578, nx583, nx585, nx590, nx592, nx597, 
         nx599, nx604, nx606, nx611, nx613, nx618, nx620, nx625, nx627, nx632, 
         nx634, nx639, nx641, nx649, nx651, nx653, nx655, nx657, nx663, nx665, 
         nx667, nx669, nx671, nx673, nx675, nx677, nx679, nx681, nx683, nx685;
    wire [30:0] \$dummy ;




    assign Q[31] = Q[32] ;
    fake_gnd ix43 (.Y (Q[32])) ;
    dffr reg_Q_0 (.Q (Q[0]), .QB (\$dummy [0]), .D (nx115), .CLK (nx665), .R (
         rst)) ;
    nand02 ix116 (.Y (nx115), .A0 (nx427), .A1 (nx431)) ;
    nand02 ix428 (.Y (nx427), .A0 (Q[0]), .A1 (nx685)) ;
    nand02 ix432 (.Y (nx431), .A0 (D[0]), .A1 (nx675)) ;
    dffr reg_Q_1 (.Q (Q[1]), .QB (\$dummy [1]), .D (nx125), .CLK (nx665), .R (
         rst)) ;
    nand02 ix126 (.Y (nx125), .A0 (nx436), .A1 (nx438)) ;
    nand02 ix437 (.Y (nx436), .A0 (Q[1]), .A1 (nx685)) ;
    nand02 ix439 (.Y (nx438), .A0 (D[1]), .A1 (nx675)) ;
    dffr reg_Q_2 (.Q (Q[2]), .QB (\$dummy [2]), .D (nx135), .CLK (nx665), .R (
         rst)) ;
    nand02 ix136 (.Y (nx135), .A0 (nx443), .A1 (nx445)) ;
    nand02 ix444 (.Y (nx443), .A0 (Q[2]), .A1 (nx685)) ;
    nand02 ix446 (.Y (nx445), .A0 (D[2]), .A1 (nx675)) ;
    dffr reg_Q_3 (.Q (Q[3]), .QB (\$dummy [3]), .D (nx145), .CLK (nx665), .R (
         rst)) ;
    nand02 ix146 (.Y (nx145), .A0 (nx450), .A1 (nx452)) ;
    nand02 ix451 (.Y (nx450), .A0 (Q[3]), .A1 (nx685)) ;
    nand02 ix453 (.Y (nx452), .A0 (D[3]), .A1 (nx675)) ;
    dffr reg_Q_4 (.Q (Q[4]), .QB (\$dummy [4]), .D (nx155), .CLK (nx665), .R (
         rst)) ;
    nand02 ix156 (.Y (nx155), .A0 (nx457), .A1 (nx459)) ;
    nand02 ix458 (.Y (nx457), .A0 (Q[4]), .A1 (nx685)) ;
    nand02 ix460 (.Y (nx459), .A0 (D[4]), .A1 (nx675)) ;
    dffr reg_Q_5 (.Q (Q[5]), .QB (\$dummy [5]), .D (nx165), .CLK (nx665), .R (
         rst)) ;
    nand02 ix166 (.Y (nx165), .A0 (nx464), .A1 (nx466)) ;
    nand02 ix465 (.Y (nx464), .A0 (Q[5]), .A1 (nx685)) ;
    nand02 ix467 (.Y (nx466), .A0 (D[5]), .A1 (nx675)) ;
    dffr reg_Q_6 (.Q (Q[6]), .QB (\$dummy [6]), .D (nx175), .CLK (nx665), .R (
         rst)) ;
    nand02 ix176 (.Y (nx175), .A0 (nx471), .A1 (nx473)) ;
    nand02 ix472 (.Y (nx471), .A0 (Q[6]), .A1 (nx685)) ;
    nand02 ix474 (.Y (nx473), .A0 (D[6]), .A1 (nx675)) ;
    dffr reg_Q_7 (.Q (Q[7]), .QB (\$dummy [7]), .D (nx185), .CLK (nx667), .R (
         rst)) ;
    nand02 ix186 (.Y (nx185), .A0 (nx478), .A1 (nx480)) ;
    nand02 ix479 (.Y (nx478), .A0 (Q[7]), .A1 (nx651)) ;
    nand02 ix481 (.Y (nx480), .A0 (D[7]), .A1 (nx677)) ;
    dffr reg_Q_8 (.Q (Q[8]), .QB (\$dummy [8]), .D (nx195), .CLK (nx667), .R (
         rst)) ;
    nand02 ix196 (.Y (nx195), .A0 (nx485), .A1 (nx487)) ;
    nand02 ix486 (.Y (nx485), .A0 (Q[8]), .A1 (nx651)) ;
    nand02 ix488 (.Y (nx487), .A0 (D[8]), .A1 (nx677)) ;
    dffr reg_Q_9 (.Q (Q[9]), .QB (\$dummy [9]), .D (nx205), .CLK (nx667), .R (
         rst)) ;
    nand02 ix206 (.Y (nx205), .A0 (nx492), .A1 (nx494)) ;
    nand02 ix493 (.Y (nx492), .A0 (Q[9]), .A1 (nx651)) ;
    nand02 ix495 (.Y (nx494), .A0 (D[9]), .A1 (nx677)) ;
    dffr reg_Q_10 (.Q (Q[10]), .QB (\$dummy [10]), .D (nx215), .CLK (nx667), .R (
         rst)) ;
    nand02 ix216 (.Y (nx215), .A0 (nx499), .A1 (nx501)) ;
    nand02 ix500 (.Y (nx499), .A0 (Q[10]), .A1 (nx651)) ;
    nand02 ix502 (.Y (nx501), .A0 (D[10]), .A1 (nx677)) ;
    dffr reg_Q_11 (.Q (Q[11]), .QB (\$dummy [11]), .D (nx225), .CLK (nx667), .R (
         rst)) ;
    nand02 ix226 (.Y (nx225), .A0 (nx506), .A1 (nx508)) ;
    nand02 ix507 (.Y (nx506), .A0 (Q[11]), .A1 (nx651)) ;
    nand02 ix509 (.Y (nx508), .A0 (D[11]), .A1 (nx677)) ;
    dffr reg_Q_12 (.Q (Q[12]), .QB (\$dummy [12]), .D (nx235), .CLK (nx667), .R (
         rst)) ;
    nand02 ix236 (.Y (nx235), .A0 (nx513), .A1 (nx515)) ;
    nand02 ix514 (.Y (nx513), .A0 (Q[12]), .A1 (nx651)) ;
    nand02 ix516 (.Y (nx515), .A0 (D[12]), .A1 (nx677)) ;
    dffr reg_Q_13 (.Q (Q[13]), .QB (\$dummy [13]), .D (nx245), .CLK (nx667), .R (
         rst)) ;
    nand02 ix246 (.Y (nx245), .A0 (nx520), .A1 (nx522)) ;
    nand02 ix521 (.Y (nx520), .A0 (Q[13]), .A1 (nx651)) ;
    nand02 ix523 (.Y (nx522), .A0 (D[13]), .A1 (nx677)) ;
    dffr reg_Q_14 (.Q (Q[14]), .QB (\$dummy [14]), .D (nx255), .CLK (nx669), .R (
         rst)) ;
    nand02 ix256 (.Y (nx255), .A0 (nx527), .A1 (nx529)) ;
    nand02 ix528 (.Y (nx527), .A0 (Q[14]), .A1 (nx653)) ;
    nand02 ix530 (.Y (nx529), .A0 (D[14]), .A1 (nx679)) ;
    dffr reg_Q_15 (.Q (Q[15]), .QB (\$dummy [15]), .D (nx265), .CLK (nx669), .R (
         rst)) ;
    nand02 ix266 (.Y (nx265), .A0 (nx534), .A1 (nx536)) ;
    nand02 ix535 (.Y (nx534), .A0 (Q[15]), .A1 (nx653)) ;
    nand02 ix537 (.Y (nx536), .A0 (D[15]), .A1 (nx679)) ;
    dffr reg_Q_16 (.Q (Q[16]), .QB (\$dummy [16]), .D (nx275), .CLK (nx669), .R (
         rst)) ;
    nand02 ix276 (.Y (nx275), .A0 (nx541), .A1 (nx543)) ;
    nand02 ix542 (.Y (nx541), .A0 (Q[16]), .A1 (nx653)) ;
    nand02 ix544 (.Y (nx543), .A0 (D[16]), .A1 (nx679)) ;
    dffr reg_Q_17 (.Q (Q[17]), .QB (\$dummy [17]), .D (nx285), .CLK (nx669), .R (
         rst)) ;
    nand02 ix286 (.Y (nx285), .A0 (nx548), .A1 (nx550)) ;
    nand02 ix549 (.Y (nx548), .A0 (Q[17]), .A1 (nx653)) ;
    nand02 ix551 (.Y (nx550), .A0 (D[17]), .A1 (nx679)) ;
    dffr reg_Q_18 (.Q (Q[18]), .QB (\$dummy [18]), .D (nx295), .CLK (nx669), .R (
         rst)) ;
    nand02 ix296 (.Y (nx295), .A0 (nx555), .A1 (nx557)) ;
    nand02 ix556 (.Y (nx555), .A0 (Q[18]), .A1 (nx653)) ;
    nand02 ix558 (.Y (nx557), .A0 (D[18]), .A1 (nx679)) ;
    dffr reg_Q_19 (.Q (Q[19]), .QB (\$dummy [19]), .D (nx305), .CLK (nx669), .R (
         rst)) ;
    nand02 ix306 (.Y (nx305), .A0 (nx562), .A1 (nx564)) ;
    nand02 ix563 (.Y (nx562), .A0 (Q[19]), .A1 (nx653)) ;
    nand02 ix565 (.Y (nx564), .A0 (D[19]), .A1 (nx679)) ;
    dffr reg_Q_20 (.Q (Q[20]), .QB (\$dummy [20]), .D (nx315), .CLK (nx669), .R (
         rst)) ;
    nand02 ix316 (.Y (nx315), .A0 (nx569), .A1 (nx571)) ;
    nand02 ix570 (.Y (nx569), .A0 (Q[20]), .A1 (nx653)) ;
    nand02 ix572 (.Y (nx571), .A0 (D[20]), .A1 (nx679)) ;
    dffr reg_Q_21 (.Q (Q[21]), .QB (\$dummy [21]), .D (nx325), .CLK (nx671), .R (
         rst)) ;
    nand02 ix326 (.Y (nx325), .A0 (nx576), .A1 (nx578)) ;
    nand02 ix577 (.Y (nx576), .A0 (Q[21]), .A1 (nx655)) ;
    nand02 ix579 (.Y (nx578), .A0 (D[21]), .A1 (nx681)) ;
    dffr reg_Q_22 (.Q (Q[22]), .QB (\$dummy [22]), .D (nx335), .CLK (nx671), .R (
         rst)) ;
    nand02 ix336 (.Y (nx335), .A0 (nx583), .A1 (nx585)) ;
    nand02 ix584 (.Y (nx583), .A0 (Q[22]), .A1 (nx655)) ;
    nand02 ix586 (.Y (nx585), .A0 (D[22]), .A1 (nx681)) ;
    dffr reg_Q_23 (.Q (Q[23]), .QB (\$dummy [23]), .D (nx345), .CLK (nx671), .R (
         rst)) ;
    nand02 ix346 (.Y (nx345), .A0 (nx590), .A1 (nx592)) ;
    nand02 ix591 (.Y (nx590), .A0 (Q[23]), .A1 (nx655)) ;
    nand02 ix593 (.Y (nx592), .A0 (D[23]), .A1 (nx681)) ;
    dffr reg_Q_24 (.Q (Q[24]), .QB (\$dummy [24]), .D (nx355), .CLK (nx671), .R (
         rst)) ;
    nand02 ix356 (.Y (nx355), .A0 (nx597), .A1 (nx599)) ;
    nand02 ix598 (.Y (nx597), .A0 (Q[24]), .A1 (nx655)) ;
    nand02 ix600 (.Y (nx599), .A0 (D[24]), .A1 (nx681)) ;
    dffr reg_Q_25 (.Q (Q[25]), .QB (\$dummy [25]), .D (nx365), .CLK (nx671), .R (
         rst)) ;
    nand02 ix366 (.Y (nx365), .A0 (nx604), .A1 (nx606)) ;
    nand02 ix605 (.Y (nx604), .A0 (Q[25]), .A1 (nx655)) ;
    nand02 ix607 (.Y (nx606), .A0 (D[25]), .A1 (nx681)) ;
    dffr reg_Q_26 (.Q (Q[26]), .QB (\$dummy [26]), .D (nx375), .CLK (nx671), .R (
         rst)) ;
    nand02 ix376 (.Y (nx375), .A0 (nx611), .A1 (nx613)) ;
    nand02 ix612 (.Y (nx611), .A0 (Q[26]), .A1 (nx655)) ;
    nand02 ix614 (.Y (nx613), .A0 (D[26]), .A1 (nx681)) ;
    dffr reg_Q_27 (.Q (Q[27]), .QB (\$dummy [27]), .D (nx385), .CLK (nx671), .R (
         rst)) ;
    nand02 ix386 (.Y (nx385), .A0 (nx618), .A1 (nx620)) ;
    nand02 ix619 (.Y (nx618), .A0 (Q[27]), .A1 (nx655)) ;
    nand02 ix621 (.Y (nx620), .A0 (D[27]), .A1 (nx681)) ;
    dffr reg_Q_28 (.Q (Q[28]), .QB (\$dummy [28]), .D (nx395), .CLK (nx673), .R (
         rst)) ;
    nand02 ix396 (.Y (nx395), .A0 (nx625), .A1 (nx627)) ;
    nand02 ix626 (.Y (nx625), .A0 (Q[28]), .A1 (nx657)) ;
    nand02 ix628 (.Y (nx627), .A0 (D[28]), .A1 (nx683)) ;
    dffr reg_Q_29 (.Q (Q[29]), .QB (\$dummy [29]), .D (nx405), .CLK (nx673), .R (
         rst)) ;
    nand02 ix406 (.Y (nx405), .A0 (nx632), .A1 (nx634)) ;
    nand02 ix633 (.Y (nx632), .A0 (Q[29]), .A1 (nx657)) ;
    nand02 ix635 (.Y (nx634), .A0 (D[29]), .A1 (nx683)) ;
    dffr reg_Q_30 (.Q (Q[30]), .QB (\$dummy [30]), .D (nx415), .CLK (nx673), .R (
         rst)) ;
    nand02 ix416 (.Y (nx415), .A0 (nx639), .A1 (nx641)) ;
    nand02 ix640 (.Y (nx639), .A0 (Q[30]), .A1 (nx657)) ;
    nand02 ix642 (.Y (nx641), .A0 (D[30]), .A1 (nx683)) ;
    inv02 ix648 (.Y (nx649), .A (en)) ;
    inv02 ix650 (.Y (nx651), .A (nx683)) ;
    inv02 ix652 (.Y (nx653), .A (nx683)) ;
    inv02 ix654 (.Y (nx655), .A (nx683)) ;
    inv02 ix656 (.Y (nx657), .A (nx683)) ;
    inv01 ix662 (.Y (nx663), .A (clk)) ;
    inv02 ix664 (.Y (nx665), .A (nx663)) ;
    inv02 ix666 (.Y (nx667), .A (nx663)) ;
    inv02 ix668 (.Y (nx669), .A (nx663)) ;
    inv02 ix670 (.Y (nx671), .A (nx663)) ;
    inv02 ix672 (.Y (nx673), .A (nx663)) ;
    inv02 ix674 (.Y (nx675), .A (nx649)) ;
    inv02 ix676 (.Y (nx677), .A (nx649)) ;
    inv02 ix678 (.Y (nx679), .A (nx649)) ;
    inv02 ix680 (.Y (nx681), .A (nx649)) ;
    inv02 ix682 (.Y (nx683), .A (nx649)) ;
    inv02 ix684 (.Y (nx685), .A (en)) ;
endmodule

