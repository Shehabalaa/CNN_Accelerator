library ieee;
use ieee.std_logic_1164.all;

package utiles is
	
	type genericarrayofvector16bit is array (natural range <>) of std_logic_vector(15 downto 0);
	type genericarrayofvector8bit is array (natural range <>) of std_logic_vector(7 downto 0);


end utiles;


-- package body section
package body utiles is

	
end utiles;


