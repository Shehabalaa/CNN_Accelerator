//
// Verilog description for cell CNNWithRAM, 
// Tue Apr 23 11:28:52 2019
//
// LeonardoSpectrum Level 3, 2018a.2 
//


module CNNWithRAM ( clk, rst, start, finishCNN ) ;

    input clk ;
    input rst ;
    input start ;
    output finishCNN ;

    wire weightsRamDataInBus_39, windowRamDataInBus_79, MFCWindowRam, 
         MFCWeightsRam, MFCWrite, weightsRamAddress_11, weightsRamAddress_10, 
         weightsRamAddress_9, weightsRamAddress_8, weightsRamAddress_7, 
         weightsRamAddress_6, weightsRamAddress_5, weightsRamAddress_4, 
         weightsRamAddress_3, weightsRamAddress_2, weightsRamAddress_1, 
         weightsRamAddress_0, windowRamAddressRead_12, windowRamAddressRead_11, 
         windowRamAddressRead_10, windowRamAddressRead_9, windowRamAddressRead_8, 
         windowRamAddressRead_7, windowRamAddressRead_6, windowRamAddressRead_5, 
         windowRamAddressRead_4, windowRamAddressRead_3, windowRamAddressRead_2, 
         windowRamAddressRead_1, windowRamAddressRead_0, 
         windowRamAddressWrite_12, windowRamAddressWrite_11, 
         windowRamAddressWrite_10, windowRamAddressWrite_9, 
         windowRamAddressWrite_8, windowRamAddressWrite_7, 
         windowRamAddressWrite_6, windowRamAddressWrite_5, 
         windowRamAddressWrite_4, windowRamAddressWrite_3, 
         windowRamAddressWrite_2, windowRamAddressWrite_1, 
         windowRamAddressWrite_0, weightsRamRead, windowRamRead, windowRamWrite, 
         GND;
    wire [134:0] \$dummy ;




    CNNModule_8_16_5_5_3_12_13 CNNMap (.startCNN (start), .clk (clk), .rst (rst)
                               , .weightsRamDataInBus ({weightsRamDataInBus_39,
                               weightsRamDataInBus_39,weightsRamDataInBus_39,
                               weightsRamDataInBus_39,weightsRamDataInBus_39,
                               weightsRamDataInBus_39,weightsRamDataInBus_39,
                               weightsRamDataInBus_39,weightsRamDataInBus_39,
                               weightsRamDataInBus_39,weightsRamDataInBus_39,
                               weightsRamDataInBus_39,weightsRamDataInBus_39,
                               weightsRamDataInBus_39,weightsRamDataInBus_39,
                               weightsRamDataInBus_39,weightsRamDataInBus_39,
                               weightsRamDataInBus_39,weightsRamDataInBus_39,
                               weightsRamDataInBus_39,weightsRamDataInBus_39,
                               weightsRamDataInBus_39,weightsRamDataInBus_39,
                               weightsRamDataInBus_39,weightsRamDataInBus_39,
                               weightsRamDataInBus_39,weightsRamDataInBus_39,
                               weightsRamDataInBus_39,weightsRamDataInBus_39,
                               weightsRamDataInBus_39,weightsRamDataInBus_39,
                               weightsRamDataInBus_39,weightsRamDataInBus_39,
                               weightsRamDataInBus_39,weightsRamDataInBus_39,
                               weightsRamDataInBus_39,weightsRamDataInBus_39,
                               weightsRamDataInBus_39,weightsRamDataInBus_39,
                               weightsRamDataInBus_39}), .windowRamDataInBus ({
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79,
                               windowRamDataInBus_79,windowRamDataInBus_79}), .MFCWindowRam (
                               MFCWindowRam), .MFCWeightsRam (MFCWeightsRam), .MFCWrite (
                               MFCWrite), .weightsRamAddress ({
                               weightsRamAddress_11,weightsRamAddress_10,
                               weightsRamAddress_9,weightsRamAddress_8,
                               weightsRamAddress_7,weightsRamAddress_6,
                               weightsRamAddress_5,weightsRamAddress_4,
                               weightsRamAddress_3,weightsRamAddress_2,
                               weightsRamAddress_1,weightsRamAddress_0}), .windowRamAddressRead (
                               {windowRamAddressRead_12,windowRamAddressRead_11,
                               windowRamAddressRead_10,windowRamAddressRead_9,
                               windowRamAddressRead_8,windowRamAddressRead_7,
                               windowRamAddressRead_6,windowRamAddressRead_5,
                               windowRamAddressRead_4,windowRamAddressRead_3,
                               windowRamAddressRead_2,windowRamAddressRead_1,
                               windowRamAddressRead_0}), .windowRamAddressWrite (
                               {windowRamAddressWrite_12,
                               windowRamAddressWrite_11,windowRamAddressWrite_10
                               ,windowRamAddressWrite_9,windowRamAddressWrite_8,
                               windowRamAddressWrite_7,windowRamAddressWrite_6,
                               windowRamAddressWrite_5,windowRamAddressWrite_4,
                               windowRamAddressWrite_3,windowRamAddressWrite_2,
                               windowRamAddressWrite_1,windowRamAddressWrite_0})
                               , .weightsRamRead (weightsRamRead), .windowRamRead (
                               windowRamRead), .windowRamWrite (windowRamWrite)
                               , .windowRamDataOutBus ({\$dummy [0],\$dummy [1],
                               \$dummy [2],\$dummy [3],\$dummy [4],\$dummy [5],
                               \$dummy [6],\$dummy [7],\$dummy [8],\$dummy [9],
                               \$dummy [10],\$dummy [11],\$dummy [12],
                               \$dummy [13],\$dummy [14],\$dummy [15]}), .finishNetwork (
                               finishCNN)) ;
    RAM_12_8_40 weightsRam (.clk (clk), .rd (weightsRamRead), .we (GND), .reset (
                rst), .addressRead ({weightsRamAddress_11,weightsRamAddress_10,
                weightsRamAddress_9,weightsRamAddress_8,weightsRamAddress_7,
                weightsRamAddress_6,weightsRamAddress_5,weightsRamAddress_4,
                weightsRamAddress_3,weightsRamAddress_2,weightsRamAddress_1,
                weightsRamAddress_0}), .addressWrite ({weightsRamAddress_11,
                weightsRamAddress_10,weightsRamAddress_9,weightsRamAddress_8,
                weightsRamAddress_7,weightsRamAddress_6,weightsRamAddress_5,
                weightsRamAddress_4,weightsRamAddress_3,weightsRamAddress_2,
                weightsRamAddress_1,weightsRamAddress_0}), .dataIn ({GND,GND,GND
                ,GND,GND,GND,GND,GND}), .dataOut ({weightsRamDataInBus_39,
                \$dummy [16],\$dummy [17],\$dummy [18],\$dummy [19],\$dummy [20]
                ,\$dummy [21],\$dummy [22],\$dummy [23],\$dummy [24],
                \$dummy [25],\$dummy [26],\$dummy [27],\$dummy [28],\$dummy [29]
                ,\$dummy [30],\$dummy [31],\$dummy [32],\$dummy [33],
                \$dummy [34],\$dummy [35],\$dummy [36],\$dummy [37],\$dummy [38]
                ,\$dummy [39],\$dummy [40],\$dummy [41],\$dummy [42],
                \$dummy [43],\$dummy [44],\$dummy [45],\$dummy [46],\$dummy [47]
                ,\$dummy [48],\$dummy [49],\$dummy [50],\$dummy [51],
                \$dummy [52],\$dummy [53],\$dummy [54]}), .MFCReadOut (
                MFCWeightsRam), .MFCWriteOut (\$dummy [55])) ;
    RAM_13_16_80 windowRam (.clk (clk), .rd (windowRamRead), .we (windowRamWrite
                 ), .reset (rst), .addressRead ({windowRamAddressRead_12,
                 windowRamAddressRead_11,windowRamAddressRead_10,
                 windowRamAddressRead_9,windowRamAddressRead_8,
                 windowRamAddressRead_7,windowRamAddressRead_6,
                 windowRamAddressRead_5,windowRamAddressRead_4,
                 windowRamAddressRead_3,windowRamAddressRead_2,
                 windowRamAddressRead_1,windowRamAddressRead_0}), .addressWrite (
                 {windowRamAddressWrite_12,windowRamAddressWrite_11,
                 windowRamAddressWrite_10,windowRamAddressWrite_9,
                 windowRamAddressWrite_8,windowRamAddressWrite_7,
                 windowRamAddressWrite_6,windowRamAddressWrite_5,
                 windowRamAddressWrite_4,windowRamAddressWrite_3,
                 windowRamAddressWrite_2,windowRamAddressWrite_1,
                 windowRamAddressWrite_0}), .dataIn ({GND,GND,GND,GND,GND,GND,
                 GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}), .dataOut ({
                 windowRamDataInBus_79,\$dummy [56],\$dummy [57],\$dummy [58],
                 \$dummy [59],\$dummy [60],\$dummy [61],\$dummy [62],
                 \$dummy [63],\$dummy [64],\$dummy [65],\$dummy [66],
                 \$dummy [67],\$dummy [68],\$dummy [69],\$dummy [70],
                 \$dummy [71],\$dummy [72],\$dummy [73],\$dummy [74],
                 \$dummy [75],\$dummy [76],\$dummy [77],\$dummy [78],
                 \$dummy [79],\$dummy [80],\$dummy [81],\$dummy [82],
                 \$dummy [83],\$dummy [84],\$dummy [85],\$dummy [86],
                 \$dummy [87],\$dummy [88],\$dummy [89],\$dummy [90],
                 \$dummy [91],\$dummy [92],\$dummy [93],\$dummy [94],
                 \$dummy [95],\$dummy [96],\$dummy [97],\$dummy [98],
                 \$dummy [99],\$dummy [100],\$dummy [101],\$dummy [102],
                 \$dummy [103],\$dummy [104],\$dummy [105],\$dummy [106],
                 \$dummy [107],\$dummy [108],\$dummy [109],\$dummy [110],
                 \$dummy [111],\$dummy [112],\$dummy [113],\$dummy [114],
                 \$dummy [115],\$dummy [116],\$dummy [117],\$dummy [118],
                 \$dummy [119],\$dummy [120],\$dummy [121],\$dummy [122],
                 \$dummy [123],\$dummy [124],\$dummy [125],\$dummy [126],
                 \$dummy [127],\$dummy [128],\$dummy [129],\$dummy [130],
                 \$dummy [131],\$dummy [132],\$dummy [133],\$dummy [134]}), .MFCReadOut (
                 MFCWindowRam), .MFCWriteOut (MFCWrite)) ;
    fake_gnd ix305 (.Y (GND)) ;
endmodule


module RAM_13_16_80 ( clk, rd, we, reset, addressRead, addressWrite, dataIn, 
                      dataOut, MFCReadOut, MFCWriteOut ) ;

    input clk ;
    input rd ;
    input we ;
    input reset ;
    input [12:0]addressRead ;
    input [12:0]addressWrite ;
    input [15:0]dataIn ;
    output [79:0]dataOut ;
    output MFCReadOut ;
    output MFCWriteOut ;

    wire NOT_clk, nx84, NOT_nx84, nx255, nx257, nx259, nx261, nx263, nx265, 
         nx267, nx269, nx271, nx273, nx275, nx277, nx279, nx281, nx283, nx285, 
         nx287, nx289;
    wire [1:0] \$dummy ;




    assign dataOut[78] = dataOut[79] ;
    assign dataOut[77] = dataOut[79] ;
    assign dataOut[76] = dataOut[79] ;
    assign dataOut[75] = dataOut[79] ;
    assign dataOut[74] = dataOut[79] ;
    assign dataOut[73] = dataOut[79] ;
    assign dataOut[72] = dataOut[79] ;
    assign dataOut[71] = dataOut[79] ;
    assign dataOut[70] = dataOut[79] ;
    assign dataOut[69] = dataOut[79] ;
    assign dataOut[68] = dataOut[79] ;
    assign dataOut[67] = dataOut[79] ;
    assign dataOut[66] = dataOut[79] ;
    assign dataOut[65] = dataOut[79] ;
    assign dataOut[64] = dataOut[79] ;
    assign dataOut[63] = dataOut[79] ;
    assign dataOut[62] = dataOut[79] ;
    assign dataOut[61] = dataOut[79] ;
    assign dataOut[60] = dataOut[79] ;
    assign dataOut[59] = dataOut[79] ;
    assign dataOut[58] = dataOut[79] ;
    assign dataOut[57] = dataOut[79] ;
    assign dataOut[56] = dataOut[79] ;
    assign dataOut[55] = dataOut[79] ;
    assign dataOut[54] = dataOut[79] ;
    assign dataOut[53] = dataOut[79] ;
    assign dataOut[52] = dataOut[79] ;
    assign dataOut[51] = dataOut[79] ;
    assign dataOut[50] = dataOut[79] ;
    assign dataOut[49] = dataOut[79] ;
    assign dataOut[48] = dataOut[79] ;
    assign dataOut[47] = dataOut[79] ;
    assign dataOut[46] = dataOut[79] ;
    assign dataOut[45] = dataOut[79] ;
    assign dataOut[44] = dataOut[79] ;
    assign dataOut[43] = dataOut[79] ;
    assign dataOut[42] = dataOut[79] ;
    assign dataOut[41] = dataOut[79] ;
    assign dataOut[40] = dataOut[79] ;
    assign dataOut[39] = dataOut[79] ;
    assign dataOut[38] = dataOut[79] ;
    assign dataOut[37] = dataOut[79] ;
    assign dataOut[36] = dataOut[79] ;
    assign dataOut[35] = dataOut[79] ;
    assign dataOut[34] = dataOut[79] ;
    assign dataOut[33] = dataOut[79] ;
    assign dataOut[32] = dataOut[79] ;
    assign dataOut[31] = dataOut[79] ;
    assign dataOut[30] = dataOut[79] ;
    assign dataOut[29] = dataOut[79] ;
    assign dataOut[28] = dataOut[79] ;
    assign dataOut[27] = dataOut[79] ;
    assign dataOut[26] = dataOut[79] ;
    assign dataOut[25] = dataOut[79] ;
    assign dataOut[24] = dataOut[79] ;
    assign dataOut[23] = dataOut[79] ;
    assign dataOut[22] = dataOut[79] ;
    assign dataOut[21] = dataOut[79] ;
    assign dataOut[20] = dataOut[79] ;
    assign dataOut[19] = dataOut[79] ;
    assign dataOut[18] = dataOut[79] ;
    assign dataOut[17] = dataOut[79] ;
    assign dataOut[16] = dataOut[79] ;
    assign dataOut[15] = dataOut[79] ;
    assign dataOut[14] = dataOut[79] ;
    assign dataOut[13] = dataOut[79] ;
    assign dataOut[12] = dataOut[79] ;
    assign dataOut[11] = dataOut[79] ;
    assign dataOut[10] = dataOut[79] ;
    assign dataOut[9] = dataOut[79] ;
    assign dataOut[8] = dataOut[79] ;
    assign dataOut[7] = dataOut[79] ;
    assign dataOut[6] = dataOut[79] ;
    assign dataOut[5] = dataOut[79] ;
    assign dataOut[4] = dataOut[79] ;
    assign dataOut[3] = dataOut[79] ;
    assign dataOut[2] = dataOut[79] ;
    assign dataOut[1] = dataOut[79] ;
    assign dataOut[0] = dataOut[79] ;
    fake_gnd ix213 (.Y (dataOut[79])) ;
    dff reg_MFCWriteOut (.Q (MFCWriteOut), .QB (\$dummy [0]), .D (NOT_nx84), .CLK (
        NOT_clk)) ;
    nand04 ix256 (.Y (nx255), .A0 (nx257), .A1 (we), .A2 (rd), .A3 (nx259)) ;
    inv01 ix258 (.Y (nx257), .A (reset)) ;
    xnor2 ix260 (.Y (nx259), .A0 (addressRead[0]), .A1 (addressWrite[0])) ;
    nand04 ix262 (.Y (nx261), .A0 (nx263), .A1 (nx265), .A2 (nx267), .A3 (nx269)
           ) ;
    xnor2 ix264 (.Y (nx263), .A0 (addressRead[1]), .A1 (addressWrite[1])) ;
    xnor2 ix266 (.Y (nx265), .A0 (addressRead[2]), .A1 (addressWrite[2])) ;
    xnor2 ix268 (.Y (nx267), .A0 (addressRead[3]), .A1 (addressWrite[3])) ;
    xnor2 ix270 (.Y (nx269), .A0 (addressRead[4]), .A1 (addressWrite[4])) ;
    nand04 ix272 (.Y (nx271), .A0 (nx273), .A1 (nx275), .A2 (nx277), .A3 (nx279)
           ) ;
    xnor2 ix274 (.Y (nx273), .A0 (addressRead[5]), .A1 (addressWrite[5])) ;
    xnor2 ix276 (.Y (nx275), .A0 (addressRead[6]), .A1 (addressWrite[6])) ;
    xnor2 ix278 (.Y (nx277), .A0 (addressRead[7]), .A1 (addressWrite[7])) ;
    xnor2 ix280 (.Y (nx279), .A0 (addressRead[12]), .A1 (addressWrite[12])) ;
    nand04 ix282 (.Y (nx281), .A0 (nx283), .A1 (nx285), .A2 (nx287), .A3 (nx289)
           ) ;
    xnor2 ix284 (.Y (nx283), .A0 (addressRead[8]), .A1 (addressWrite[8])) ;
    xnor2 ix286 (.Y (nx285), .A0 (addressRead[9]), .A1 (addressWrite[9])) ;
    xnor2 ix288 (.Y (nx287), .A0 (addressRead[10]), .A1 (addressWrite[10])) ;
    xnor2 ix290 (.Y (nx289), .A0 (addressRead[11]), .A1 (addressWrite[11])) ;
    inv01 ix292 (.Y (NOT_clk), .A (clk)) ;
    dff reg_MFCReadOut (.Q (MFCReadOut), .QB (\$dummy [1]), .D (nx84), .CLK (
        NOT_clk)) ;
    nor04 ix85 (.Y (nx84), .A0 (nx255), .A1 (nx261), .A2 (nx271), .A3 (nx281)) ;
    inv01 ix254 (.Y (NOT_nx84), .A (nx84)) ;
endmodule


module RAM_12_8_40 ( clk, rd, we, reset, addressRead, addressWrite, dataIn, 
                     dataOut, MFCReadOut, MFCWriteOut ) ;

    input clk ;
    input rd ;
    input we ;
    input reset ;
    input [11:0]addressRead ;
    input [11:0]addressWrite ;
    input [7:0]dataIn ;
    output [39:0]dataOut ;
    output MFCReadOut ;
    output MFCWriteOut ;

    wire NOT_clk, nx78, NOT_nx78, nx173, nx175, nx177, nx179, nx181, nx183, 
         nx185, nx187, nx189, nx191, nx193, nx195, nx197, nx199, nx201, nx203, 
         nx205;
    wire [1:0] \$dummy ;




    assign dataOut[38] = dataOut[39] ;
    assign dataOut[37] = dataOut[39] ;
    assign dataOut[36] = dataOut[39] ;
    assign dataOut[35] = dataOut[39] ;
    assign dataOut[34] = dataOut[39] ;
    assign dataOut[33] = dataOut[39] ;
    assign dataOut[32] = dataOut[39] ;
    assign dataOut[31] = dataOut[39] ;
    assign dataOut[30] = dataOut[39] ;
    assign dataOut[29] = dataOut[39] ;
    assign dataOut[28] = dataOut[39] ;
    assign dataOut[27] = dataOut[39] ;
    assign dataOut[26] = dataOut[39] ;
    assign dataOut[25] = dataOut[39] ;
    assign dataOut[24] = dataOut[39] ;
    assign dataOut[23] = dataOut[39] ;
    assign dataOut[22] = dataOut[39] ;
    assign dataOut[21] = dataOut[39] ;
    assign dataOut[20] = dataOut[39] ;
    assign dataOut[19] = dataOut[39] ;
    assign dataOut[18] = dataOut[39] ;
    assign dataOut[17] = dataOut[39] ;
    assign dataOut[16] = dataOut[39] ;
    assign dataOut[15] = dataOut[39] ;
    assign dataOut[14] = dataOut[39] ;
    assign dataOut[13] = dataOut[39] ;
    assign dataOut[12] = dataOut[39] ;
    assign dataOut[11] = dataOut[39] ;
    assign dataOut[10] = dataOut[39] ;
    assign dataOut[9] = dataOut[39] ;
    assign dataOut[8] = dataOut[39] ;
    assign dataOut[7] = dataOut[39] ;
    assign dataOut[6] = dataOut[39] ;
    assign dataOut[5] = dataOut[39] ;
    assign dataOut[4] = dataOut[39] ;
    assign dataOut[3] = dataOut[39] ;
    assign dataOut[2] = dataOut[39] ;
    assign dataOut[1] = dataOut[39] ;
    assign dataOut[0] = dataOut[39] ;
    fake_gnd ix133 (.Y (dataOut[39])) ;
    dff reg_MFCWriteOut (.Q (MFCWriteOut), .QB (\$dummy [0]), .D (NOT_nx78), .CLK (
        NOT_clk)) ;
    nand04 ix174 (.Y (nx173), .A0 (nx175), .A1 (we), .A2 (rd), .A3 (nx177)) ;
    inv01 ix176 (.Y (nx175), .A (reset)) ;
    xnor2 ix178 (.Y (nx177), .A0 (addressRead[0]), .A1 (addressWrite[0])) ;
    nand04 ix180 (.Y (nx179), .A0 (nx181), .A1 (nx183), .A2 (nx185), .A3 (nx187)
           ) ;
    xnor2 ix182 (.Y (nx181), .A0 (addressRead[1]), .A1 (addressWrite[1])) ;
    xnor2 ix184 (.Y (nx183), .A0 (addressRead[2]), .A1 (addressWrite[2])) ;
    xnor2 ix186 (.Y (nx185), .A0 (addressRead[3]), .A1 (addressWrite[3])) ;
    xnor2 ix188 (.Y (nx187), .A0 (addressRead[4]), .A1 (addressWrite[4])) ;
    nand04 ix190 (.Y (nx189), .A0 (nx191), .A1 (nx193), .A2 (nx195), .A3 (nx197)
           ) ;
    xnor2 ix192 (.Y (nx191), .A0 (addressRead[5]), .A1 (addressWrite[5])) ;
    xnor2 ix194 (.Y (nx193), .A0 (addressRead[6]), .A1 (addressWrite[6])) ;
    xnor2 ix196 (.Y (nx195), .A0 (addressRead[7]), .A1 (addressWrite[7])) ;
    xnor2 ix198 (.Y (nx197), .A0 (addressRead[8]), .A1 (addressWrite[8])) ;
    nand03 ix200 (.Y (nx199), .A0 (nx201), .A1 (nx203), .A2 (nx205)) ;
    xnor2 ix202 (.Y (nx201), .A0 (addressRead[11]), .A1 (addressWrite[11])) ;
    xnor2 ix204 (.Y (nx203), .A0 (addressRead[9]), .A1 (addressWrite[9])) ;
    xnor2 ix206 (.Y (nx205), .A0 (addressRead[10]), .A1 (addressWrite[10])) ;
    inv01 ix208 (.Y (NOT_clk), .A (clk)) ;
    dff reg_MFCReadOut (.Q (MFCReadOut), .QB (\$dummy [1]), .D (nx78), .CLK (
        NOT_clk)) ;
    nor04 ix79 (.Y (nx78), .A0 (nx173), .A1 (nx179), .A2 (nx189), .A3 (nx199)) ;
    inv01 ix172 (.Y (NOT_nx78), .A (nx78)) ;
endmodule


module CNNModule_8_16_5_5_3_12_13 ( startCNN, clk, rst, weightsRamDataInBus, 
                                    windowRamDataInBus, MFCWindowRam, 
                                    MFCWeightsRam, MFCWrite, weightsRamAddress, 
                                    windowRamAddressRead, windowRamAddressWrite, 
                                    weightsRamRead, windowRamRead, 
                                    windowRamWrite, windowRamDataOutBus, 
                                    finishNetwork ) ;

    input startCNN ;
    input clk ;
    input rst ;
    input [39:0]weightsRamDataInBus ;
    input [79:0]windowRamDataInBus ;
    input MFCWindowRam ;
    input MFCWeightsRam ;
    input MFCWrite ;
    output [11:0]weightsRamAddress ;
    output [12:0]windowRamAddressRead ;
    output [12:0]windowRamAddressWrite ;
    output weightsRamRead ;
    output windowRamRead ;
    output windowRamWrite ;
    output [15:0]windowRamDataOutBus ;
    output finishNetwork ;

    wire conv, pool, layerType, filterType, currentPage_0, filterBus_39, 
         filterBus_38, filterBus_37, filterBus_36, filterBus_35, filterBus_34, 
         filterBus_33, filterBus_32, filterBus_31, filterBus_30, filterBus_29, 
         filterBus_28, filterBus_27, filterBus_26, filterBus_25, filterBus_24, 
         filterBus_23, filterBus_22, filterBus_21, filterBus_20, filterBus_19, 
         filterBus_18, filterBus_17, filterBus_16, filterBus_15, filterBus_14, 
         filterBus_13, filterBus_12, filterBus_11, filterBus_10, filterBus_9, 
         filterBus_8, filterBus_7, filterBus_6, filterBus_5, filterBus_4, 
         filterBus_3, filterBus_2, filterBus_1, filterBus_0, windowBus_79, 
         windowBus_78, windowBus_77, windowBus_76, windowBus_75, windowBus_74, 
         windowBus_73, windowBus_72, windowBus_71, windowBus_70, windowBus_69, 
         windowBus_68, windowBus_67, windowBus_66, windowBus_65, windowBus_64, 
         windowBus_63, windowBus_62, windowBus_61, windowBus_60, windowBus_59, 
         windowBus_58, windowBus_57, windowBus_56, windowBus_55, windowBus_54, 
         windowBus_53, windowBus_52, windowBus_51, windowBus_50, windowBus_49, 
         windowBus_48, windowBus_47, windowBus_46, windowBus_45, windowBus_44, 
         windowBus_43, windowBus_42, windowBus_41, windowBus_40, windowBus_39, 
         windowBus_38, windowBus_37, windowBus_36, windowBus_35, windowBus_34, 
         windowBus_33, windowBus_32, windowBus_31, windowBus_30, windowBus_29, 
         windowBus_28, windowBus_27, windowBus_26, windowBus_25, windowBus_24, 
         windowBus_23, windowBus_22, windowBus_21, windowBus_20, windowBus_19, 
         windowBus_18, windowBus_17, windowBus_16, windowBus_15, windowBus_14, 
         windowBus_13, windowBus_12, windowBus_11, windowBus_10, windowBus_9, 
         windowBus_8, windowBus_7, windowBus_6, windowBus_5, windowBus_4, 
         windowBus_3, windowBus_2, windowBus_1, windowBus_0, writeBus_15, 
         writeBus_14, writeBus_13, writeBus_12, writeBus_11, writeBus_10, 
         writeBus_9, writeBus_8, writeBus_7, writeBus_6, writeBus_5, writeBus_4, 
         writeBus_3, writeBus_2, writeBus_1, writeBus_0, decoderRow_2, 
         decoderRow_1, decoderRow_0, writePage1, writePage2, writeFilter, 
         shift2To1, shift1To2, doneCores, startConv, dmaFilterFinish, 
         loadOneWord, loadTwoWord, readAllFinish, writeOneFinish, sumOutCores_15, 
         sumOutCores_14, sumOutCores_13, sumOutCores_12, sumOutCores_11, 
         sumOutCores_10, sumOutCores_9, sumOutCores_8, sumOutCores_7, 
         sumOutCores_6, sumOutCores_5, sumOutCores_4, sumOutCores_3, 
         sumOutCores_2, sumOutCores_1, sumOutCores_0, loadNetworkConfig, 
         loadFilterConfig, loadWindow, loadFilter, readNextCol, finishLayer, 
         finishSlice, inputSizeAddress_4, inputSizeAddress_3, inputSizeAddress_2, 
         inputSizeAddress_1, inputSizeAddress_0, outputSizeAddress_4, 
         outputSizeAddress_3, outputSizeAddress_2, outputSizeAddress_1, 
         outputSizeAddress_0, outputSizeAddressForDMA_12, 
         outputSizeAddressForDMA_11, outputSizeAddressForDMA_10, 
         outputSizeAddressForDMA_9, outputSizeAddressForDMA_8, 
         outputSizeAddressForDMA_7, outputSizeAddressForDMA_6, 
         outputSizeAddressForDMA_5, outputSizeAddressForDMA_4, 
         outputSizeAddressForDMA_3, outputSizeAddressForDMA_2, 
         outputSizeAddressForDMA_1, outputSizeAddressForDMA_0, 
         finishReadRowWindow, finishReadRowFilter, aluNumberWindow_2, 
         aluNumberWindow_1, aluNumberWindow_0, layersNumber_1, layersNumber_0, 
         filtersNumber_2, filtersNumber_1, filtersNumber_0, filterDepth_2, 
         filterDepth_1, filterDepth_0, outputBufferEn, saveToRAM, allRead, 
         currentRegFromOutBuffer_15, currentRegFromOutBuffer_14, 
         currentRegFromOutBuffer_13, currentRegFromOutBuffer_12, 
         currentRegFromOutBuffer_11, currentRegFromOutBuffer_10, 
         currentRegFromOutBuffer_9, currentRegFromOutBuffer_8, 
         currentRegFromOutBuffer_7, currentRegFromOutBuffer_6, 
         currentRegFromOutBuffer_5, currentRegFromOutBuffer_4, 
         currentRegFromOutBuffer_3, currentRegFromOutBuffer_2, 
         currentRegFromOutBuffer_1, currentRegFromOutBuffer_0, finalAdderOut_15, 
         finalAdderOut_14, finalAdderOut_13, finalAdderOut_12, finalAdderOut_11, 
         finalAdderOut_10, finalAdderOut_9, finalAdderOut_8, finalAdderOut_7, 
         finalAdderOut_6, finalAdderOut_5, finalAdderOut_4, finalAdderOut_3, 
         finalAdderOut_2, finalAdderOut_1, finalAdderOut_0, inputToFinalAdder_15, 
         inputToFinalAdder_14, inputToFinalAdder_13, inputToFinalAdder_12, 
         inputToFinalAdder_11, inputToFinalAdder_10, inputToFinalAdder_9, 
         inputToFinalAdder_8, inputToFinalAdder_7, inputToFinalAdder_6, 
         inputToFinalAdder_5, inputToFinalAdder_4, inputToFinalAdder_3, 
         inputToFinalAdder_2, inputToFinalAdder_1, inputToFinalAdder_0, 
         readNumLayers, readLayerConfig, finishFilter, baseAddressTwo_11, 
         inputSizeAddress_12, nx0, nx2, nx12, nx20, nx38, nx64, nx619, nx621, 
         nx624, nx626, nx628, nx638, nx645, nx647, nx649, nx651, nx653, nx655, 
         nx657, nx659, nx661, nx663, nx665, nx667, nx669;
    wire [6:0] \$dummy ;




    CNNCores_8_16_5_5_3 coresMap (.filterBus ({filterBus_39,filterBus_38,
                        filterBus_37,filterBus_36,filterBus_35,filterBus_34,
                        filterBus_33,filterBus_32,filterBus_31,filterBus_30,
                        filterBus_29,filterBus_28,filterBus_27,filterBus_26,
                        filterBus_25,filterBus_24,filterBus_23,filterBus_22,
                        filterBus_21,filterBus_20,filterBus_19,filterBus_18,
                        filterBus_17,filterBus_16,filterBus_15,filterBus_14,
                        filterBus_13,filterBus_12,filterBus_11,filterBus_10,
                        filterBus_9,filterBus_8,nx653,nx657,filterBus_5,
                        filterBus_4,filterBus_3,filterBus_2,filterBus_1,
                        filterBus_0}), .windowBus ({windowBus_79,windowBus_78,
                        windowBus_77,windowBus_76,windowBus_75,windowBus_74,
                        windowBus_73,windowBus_72,windowBus_71,windowBus_70,
                        windowBus_69,windowBus_68,windowBus_67,windowBus_66,
                        windowBus_65,windowBus_64,windowBus_63,windowBus_62,
                        windowBus_61,windowBus_60,windowBus_59,windowBus_58,
                        windowBus_57,windowBus_56,windowBus_55,windowBus_54,
                        windowBus_53,windowBus_52,windowBus_51,windowBus_50,
                        windowBus_49,windowBus_48,windowBus_47,windowBus_46,
                        windowBus_45,windowBus_44,windowBus_43,windowBus_42,
                        windowBus_41,windowBus_40,windowBus_39,windowBus_38,
                        windowBus_37,windowBus_36,windowBus_35,windowBus_34,
                        windowBus_33,windowBus_32,windowBus_31,windowBus_30,
                        windowBus_29,windowBus_28,windowBus_27,windowBus_26,
                        windowBus_25,windowBus_24,windowBus_23,windowBus_22,
                        windowBus_21,windowBus_20,windowBus_19,windowBus_18,
                        windowBus_17,windowBus_16,windowBus_15,windowBus_14,
                        windowBus_13,windowBus_12,windowBus_11,windowBus_10,
                        windowBus_9,windowBus_8,windowBus_7,windowBus_6,
                        windowBus_5,windowBus_4,windowBus_3,windowBus_2,
                        windowBus_1,windowBus_0}), .decoderRow ({decoderRow_2,
                        decoderRow_1,decoderRow_0}), .clk (clk), .rst (rst), .writePage1 (
                        nx661), .writePage2 (writePage2), .writeFilter (
                        writeFilter), .shift2To1 (shift2To1), .shift1To2 (
                        shift1To2), .pageTurn (currentPage_0), .start (startConv
                        ), .layerType (nx645), .filterType (nx649), .doneCores (
                        doneCores), .finalSumConv ({sumOutCores_15,
                        sumOutCores_14,sumOutCores_13,sumOutCores_12,
                        sumOutCores_11,sumOutCores_10,sumOutCores_9,
                        sumOutCores_8,sumOutCores_7,sumOutCores_6,sumOutCores_5,
                        sumOutCores_4,sumOutCores_3,sumOutCores_2,sumOutCores_1,
                        sumOutCores_0})) ;
    ControlUnit controlUnitMap (.clk (clk), .layersNumber ({layersNumber_1,
                layersNumber_0}), .filtersNumber ({filtersNumber_2,
                filtersNumber_1,filtersNumber_0}), .filterDepth ({filterDepth_2,
                filterDepth_1,filterDepth_0}), .filterOutputSize ({
                outputSizeAddress_4,outputSizeAddress_3,outputSizeAddress_2,
                outputSizeAddress_1,outputSizeAddress_0}), .startNetwork (
                startCNN), .layerType (nx645), .convFinish (doneCores), .dmaAFinish (
                dmaFilterFinish), .dmaBFinish (readAllFinish), .dmaCFinish (
                writeOneFinish), .resetNetwork (rst), .loadLayerConfig (
                loadTwoWord), .loadNetworkConfig (loadNetworkConfig), .loadFilterConfig (
                loadFilterConfig), .loadWindow (loadWindow), .loadFilter (
                loadFilter), .conv (conv), .pool (pool), .shift12 (shift1To2), .shift21 (
                shift2To1), .readNextCol (readNextCol), .addToOutputBuffer (
                \$dummy [0]), .outputBufferEn (outputBufferEn), .saveToRAM (
                saveToRAM), .currentPage ({currentPage_0}), .finishCurrentSlice (
                finishSlice), .finishFilter (finishFilter), .finishOneLayer (
                finishLayer), .finishNetwork (finishNetwork)) ;
    NBitAdder_13 outputSizeAddMap (.a ({inputSizeAddress_12,inputSizeAddress_12,
                 inputSizeAddress_12,inputSizeAddress_12,inputSizeAddress_12,
                 inputSizeAddress_12,inputSizeAddress_12,inputSizeAddress_12,
                 outputSizeAddress_4,outputSizeAddress_3,outputSizeAddress_2,
                 outputSizeAddress_1,outputSizeAddress_0}), .b ({
                 inputSizeAddress_12,inputSizeAddress_12,inputSizeAddress_12,
                 inputSizeAddress_12,inputSizeAddress_12,inputSizeAddress_12,
                 inputSizeAddress_12,inputSizeAddress_12,inputSizeAddress_12,
                 inputSizeAddress_12,inputSizeAddress_12,inputSizeAddress_12,
                 inputSizeAddress_12}), .carryIn (baseAddressTwo_11), .sum ({
                 outputSizeAddressForDMA_12,outputSizeAddressForDMA_11,
                 outputSizeAddressForDMA_10,outputSizeAddressForDMA_9,
                 outputSizeAddressForDMA_8,outputSizeAddressForDMA_7,
                 outputSizeAddressForDMA_6,outputSizeAddressForDMA_5,
                 outputSizeAddressForDMA_4,outputSizeAddressForDMA_3,
                 outputSizeAddressForDMA_2,outputSizeAddressForDMA_1,
                 outputSizeAddressForDMA_0}), .carryOut (\$dummy [1])) ;
    DMAController_12_13_8_16_5 DMAControllerMap (.clk (clk), .reset (rst), .weightsInternalBus (
                               {filterBus_39,filterBus_38,filterBus_37,
                               filterBus_36,filterBus_35,filterBus_34,
                               filterBus_33,filterBus_32,filterBus_31,
                               filterBus_30,filterBus_29,filterBus_28,
                               filterBus_27,filterBus_26,filterBus_25,
                               filterBus_24,filterBus_23,filterBus_22,
                               filterBus_21,filterBus_20,filterBus_19,
                               filterBus_18,filterBus_17,filterBus_16,
                               filterBus_15,filterBus_14,filterBus_13,
                               filterBus_12,filterBus_11,filterBus_10,
                               filterBus_9,filterBus_8,filterBus_7,filterBus_6,
                               filterBus_5,filterBus_4,filterBus_3,filterBus_2,
                               filterBus_1,filterBus_0}), .windowInternalBus ({
                               windowBus_79,windowBus_78,windowBus_77,
                               windowBus_76,windowBus_75,windowBus_74,
                               windowBus_73,windowBus_72,windowBus_71,
                               windowBus_70,windowBus_69,windowBus_68,
                               windowBus_67,windowBus_66,windowBus_65,
                               windowBus_64,windowBus_63,windowBus_62,
                               windowBus_61,windowBus_60,windowBus_59,
                               windowBus_58,windowBus_57,windowBus_56,
                               windowBus_55,windowBus_54,windowBus_53,
                               windowBus_52,windowBus_51,windowBus_50,
                               windowBus_49,windowBus_48,windowBus_47,
                               windowBus_46,windowBus_45,windowBus_44,
                               windowBus_43,windowBus_42,windowBus_41,
                               windowBus_40,windowBus_39,windowBus_38,
                               windowBus_37,windowBus_36,windowBus_35,
                               windowBus_34,windowBus_33,windowBus_32,
                               windowBus_31,windowBus_30,windowBus_29,
                               windowBus_28,windowBus_27,windowBus_26,
                               windowBus_25,windowBus_24,windowBus_23,
                               windowBus_22,windowBus_21,windowBus_20,
                               windowBus_19,windowBus_18,windowBus_17,
                               windowBus_16,windowBus_15,windowBus_14,
                               windowBus_13,windowBus_12,windowBus_11,
                               windowBus_10,windowBus_9,windowBus_8,windowBus_7,
                               windowBus_6,windowBus_5,windowBus_4,windowBus_3,
                               windowBus_2,windowBus_1,windowBus_0}), .writeInternalBus (
                               {writeBus_15,writeBus_14,writeBus_13,writeBus_12,
                               writeBus_11,writeBus_10,writeBus_9,writeBus_8,
                               writeBus_7,writeBus_6,writeBus_5,writeBus_4,
                               writeBus_3,writeBus_2,writeBus_1,writeBus_0}), .weightsRamAddress (
                               {weightsRamAddress[11],weightsRamAddress[10],
                               weightsRamAddress[9],weightsRamAddress[8],
                               weightsRamAddress[7],weightsRamAddress[6],
                               weightsRamAddress[5],weightsRamAddress[4],
                               weightsRamAddress[3],weightsRamAddress[2],
                               weightsRamAddress[1],weightsRamAddress[0]}), .windowRamAddressRead (
                               {windowRamAddressRead[12],
                               windowRamAddressRead[11],windowRamAddressRead[10]
                               ,windowRamAddressRead[9],windowRamAddressRead[8],
                               windowRamAddressRead[7],windowRamAddressRead[6],
                               windowRamAddressRead[5],windowRamAddressRead[4],
                               windowRamAddressRead[3],windowRamAddressRead[2],
                               windowRamAddressRead[1],windowRamAddressRead[0]})
                               , .windowRamAddressWrite ({
                               windowRamAddressWrite[12],
                               windowRamAddressWrite[11],
                               windowRamAddressWrite[10],
                               windowRamAddressWrite[9],windowRamAddressWrite[8]
                               ,windowRamAddressWrite[7],
                               windowRamAddressWrite[6],windowRamAddressWrite[5]
                               ,windowRamAddressWrite[4],
                               windowRamAddressWrite[3],windowRamAddressWrite[2]
                               ,windowRamAddressWrite[1],
                               windowRamAddressWrite[0]}), .weightsRamDataInBus (
                               {weightsRamDataInBus[39],weightsRamDataInBus[38],
                               weightsRamDataInBus[37],weightsRamDataInBus[36],
                               weightsRamDataInBus[35],weightsRamDataInBus[34],
                               weightsRamDataInBus[33],weightsRamDataInBus[32],
                               weightsRamDataInBus[31],weightsRamDataInBus[30],
                               weightsRamDataInBus[29],weightsRamDataInBus[28],
                               weightsRamDataInBus[27],weightsRamDataInBus[26],
                               weightsRamDataInBus[25],weightsRamDataInBus[24],
                               weightsRamDataInBus[23],weightsRamDataInBus[22],
                               weightsRamDataInBus[21],weightsRamDataInBus[20],
                               weightsRamDataInBus[19],weightsRamDataInBus[18],
                               weightsRamDataInBus[17],weightsRamDataInBus[16],
                               weightsRamDataInBus[15],weightsRamDataInBus[14],
                               weightsRamDataInBus[13],weightsRamDataInBus[12],
                               weightsRamDataInBus[11],weightsRamDataInBus[10],
                               weightsRamDataInBus[9],weightsRamDataInBus[8],
                               weightsRamDataInBus[7],weightsRamDataInBus[6],
                               weightsRamDataInBus[5],weightsRamDataInBus[4],
                               weightsRamDataInBus[3],weightsRamDataInBus[2],
                               weightsRamDataInBus[1],weightsRamDataInBus[0]}), 
                               .windowRamDataInBus ({windowRamDataInBus[79],
                               windowRamDataInBus[78],windowRamDataInBus[77],
                               windowRamDataInBus[76],windowRamDataInBus[75],
                               windowRamDataInBus[74],windowRamDataInBus[73],
                               windowRamDataInBus[72],windowRamDataInBus[71],
                               windowRamDataInBus[70],windowRamDataInBus[69],
                               windowRamDataInBus[68],windowRamDataInBus[67],
                               windowRamDataInBus[66],windowRamDataInBus[65],
                               windowRamDataInBus[64],windowRamDataInBus[63],
                               windowRamDataInBus[62],windowRamDataInBus[61],
                               windowRamDataInBus[60],windowRamDataInBus[59],
                               windowRamDataInBus[58],windowRamDataInBus[57],
                               windowRamDataInBus[56],windowRamDataInBus[55],
                               windowRamDataInBus[54],windowRamDataInBus[53],
                               windowRamDataInBus[52],windowRamDataInBus[51],
                               windowRamDataInBus[50],windowRamDataInBus[49],
                               windowRamDataInBus[48],windowRamDataInBus[47],
                               windowRamDataInBus[46],windowRamDataInBus[45],
                               windowRamDataInBus[44],windowRamDataInBus[43],
                               windowRamDataInBus[42],windowRamDataInBus[41],
                               windowRamDataInBus[40],windowRamDataInBus[39],
                               windowRamDataInBus[38],windowRamDataInBus[37],
                               windowRamDataInBus[36],windowRamDataInBus[35],
                               windowRamDataInBus[34],windowRamDataInBus[33],
                               windowRamDataInBus[32],windowRamDataInBus[31],
                               windowRamDataInBus[30],windowRamDataInBus[29],
                               windowRamDataInBus[28],windowRamDataInBus[27],
                               windowRamDataInBus[26],windowRamDataInBus[25],
                               windowRamDataInBus[24],windowRamDataInBus[23],
                               windowRamDataInBus[22],windowRamDataInBus[21],
                               windowRamDataInBus[20],windowRamDataInBus[19],
                               windowRamDataInBus[18],windowRamDataInBus[17],
                               windowRamDataInBus[16],windowRamDataInBus[15],
                               windowRamDataInBus[14],windowRamDataInBus[13],
                               windowRamDataInBus[12],windowRamDataInBus[11],
                               windowRamDataInBus[10],windowRamDataInBus[9],
                               windowRamDataInBus[8],windowRamDataInBus[7],
                               windowRamDataInBus[6],windowRamDataInBus[5],
                               windowRamDataInBus[4],windowRamDataInBus[3],
                               windowRamDataInBus[2],windowRamDataInBus[1],
                               windowRamDataInBus[0]}), .weightsRamRead (
                               weightsRamRead), .windowRamRead (windowRamRead), 
                               .windowRamWrite (windowRamWrite), .windowRamDataOutBus (
                               {windowRamDataOutBus[15],windowRamDataOutBus[14],
                               windowRamDataOutBus[13],windowRamDataOutBus[12],
                               windowRamDataOutBus[11],windowRamDataOutBus[10],
                               windowRamDataOutBus[9],windowRamDataOutBus[8],
                               windowRamDataOutBus[7],windowRamDataOutBus[6],
                               windowRamDataOutBus[5],windowRamDataOutBus[4],
                               windowRamDataOutBus[3],windowRamDataOutBus[2],
                               windowRamDataOutBus[1],windowRamDataOutBus[0]}), 
                               .MFCWindowRam (MFCWindowRam), .MFCWeightsRam (
                               MFCWeightsRam), .MFCWrite (MFCWrite), .loadNextFilter (
                               loadFilter), .loadNextWindow (nx663), .loadNextRow (
                               readNextCol), .loadOneWord (loadOneWord), .loadThreeWord (
                               loadTwoWord), .filterFinished (finishFilter), .sliceFinished (
                               finishSlice), .layerFinished (finishLayer), .layerType (
                               nx645), .write (saveToRAM), .weightsSizeType (
                               nx651), .inputSize ({inputSizeAddress_12,
                               inputSizeAddress_12,inputSizeAddress_12,
                               inputSizeAddress_12,inputSizeAddress_12,
                               inputSizeAddress_12,inputSizeAddress_12,
                               inputSizeAddress_12,inputSizeAddress_4,
                               inputSizeAddress_3,inputSizeAddress_2,
                               inputSizeAddress_1,inputSizeAddress_0}), .outputSize (
                               {outputSizeAddressForDMA_12,
                               outputSizeAddressForDMA_11,
                               outputSizeAddressForDMA_10,
                               outputSizeAddressForDMA_9,
                               outputSizeAddressForDMA_8,
                               outputSizeAddressForDMA_7,
                               outputSizeAddressForDMA_6,
                               outputSizeAddressForDMA_5,
                               outputSizeAddressForDMA_4,
                               outputSizeAddressForDMA_3,
                               outputSizeAddressForDMA_2,
                               outputSizeAddressForDMA_1,
                               outputSizeAddressForDMA_0}), .windowRamBaseAddress1 (
                               {inputSizeAddress_12,inputSizeAddress_12,
                               inputSizeAddress_12,inputSizeAddress_12,
                               inputSizeAddress_12,inputSizeAddress_12,
                               inputSizeAddress_12,inputSizeAddress_12,
                               inputSizeAddress_12,inputSizeAddress_12,
                               inputSizeAddress_12,inputSizeAddress_12,
                               inputSizeAddress_12}), .windowRamBaseAddress2 ({
                               inputSizeAddress_12,baseAddressTwo_11,
                               baseAddressTwo_11,baseAddressTwo_11,
                               baseAddressTwo_11,inputSizeAddress_12,
                               inputSizeAddress_12,baseAddressTwo_11,
                               inputSizeAddress_12,inputSizeAddress_12,
                               inputSizeAddress_12,inputSizeAddress_12,
                               inputSizeAddress_12}), .filterRamBaseAddress ({
                               inputSizeAddress_12,inputSizeAddress_12,
                               inputSizeAddress_12,inputSizeAddress_12,
                               inputSizeAddress_12,inputSizeAddress_12,
                               inputSizeAddress_12,inputSizeAddress_12,
                               inputSizeAddress_12,inputSizeAddress_12,
                               inputSizeAddress_12,inputSizeAddress_12}), .windowReadOne (
                               finishReadRowWindow), .windowReadFinal (
                               readAllFinish), .weightsReadOne (
                               finishReadRowFilter), .weightsReadFinal (
                               dmaFilterFinish), .writeDoneAll (\$dummy [2]), .writeDoneOne (
                               writeOneFinish), .filterAluNumber ({\$dummy [3],
                               \$dummy [4],\$dummy [5]}), .windowAluNumber ({
                               aluNumberWindow_2,aluNumberWindow_1,
                               aluNumberWindow_0})) ;
    OutputBuffer_40_484_16_8_9_6 outbufferMap (.sumInput ({finalAdderOut_15,
                                 finalAdderOut_14,finalAdderOut_13,
                                 finalAdderOut_12,finalAdderOut_11,
                                 finalAdderOut_10,finalAdderOut_9,
                                 finalAdderOut_8,finalAdderOut_7,finalAdderOut_6
                                 ,finalAdderOut_5,finalAdderOut_4,
                                 finalAdderOut_3,finalAdderOut_2,finalAdderOut_1
                                 ,finalAdderOut_0}), .weightsBus ({
                                 inputSizeAddress_12,inputSizeAddress_12,
                                 inputSizeAddress_12,inputSizeAddress_12,
                                 inputSizeAddress_12,inputSizeAddress_12,
                                 inputSizeAddress_12,inputSizeAddress_12,
                                 inputSizeAddress_12,inputSizeAddress_12,
                                 inputSizeAddress_12,inputSizeAddress_12,
                                 inputSizeAddress_12,inputSizeAddress_12,
                                 inputSizeAddress_12,inputSizeAddress_12,
                                 inputSizeAddress_12,inputSizeAddress_12,
                                 inputSizeAddress_12,inputSizeAddress_12,
                                 inputSizeAddress_12,inputSizeAddress_12,
                                 inputSizeAddress_12,inputSizeAddress_12,
                                 inputSizeAddress_12,inputSizeAddress_12,
                                 inputSizeAddress_12,inputSizeAddress_12,
                                 inputSizeAddress_12,inputSizeAddress_12,
                                 inputSizeAddress_12,inputSizeAddress_12,nx653,
                                 nx657,filterBus_5,filterBus_4,filterBus_3,
                                 filterBus_2,filterBus_1,filterBus_0}), .writeBus (
                                 {writeBus_15,writeBus_14,writeBus_13,
                                 writeBus_12,writeBus_11,writeBus_10,writeBus_9,
                                 writeBus_8,writeBus_7,writeBus_6,writeBus_5,
                                 writeBus_4,writeBus_3,writeBus_2,writeBus_1,
                                 writeBus_0}), .AllRead (allRead), .enableDecoder (
                                 nx667), .selectedRegisterMuxOutput ({
                                 currentRegFromOutBuffer_15,
                                 currentRegFromOutBuffer_14,
                                 currentRegFromOutBuffer_13,
                                 currentRegFromOutBuffer_12,
                                 currentRegFromOutBuffer_11,
                                 currentRegFromOutBuffer_10,
                                 currentRegFromOutBuffer_9,
                                 currentRegFromOutBuffer_8,
                                 currentRegFromOutBuffer_7,
                                 currentRegFromOutBuffer_6,
                                 currentRegFromOutBuffer_5,
                                 currentRegFromOutBuffer_4,
                                 currentRegFromOutBuffer_3,
                                 currentRegFromOutBuffer_2,
                                 currentRegFromOutBuffer_1,
                                 currentRegFromOutBuffer_0}), .clk (clk), .finishSlice (
                                 finishSlice), .resetRegisters (rst), .tristateEnable (
                                 saveToRAM), .counterEnable (nx669), .isPool (
                                 nx645)) ;
    Mux2_16 convOrPoolMuxMap (.A ({currentRegFromOutBuffer_15,
            currentRegFromOutBuffer_14,currentRegFromOutBuffer_13,
            currentRegFromOutBuffer_12,currentRegFromOutBuffer_11,
            currentRegFromOutBuffer_10,currentRegFromOutBuffer_9,
            currentRegFromOutBuffer_8,currentRegFromOutBuffer_7,
            currentRegFromOutBuffer_6,currentRegFromOutBuffer_5,
            currentRegFromOutBuffer_4,currentRegFromOutBuffer_3,
            currentRegFromOutBuffer_2,currentRegFromOutBuffer_1,
            currentRegFromOutBuffer_0}), .B ({inputSizeAddress_12,
            inputSizeAddress_12,inputSizeAddress_12,inputSizeAddress_12,
            inputSizeAddress_12,inputSizeAddress_12,inputSizeAddress_12,
            inputSizeAddress_12,inputSizeAddress_12,inputSizeAddress_12,
            inputSizeAddress_12,inputSizeAddress_12,inputSizeAddress_12,
            inputSizeAddress_12,inputSizeAddress_12,inputSizeAddress_12}), .S (
            nx645), .C ({inputToFinalAdder_15,inputToFinalAdder_14,
            inputToFinalAdder_13,inputToFinalAdder_12,inputToFinalAdder_11,
            inputToFinalAdder_10,inputToFinalAdder_9,inputToFinalAdder_8,
            inputToFinalAdder_7,inputToFinalAdder_6,inputToFinalAdder_5,
            inputToFinalAdder_4,inputToFinalAdder_3,inputToFinalAdder_2,
            inputToFinalAdder_1,inputToFinalAdder_0})) ;
    NBitAdder_16 finalAdderMap (.a ({inputToFinalAdder_15,inputToFinalAdder_14,
                 inputToFinalAdder_13,inputToFinalAdder_12,inputToFinalAdder_11,
                 inputToFinalAdder_10,inputToFinalAdder_9,inputToFinalAdder_8,
                 inputToFinalAdder_7,inputToFinalAdder_6,inputToFinalAdder_5,
                 inputToFinalAdder_4,inputToFinalAdder_3,inputToFinalAdder_2,
                 inputToFinalAdder_1,inputToFinalAdder_0}), .b ({sumOutCores_15,
                 sumOutCores_14,sumOutCores_13,sumOutCores_12,sumOutCores_11,
                 sumOutCores_10,sumOutCores_9,sumOutCores_8,sumOutCores_7,
                 sumOutCores_6,sumOutCores_5,sumOutCores_4,sumOutCores_3,
                 sumOutCores_2,sumOutCores_1,sumOutCores_0}), .carryIn (
                 inputSizeAddress_12), .sum ({finalAdderOut_15,finalAdderOut_14,
                 finalAdderOut_13,finalAdderOut_12,finalAdderOut_11,
                 finalAdderOut_10,finalAdderOut_9,finalAdderOut_8,
                 finalAdderOut_7,finalAdderOut_6,finalAdderOut_5,finalAdderOut_4
                 ,finalAdderOut_3,finalAdderOut_2,finalAdderOut_1,
                 finalAdderOut_0}), .carryOut (\$dummy [6])) ;
    Config_40 configMap (.filterBus ({inputSizeAddress_12,inputSizeAddress_12,
              inputSizeAddress_12,inputSizeAddress_12,inputSizeAddress_12,
              inputSizeAddress_12,inputSizeAddress_12,inputSizeAddress_12,
              inputSizeAddress_12,inputSizeAddress_12,inputSizeAddress_12,
              inputSizeAddress_12,inputSizeAddress_12,inputSizeAddress_12,
              inputSizeAddress_12,inputSizeAddress_12,filterBus_23,filterBus_22,
              filterBus_21,filterBus_20,filterBus_19,inputSizeAddress_12,
              inputSizeAddress_12,inputSizeAddress_12,filterBus_15,filterBus_14,
              filterBus_13,filterBus_12,filterBus_11,inputSizeAddress_12,
              inputSizeAddress_12,inputSizeAddress_12,nx655,nx659,filterBus_5,
              filterBus_4,filterBus_3,filterBus_2,filterBus_1,filterBus_0}), .clk (
              clk), .rst (rst), .readNumLayers (readNumLayers), .readLayerConfig (
              readLayerConfig), .numLayers ({layersNumber_1,layersNumber_0}), .layerType (
              layerType), .filterType (filterType), .numFilters ({
              filtersNumber_2,filtersNumber_1,filtersNumber_0}), .filterDepth ({
              filterDepth_2,filterDepth_1,filterDepth_0}), .inputSize ({
              inputSizeAddress_4,inputSizeAddress_3,inputSizeAddress_2,
              inputSizeAddress_1,inputSizeAddress_0}), .outputSize ({
              outputSizeAddress_4,outputSizeAddress_3,outputSizeAddress_2,
              outputSizeAddress_1,outputSizeAddress_0})) ;
    fake_gnd ix588 (.Y (inputSizeAddress_12)) ;
    fake_vcc ix586 (.Y (baseAddressTwo_11)) ;
    and02 ix47 (.Y (readLayerConfig), .A0 (loadTwoWord), .A1 (
          finishReadRowFilter)) ;
    and02 ix49 (.Y (readNumLayers), .A0 (loadNetworkConfig), .A1 (
          finishReadRowFilter)) ;
    and02 ix51 (.Y (allRead), .A0 (dmaFilterFinish), .A1 (loadFilterConfig)) ;
    or02 ix53 (.Y (loadOneWord), .A0 (loadNetworkConfig), .A1 (loadFilterConfig)
         ) ;
    or02 ix79 (.Y (startConv), .A0 (conv), .A1 (pool)) ;
    and02 ix55 (.Y (writeFilter), .A0 (finishReadRowFilter), .A1 (loadFilter)) ;
    and02 ix67 (.Y (writePage2), .A0 (finishReadRowWindow), .A1 (nx64)) ;
    oai21 ix65 (.Y (nx64), .A0 (currentPage_0), .A1 (nx619), .B0 (nx621)) ;
    nor02_2x ix620 (.Y (nx619), .A0 (nx663), .A1 (readNextCol)) ;
    oai21 ix622 (.Y (nx621), .A0 (loadFilter), .A1 (nx645), .B0 (nx663)) ;
    aoi21 ix77 (.Y (writePage1), .A0 (nx624), .A1 (nx626), .B0 (nx628)) ;
    oai21 ix625 (.Y (nx624), .A0 (nx665), .A1 (readNextCol), .B0 (currentPage_0)
          ) ;
    oai21 ix627 (.Y (nx626), .A0 (loadFilter), .A1 (nx647), .B0 (nx665)) ;
    inv01 ix629 (.Y (nx628), .A (finishReadRowWindow)) ;
    latch lat_decoderRow_0 (.Q (decoderRow_0), .D (nx2), .CLK (nx0)) ;
    and02 ix3 (.Y (nx2), .A0 (aluNumberWindow_0), .A1 (nx665)) ;
    latch lat_decoderRow_1 (.Q (decoderRow_1), .D (nx20), .CLK (nx0)) ;
    mux21_ni ix21 (.Y (nx20), .A0 (nx12), .A1 (aluNumberWindow_1), .S0 (nx665)
             ) ;
    nor02ii ix13 (.Y (nx12), .A0 (nx649), .A1 (readNextCol)) ;
    latch lat_decoderRow_2 (.Q (decoderRow_2), .D (nx38), .CLK (nx0)) ;
    oai21 ix39 (.Y (nx38), .A0 (nx665), .A1 (readNextCol), .B0 (nx638)) ;
    mux21 ix639 (.Y (nx638), .A0 (nx649), .A1 (aluNumberWindow_2), .S0 (nx665)
          ) ;
    inv01 ix1 (.Y (nx0), .A (nx619)) ;
    buf02 ix644 (.Y (nx645), .A (layerType)) ;
    buf02 ix646 (.Y (nx647), .A (layerType)) ;
    buf02 ix648 (.Y (nx649), .A (filterType)) ;
    buf02 ix650 (.Y (nx651), .A (filterType)) ;
    buf02 ix652 (.Y (nx653), .A (filterBus_7)) ;
    buf02 ix654 (.Y (nx655), .A (filterBus_7)) ;
    buf02 ix656 (.Y (nx657), .A (filterBus_6)) ;
    buf02 ix658 (.Y (nx659), .A (filterBus_6)) ;
    buf02 ix660 (.Y (nx661), .A (writePage1)) ;
    buf02 ix662 (.Y (nx663), .A (loadWindow)) ;
    buf02 ix664 (.Y (nx665), .A (loadWindow)) ;
    buf02 ix666 (.Y (nx667), .A (outputBufferEn)) ;
    buf02 ix668 (.Y (nx669), .A (outputBufferEn)) ;
endmodule


module Config_40 ( filterBus, clk, rst, readNumLayers, readLayerConfig, 
                   numLayers, layerType, filterType, numFilters, filterDepth, 
                   inputSize, outputSize ) ;

    input [39:0]filterBus ;
    input clk ;
    input rst ;
    input readNumLayers ;
    input readLayerConfig ;
    output [1:0]numLayers ;
    output layerType ;
    output filterType ;
    output [2:0]numFilters ;
    output [2:0]filterDepth ;
    output [4:0]inputSize ;
    output [4:0]outputSize ;

    wire nx90, nx92;



    Reg_2 numLayerRegMap (.D ({filterBus[7],filterBus[6]}), .en (readNumLayers)
          , .clk (clk), .rst (rst), .Q ({numLayers[1],numLayers[0]})) ;
    Reg_3 numFiltersRegMap (.D ({filterBus[5],filterBus[4],filterBus[3]}), .en (
          nx90), .clk (clk), .rst (rst), .Q ({numFilters[2],numFilters[1],
          numFilters[0]})) ;
    Reg_3 filterDepthRegMap (.D ({filterBus[2],filterBus[1],filterBus[0]}), .en (
          nx90), .clk (clk), .rst (rst), .Q ({filterDepth[2],filterDepth[1],
          filterDepth[0]})) ;
    Reg_2 layerTypeRegMap (.D ({filterBus[7],filterBus[6]}), .en (nx92), .clk (
          clk), .rst (rst), .Q ({layerType,filterType})) ;
    Reg_5 inputSizeRegMap (.D ({filterBus[15],filterBus[14],filterBus[13],
          filterBus[12],filterBus[11]}), .en (nx90), .clk (clk), .rst (rst), .Q (
          {inputSize[4],inputSize[3],inputSize[2],inputSize[1],inputSize[0]})) ;
    Reg_5 outputSizeRegMap (.D ({filterBus[23],filterBus[22],filterBus[21],
          filterBus[20],filterBus[19]}), .en (nx92), .clk (clk), .rst (rst), .Q (
          {outputSize[4],outputSize[3],outputSize[2],outputSize[1],outputSize[0]
          })) ;
    buf02 ix89 (.Y (nx90), .A (readLayerConfig)) ;
    buf02 ix91 (.Y (nx92), .A (readLayerConfig)) ;
endmodule


module OutputBuffer_40_484_16_8_9_6 ( sumInput, weightsBus, writeBus, AllRead, 
                                      enableDecoder, selectedRegisterMuxOutput, 
                                      clk, finishSlice, resetRegisters, 
                                      tristateEnable, counterEnable, isPool ) ;

    input [15:0]sumInput ;
    input [39:0]weightsBus ;
    output [15:0]writeBus ;
    input AllRead ;
    input enableDecoder ;
    output [15:0]selectedRegisterMuxOutput ;
    input clk ;
    input finishSlice ;
    input resetRegisters ;
    input tristateEnable ;
    input counterEnable ;
    input isPool ;

    wire decoderOutput_483, decoderOutput_482, decoderOutput_481, 
         decoderOutput_480, decoderOutput_479, decoderOutput_478, 
         decoderOutput_477, decoderOutput_476, decoderOutput_475, 
         decoderOutput_474, decoderOutput_473, decoderOutput_472, 
         decoderOutput_471, decoderOutput_470, decoderOutput_469, 
         decoderOutput_468, decoderOutput_467, decoderOutput_466, 
         decoderOutput_465, decoderOutput_464, decoderOutput_463, 
         decoderOutput_462, decoderOutput_461, decoderOutput_460, 
         decoderOutput_459, decoderOutput_458, decoderOutput_457, 
         decoderOutput_456, decoderOutput_455, decoderOutput_454, 
         decoderOutput_453, decoderOutput_452, decoderOutput_451, 
         decoderOutput_450, decoderOutput_449, decoderOutput_448, 
         decoderOutput_447, decoderOutput_446, decoderOutput_445, 
         decoderOutput_444, decoderOutput_443, decoderOutput_442, 
         decoderOutput_441, decoderOutput_440, decoderOutput_439, 
         decoderOutput_438, decoderOutput_437, decoderOutput_436, 
         decoderOutput_435, decoderOutput_434, decoderOutput_433, 
         decoderOutput_432, decoderOutput_431, decoderOutput_430, 
         decoderOutput_429, decoderOutput_428, decoderOutput_427, 
         decoderOutput_426, decoderOutput_425, decoderOutput_424, 
         decoderOutput_423, decoderOutput_422, decoderOutput_421, 
         decoderOutput_420, decoderOutput_419, decoderOutput_418, 
         decoderOutput_417, decoderOutput_416, decoderOutput_415, 
         decoderOutput_414, decoderOutput_413, decoderOutput_412, 
         decoderOutput_411, decoderOutput_410, decoderOutput_409, 
         decoderOutput_408, decoderOutput_407, decoderOutput_406, 
         decoderOutput_405, decoderOutput_404, decoderOutput_403, 
         decoderOutput_402, decoderOutput_401, decoderOutput_400, 
         decoderOutput_399, decoderOutput_398, decoderOutput_397, 
         decoderOutput_396, decoderOutput_395, decoderOutput_394, 
         decoderOutput_393, decoderOutput_392, decoderOutput_391, 
         decoderOutput_390, decoderOutput_389, decoderOutput_388, 
         decoderOutput_387, decoderOutput_386, decoderOutput_385, 
         decoderOutput_384, decoderOutput_383, decoderOutput_382, 
         decoderOutput_381, decoderOutput_380, decoderOutput_379, 
         decoderOutput_378, decoderOutput_377, decoderOutput_376, 
         decoderOutput_375, decoderOutput_374, decoderOutput_373, 
         decoderOutput_372, decoderOutput_371, decoderOutput_370, 
         decoderOutput_369, decoderOutput_368, decoderOutput_367, 
         decoderOutput_366, decoderOutput_365, decoderOutput_364, 
         decoderOutput_363, decoderOutput_362, decoderOutput_361, 
         decoderOutput_360, decoderOutput_359, decoderOutput_358, 
         decoderOutput_357, decoderOutput_356, decoderOutput_355, 
         decoderOutput_354, decoderOutput_353, decoderOutput_352, 
         decoderOutput_351, decoderOutput_350, decoderOutput_349, 
         decoderOutput_348, decoderOutput_347, decoderOutput_346, 
         decoderOutput_345, decoderOutput_344, decoderOutput_343, 
         decoderOutput_342, decoderOutput_341, decoderOutput_340, 
         decoderOutput_339, decoderOutput_338, decoderOutput_337, 
         decoderOutput_336, decoderOutput_335, decoderOutput_334, 
         decoderOutput_333, decoderOutput_332, decoderOutput_331, 
         decoderOutput_330, decoderOutput_329, decoderOutput_328, 
         decoderOutput_327, decoderOutput_326, decoderOutput_325, 
         decoderOutput_324, decoderOutput_323, decoderOutput_322, 
         decoderOutput_321, decoderOutput_320, decoderOutput_319, 
         decoderOutput_318, decoderOutput_317, decoderOutput_316, 
         decoderOutput_315, decoderOutput_314, decoderOutput_313, 
         decoderOutput_312, decoderOutput_311, decoderOutput_310, 
         decoderOutput_309, decoderOutput_308, decoderOutput_307, 
         decoderOutput_306, decoderOutput_305, decoderOutput_304, 
         decoderOutput_303, decoderOutput_302, decoderOutput_301, 
         decoderOutput_300, decoderOutput_299, decoderOutput_298, 
         decoderOutput_297, decoderOutput_296, decoderOutput_295, 
         decoderOutput_294, decoderOutput_293, decoderOutput_292, 
         decoderOutput_291, decoderOutput_290, decoderOutput_289, 
         decoderOutput_288, decoderOutput_287, decoderOutput_286, 
         decoderOutput_285, decoderOutput_284, decoderOutput_283, 
         decoderOutput_282, decoderOutput_281, decoderOutput_280, 
         decoderOutput_279, decoderOutput_278, decoderOutput_277, 
         decoderOutput_276, decoderOutput_275, decoderOutput_274, 
         decoderOutput_273, decoderOutput_272, decoderOutput_271, 
         decoderOutput_270, decoderOutput_269, decoderOutput_268, 
         decoderOutput_267, decoderOutput_266, decoderOutput_265, 
         decoderOutput_264, decoderOutput_263, decoderOutput_262, 
         decoderOutput_261, decoderOutput_260, decoderOutput_259, 
         decoderOutput_258, decoderOutput_257, decoderOutput_256, 
         decoderOutput_255, decoderOutput_254, decoderOutput_253, 
         decoderOutput_252, decoderOutput_251, decoderOutput_250, 
         decoderOutput_249, decoderOutput_248, decoderOutput_247, 
         decoderOutput_246, decoderOutput_245, decoderOutput_244, 
         decoderOutput_243, decoderOutput_242, decoderOutput_241, 
         decoderOutput_240, decoderOutput_239, decoderOutput_238, 
         decoderOutput_237, decoderOutput_236, decoderOutput_235, 
         decoderOutput_234, decoderOutput_233, decoderOutput_232, 
         decoderOutput_231, decoderOutput_230, decoderOutput_229, 
         decoderOutput_228, decoderOutput_227, decoderOutput_226, 
         decoderOutput_225, decoderOutput_224, decoderOutput_223, 
         decoderOutput_222, decoderOutput_221, decoderOutput_220, 
         decoderOutput_219, decoderOutput_218, decoderOutput_217, 
         decoderOutput_216, decoderOutput_215, decoderOutput_214, 
         decoderOutput_213, decoderOutput_212, decoderOutput_211, 
         decoderOutput_210, decoderOutput_209, decoderOutput_208, 
         decoderOutput_207, decoderOutput_206, decoderOutput_205, 
         decoderOutput_204, decoderOutput_203, decoderOutput_202, 
         decoderOutput_201, decoderOutput_200, decoderOutput_199, 
         decoderOutput_198, decoderOutput_197, decoderOutput_196, 
         decoderOutput_195, decoderOutput_194, decoderOutput_193, 
         decoderOutput_192, decoderOutput_191, decoderOutput_190, 
         decoderOutput_189, decoderOutput_188, decoderOutput_187, 
         decoderOutput_186, decoderOutput_185, decoderOutput_184, 
         decoderOutput_183, decoderOutput_182, decoderOutput_181, 
         decoderOutput_180, decoderOutput_179, decoderOutput_178, 
         decoderOutput_177, decoderOutput_176, decoderOutput_175, 
         decoderOutput_174, decoderOutput_173, decoderOutput_172, 
         decoderOutput_171, decoderOutput_170, decoderOutput_169, 
         decoderOutput_168, decoderOutput_167, decoderOutput_166, 
         decoderOutput_165, decoderOutput_164, decoderOutput_163, 
         decoderOutput_162, decoderOutput_161, decoderOutput_160, 
         decoderOutput_159, decoderOutput_158, decoderOutput_157, 
         decoderOutput_156, decoderOutput_155, decoderOutput_154, 
         decoderOutput_153, decoderOutput_152, decoderOutput_151, 
         decoderOutput_150, decoderOutput_149, decoderOutput_148, 
         decoderOutput_147, decoderOutput_146, decoderOutput_145, 
         decoderOutput_144, decoderOutput_143, decoderOutput_142, 
         decoderOutput_141, decoderOutput_140, decoderOutput_139, 
         decoderOutput_138, decoderOutput_137, decoderOutput_136, 
         decoderOutput_135, decoderOutput_134, decoderOutput_133, 
         decoderOutput_132, decoderOutput_131, decoderOutput_130, 
         decoderOutput_129, decoderOutput_128, decoderOutput_127, 
         decoderOutput_126, decoderOutput_125, decoderOutput_124, 
         decoderOutput_123, decoderOutput_122, decoderOutput_121, 
         decoderOutput_120, decoderOutput_119, decoderOutput_118, 
         decoderOutput_117, decoderOutput_116, decoderOutput_115, 
         decoderOutput_114, decoderOutput_113, decoderOutput_112, 
         decoderOutput_111, decoderOutput_110, decoderOutput_109, 
         decoderOutput_108, decoderOutput_107, decoderOutput_106, 
         decoderOutput_105, decoderOutput_104, decoderOutput_103, 
         decoderOutput_102, decoderOutput_101, decoderOutput_100, 
         decoderOutput_99, decoderOutput_98, decoderOutput_97, decoderOutput_96, 
         decoderOutput_95, decoderOutput_94, decoderOutput_93, decoderOutput_92, 
         decoderOutput_91, decoderOutput_90, decoderOutput_89, decoderOutput_88, 
         decoderOutput_87, decoderOutput_86, decoderOutput_85, decoderOutput_84, 
         decoderOutput_83, decoderOutput_82, decoderOutput_81, decoderOutput_80, 
         decoderOutput_79, decoderOutput_78, decoderOutput_77, decoderOutput_76, 
         decoderOutput_75, decoderOutput_74, decoderOutput_73, decoderOutput_72, 
         decoderOutput_71, decoderOutput_70, decoderOutput_69, decoderOutput_68, 
         decoderOutput_67, decoderOutput_66, decoderOutput_65, decoderOutput_64, 
         decoderOutput_63, decoderOutput_62, decoderOutput_61, decoderOutput_60, 
         decoderOutput_59, decoderOutput_58, decoderOutput_57, decoderOutput_56, 
         decoderOutput_55, decoderOutput_54, decoderOutput_53, decoderOutput_52, 
         decoderOutput_51, decoderOutput_50, decoderOutput_49, decoderOutput_48, 
         decoderOutput_47, decoderOutput_46, decoderOutput_45, decoderOutput_44, 
         decoderOutput_43, decoderOutput_42, decoderOutput_41, decoderOutput_40, 
         decoderOutput_39, decoderOutput_38, decoderOutput_37, decoderOutput_36, 
         decoderOutput_35, decoderOutput_34, decoderOutput_33, decoderOutput_32, 
         decoderOutput_31, decoderOutput_30, decoderOutput_29, decoderOutput_28, 
         decoderOutput_27, decoderOutput_26, decoderOutput_25, decoderOutput_24, 
         decoderOutput_23, decoderOutput_22, decoderOutput_21, decoderOutput_20, 
         decoderOutput_19, decoderOutput_18, decoderOutput_17, decoderOutput_16, 
         decoderOutput_15, decoderOutput_14, decoderOutput_13, decoderOutput_12, 
         decoderOutput_11, decoderOutput_10, decoderOutput_9, decoderOutput_8, 
         decoderOutput_7, decoderOutput_6, decoderOutput_5, decoderOutput_4, 
         decoderOutput_3, decoderOutput_2, decoderOutput_1, decoderOutput_0, 
         registerOutputs_0__15, registerOutputs_0__14, registerOutputs_0__13, 
         registerOutputs_0__12, registerOutputs_0__11, registerOutputs_0__10, 
         registerOutputs_0__9, registerOutputs_0__8, registerOutputs_0__7, 
         registerOutputs_0__6, registerOutputs_0__5, registerOutputs_0__4, 
         registerOutputs_0__3, registerOutputs_0__2, registerOutputs_0__1, 
         registerOutputs_0__0, registerOutputs_1__15, registerOutputs_1__14, 
         registerOutputs_1__13, registerOutputs_1__12, registerOutputs_1__11, 
         registerOutputs_1__10, registerOutputs_1__9, registerOutputs_1__8, 
         registerOutputs_1__7, registerOutputs_1__6, registerOutputs_1__5, 
         registerOutputs_1__4, registerOutputs_1__3, registerOutputs_1__2, 
         registerOutputs_1__1, registerOutputs_1__0, registerOutputs_2__15, 
         registerOutputs_2__14, registerOutputs_2__13, registerOutputs_2__12, 
         registerOutputs_2__11, registerOutputs_2__10, registerOutputs_2__9, 
         registerOutputs_2__8, registerOutputs_2__7, registerOutputs_2__6, 
         registerOutputs_2__5, registerOutputs_2__4, registerOutputs_2__3, 
         registerOutputs_2__2, registerOutputs_2__1, registerOutputs_2__0, 
         registerOutputs_3__15, registerOutputs_3__14, registerOutputs_3__13, 
         registerOutputs_3__12, registerOutputs_3__11, registerOutputs_3__10, 
         registerOutputs_3__9, registerOutputs_3__8, registerOutputs_3__7, 
         registerOutputs_3__6, registerOutputs_3__5, registerOutputs_3__4, 
         registerOutputs_3__3, registerOutputs_3__2, registerOutputs_3__1, 
         registerOutputs_3__0, registerOutputs_4__15, registerOutputs_4__14, 
         registerOutputs_4__13, registerOutputs_4__12, registerOutputs_4__11, 
         registerOutputs_4__10, registerOutputs_4__9, registerOutputs_4__8, 
         registerOutputs_4__7, registerOutputs_4__6, registerOutputs_4__5, 
         registerOutputs_4__4, registerOutputs_4__3, registerOutputs_4__2, 
         registerOutputs_4__1, registerOutputs_4__0, registerOutputs_5__15, 
         registerOutputs_5__14, registerOutputs_5__13, registerOutputs_5__12, 
         registerOutputs_5__11, registerOutputs_5__10, registerOutputs_5__9, 
         registerOutputs_5__8, registerOutputs_5__7, registerOutputs_5__6, 
         registerOutputs_5__5, registerOutputs_5__4, registerOutputs_5__3, 
         registerOutputs_5__2, registerOutputs_5__1, registerOutputs_5__0, 
         registerOutputs_6__15, registerOutputs_6__14, registerOutputs_6__13, 
         registerOutputs_6__12, registerOutputs_6__11, registerOutputs_6__10, 
         registerOutputs_6__9, registerOutputs_6__8, registerOutputs_6__7, 
         registerOutputs_6__6, registerOutputs_6__5, registerOutputs_6__4, 
         registerOutputs_6__3, registerOutputs_6__2, registerOutputs_6__1, 
         registerOutputs_6__0, registerOutputs_7__15, registerOutputs_7__14, 
         registerOutputs_7__13, registerOutputs_7__12, registerOutputs_7__11, 
         registerOutputs_7__10, registerOutputs_7__9, registerOutputs_7__8, 
         registerOutputs_7__7, registerOutputs_7__6, registerOutputs_7__5, 
         registerOutputs_7__4, registerOutputs_7__3, registerOutputs_7__2, 
         registerOutputs_7__1, registerOutputs_7__0, registerOutputs_8__15, 
         registerOutputs_8__14, registerOutputs_8__13, registerOutputs_8__12, 
         registerOutputs_8__11, registerOutputs_8__10, registerOutputs_8__9, 
         registerOutputs_8__8, registerOutputs_8__7, registerOutputs_8__6, 
         registerOutputs_8__5, registerOutputs_8__4, registerOutputs_8__3, 
         registerOutputs_8__2, registerOutputs_8__1, registerOutputs_8__0, 
         registerOutputs_9__15, registerOutputs_9__14, registerOutputs_9__13, 
         registerOutputs_9__12, registerOutputs_9__11, registerOutputs_9__10, 
         registerOutputs_9__9, registerOutputs_9__8, registerOutputs_9__7, 
         registerOutputs_9__6, registerOutputs_9__5, registerOutputs_9__4, 
         registerOutputs_9__3, registerOutputs_9__2, registerOutputs_9__1, 
         registerOutputs_9__0, registerOutputs_10__15, registerOutputs_10__14, 
         registerOutputs_10__13, registerOutputs_10__12, registerOutputs_10__11, 
         registerOutputs_10__10, registerOutputs_10__9, registerOutputs_10__8, 
         registerOutputs_10__7, registerOutputs_10__6, registerOutputs_10__5, 
         registerOutputs_10__4, registerOutputs_10__3, registerOutputs_10__2, 
         registerOutputs_10__1, registerOutputs_10__0, registerOutputs_11__15, 
         registerOutputs_11__14, registerOutputs_11__13, registerOutputs_11__12, 
         registerOutputs_11__11, registerOutputs_11__10, registerOutputs_11__9, 
         registerOutputs_11__8, registerOutputs_11__7, registerOutputs_11__6, 
         registerOutputs_11__5, registerOutputs_11__4, registerOutputs_11__3, 
         registerOutputs_11__2, registerOutputs_11__1, registerOutputs_11__0, 
         registerOutputs_12__15, registerOutputs_12__14, registerOutputs_12__13, 
         registerOutputs_12__12, registerOutputs_12__11, registerOutputs_12__10, 
         registerOutputs_12__9, registerOutputs_12__8, registerOutputs_12__7, 
         registerOutputs_12__6, registerOutputs_12__5, registerOutputs_12__4, 
         registerOutputs_12__3, registerOutputs_12__2, registerOutputs_12__1, 
         registerOutputs_12__0, registerOutputs_13__15, registerOutputs_13__14, 
         registerOutputs_13__13, registerOutputs_13__12, registerOutputs_13__11, 
         registerOutputs_13__10, registerOutputs_13__9, registerOutputs_13__8, 
         registerOutputs_13__7, registerOutputs_13__6, registerOutputs_13__5, 
         registerOutputs_13__4, registerOutputs_13__3, registerOutputs_13__2, 
         registerOutputs_13__1, registerOutputs_13__0, registerOutputs_14__15, 
         registerOutputs_14__14, registerOutputs_14__13, registerOutputs_14__12, 
         registerOutputs_14__11, registerOutputs_14__10, registerOutputs_14__9, 
         registerOutputs_14__8, registerOutputs_14__7, registerOutputs_14__6, 
         registerOutputs_14__5, registerOutputs_14__4, registerOutputs_14__3, 
         registerOutputs_14__2, registerOutputs_14__1, registerOutputs_14__0, 
         registerOutputs_15__15, registerOutputs_15__14, registerOutputs_15__13, 
         registerOutputs_15__12, registerOutputs_15__11, registerOutputs_15__10, 
         registerOutputs_15__9, registerOutputs_15__8, registerOutputs_15__7, 
         registerOutputs_15__6, registerOutputs_15__5, registerOutputs_15__4, 
         registerOutputs_15__3, registerOutputs_15__2, registerOutputs_15__1, 
         registerOutputs_15__0, registerOutputs_16__15, registerOutputs_16__14, 
         registerOutputs_16__13, registerOutputs_16__12, registerOutputs_16__11, 
         registerOutputs_16__10, registerOutputs_16__9, registerOutputs_16__8, 
         registerOutputs_16__7, registerOutputs_16__6, registerOutputs_16__5, 
         registerOutputs_16__4, registerOutputs_16__3, registerOutputs_16__2, 
         registerOutputs_16__1, registerOutputs_16__0, registerOutputs_17__15, 
         registerOutputs_17__14, registerOutputs_17__13, registerOutputs_17__12, 
         registerOutputs_17__11, registerOutputs_17__10, registerOutputs_17__9, 
         registerOutputs_17__8, registerOutputs_17__7, registerOutputs_17__6, 
         registerOutputs_17__5, registerOutputs_17__4, registerOutputs_17__3, 
         registerOutputs_17__2, registerOutputs_17__1, registerOutputs_17__0, 
         registerOutputs_18__15, registerOutputs_18__14, registerOutputs_18__13, 
         registerOutputs_18__12, registerOutputs_18__11, registerOutputs_18__10, 
         registerOutputs_18__9, registerOutputs_18__8, registerOutputs_18__7, 
         registerOutputs_18__6, registerOutputs_18__5, registerOutputs_18__4, 
         registerOutputs_18__3, registerOutputs_18__2, registerOutputs_18__1, 
         registerOutputs_18__0, registerOutputs_19__15, registerOutputs_19__14, 
         registerOutputs_19__13, registerOutputs_19__12, registerOutputs_19__11, 
         registerOutputs_19__10, registerOutputs_19__9, registerOutputs_19__8, 
         registerOutputs_19__7, registerOutputs_19__6, registerOutputs_19__5, 
         registerOutputs_19__4, registerOutputs_19__3, registerOutputs_19__2, 
         registerOutputs_19__1, registerOutputs_19__0, registerOutputs_20__15, 
         registerOutputs_20__14, registerOutputs_20__13, registerOutputs_20__12, 
         registerOutputs_20__11, registerOutputs_20__10, registerOutputs_20__9, 
         registerOutputs_20__8, registerOutputs_20__7, registerOutputs_20__6, 
         registerOutputs_20__5, registerOutputs_20__4, registerOutputs_20__3, 
         registerOutputs_20__2, registerOutputs_20__1, registerOutputs_20__0, 
         registerOutputs_21__15, registerOutputs_21__14, registerOutputs_21__13, 
         registerOutputs_21__12, registerOutputs_21__11, registerOutputs_21__10, 
         registerOutputs_21__9, registerOutputs_21__8, registerOutputs_21__7, 
         registerOutputs_21__6, registerOutputs_21__5, registerOutputs_21__4, 
         registerOutputs_21__3, registerOutputs_21__2, registerOutputs_21__1, 
         registerOutputs_21__0, registerOutputs_22__15, registerOutputs_22__14, 
         registerOutputs_22__13, registerOutputs_22__12, registerOutputs_22__11, 
         registerOutputs_22__10, registerOutputs_22__9, registerOutputs_22__8, 
         registerOutputs_22__7, registerOutputs_22__6, registerOutputs_22__5, 
         registerOutputs_22__4, registerOutputs_22__3, registerOutputs_22__2, 
         registerOutputs_22__1, registerOutputs_22__0, registerOutputs_23__15, 
         registerOutputs_23__14, registerOutputs_23__13, registerOutputs_23__12, 
         registerOutputs_23__11, registerOutputs_23__10, registerOutputs_23__9, 
         registerOutputs_23__8, registerOutputs_23__7, registerOutputs_23__6, 
         registerOutputs_23__5, registerOutputs_23__4, registerOutputs_23__3, 
         registerOutputs_23__2, registerOutputs_23__1, registerOutputs_23__0, 
         registerOutputs_24__15, registerOutputs_24__14, registerOutputs_24__13, 
         registerOutputs_24__12, registerOutputs_24__11, registerOutputs_24__10, 
         registerOutputs_24__9, registerOutputs_24__8, registerOutputs_24__7, 
         registerOutputs_24__6, registerOutputs_24__5, registerOutputs_24__4, 
         registerOutputs_24__3, registerOutputs_24__2, registerOutputs_24__1, 
         registerOutputs_24__0, registerOutputs_25__15, registerOutputs_25__14, 
         registerOutputs_25__13, registerOutputs_25__12, registerOutputs_25__11, 
         registerOutputs_25__10, registerOutputs_25__9, registerOutputs_25__8, 
         registerOutputs_25__7, registerOutputs_25__6, registerOutputs_25__5, 
         registerOutputs_25__4, registerOutputs_25__3, registerOutputs_25__2, 
         registerOutputs_25__1, registerOutputs_25__0, registerOutputs_26__15, 
         registerOutputs_26__14, registerOutputs_26__13, registerOutputs_26__12, 
         registerOutputs_26__11, registerOutputs_26__10, registerOutputs_26__9, 
         registerOutputs_26__8, registerOutputs_26__7, registerOutputs_26__6, 
         registerOutputs_26__5, registerOutputs_26__4, registerOutputs_26__3, 
         registerOutputs_26__2, registerOutputs_26__1, registerOutputs_26__0, 
         registerOutputs_27__15, registerOutputs_27__14, registerOutputs_27__13, 
         registerOutputs_27__12, registerOutputs_27__11, registerOutputs_27__10, 
         registerOutputs_27__9, registerOutputs_27__8, registerOutputs_27__7, 
         registerOutputs_27__6, registerOutputs_27__5, registerOutputs_27__4, 
         registerOutputs_27__3, registerOutputs_27__2, registerOutputs_27__1, 
         registerOutputs_27__0, registerOutputs_28__15, registerOutputs_28__14, 
         registerOutputs_28__13, registerOutputs_28__12, registerOutputs_28__11, 
         registerOutputs_28__10, registerOutputs_28__9, registerOutputs_28__8, 
         registerOutputs_28__7, registerOutputs_28__6, registerOutputs_28__5, 
         registerOutputs_28__4, registerOutputs_28__3, registerOutputs_28__2, 
         registerOutputs_28__1, registerOutputs_28__0, registerOutputs_29__15, 
         registerOutputs_29__14, registerOutputs_29__13, registerOutputs_29__12, 
         registerOutputs_29__11, registerOutputs_29__10, registerOutputs_29__9, 
         registerOutputs_29__8, registerOutputs_29__7, registerOutputs_29__6, 
         registerOutputs_29__5, registerOutputs_29__4, registerOutputs_29__3, 
         registerOutputs_29__2, registerOutputs_29__1, registerOutputs_29__0, 
         registerOutputs_30__15, registerOutputs_30__14, registerOutputs_30__13, 
         registerOutputs_30__12, registerOutputs_30__11, registerOutputs_30__10, 
         registerOutputs_30__9, registerOutputs_30__8, registerOutputs_30__7, 
         registerOutputs_30__6, registerOutputs_30__5, registerOutputs_30__4, 
         registerOutputs_30__3, registerOutputs_30__2, registerOutputs_30__1, 
         registerOutputs_30__0, registerOutputs_31__15, registerOutputs_31__14, 
         registerOutputs_31__13, registerOutputs_31__12, registerOutputs_31__11, 
         registerOutputs_31__10, registerOutputs_31__9, registerOutputs_31__8, 
         registerOutputs_31__7, registerOutputs_31__6, registerOutputs_31__5, 
         registerOutputs_31__4, registerOutputs_31__3, registerOutputs_31__2, 
         registerOutputs_31__1, registerOutputs_31__0, registerOutputs_32__15, 
         registerOutputs_32__14, registerOutputs_32__13, registerOutputs_32__12, 
         registerOutputs_32__11, registerOutputs_32__10, registerOutputs_32__9, 
         registerOutputs_32__8, registerOutputs_32__7, registerOutputs_32__6, 
         registerOutputs_32__5, registerOutputs_32__4, registerOutputs_32__3, 
         registerOutputs_32__2, registerOutputs_32__1, registerOutputs_32__0, 
         registerOutputs_33__15, registerOutputs_33__14, registerOutputs_33__13, 
         registerOutputs_33__12, registerOutputs_33__11, registerOutputs_33__10, 
         registerOutputs_33__9, registerOutputs_33__8, registerOutputs_33__7, 
         registerOutputs_33__6, registerOutputs_33__5, registerOutputs_33__4, 
         registerOutputs_33__3, registerOutputs_33__2, registerOutputs_33__1, 
         registerOutputs_33__0, registerOutputs_34__15, registerOutputs_34__14, 
         registerOutputs_34__13, registerOutputs_34__12, registerOutputs_34__11, 
         registerOutputs_34__10, registerOutputs_34__9, registerOutputs_34__8, 
         registerOutputs_34__7, registerOutputs_34__6, registerOutputs_34__5, 
         registerOutputs_34__4, registerOutputs_34__3, registerOutputs_34__2, 
         registerOutputs_34__1, registerOutputs_34__0, registerOutputs_35__15, 
         registerOutputs_35__14, registerOutputs_35__13, registerOutputs_35__12, 
         registerOutputs_35__11, registerOutputs_35__10, registerOutputs_35__9, 
         registerOutputs_35__8, registerOutputs_35__7, registerOutputs_35__6, 
         registerOutputs_35__5, registerOutputs_35__4, registerOutputs_35__3, 
         registerOutputs_35__2, registerOutputs_35__1, registerOutputs_35__0, 
         registerOutputs_36__15, registerOutputs_36__14, registerOutputs_36__13, 
         registerOutputs_36__12, registerOutputs_36__11, registerOutputs_36__10, 
         registerOutputs_36__9, registerOutputs_36__8, registerOutputs_36__7, 
         registerOutputs_36__6, registerOutputs_36__5, registerOutputs_36__4, 
         registerOutputs_36__3, registerOutputs_36__2, registerOutputs_36__1, 
         registerOutputs_36__0, registerOutputs_37__15, registerOutputs_37__14, 
         registerOutputs_37__13, registerOutputs_37__12, registerOutputs_37__11, 
         registerOutputs_37__10, registerOutputs_37__9, registerOutputs_37__8, 
         registerOutputs_37__7, registerOutputs_37__6, registerOutputs_37__5, 
         registerOutputs_37__4, registerOutputs_37__3, registerOutputs_37__2, 
         registerOutputs_37__1, registerOutputs_37__0, registerOutputs_38__15, 
         registerOutputs_38__14, registerOutputs_38__13, registerOutputs_38__12, 
         registerOutputs_38__11, registerOutputs_38__10, registerOutputs_38__9, 
         registerOutputs_38__8, registerOutputs_38__7, registerOutputs_38__6, 
         registerOutputs_38__5, registerOutputs_38__4, registerOutputs_38__3, 
         registerOutputs_38__2, registerOutputs_38__1, registerOutputs_38__0, 
         registerOutputs_39__15, registerOutputs_39__14, registerOutputs_39__13, 
         registerOutputs_39__12, registerOutputs_39__11, registerOutputs_39__10, 
         registerOutputs_39__9, registerOutputs_39__8, registerOutputs_39__7, 
         registerOutputs_39__6, registerOutputs_39__5, registerOutputs_39__4, 
         registerOutputs_39__3, registerOutputs_39__2, registerOutputs_39__1, 
         registerOutputs_39__0, registerOutputs_40__15, registerOutputs_40__14, 
         registerOutputs_40__13, registerOutputs_40__12, registerOutputs_40__11, 
         registerOutputs_40__10, registerOutputs_40__9, registerOutputs_40__8, 
         registerOutputs_40__7, registerOutputs_40__6, registerOutputs_40__5, 
         registerOutputs_40__4, registerOutputs_40__3, registerOutputs_40__2, 
         registerOutputs_40__1, registerOutputs_40__0, registerOutputs_41__15, 
         registerOutputs_41__14, registerOutputs_41__13, registerOutputs_41__12, 
         registerOutputs_41__11, registerOutputs_41__10, registerOutputs_41__9, 
         registerOutputs_41__8, registerOutputs_41__7, registerOutputs_41__6, 
         registerOutputs_41__5, registerOutputs_41__4, registerOutputs_41__3, 
         registerOutputs_41__2, registerOutputs_41__1, registerOutputs_41__0, 
         registerOutputs_42__15, registerOutputs_42__14, registerOutputs_42__13, 
         registerOutputs_42__12, registerOutputs_42__11, registerOutputs_42__10, 
         registerOutputs_42__9, registerOutputs_42__8, registerOutputs_42__7, 
         registerOutputs_42__6, registerOutputs_42__5, registerOutputs_42__4, 
         registerOutputs_42__3, registerOutputs_42__2, registerOutputs_42__1, 
         registerOutputs_42__0, registerOutputs_43__15, registerOutputs_43__14, 
         registerOutputs_43__13, registerOutputs_43__12, registerOutputs_43__11, 
         registerOutputs_43__10, registerOutputs_43__9, registerOutputs_43__8, 
         registerOutputs_43__7, registerOutputs_43__6, registerOutputs_43__5, 
         registerOutputs_43__4, registerOutputs_43__3, registerOutputs_43__2, 
         registerOutputs_43__1, registerOutputs_43__0, registerOutputs_44__15, 
         registerOutputs_44__14, registerOutputs_44__13, registerOutputs_44__12, 
         registerOutputs_44__11, registerOutputs_44__10, registerOutputs_44__9, 
         registerOutputs_44__8, registerOutputs_44__7, registerOutputs_44__6, 
         registerOutputs_44__5, registerOutputs_44__4, registerOutputs_44__3, 
         registerOutputs_44__2, registerOutputs_44__1, registerOutputs_44__0, 
         registerOutputs_45__15, registerOutputs_45__14, registerOutputs_45__13, 
         registerOutputs_45__12, registerOutputs_45__11, registerOutputs_45__10, 
         registerOutputs_45__9, registerOutputs_45__8, registerOutputs_45__7, 
         registerOutputs_45__6, registerOutputs_45__5, registerOutputs_45__4, 
         registerOutputs_45__3, registerOutputs_45__2, registerOutputs_45__1, 
         registerOutputs_45__0, registerOutputs_46__15, registerOutputs_46__14, 
         registerOutputs_46__13, registerOutputs_46__12, registerOutputs_46__11, 
         registerOutputs_46__10, registerOutputs_46__9, registerOutputs_46__8, 
         registerOutputs_46__7, registerOutputs_46__6, registerOutputs_46__5, 
         registerOutputs_46__4, registerOutputs_46__3, registerOutputs_46__2, 
         registerOutputs_46__1, registerOutputs_46__0, registerOutputs_47__15, 
         registerOutputs_47__14, registerOutputs_47__13, registerOutputs_47__12, 
         registerOutputs_47__11, registerOutputs_47__10, registerOutputs_47__9, 
         registerOutputs_47__8, registerOutputs_47__7, registerOutputs_47__6, 
         registerOutputs_47__5, registerOutputs_47__4, registerOutputs_47__3, 
         registerOutputs_47__2, registerOutputs_47__1, registerOutputs_47__0, 
         registerOutputs_48__15, registerOutputs_48__14, registerOutputs_48__13, 
         registerOutputs_48__12, registerOutputs_48__11, registerOutputs_48__10, 
         registerOutputs_48__9, registerOutputs_48__8, registerOutputs_48__7, 
         registerOutputs_48__6, registerOutputs_48__5, registerOutputs_48__4, 
         registerOutputs_48__3, registerOutputs_48__2, registerOutputs_48__1, 
         registerOutputs_48__0, registerOutputs_49__15, registerOutputs_49__14, 
         registerOutputs_49__13, registerOutputs_49__12, registerOutputs_49__11, 
         registerOutputs_49__10, registerOutputs_49__9, registerOutputs_49__8, 
         registerOutputs_49__7, registerOutputs_49__6, registerOutputs_49__5, 
         registerOutputs_49__4, registerOutputs_49__3, registerOutputs_49__2, 
         registerOutputs_49__1, registerOutputs_49__0, registerOutputs_50__15, 
         registerOutputs_50__14, registerOutputs_50__13, registerOutputs_50__12, 
         registerOutputs_50__11, registerOutputs_50__10, registerOutputs_50__9, 
         registerOutputs_50__8, registerOutputs_50__7, registerOutputs_50__6, 
         registerOutputs_50__5, registerOutputs_50__4, registerOutputs_50__3, 
         registerOutputs_50__2, registerOutputs_50__1, registerOutputs_50__0, 
         registerOutputs_51__15, registerOutputs_51__14, registerOutputs_51__13, 
         registerOutputs_51__12, registerOutputs_51__11, registerOutputs_51__10, 
         registerOutputs_51__9, registerOutputs_51__8, registerOutputs_51__7, 
         registerOutputs_51__6, registerOutputs_51__5, registerOutputs_51__4, 
         registerOutputs_51__3, registerOutputs_51__2, registerOutputs_51__1, 
         registerOutputs_51__0, registerOutputs_52__15, registerOutputs_52__14, 
         registerOutputs_52__13, registerOutputs_52__12, registerOutputs_52__11, 
         registerOutputs_52__10, registerOutputs_52__9, registerOutputs_52__8, 
         registerOutputs_52__7, registerOutputs_52__6, registerOutputs_52__5, 
         registerOutputs_52__4, registerOutputs_52__3, registerOutputs_52__2, 
         registerOutputs_52__1, registerOutputs_52__0, registerOutputs_53__15, 
         registerOutputs_53__14, registerOutputs_53__13, registerOutputs_53__12, 
         registerOutputs_53__11, registerOutputs_53__10, registerOutputs_53__9, 
         registerOutputs_53__8, registerOutputs_53__7, registerOutputs_53__6, 
         registerOutputs_53__5, registerOutputs_53__4, registerOutputs_53__3, 
         registerOutputs_53__2, registerOutputs_53__1, registerOutputs_53__0, 
         registerOutputs_54__15, registerOutputs_54__14, registerOutputs_54__13, 
         registerOutputs_54__12, registerOutputs_54__11, registerOutputs_54__10, 
         registerOutputs_54__9, registerOutputs_54__8, registerOutputs_54__7, 
         registerOutputs_54__6, registerOutputs_54__5, registerOutputs_54__4, 
         registerOutputs_54__3, registerOutputs_54__2, registerOutputs_54__1, 
         registerOutputs_54__0, registerOutputs_55__15, registerOutputs_55__14, 
         registerOutputs_55__13, registerOutputs_55__12, registerOutputs_55__11, 
         registerOutputs_55__10, registerOutputs_55__9, registerOutputs_55__8, 
         registerOutputs_55__7, registerOutputs_55__6, registerOutputs_55__5, 
         registerOutputs_55__4, registerOutputs_55__3, registerOutputs_55__2, 
         registerOutputs_55__1, registerOutputs_55__0, registerOutputs_56__15, 
         registerOutputs_56__14, registerOutputs_56__13, registerOutputs_56__12, 
         registerOutputs_56__11, registerOutputs_56__10, registerOutputs_56__9, 
         registerOutputs_56__8, registerOutputs_56__7, registerOutputs_56__6, 
         registerOutputs_56__5, registerOutputs_56__4, registerOutputs_56__3, 
         registerOutputs_56__2, registerOutputs_56__1, registerOutputs_56__0, 
         registerOutputs_57__15, registerOutputs_57__14, registerOutputs_57__13, 
         registerOutputs_57__12, registerOutputs_57__11, registerOutputs_57__10, 
         registerOutputs_57__9, registerOutputs_57__8, registerOutputs_57__7, 
         registerOutputs_57__6, registerOutputs_57__5, registerOutputs_57__4, 
         registerOutputs_57__3, registerOutputs_57__2, registerOutputs_57__1, 
         registerOutputs_57__0, registerOutputs_58__15, registerOutputs_58__14, 
         registerOutputs_58__13, registerOutputs_58__12, registerOutputs_58__11, 
         registerOutputs_58__10, registerOutputs_58__9, registerOutputs_58__8, 
         registerOutputs_58__7, registerOutputs_58__6, registerOutputs_58__5, 
         registerOutputs_58__4, registerOutputs_58__3, registerOutputs_58__2, 
         registerOutputs_58__1, registerOutputs_58__0, registerOutputs_59__15, 
         registerOutputs_59__14, registerOutputs_59__13, registerOutputs_59__12, 
         registerOutputs_59__11, registerOutputs_59__10, registerOutputs_59__9, 
         registerOutputs_59__8, registerOutputs_59__7, registerOutputs_59__6, 
         registerOutputs_59__5, registerOutputs_59__4, registerOutputs_59__3, 
         registerOutputs_59__2, registerOutputs_59__1, registerOutputs_59__0, 
         registerOutputs_60__15, registerOutputs_60__14, registerOutputs_60__13, 
         registerOutputs_60__12, registerOutputs_60__11, registerOutputs_60__10, 
         registerOutputs_60__9, registerOutputs_60__8, registerOutputs_60__7, 
         registerOutputs_60__6, registerOutputs_60__5, registerOutputs_60__4, 
         registerOutputs_60__3, registerOutputs_60__2, registerOutputs_60__1, 
         registerOutputs_60__0, registerOutputs_61__15, registerOutputs_61__14, 
         registerOutputs_61__13, registerOutputs_61__12, registerOutputs_61__11, 
         registerOutputs_61__10, registerOutputs_61__9, registerOutputs_61__8, 
         registerOutputs_61__7, registerOutputs_61__6, registerOutputs_61__5, 
         registerOutputs_61__4, registerOutputs_61__3, registerOutputs_61__2, 
         registerOutputs_61__1, registerOutputs_61__0, registerOutputs_62__15, 
         registerOutputs_62__14, registerOutputs_62__13, registerOutputs_62__12, 
         registerOutputs_62__11, registerOutputs_62__10, registerOutputs_62__9, 
         registerOutputs_62__8, registerOutputs_62__7, registerOutputs_62__6, 
         registerOutputs_62__5, registerOutputs_62__4, registerOutputs_62__3, 
         registerOutputs_62__2, registerOutputs_62__1, registerOutputs_62__0, 
         registerOutputs_63__15, registerOutputs_63__14, registerOutputs_63__13, 
         registerOutputs_63__12, registerOutputs_63__11, registerOutputs_63__10, 
         registerOutputs_63__9, registerOutputs_63__8, registerOutputs_63__7, 
         registerOutputs_63__6, registerOutputs_63__5, registerOutputs_63__4, 
         registerOutputs_63__3, registerOutputs_63__2, registerOutputs_63__1, 
         registerOutputs_63__0, registerOutputs_64__15, registerOutputs_64__14, 
         registerOutputs_64__13, registerOutputs_64__12, registerOutputs_64__11, 
         registerOutputs_64__10, registerOutputs_64__9, registerOutputs_64__8, 
         registerOutputs_64__7, registerOutputs_64__6, registerOutputs_64__5, 
         registerOutputs_64__4, registerOutputs_64__3, registerOutputs_64__2, 
         registerOutputs_64__1, registerOutputs_64__0, registerOutputs_65__15, 
         registerOutputs_65__14, registerOutputs_65__13, registerOutputs_65__12, 
         registerOutputs_65__11, registerOutputs_65__10, registerOutputs_65__9, 
         registerOutputs_65__8, registerOutputs_65__7, registerOutputs_65__6, 
         registerOutputs_65__5, registerOutputs_65__4, registerOutputs_65__3, 
         registerOutputs_65__2, registerOutputs_65__1, registerOutputs_65__0, 
         registerOutputs_66__15, registerOutputs_66__14, registerOutputs_66__13, 
         registerOutputs_66__12, registerOutputs_66__11, registerOutputs_66__10, 
         registerOutputs_66__9, registerOutputs_66__8, registerOutputs_66__7, 
         registerOutputs_66__6, registerOutputs_66__5, registerOutputs_66__4, 
         registerOutputs_66__3, registerOutputs_66__2, registerOutputs_66__1, 
         registerOutputs_66__0, registerOutputs_67__15, registerOutputs_67__14, 
         registerOutputs_67__13, registerOutputs_67__12, registerOutputs_67__11, 
         registerOutputs_67__10, registerOutputs_67__9, registerOutputs_67__8, 
         registerOutputs_67__7, registerOutputs_67__6, registerOutputs_67__5, 
         registerOutputs_67__4, registerOutputs_67__3, registerOutputs_67__2, 
         registerOutputs_67__1, registerOutputs_67__0, registerOutputs_68__15, 
         registerOutputs_68__14, registerOutputs_68__13, registerOutputs_68__12, 
         registerOutputs_68__11, registerOutputs_68__10, registerOutputs_68__9, 
         registerOutputs_68__8, registerOutputs_68__7, registerOutputs_68__6, 
         registerOutputs_68__5, registerOutputs_68__4, registerOutputs_68__3, 
         registerOutputs_68__2, registerOutputs_68__1, registerOutputs_68__0, 
         registerOutputs_69__15, registerOutputs_69__14, registerOutputs_69__13, 
         registerOutputs_69__12, registerOutputs_69__11, registerOutputs_69__10, 
         registerOutputs_69__9, registerOutputs_69__8, registerOutputs_69__7, 
         registerOutputs_69__6, registerOutputs_69__5, registerOutputs_69__4, 
         registerOutputs_69__3, registerOutputs_69__2, registerOutputs_69__1, 
         registerOutputs_69__0, registerOutputs_70__15, registerOutputs_70__14, 
         registerOutputs_70__13, registerOutputs_70__12, registerOutputs_70__11, 
         registerOutputs_70__10, registerOutputs_70__9, registerOutputs_70__8, 
         registerOutputs_70__7, registerOutputs_70__6, registerOutputs_70__5, 
         registerOutputs_70__4, registerOutputs_70__3, registerOutputs_70__2, 
         registerOutputs_70__1, registerOutputs_70__0, registerOutputs_71__15, 
         registerOutputs_71__14, registerOutputs_71__13, registerOutputs_71__12, 
         registerOutputs_71__11, registerOutputs_71__10, registerOutputs_71__9, 
         registerOutputs_71__8, registerOutputs_71__7, registerOutputs_71__6, 
         registerOutputs_71__5, registerOutputs_71__4, registerOutputs_71__3, 
         registerOutputs_71__2, registerOutputs_71__1, registerOutputs_71__0, 
         registerOutputs_72__15, registerOutputs_72__14, registerOutputs_72__13, 
         registerOutputs_72__12, registerOutputs_72__11, registerOutputs_72__10, 
         registerOutputs_72__9, registerOutputs_72__8, registerOutputs_72__7, 
         registerOutputs_72__6, registerOutputs_72__5, registerOutputs_72__4, 
         registerOutputs_72__3, registerOutputs_72__2, registerOutputs_72__1, 
         registerOutputs_72__0, registerOutputs_73__15, registerOutputs_73__14, 
         registerOutputs_73__13, registerOutputs_73__12, registerOutputs_73__11, 
         registerOutputs_73__10, registerOutputs_73__9, registerOutputs_73__8, 
         registerOutputs_73__7, registerOutputs_73__6, registerOutputs_73__5, 
         registerOutputs_73__4, registerOutputs_73__3, registerOutputs_73__2, 
         registerOutputs_73__1, registerOutputs_73__0, registerOutputs_74__15, 
         registerOutputs_74__14, registerOutputs_74__13, registerOutputs_74__12, 
         registerOutputs_74__11, registerOutputs_74__10, registerOutputs_74__9, 
         registerOutputs_74__8, registerOutputs_74__7, registerOutputs_74__6, 
         registerOutputs_74__5, registerOutputs_74__4, registerOutputs_74__3, 
         registerOutputs_74__2, registerOutputs_74__1, registerOutputs_74__0, 
         registerOutputs_75__15, registerOutputs_75__14, registerOutputs_75__13, 
         registerOutputs_75__12, registerOutputs_75__11, registerOutputs_75__10, 
         registerOutputs_75__9, registerOutputs_75__8, registerOutputs_75__7, 
         registerOutputs_75__6, registerOutputs_75__5, registerOutputs_75__4, 
         registerOutputs_75__3, registerOutputs_75__2, registerOutputs_75__1, 
         registerOutputs_75__0, registerOutputs_76__15, registerOutputs_76__14, 
         registerOutputs_76__13, registerOutputs_76__12, registerOutputs_76__11, 
         registerOutputs_76__10, registerOutputs_76__9, registerOutputs_76__8, 
         registerOutputs_76__7, registerOutputs_76__6, registerOutputs_76__5, 
         registerOutputs_76__4, registerOutputs_76__3, registerOutputs_76__2, 
         registerOutputs_76__1, registerOutputs_76__0, registerOutputs_77__15, 
         registerOutputs_77__14, registerOutputs_77__13, registerOutputs_77__12, 
         registerOutputs_77__11, registerOutputs_77__10, registerOutputs_77__9, 
         registerOutputs_77__8, registerOutputs_77__7, registerOutputs_77__6, 
         registerOutputs_77__5, registerOutputs_77__4, registerOutputs_77__3, 
         registerOutputs_77__2, registerOutputs_77__1, registerOutputs_77__0, 
         registerOutputs_78__15, registerOutputs_78__14, registerOutputs_78__13, 
         registerOutputs_78__12, registerOutputs_78__11, registerOutputs_78__10, 
         registerOutputs_78__9, registerOutputs_78__8, registerOutputs_78__7, 
         registerOutputs_78__6, registerOutputs_78__5, registerOutputs_78__4, 
         registerOutputs_78__3, registerOutputs_78__2, registerOutputs_78__1, 
         registerOutputs_78__0, registerOutputs_79__15, registerOutputs_79__14, 
         registerOutputs_79__13, registerOutputs_79__12, registerOutputs_79__11, 
         registerOutputs_79__10, registerOutputs_79__9, registerOutputs_79__8, 
         registerOutputs_79__7, registerOutputs_79__6, registerOutputs_79__5, 
         registerOutputs_79__4, registerOutputs_79__3, registerOutputs_79__2, 
         registerOutputs_79__1, registerOutputs_79__0, registerOutputs_80__15, 
         registerOutputs_80__14, registerOutputs_80__13, registerOutputs_80__12, 
         registerOutputs_80__11, registerOutputs_80__10, registerOutputs_80__9, 
         registerOutputs_80__8, registerOutputs_80__7, registerOutputs_80__6, 
         registerOutputs_80__5, registerOutputs_80__4, registerOutputs_80__3, 
         registerOutputs_80__2, registerOutputs_80__1, registerOutputs_80__0, 
         registerOutputs_81__15, registerOutputs_81__14, registerOutputs_81__13, 
         registerOutputs_81__12, registerOutputs_81__11, registerOutputs_81__10, 
         registerOutputs_81__9, registerOutputs_81__8, registerOutputs_81__7, 
         registerOutputs_81__6, registerOutputs_81__5, registerOutputs_81__4, 
         registerOutputs_81__3, registerOutputs_81__2, registerOutputs_81__1, 
         registerOutputs_81__0, registerOutputs_82__15, registerOutputs_82__14, 
         registerOutputs_82__13, registerOutputs_82__12, registerOutputs_82__11, 
         registerOutputs_82__10, registerOutputs_82__9, registerOutputs_82__8, 
         registerOutputs_82__7, registerOutputs_82__6, registerOutputs_82__5, 
         registerOutputs_82__4, registerOutputs_82__3, registerOutputs_82__2, 
         registerOutputs_82__1, registerOutputs_82__0, registerOutputs_83__15, 
         registerOutputs_83__14, registerOutputs_83__13, registerOutputs_83__12, 
         registerOutputs_83__11, registerOutputs_83__10, registerOutputs_83__9, 
         registerOutputs_83__8, registerOutputs_83__7, registerOutputs_83__6, 
         registerOutputs_83__5, registerOutputs_83__4, registerOutputs_83__3, 
         registerOutputs_83__2, registerOutputs_83__1, registerOutputs_83__0, 
         registerOutputs_84__15, registerOutputs_84__14, registerOutputs_84__13, 
         registerOutputs_84__12, registerOutputs_84__11, registerOutputs_84__10, 
         registerOutputs_84__9, registerOutputs_84__8, registerOutputs_84__7, 
         registerOutputs_84__6, registerOutputs_84__5, registerOutputs_84__4, 
         registerOutputs_84__3, registerOutputs_84__2, registerOutputs_84__1, 
         registerOutputs_84__0, registerOutputs_85__15, registerOutputs_85__14, 
         registerOutputs_85__13, registerOutputs_85__12, registerOutputs_85__11, 
         registerOutputs_85__10, registerOutputs_85__9, registerOutputs_85__8, 
         registerOutputs_85__7, registerOutputs_85__6, registerOutputs_85__5, 
         registerOutputs_85__4, registerOutputs_85__3, registerOutputs_85__2, 
         registerOutputs_85__1, registerOutputs_85__0, registerOutputs_86__15, 
         registerOutputs_86__14, registerOutputs_86__13, registerOutputs_86__12, 
         registerOutputs_86__11, registerOutputs_86__10, registerOutputs_86__9, 
         registerOutputs_86__8, registerOutputs_86__7, registerOutputs_86__6, 
         registerOutputs_86__5, registerOutputs_86__4, registerOutputs_86__3, 
         registerOutputs_86__2, registerOutputs_86__1, registerOutputs_86__0, 
         registerOutputs_87__15, registerOutputs_87__14, registerOutputs_87__13, 
         registerOutputs_87__12, registerOutputs_87__11, registerOutputs_87__10, 
         registerOutputs_87__9, registerOutputs_87__8, registerOutputs_87__7, 
         registerOutputs_87__6, registerOutputs_87__5, registerOutputs_87__4, 
         registerOutputs_87__3, registerOutputs_87__2, registerOutputs_87__1, 
         registerOutputs_87__0, registerOutputs_88__15, registerOutputs_88__14, 
         registerOutputs_88__13, registerOutputs_88__12, registerOutputs_88__11, 
         registerOutputs_88__10, registerOutputs_88__9, registerOutputs_88__8, 
         registerOutputs_88__7, registerOutputs_88__6, registerOutputs_88__5, 
         registerOutputs_88__4, registerOutputs_88__3, registerOutputs_88__2, 
         registerOutputs_88__1, registerOutputs_88__0, registerOutputs_89__15, 
         registerOutputs_89__14, registerOutputs_89__13, registerOutputs_89__12, 
         registerOutputs_89__11, registerOutputs_89__10, registerOutputs_89__9, 
         registerOutputs_89__8, registerOutputs_89__7, registerOutputs_89__6, 
         registerOutputs_89__5, registerOutputs_89__4, registerOutputs_89__3, 
         registerOutputs_89__2, registerOutputs_89__1, registerOutputs_89__0, 
         registerOutputs_90__15, registerOutputs_90__14, registerOutputs_90__13, 
         registerOutputs_90__12, registerOutputs_90__11, registerOutputs_90__10, 
         registerOutputs_90__9, registerOutputs_90__8, registerOutputs_90__7, 
         registerOutputs_90__6, registerOutputs_90__5, registerOutputs_90__4, 
         registerOutputs_90__3, registerOutputs_90__2, registerOutputs_90__1, 
         registerOutputs_90__0, registerOutputs_91__15, registerOutputs_91__14, 
         registerOutputs_91__13, registerOutputs_91__12, registerOutputs_91__11, 
         registerOutputs_91__10, registerOutputs_91__9, registerOutputs_91__8, 
         registerOutputs_91__7, registerOutputs_91__6, registerOutputs_91__5, 
         registerOutputs_91__4, registerOutputs_91__3, registerOutputs_91__2, 
         registerOutputs_91__1, registerOutputs_91__0, registerOutputs_92__15, 
         registerOutputs_92__14, registerOutputs_92__13, registerOutputs_92__12, 
         registerOutputs_92__11, registerOutputs_92__10, registerOutputs_92__9, 
         registerOutputs_92__8, registerOutputs_92__7, registerOutputs_92__6, 
         registerOutputs_92__5, registerOutputs_92__4, registerOutputs_92__3, 
         registerOutputs_92__2, registerOutputs_92__1, registerOutputs_92__0, 
         registerOutputs_93__15, registerOutputs_93__14, registerOutputs_93__13, 
         registerOutputs_93__12, registerOutputs_93__11, registerOutputs_93__10, 
         registerOutputs_93__9, registerOutputs_93__8, registerOutputs_93__7, 
         registerOutputs_93__6, registerOutputs_93__5, registerOutputs_93__4, 
         registerOutputs_93__3, registerOutputs_93__2, registerOutputs_93__1, 
         registerOutputs_93__0, registerOutputs_94__15, registerOutputs_94__14, 
         registerOutputs_94__13, registerOutputs_94__12, registerOutputs_94__11, 
         registerOutputs_94__10, registerOutputs_94__9, registerOutputs_94__8, 
         registerOutputs_94__7, registerOutputs_94__6, registerOutputs_94__5, 
         registerOutputs_94__4, registerOutputs_94__3, registerOutputs_94__2, 
         registerOutputs_94__1, registerOutputs_94__0, registerOutputs_95__15, 
         registerOutputs_95__14, registerOutputs_95__13, registerOutputs_95__12, 
         registerOutputs_95__11, registerOutputs_95__10, registerOutputs_95__9, 
         registerOutputs_95__8, registerOutputs_95__7, registerOutputs_95__6, 
         registerOutputs_95__5, registerOutputs_95__4, registerOutputs_95__3, 
         registerOutputs_95__2, registerOutputs_95__1, registerOutputs_95__0, 
         registerOutputs_96__15, registerOutputs_96__14, registerOutputs_96__13, 
         registerOutputs_96__12, registerOutputs_96__11, registerOutputs_96__10, 
         registerOutputs_96__9, registerOutputs_96__8, registerOutputs_96__7, 
         registerOutputs_96__6, registerOutputs_96__5, registerOutputs_96__4, 
         registerOutputs_96__3, registerOutputs_96__2, registerOutputs_96__1, 
         registerOutputs_96__0, registerOutputs_97__15, registerOutputs_97__14, 
         registerOutputs_97__13, registerOutputs_97__12, registerOutputs_97__11, 
         registerOutputs_97__10, registerOutputs_97__9, registerOutputs_97__8, 
         registerOutputs_97__7, registerOutputs_97__6, registerOutputs_97__5, 
         registerOutputs_97__4, registerOutputs_97__3, registerOutputs_97__2, 
         registerOutputs_97__1, registerOutputs_97__0, registerOutputs_98__15, 
         registerOutputs_98__14, registerOutputs_98__13, registerOutputs_98__12, 
         registerOutputs_98__11, registerOutputs_98__10, registerOutputs_98__9, 
         registerOutputs_98__8, registerOutputs_98__7, registerOutputs_98__6, 
         registerOutputs_98__5, registerOutputs_98__4, registerOutputs_98__3, 
         registerOutputs_98__2, registerOutputs_98__1, registerOutputs_98__0, 
         registerOutputs_99__15, registerOutputs_99__14, registerOutputs_99__13, 
         registerOutputs_99__12, registerOutputs_99__11, registerOutputs_99__10, 
         registerOutputs_99__9, registerOutputs_99__8, registerOutputs_99__7, 
         registerOutputs_99__6, registerOutputs_99__5, registerOutputs_99__4, 
         registerOutputs_99__3, registerOutputs_99__2, registerOutputs_99__1, 
         registerOutputs_99__0, registerOutputs_100__15, registerOutputs_100__14, 
         registerOutputs_100__13, registerOutputs_100__12, 
         registerOutputs_100__11, registerOutputs_100__10, 
         registerOutputs_100__9, registerOutputs_100__8, registerOutputs_100__7, 
         registerOutputs_100__6, registerOutputs_100__5, registerOutputs_100__4, 
         registerOutputs_100__3, registerOutputs_100__2, registerOutputs_100__1, 
         registerOutputs_100__0, registerOutputs_101__15, 
         registerOutputs_101__14, registerOutputs_101__13, 
         registerOutputs_101__12, registerOutputs_101__11, 
         registerOutputs_101__10, registerOutputs_101__9, registerOutputs_101__8, 
         registerOutputs_101__7, registerOutputs_101__6, registerOutputs_101__5, 
         registerOutputs_101__4, registerOutputs_101__3, registerOutputs_101__2, 
         registerOutputs_101__1, registerOutputs_101__0, registerOutputs_102__15, 
         registerOutputs_102__14, registerOutputs_102__13, 
         registerOutputs_102__12, registerOutputs_102__11, 
         registerOutputs_102__10, registerOutputs_102__9, registerOutputs_102__8, 
         registerOutputs_102__7, registerOutputs_102__6, registerOutputs_102__5, 
         registerOutputs_102__4, registerOutputs_102__3, registerOutputs_102__2, 
         registerOutputs_102__1, registerOutputs_102__0, registerOutputs_103__15, 
         registerOutputs_103__14, registerOutputs_103__13, 
         registerOutputs_103__12, registerOutputs_103__11, 
         registerOutputs_103__10, registerOutputs_103__9, registerOutputs_103__8, 
         registerOutputs_103__7, registerOutputs_103__6, registerOutputs_103__5, 
         registerOutputs_103__4, registerOutputs_103__3, registerOutputs_103__2, 
         registerOutputs_103__1, registerOutputs_103__0, registerOutputs_104__15, 
         registerOutputs_104__14, registerOutputs_104__13, 
         registerOutputs_104__12, registerOutputs_104__11, 
         registerOutputs_104__10, registerOutputs_104__9, registerOutputs_104__8, 
         registerOutputs_104__7, registerOutputs_104__6, registerOutputs_104__5, 
         registerOutputs_104__4, registerOutputs_104__3, registerOutputs_104__2, 
         registerOutputs_104__1, registerOutputs_104__0, registerOutputs_105__15, 
         registerOutputs_105__14, registerOutputs_105__13, 
         registerOutputs_105__12, registerOutputs_105__11, 
         registerOutputs_105__10, registerOutputs_105__9, registerOutputs_105__8, 
         registerOutputs_105__7, registerOutputs_105__6, registerOutputs_105__5, 
         registerOutputs_105__4, registerOutputs_105__3, registerOutputs_105__2, 
         registerOutputs_105__1, registerOutputs_105__0, registerOutputs_106__15, 
         registerOutputs_106__14, registerOutputs_106__13, 
         registerOutputs_106__12, registerOutputs_106__11, 
         registerOutputs_106__10, registerOutputs_106__9, registerOutputs_106__8, 
         registerOutputs_106__7, registerOutputs_106__6, registerOutputs_106__5, 
         registerOutputs_106__4, registerOutputs_106__3, registerOutputs_106__2, 
         registerOutputs_106__1, registerOutputs_106__0, registerOutputs_107__15, 
         registerOutputs_107__14, registerOutputs_107__13, 
         registerOutputs_107__12, registerOutputs_107__11, 
         registerOutputs_107__10, registerOutputs_107__9, registerOutputs_107__8, 
         registerOutputs_107__7, registerOutputs_107__6, registerOutputs_107__5, 
         registerOutputs_107__4, registerOutputs_107__3, registerOutputs_107__2, 
         registerOutputs_107__1, registerOutputs_107__0, registerOutputs_108__15, 
         registerOutputs_108__14, registerOutputs_108__13, 
         registerOutputs_108__12, registerOutputs_108__11, 
         registerOutputs_108__10, registerOutputs_108__9, registerOutputs_108__8, 
         registerOutputs_108__7, registerOutputs_108__6, registerOutputs_108__5, 
         registerOutputs_108__4, registerOutputs_108__3, registerOutputs_108__2, 
         registerOutputs_108__1, registerOutputs_108__0, registerOutputs_109__15, 
         registerOutputs_109__14, registerOutputs_109__13, 
         registerOutputs_109__12, registerOutputs_109__11, 
         registerOutputs_109__10, registerOutputs_109__9, registerOutputs_109__8, 
         registerOutputs_109__7, registerOutputs_109__6, registerOutputs_109__5, 
         registerOutputs_109__4, registerOutputs_109__3, registerOutputs_109__2, 
         registerOutputs_109__1, registerOutputs_109__0, registerOutputs_110__15, 
         registerOutputs_110__14, registerOutputs_110__13, 
         registerOutputs_110__12, registerOutputs_110__11, 
         registerOutputs_110__10, registerOutputs_110__9, registerOutputs_110__8, 
         registerOutputs_110__7, registerOutputs_110__6, registerOutputs_110__5, 
         registerOutputs_110__4, registerOutputs_110__3, registerOutputs_110__2, 
         registerOutputs_110__1, registerOutputs_110__0, registerOutputs_111__15, 
         registerOutputs_111__14, registerOutputs_111__13, 
         registerOutputs_111__12, registerOutputs_111__11, 
         registerOutputs_111__10, registerOutputs_111__9, registerOutputs_111__8, 
         registerOutputs_111__7, registerOutputs_111__6, registerOutputs_111__5, 
         registerOutputs_111__4, registerOutputs_111__3, registerOutputs_111__2, 
         registerOutputs_111__1, registerOutputs_111__0, registerOutputs_112__15, 
         registerOutputs_112__14, registerOutputs_112__13, 
         registerOutputs_112__12, registerOutputs_112__11, 
         registerOutputs_112__10, registerOutputs_112__9, registerOutputs_112__8, 
         registerOutputs_112__7, registerOutputs_112__6, registerOutputs_112__5, 
         registerOutputs_112__4, registerOutputs_112__3, registerOutputs_112__2, 
         registerOutputs_112__1, registerOutputs_112__0, registerOutputs_113__15, 
         registerOutputs_113__14, registerOutputs_113__13, 
         registerOutputs_113__12, registerOutputs_113__11, 
         registerOutputs_113__10, registerOutputs_113__9, registerOutputs_113__8, 
         registerOutputs_113__7, registerOutputs_113__6, registerOutputs_113__5, 
         registerOutputs_113__4, registerOutputs_113__3, registerOutputs_113__2, 
         registerOutputs_113__1, registerOutputs_113__0, registerOutputs_114__15, 
         registerOutputs_114__14, registerOutputs_114__13, 
         registerOutputs_114__12, registerOutputs_114__11, 
         registerOutputs_114__10, registerOutputs_114__9, registerOutputs_114__8, 
         registerOutputs_114__7, registerOutputs_114__6, registerOutputs_114__5, 
         registerOutputs_114__4, registerOutputs_114__3, registerOutputs_114__2, 
         registerOutputs_114__1, registerOutputs_114__0, registerOutputs_115__15, 
         registerOutputs_115__14, registerOutputs_115__13, 
         registerOutputs_115__12, registerOutputs_115__11, 
         registerOutputs_115__10, registerOutputs_115__9, registerOutputs_115__8, 
         registerOutputs_115__7, registerOutputs_115__6, registerOutputs_115__5, 
         registerOutputs_115__4, registerOutputs_115__3, registerOutputs_115__2, 
         registerOutputs_115__1, registerOutputs_115__0, registerOutputs_116__15, 
         registerOutputs_116__14, registerOutputs_116__13, 
         registerOutputs_116__12, registerOutputs_116__11, 
         registerOutputs_116__10, registerOutputs_116__9, registerOutputs_116__8, 
         registerOutputs_116__7, registerOutputs_116__6, registerOutputs_116__5, 
         registerOutputs_116__4, registerOutputs_116__3, registerOutputs_116__2, 
         registerOutputs_116__1, registerOutputs_116__0, registerOutputs_117__15, 
         registerOutputs_117__14, registerOutputs_117__13, 
         registerOutputs_117__12, registerOutputs_117__11, 
         registerOutputs_117__10, registerOutputs_117__9, registerOutputs_117__8, 
         registerOutputs_117__7, registerOutputs_117__6, registerOutputs_117__5, 
         registerOutputs_117__4, registerOutputs_117__3, registerOutputs_117__2, 
         registerOutputs_117__1, registerOutputs_117__0, registerOutputs_118__15, 
         registerOutputs_118__14, registerOutputs_118__13, 
         registerOutputs_118__12, registerOutputs_118__11, 
         registerOutputs_118__10, registerOutputs_118__9, registerOutputs_118__8, 
         registerOutputs_118__7, registerOutputs_118__6, registerOutputs_118__5, 
         registerOutputs_118__4, registerOutputs_118__3, registerOutputs_118__2, 
         registerOutputs_118__1, registerOutputs_118__0, registerOutputs_119__15, 
         registerOutputs_119__14, registerOutputs_119__13, 
         registerOutputs_119__12, registerOutputs_119__11, 
         registerOutputs_119__10, registerOutputs_119__9, registerOutputs_119__8, 
         registerOutputs_119__7, registerOutputs_119__6, registerOutputs_119__5, 
         registerOutputs_119__4, registerOutputs_119__3, registerOutputs_119__2, 
         registerOutputs_119__1, registerOutputs_119__0, registerOutputs_120__15, 
         registerOutputs_120__14, registerOutputs_120__13, 
         registerOutputs_120__12, registerOutputs_120__11, 
         registerOutputs_120__10, registerOutputs_120__9, registerOutputs_120__8, 
         registerOutputs_120__7, registerOutputs_120__6, registerOutputs_120__5, 
         registerOutputs_120__4, registerOutputs_120__3, registerOutputs_120__2, 
         registerOutputs_120__1, registerOutputs_120__0, registerOutputs_121__15, 
         registerOutputs_121__14, registerOutputs_121__13, 
         registerOutputs_121__12, registerOutputs_121__11, 
         registerOutputs_121__10, registerOutputs_121__9, registerOutputs_121__8, 
         registerOutputs_121__7, registerOutputs_121__6, registerOutputs_121__5, 
         registerOutputs_121__4, registerOutputs_121__3, registerOutputs_121__2, 
         registerOutputs_121__1, registerOutputs_121__0, registerOutputs_122__15, 
         registerOutputs_122__14, registerOutputs_122__13, 
         registerOutputs_122__12, registerOutputs_122__11, 
         registerOutputs_122__10, registerOutputs_122__9, registerOutputs_122__8, 
         registerOutputs_122__7, registerOutputs_122__6, registerOutputs_122__5, 
         registerOutputs_122__4, registerOutputs_122__3, registerOutputs_122__2, 
         registerOutputs_122__1, registerOutputs_122__0, registerOutputs_123__15, 
         registerOutputs_123__14, registerOutputs_123__13, 
         registerOutputs_123__12, registerOutputs_123__11, 
         registerOutputs_123__10, registerOutputs_123__9, registerOutputs_123__8, 
         registerOutputs_123__7, registerOutputs_123__6, registerOutputs_123__5, 
         registerOutputs_123__4, registerOutputs_123__3, registerOutputs_123__2, 
         registerOutputs_123__1, registerOutputs_123__0, registerOutputs_124__15, 
         registerOutputs_124__14, registerOutputs_124__13, 
         registerOutputs_124__12, registerOutputs_124__11, 
         registerOutputs_124__10, registerOutputs_124__9, registerOutputs_124__8, 
         registerOutputs_124__7, registerOutputs_124__6, registerOutputs_124__5, 
         registerOutputs_124__4, registerOutputs_124__3, registerOutputs_124__2, 
         registerOutputs_124__1, registerOutputs_124__0, registerOutputs_125__15, 
         registerOutputs_125__14, registerOutputs_125__13, 
         registerOutputs_125__12, registerOutputs_125__11, 
         registerOutputs_125__10, registerOutputs_125__9, registerOutputs_125__8, 
         registerOutputs_125__7, registerOutputs_125__6, registerOutputs_125__5, 
         registerOutputs_125__4, registerOutputs_125__3, registerOutputs_125__2, 
         registerOutputs_125__1, registerOutputs_125__0, registerOutputs_126__15, 
         registerOutputs_126__14, registerOutputs_126__13, 
         registerOutputs_126__12, registerOutputs_126__11, 
         registerOutputs_126__10, registerOutputs_126__9, registerOutputs_126__8, 
         registerOutputs_126__7, registerOutputs_126__6, registerOutputs_126__5, 
         registerOutputs_126__4, registerOutputs_126__3, registerOutputs_126__2, 
         registerOutputs_126__1, registerOutputs_126__0, registerOutputs_127__15, 
         registerOutputs_127__14, registerOutputs_127__13, 
         registerOutputs_127__12, registerOutputs_127__11, 
         registerOutputs_127__10, registerOutputs_127__9, registerOutputs_127__8, 
         registerOutputs_127__7, registerOutputs_127__6, registerOutputs_127__5, 
         registerOutputs_127__4, registerOutputs_127__3, registerOutputs_127__2, 
         registerOutputs_127__1, registerOutputs_127__0, registerOutputs_128__15, 
         registerOutputs_128__14, registerOutputs_128__13, 
         registerOutputs_128__12, registerOutputs_128__11, 
         registerOutputs_128__10, registerOutputs_128__9, registerOutputs_128__8, 
         registerOutputs_128__7, registerOutputs_128__6, registerOutputs_128__5, 
         registerOutputs_128__4, registerOutputs_128__3, registerOutputs_128__2, 
         registerOutputs_128__1, registerOutputs_128__0, registerOutputs_129__15, 
         registerOutputs_129__14, registerOutputs_129__13, 
         registerOutputs_129__12, registerOutputs_129__11, 
         registerOutputs_129__10, registerOutputs_129__9, registerOutputs_129__8, 
         registerOutputs_129__7, registerOutputs_129__6, registerOutputs_129__5, 
         registerOutputs_129__4, registerOutputs_129__3, registerOutputs_129__2, 
         registerOutputs_129__1, registerOutputs_129__0, registerOutputs_130__15, 
         registerOutputs_130__14, registerOutputs_130__13, 
         registerOutputs_130__12, registerOutputs_130__11, 
         registerOutputs_130__10, registerOutputs_130__9, registerOutputs_130__8, 
         registerOutputs_130__7, registerOutputs_130__6, registerOutputs_130__5, 
         registerOutputs_130__4, registerOutputs_130__3, registerOutputs_130__2, 
         registerOutputs_130__1, registerOutputs_130__0, registerOutputs_131__15, 
         registerOutputs_131__14, registerOutputs_131__13, 
         registerOutputs_131__12, registerOutputs_131__11, 
         registerOutputs_131__10, registerOutputs_131__9, registerOutputs_131__8, 
         registerOutputs_131__7, registerOutputs_131__6, registerOutputs_131__5, 
         registerOutputs_131__4, registerOutputs_131__3, registerOutputs_131__2, 
         registerOutputs_131__1, registerOutputs_131__0, registerOutputs_132__15, 
         registerOutputs_132__14, registerOutputs_132__13, 
         registerOutputs_132__12, registerOutputs_132__11, 
         registerOutputs_132__10, registerOutputs_132__9, registerOutputs_132__8, 
         registerOutputs_132__7, registerOutputs_132__6, registerOutputs_132__5, 
         registerOutputs_132__4, registerOutputs_132__3, registerOutputs_132__2, 
         registerOutputs_132__1, registerOutputs_132__0, registerOutputs_133__15, 
         registerOutputs_133__14, registerOutputs_133__13, 
         registerOutputs_133__12, registerOutputs_133__11, 
         registerOutputs_133__10, registerOutputs_133__9, registerOutputs_133__8, 
         registerOutputs_133__7, registerOutputs_133__6, registerOutputs_133__5, 
         registerOutputs_133__4, registerOutputs_133__3, registerOutputs_133__2, 
         registerOutputs_133__1, registerOutputs_133__0, registerOutputs_134__15, 
         registerOutputs_134__14, registerOutputs_134__13, 
         registerOutputs_134__12, registerOutputs_134__11, 
         registerOutputs_134__10, registerOutputs_134__9, registerOutputs_134__8, 
         registerOutputs_134__7, registerOutputs_134__6, registerOutputs_134__5, 
         registerOutputs_134__4, registerOutputs_134__3, registerOutputs_134__2, 
         registerOutputs_134__1, registerOutputs_134__0, registerOutputs_135__15, 
         registerOutputs_135__14, registerOutputs_135__13, 
         registerOutputs_135__12, registerOutputs_135__11, 
         registerOutputs_135__10, registerOutputs_135__9, registerOutputs_135__8, 
         registerOutputs_135__7, registerOutputs_135__6, registerOutputs_135__5, 
         registerOutputs_135__4, registerOutputs_135__3, registerOutputs_135__2, 
         registerOutputs_135__1, registerOutputs_135__0, registerOutputs_136__15, 
         registerOutputs_136__14, registerOutputs_136__13, 
         registerOutputs_136__12, registerOutputs_136__11, 
         registerOutputs_136__10, registerOutputs_136__9, registerOutputs_136__8, 
         registerOutputs_136__7, registerOutputs_136__6, registerOutputs_136__5, 
         registerOutputs_136__4, registerOutputs_136__3, registerOutputs_136__2, 
         registerOutputs_136__1, registerOutputs_136__0, registerOutputs_137__15, 
         registerOutputs_137__14, registerOutputs_137__13, 
         registerOutputs_137__12, registerOutputs_137__11, 
         registerOutputs_137__10, registerOutputs_137__9, registerOutputs_137__8, 
         registerOutputs_137__7, registerOutputs_137__6, registerOutputs_137__5, 
         registerOutputs_137__4, registerOutputs_137__3, registerOutputs_137__2, 
         registerOutputs_137__1, registerOutputs_137__0, registerOutputs_138__15, 
         registerOutputs_138__14, registerOutputs_138__13, 
         registerOutputs_138__12, registerOutputs_138__11, 
         registerOutputs_138__10, registerOutputs_138__9, registerOutputs_138__8, 
         registerOutputs_138__7, registerOutputs_138__6, registerOutputs_138__5, 
         registerOutputs_138__4, registerOutputs_138__3, registerOutputs_138__2, 
         registerOutputs_138__1, registerOutputs_138__0, registerOutputs_139__15, 
         registerOutputs_139__14, registerOutputs_139__13, 
         registerOutputs_139__12, registerOutputs_139__11, 
         registerOutputs_139__10, registerOutputs_139__9, registerOutputs_139__8, 
         registerOutputs_139__7, registerOutputs_139__6, registerOutputs_139__5, 
         registerOutputs_139__4, registerOutputs_139__3, registerOutputs_139__2, 
         registerOutputs_139__1, registerOutputs_139__0, registerOutputs_140__15, 
         registerOutputs_140__14, registerOutputs_140__13, 
         registerOutputs_140__12, registerOutputs_140__11, 
         registerOutputs_140__10, registerOutputs_140__9, registerOutputs_140__8, 
         registerOutputs_140__7, registerOutputs_140__6, registerOutputs_140__5, 
         registerOutputs_140__4, registerOutputs_140__3, registerOutputs_140__2, 
         registerOutputs_140__1, registerOutputs_140__0, registerOutputs_141__15, 
         registerOutputs_141__14, registerOutputs_141__13, 
         registerOutputs_141__12, registerOutputs_141__11, 
         registerOutputs_141__10, registerOutputs_141__9, registerOutputs_141__8, 
         registerOutputs_141__7, registerOutputs_141__6, registerOutputs_141__5, 
         registerOutputs_141__4, registerOutputs_141__3, registerOutputs_141__2, 
         registerOutputs_141__1, registerOutputs_141__0, registerOutputs_142__15, 
         registerOutputs_142__14, registerOutputs_142__13, 
         registerOutputs_142__12, registerOutputs_142__11, 
         registerOutputs_142__10, registerOutputs_142__9, registerOutputs_142__8, 
         registerOutputs_142__7, registerOutputs_142__6, registerOutputs_142__5, 
         registerOutputs_142__4, registerOutputs_142__3, registerOutputs_142__2, 
         registerOutputs_142__1, registerOutputs_142__0, registerOutputs_143__15, 
         registerOutputs_143__14, registerOutputs_143__13, 
         registerOutputs_143__12, registerOutputs_143__11, 
         registerOutputs_143__10, registerOutputs_143__9, registerOutputs_143__8, 
         registerOutputs_143__7, registerOutputs_143__6, registerOutputs_143__5, 
         registerOutputs_143__4, registerOutputs_143__3, registerOutputs_143__2, 
         registerOutputs_143__1, registerOutputs_143__0, registerOutputs_144__15, 
         registerOutputs_144__14, registerOutputs_144__13, 
         registerOutputs_144__12, registerOutputs_144__11, 
         registerOutputs_144__10, registerOutputs_144__9, registerOutputs_144__8, 
         registerOutputs_144__7, registerOutputs_144__6, registerOutputs_144__5, 
         registerOutputs_144__4, registerOutputs_144__3, registerOutputs_144__2, 
         registerOutputs_144__1, registerOutputs_144__0, registerOutputs_145__15, 
         registerOutputs_145__14, registerOutputs_145__13, 
         registerOutputs_145__12, registerOutputs_145__11, 
         registerOutputs_145__10, registerOutputs_145__9, registerOutputs_145__8, 
         registerOutputs_145__7, registerOutputs_145__6, registerOutputs_145__5, 
         registerOutputs_145__4, registerOutputs_145__3, registerOutputs_145__2, 
         registerOutputs_145__1, registerOutputs_145__0, registerOutputs_146__15, 
         registerOutputs_146__14, registerOutputs_146__13, 
         registerOutputs_146__12, registerOutputs_146__11, 
         registerOutputs_146__10, registerOutputs_146__9, registerOutputs_146__8, 
         registerOutputs_146__7, registerOutputs_146__6, registerOutputs_146__5, 
         registerOutputs_146__4, registerOutputs_146__3, registerOutputs_146__2, 
         registerOutputs_146__1, registerOutputs_146__0, registerOutputs_147__15, 
         registerOutputs_147__14, registerOutputs_147__13, 
         registerOutputs_147__12, registerOutputs_147__11, 
         registerOutputs_147__10, registerOutputs_147__9, registerOutputs_147__8, 
         registerOutputs_147__7, registerOutputs_147__6, registerOutputs_147__5, 
         registerOutputs_147__4, registerOutputs_147__3, registerOutputs_147__2, 
         registerOutputs_147__1, registerOutputs_147__0, registerOutputs_148__15, 
         registerOutputs_148__14, registerOutputs_148__13, 
         registerOutputs_148__12, registerOutputs_148__11, 
         registerOutputs_148__10, registerOutputs_148__9, registerOutputs_148__8, 
         registerOutputs_148__7, registerOutputs_148__6, registerOutputs_148__5, 
         registerOutputs_148__4, registerOutputs_148__3, registerOutputs_148__2, 
         registerOutputs_148__1, registerOutputs_148__0, registerOutputs_149__15, 
         registerOutputs_149__14, registerOutputs_149__13, 
         registerOutputs_149__12, registerOutputs_149__11, 
         registerOutputs_149__10, registerOutputs_149__9, registerOutputs_149__8, 
         registerOutputs_149__7, registerOutputs_149__6, registerOutputs_149__5, 
         registerOutputs_149__4, registerOutputs_149__3, registerOutputs_149__2, 
         registerOutputs_149__1, registerOutputs_149__0, registerOutputs_150__15, 
         registerOutputs_150__14, registerOutputs_150__13, 
         registerOutputs_150__12, registerOutputs_150__11, 
         registerOutputs_150__10, registerOutputs_150__9, registerOutputs_150__8, 
         registerOutputs_150__7, registerOutputs_150__6, registerOutputs_150__5, 
         registerOutputs_150__4, registerOutputs_150__3, registerOutputs_150__2, 
         registerOutputs_150__1, registerOutputs_150__0, registerOutputs_151__15, 
         registerOutputs_151__14, registerOutputs_151__13, 
         registerOutputs_151__12, registerOutputs_151__11, 
         registerOutputs_151__10, registerOutputs_151__9, registerOutputs_151__8, 
         registerOutputs_151__7, registerOutputs_151__6, registerOutputs_151__5, 
         registerOutputs_151__4, registerOutputs_151__3, registerOutputs_151__2, 
         registerOutputs_151__1, registerOutputs_151__0, registerOutputs_152__15, 
         registerOutputs_152__14, registerOutputs_152__13, 
         registerOutputs_152__12, registerOutputs_152__11, 
         registerOutputs_152__10, registerOutputs_152__9, registerOutputs_152__8, 
         registerOutputs_152__7, registerOutputs_152__6, registerOutputs_152__5, 
         registerOutputs_152__4, registerOutputs_152__3, registerOutputs_152__2, 
         registerOutputs_152__1, registerOutputs_152__0, registerOutputs_153__15, 
         registerOutputs_153__14, registerOutputs_153__13, 
         registerOutputs_153__12, registerOutputs_153__11, 
         registerOutputs_153__10, registerOutputs_153__9, registerOutputs_153__8, 
         registerOutputs_153__7, registerOutputs_153__6, registerOutputs_153__5, 
         registerOutputs_153__4, registerOutputs_153__3, registerOutputs_153__2, 
         registerOutputs_153__1, registerOutputs_153__0, registerOutputs_154__15, 
         registerOutputs_154__14, registerOutputs_154__13, 
         registerOutputs_154__12, registerOutputs_154__11, 
         registerOutputs_154__10, registerOutputs_154__9, registerOutputs_154__8, 
         registerOutputs_154__7, registerOutputs_154__6, registerOutputs_154__5, 
         registerOutputs_154__4, registerOutputs_154__3, registerOutputs_154__2, 
         registerOutputs_154__1, registerOutputs_154__0, registerOutputs_155__15, 
         registerOutputs_155__14, registerOutputs_155__13, 
         registerOutputs_155__12, registerOutputs_155__11, 
         registerOutputs_155__10, registerOutputs_155__9, registerOutputs_155__8, 
         registerOutputs_155__7, registerOutputs_155__6, registerOutputs_155__5, 
         registerOutputs_155__4, registerOutputs_155__3, registerOutputs_155__2, 
         registerOutputs_155__1, registerOutputs_155__0, registerOutputs_156__15, 
         registerOutputs_156__14, registerOutputs_156__13, 
         registerOutputs_156__12, registerOutputs_156__11, 
         registerOutputs_156__10, registerOutputs_156__9, registerOutputs_156__8, 
         registerOutputs_156__7, registerOutputs_156__6, registerOutputs_156__5, 
         registerOutputs_156__4, registerOutputs_156__3, registerOutputs_156__2, 
         registerOutputs_156__1, registerOutputs_156__0, registerOutputs_157__15, 
         registerOutputs_157__14, registerOutputs_157__13, 
         registerOutputs_157__12, registerOutputs_157__11, 
         registerOutputs_157__10, registerOutputs_157__9, registerOutputs_157__8, 
         registerOutputs_157__7, registerOutputs_157__6, registerOutputs_157__5, 
         registerOutputs_157__4, registerOutputs_157__3, registerOutputs_157__2, 
         registerOutputs_157__1, registerOutputs_157__0, registerOutputs_158__15, 
         registerOutputs_158__14, registerOutputs_158__13, 
         registerOutputs_158__12, registerOutputs_158__11, 
         registerOutputs_158__10, registerOutputs_158__9, registerOutputs_158__8, 
         registerOutputs_158__7, registerOutputs_158__6, registerOutputs_158__5, 
         registerOutputs_158__4, registerOutputs_158__3, registerOutputs_158__2, 
         registerOutputs_158__1, registerOutputs_158__0, registerOutputs_159__15, 
         registerOutputs_159__14, registerOutputs_159__13, 
         registerOutputs_159__12, registerOutputs_159__11, 
         registerOutputs_159__10, registerOutputs_159__9, registerOutputs_159__8, 
         registerOutputs_159__7, registerOutputs_159__6, registerOutputs_159__5, 
         registerOutputs_159__4, registerOutputs_159__3, registerOutputs_159__2, 
         registerOutputs_159__1, registerOutputs_159__0, registerOutputs_160__15, 
         registerOutputs_160__14, registerOutputs_160__13, 
         registerOutputs_160__12, registerOutputs_160__11, 
         registerOutputs_160__10, registerOutputs_160__9, registerOutputs_160__8, 
         registerOutputs_160__7, registerOutputs_160__6, registerOutputs_160__5, 
         registerOutputs_160__4, registerOutputs_160__3, registerOutputs_160__2, 
         registerOutputs_160__1, registerOutputs_160__0, registerOutputs_161__15, 
         registerOutputs_161__14, registerOutputs_161__13, 
         registerOutputs_161__12, registerOutputs_161__11, 
         registerOutputs_161__10, registerOutputs_161__9, registerOutputs_161__8, 
         registerOutputs_161__7, registerOutputs_161__6, registerOutputs_161__5, 
         registerOutputs_161__4, registerOutputs_161__3, registerOutputs_161__2, 
         registerOutputs_161__1, registerOutputs_161__0, registerOutputs_162__15, 
         registerOutputs_162__14, registerOutputs_162__13, 
         registerOutputs_162__12, registerOutputs_162__11, 
         registerOutputs_162__10, registerOutputs_162__9, registerOutputs_162__8, 
         registerOutputs_162__7, registerOutputs_162__6, registerOutputs_162__5, 
         registerOutputs_162__4, registerOutputs_162__3, registerOutputs_162__2, 
         registerOutputs_162__1, registerOutputs_162__0, registerOutputs_163__15, 
         registerOutputs_163__14, registerOutputs_163__13, 
         registerOutputs_163__12, registerOutputs_163__11, 
         registerOutputs_163__10, registerOutputs_163__9, registerOutputs_163__8, 
         registerOutputs_163__7, registerOutputs_163__6, registerOutputs_163__5, 
         registerOutputs_163__4, registerOutputs_163__3, registerOutputs_163__2, 
         registerOutputs_163__1, registerOutputs_163__0, registerOutputs_164__15, 
         registerOutputs_164__14, registerOutputs_164__13, 
         registerOutputs_164__12, registerOutputs_164__11, 
         registerOutputs_164__10, registerOutputs_164__9, registerOutputs_164__8, 
         registerOutputs_164__7, registerOutputs_164__6, registerOutputs_164__5, 
         registerOutputs_164__4, registerOutputs_164__3, registerOutputs_164__2, 
         registerOutputs_164__1, registerOutputs_164__0, registerOutputs_165__15, 
         registerOutputs_165__14, registerOutputs_165__13, 
         registerOutputs_165__12, registerOutputs_165__11, 
         registerOutputs_165__10, registerOutputs_165__9, registerOutputs_165__8, 
         registerOutputs_165__7, registerOutputs_165__6, registerOutputs_165__5, 
         registerOutputs_165__4, registerOutputs_165__3, registerOutputs_165__2, 
         registerOutputs_165__1, registerOutputs_165__0, registerOutputs_166__15, 
         registerOutputs_166__14, registerOutputs_166__13, 
         registerOutputs_166__12, registerOutputs_166__11, 
         registerOutputs_166__10, registerOutputs_166__9, registerOutputs_166__8, 
         registerOutputs_166__7, registerOutputs_166__6, registerOutputs_166__5, 
         registerOutputs_166__4, registerOutputs_166__3, registerOutputs_166__2, 
         registerOutputs_166__1, registerOutputs_166__0, registerOutputs_167__15, 
         registerOutputs_167__14, registerOutputs_167__13, 
         registerOutputs_167__12, registerOutputs_167__11, 
         registerOutputs_167__10, registerOutputs_167__9, registerOutputs_167__8, 
         registerOutputs_167__7, registerOutputs_167__6, registerOutputs_167__5, 
         registerOutputs_167__4, registerOutputs_167__3, registerOutputs_167__2, 
         registerOutputs_167__1, registerOutputs_167__0, registerOutputs_168__15, 
         registerOutputs_168__14, registerOutputs_168__13, 
         registerOutputs_168__12, registerOutputs_168__11, 
         registerOutputs_168__10, registerOutputs_168__9, registerOutputs_168__8, 
         registerOutputs_168__7, registerOutputs_168__6, registerOutputs_168__5, 
         registerOutputs_168__4, registerOutputs_168__3, registerOutputs_168__2, 
         registerOutputs_168__1, registerOutputs_168__0, registerOutputs_169__15, 
         registerOutputs_169__14, registerOutputs_169__13, 
         registerOutputs_169__12, registerOutputs_169__11, 
         registerOutputs_169__10, registerOutputs_169__9, registerOutputs_169__8, 
         registerOutputs_169__7, registerOutputs_169__6, registerOutputs_169__5, 
         registerOutputs_169__4, registerOutputs_169__3, registerOutputs_169__2, 
         registerOutputs_169__1, registerOutputs_169__0, registerOutputs_170__15, 
         registerOutputs_170__14, registerOutputs_170__13, 
         registerOutputs_170__12, registerOutputs_170__11, 
         registerOutputs_170__10, registerOutputs_170__9, registerOutputs_170__8, 
         registerOutputs_170__7, registerOutputs_170__6, registerOutputs_170__5, 
         registerOutputs_170__4, registerOutputs_170__3, registerOutputs_170__2, 
         registerOutputs_170__1, registerOutputs_170__0, registerOutputs_171__15, 
         registerOutputs_171__14, registerOutputs_171__13, 
         registerOutputs_171__12, registerOutputs_171__11, 
         registerOutputs_171__10, registerOutputs_171__9, registerOutputs_171__8, 
         registerOutputs_171__7, registerOutputs_171__6, registerOutputs_171__5, 
         registerOutputs_171__4, registerOutputs_171__3, registerOutputs_171__2, 
         registerOutputs_171__1, registerOutputs_171__0, registerOutputs_172__15, 
         registerOutputs_172__14, registerOutputs_172__13, 
         registerOutputs_172__12, registerOutputs_172__11, 
         registerOutputs_172__10, registerOutputs_172__9, registerOutputs_172__8, 
         registerOutputs_172__7, registerOutputs_172__6, registerOutputs_172__5, 
         registerOutputs_172__4, registerOutputs_172__3, registerOutputs_172__2, 
         registerOutputs_172__1, registerOutputs_172__0, registerOutputs_173__15, 
         registerOutputs_173__14, registerOutputs_173__13, 
         registerOutputs_173__12, registerOutputs_173__11, 
         registerOutputs_173__10, registerOutputs_173__9, registerOutputs_173__8, 
         registerOutputs_173__7, registerOutputs_173__6, registerOutputs_173__5, 
         registerOutputs_173__4, registerOutputs_173__3, registerOutputs_173__2, 
         registerOutputs_173__1, registerOutputs_173__0, registerOutputs_174__15, 
         registerOutputs_174__14, registerOutputs_174__13, 
         registerOutputs_174__12, registerOutputs_174__11, 
         registerOutputs_174__10, registerOutputs_174__9, registerOutputs_174__8, 
         registerOutputs_174__7, registerOutputs_174__6, registerOutputs_174__5, 
         registerOutputs_174__4, registerOutputs_174__3, registerOutputs_174__2, 
         registerOutputs_174__1, registerOutputs_174__0, registerOutputs_175__15, 
         registerOutputs_175__14, registerOutputs_175__13, 
         registerOutputs_175__12, registerOutputs_175__11, 
         registerOutputs_175__10, registerOutputs_175__9, registerOutputs_175__8, 
         registerOutputs_175__7, registerOutputs_175__6, registerOutputs_175__5, 
         registerOutputs_175__4, registerOutputs_175__3, registerOutputs_175__2, 
         registerOutputs_175__1, registerOutputs_175__0, registerOutputs_176__15, 
         registerOutputs_176__14, registerOutputs_176__13, 
         registerOutputs_176__12, registerOutputs_176__11, 
         registerOutputs_176__10, registerOutputs_176__9, registerOutputs_176__8, 
         registerOutputs_176__7, registerOutputs_176__6, registerOutputs_176__5, 
         registerOutputs_176__4, registerOutputs_176__3, registerOutputs_176__2, 
         registerOutputs_176__1, registerOutputs_176__0, registerOutputs_177__15, 
         registerOutputs_177__14, registerOutputs_177__13, 
         registerOutputs_177__12, registerOutputs_177__11, 
         registerOutputs_177__10, registerOutputs_177__9, registerOutputs_177__8, 
         registerOutputs_177__7, registerOutputs_177__6, registerOutputs_177__5, 
         registerOutputs_177__4, registerOutputs_177__3, registerOutputs_177__2, 
         registerOutputs_177__1, registerOutputs_177__0, registerOutputs_178__15, 
         registerOutputs_178__14, registerOutputs_178__13, 
         registerOutputs_178__12, registerOutputs_178__11, 
         registerOutputs_178__10, registerOutputs_178__9, registerOutputs_178__8, 
         registerOutputs_178__7, registerOutputs_178__6, registerOutputs_178__5, 
         registerOutputs_178__4, registerOutputs_178__3, registerOutputs_178__2, 
         registerOutputs_178__1, registerOutputs_178__0, registerOutputs_179__15, 
         registerOutputs_179__14, registerOutputs_179__13, 
         registerOutputs_179__12, registerOutputs_179__11, 
         registerOutputs_179__10, registerOutputs_179__9, registerOutputs_179__8, 
         registerOutputs_179__7, registerOutputs_179__6, registerOutputs_179__5, 
         registerOutputs_179__4, registerOutputs_179__3, registerOutputs_179__2, 
         registerOutputs_179__1, registerOutputs_179__0, registerOutputs_180__15, 
         registerOutputs_180__14, registerOutputs_180__13, 
         registerOutputs_180__12, registerOutputs_180__11, 
         registerOutputs_180__10, registerOutputs_180__9, registerOutputs_180__8, 
         registerOutputs_180__7, registerOutputs_180__6, registerOutputs_180__5, 
         registerOutputs_180__4, registerOutputs_180__3, registerOutputs_180__2, 
         registerOutputs_180__1, registerOutputs_180__0, registerOutputs_181__15, 
         registerOutputs_181__14, registerOutputs_181__13, 
         registerOutputs_181__12, registerOutputs_181__11, 
         registerOutputs_181__10, registerOutputs_181__9, registerOutputs_181__8, 
         registerOutputs_181__7, registerOutputs_181__6, registerOutputs_181__5, 
         registerOutputs_181__4, registerOutputs_181__3, registerOutputs_181__2, 
         registerOutputs_181__1, registerOutputs_181__0, registerOutputs_182__15, 
         registerOutputs_182__14, registerOutputs_182__13, 
         registerOutputs_182__12, registerOutputs_182__11, 
         registerOutputs_182__10, registerOutputs_182__9, registerOutputs_182__8, 
         registerOutputs_182__7, registerOutputs_182__6, registerOutputs_182__5, 
         registerOutputs_182__4, registerOutputs_182__3, registerOutputs_182__2, 
         registerOutputs_182__1, registerOutputs_182__0, registerOutputs_183__15, 
         registerOutputs_183__14, registerOutputs_183__13, 
         registerOutputs_183__12, registerOutputs_183__11, 
         registerOutputs_183__10, registerOutputs_183__9, registerOutputs_183__8, 
         registerOutputs_183__7, registerOutputs_183__6, registerOutputs_183__5, 
         registerOutputs_183__4, registerOutputs_183__3, registerOutputs_183__2, 
         registerOutputs_183__1, registerOutputs_183__0, registerOutputs_184__15, 
         registerOutputs_184__14, registerOutputs_184__13, 
         registerOutputs_184__12, registerOutputs_184__11, 
         registerOutputs_184__10, registerOutputs_184__9, registerOutputs_184__8, 
         registerOutputs_184__7, registerOutputs_184__6, registerOutputs_184__5, 
         registerOutputs_184__4, registerOutputs_184__3, registerOutputs_184__2, 
         registerOutputs_184__1, registerOutputs_184__0, registerOutputs_185__15, 
         registerOutputs_185__14, registerOutputs_185__13, 
         registerOutputs_185__12, registerOutputs_185__11, 
         registerOutputs_185__10, registerOutputs_185__9, registerOutputs_185__8, 
         registerOutputs_185__7, registerOutputs_185__6, registerOutputs_185__5, 
         registerOutputs_185__4, registerOutputs_185__3, registerOutputs_185__2, 
         registerOutputs_185__1, registerOutputs_185__0, registerOutputs_186__15, 
         registerOutputs_186__14, registerOutputs_186__13, 
         registerOutputs_186__12, registerOutputs_186__11, 
         registerOutputs_186__10, registerOutputs_186__9, registerOutputs_186__8, 
         registerOutputs_186__7, registerOutputs_186__6, registerOutputs_186__5, 
         registerOutputs_186__4, registerOutputs_186__3, registerOutputs_186__2, 
         registerOutputs_186__1, registerOutputs_186__0, registerOutputs_187__15, 
         registerOutputs_187__14, registerOutputs_187__13, 
         registerOutputs_187__12, registerOutputs_187__11, 
         registerOutputs_187__10, registerOutputs_187__9, registerOutputs_187__8, 
         registerOutputs_187__7, registerOutputs_187__6, registerOutputs_187__5, 
         registerOutputs_187__4, registerOutputs_187__3, registerOutputs_187__2, 
         registerOutputs_187__1, registerOutputs_187__0, registerOutputs_188__15, 
         registerOutputs_188__14, registerOutputs_188__13, 
         registerOutputs_188__12, registerOutputs_188__11, 
         registerOutputs_188__10, registerOutputs_188__9, registerOutputs_188__8, 
         registerOutputs_188__7, registerOutputs_188__6, registerOutputs_188__5, 
         registerOutputs_188__4, registerOutputs_188__3, registerOutputs_188__2, 
         registerOutputs_188__1, registerOutputs_188__0, registerOutputs_189__15, 
         registerOutputs_189__14, registerOutputs_189__13, 
         registerOutputs_189__12, registerOutputs_189__11, 
         registerOutputs_189__10, registerOutputs_189__9, registerOutputs_189__8, 
         registerOutputs_189__7, registerOutputs_189__6, registerOutputs_189__5, 
         registerOutputs_189__4, registerOutputs_189__3, registerOutputs_189__2, 
         registerOutputs_189__1, registerOutputs_189__0, registerOutputs_190__15, 
         registerOutputs_190__14, registerOutputs_190__13, 
         registerOutputs_190__12, registerOutputs_190__11, 
         registerOutputs_190__10, registerOutputs_190__9, registerOutputs_190__8, 
         registerOutputs_190__7, registerOutputs_190__6, registerOutputs_190__5, 
         registerOutputs_190__4, registerOutputs_190__3, registerOutputs_190__2, 
         registerOutputs_190__1, registerOutputs_190__0, registerOutputs_191__15, 
         registerOutputs_191__14, registerOutputs_191__13, 
         registerOutputs_191__12, registerOutputs_191__11, 
         registerOutputs_191__10, registerOutputs_191__9, registerOutputs_191__8, 
         registerOutputs_191__7, registerOutputs_191__6, registerOutputs_191__5, 
         registerOutputs_191__4, registerOutputs_191__3, registerOutputs_191__2, 
         registerOutputs_191__1, registerOutputs_191__0, registerOutputs_192__15, 
         registerOutputs_192__14, registerOutputs_192__13, 
         registerOutputs_192__12, registerOutputs_192__11, 
         registerOutputs_192__10, registerOutputs_192__9, registerOutputs_192__8, 
         registerOutputs_192__7, registerOutputs_192__6, registerOutputs_192__5, 
         registerOutputs_192__4, registerOutputs_192__3, registerOutputs_192__2, 
         registerOutputs_192__1, registerOutputs_192__0, registerOutputs_193__15, 
         registerOutputs_193__14, registerOutputs_193__13, 
         registerOutputs_193__12, registerOutputs_193__11, 
         registerOutputs_193__10, registerOutputs_193__9, registerOutputs_193__8, 
         registerOutputs_193__7, registerOutputs_193__6, registerOutputs_193__5, 
         registerOutputs_193__4, registerOutputs_193__3, registerOutputs_193__2, 
         registerOutputs_193__1, registerOutputs_193__0, registerOutputs_194__15, 
         registerOutputs_194__14, registerOutputs_194__13, 
         registerOutputs_194__12, registerOutputs_194__11, 
         registerOutputs_194__10, registerOutputs_194__9, registerOutputs_194__8, 
         registerOutputs_194__7, registerOutputs_194__6, registerOutputs_194__5, 
         registerOutputs_194__4, registerOutputs_194__3, registerOutputs_194__2, 
         registerOutputs_194__1, registerOutputs_194__0, registerOutputs_195__15, 
         registerOutputs_195__14, registerOutputs_195__13, 
         registerOutputs_195__12, registerOutputs_195__11, 
         registerOutputs_195__10, registerOutputs_195__9, registerOutputs_195__8, 
         registerOutputs_195__7, registerOutputs_195__6, registerOutputs_195__5, 
         registerOutputs_195__4, registerOutputs_195__3, registerOutputs_195__2, 
         registerOutputs_195__1, registerOutputs_195__0, registerOutputs_196__15, 
         registerOutputs_196__14, registerOutputs_196__13, 
         registerOutputs_196__12, registerOutputs_196__11, 
         registerOutputs_196__10, registerOutputs_196__9, registerOutputs_196__8, 
         registerOutputs_196__7, registerOutputs_196__6, registerOutputs_196__5, 
         registerOutputs_196__4, registerOutputs_196__3, registerOutputs_196__2, 
         registerOutputs_196__1, registerOutputs_196__0, registerOutputs_197__15, 
         registerOutputs_197__14, registerOutputs_197__13, 
         registerOutputs_197__12, registerOutputs_197__11, 
         registerOutputs_197__10, registerOutputs_197__9, registerOutputs_197__8, 
         registerOutputs_197__7, registerOutputs_197__6, registerOutputs_197__5, 
         registerOutputs_197__4, registerOutputs_197__3, registerOutputs_197__2, 
         registerOutputs_197__1, registerOutputs_197__0, registerOutputs_198__15, 
         registerOutputs_198__14, registerOutputs_198__13, 
         registerOutputs_198__12, registerOutputs_198__11, 
         registerOutputs_198__10, registerOutputs_198__9, registerOutputs_198__8, 
         registerOutputs_198__7, registerOutputs_198__6, registerOutputs_198__5, 
         registerOutputs_198__4, registerOutputs_198__3, registerOutputs_198__2, 
         registerOutputs_198__1, registerOutputs_198__0, registerOutputs_199__15, 
         registerOutputs_199__14, registerOutputs_199__13, 
         registerOutputs_199__12, registerOutputs_199__11, 
         registerOutputs_199__10, registerOutputs_199__9, registerOutputs_199__8, 
         registerOutputs_199__7, registerOutputs_199__6, registerOutputs_199__5, 
         registerOutputs_199__4, registerOutputs_199__3, registerOutputs_199__2, 
         registerOutputs_199__1, registerOutputs_199__0, registerOutputs_200__15, 
         registerOutputs_200__14, registerOutputs_200__13, 
         registerOutputs_200__12, registerOutputs_200__11, 
         registerOutputs_200__10, registerOutputs_200__9, registerOutputs_200__8, 
         registerOutputs_200__7, registerOutputs_200__6, registerOutputs_200__5, 
         registerOutputs_200__4, registerOutputs_200__3, registerOutputs_200__2, 
         registerOutputs_200__1, registerOutputs_200__0, registerOutputs_201__15, 
         registerOutputs_201__14, registerOutputs_201__13, 
         registerOutputs_201__12, registerOutputs_201__11, 
         registerOutputs_201__10, registerOutputs_201__9, registerOutputs_201__8, 
         registerOutputs_201__7, registerOutputs_201__6, registerOutputs_201__5, 
         registerOutputs_201__4, registerOutputs_201__3, registerOutputs_201__2, 
         registerOutputs_201__1, registerOutputs_201__0, registerOutputs_202__15, 
         registerOutputs_202__14, registerOutputs_202__13, 
         registerOutputs_202__12, registerOutputs_202__11, 
         registerOutputs_202__10, registerOutputs_202__9, registerOutputs_202__8, 
         registerOutputs_202__7, registerOutputs_202__6, registerOutputs_202__5, 
         registerOutputs_202__4, registerOutputs_202__3, registerOutputs_202__2, 
         registerOutputs_202__1, registerOutputs_202__0, registerOutputs_203__15, 
         registerOutputs_203__14, registerOutputs_203__13, 
         registerOutputs_203__12, registerOutputs_203__11, 
         registerOutputs_203__10, registerOutputs_203__9, registerOutputs_203__8, 
         registerOutputs_203__7, registerOutputs_203__6, registerOutputs_203__5, 
         registerOutputs_203__4, registerOutputs_203__3, registerOutputs_203__2, 
         registerOutputs_203__1, registerOutputs_203__0, registerOutputs_204__15, 
         registerOutputs_204__14, registerOutputs_204__13, 
         registerOutputs_204__12, registerOutputs_204__11, 
         registerOutputs_204__10, registerOutputs_204__9, registerOutputs_204__8, 
         registerOutputs_204__7, registerOutputs_204__6, registerOutputs_204__5, 
         registerOutputs_204__4, registerOutputs_204__3, registerOutputs_204__2, 
         registerOutputs_204__1, registerOutputs_204__0, registerOutputs_205__15, 
         registerOutputs_205__14, registerOutputs_205__13, 
         registerOutputs_205__12, registerOutputs_205__11, 
         registerOutputs_205__10, registerOutputs_205__9, registerOutputs_205__8, 
         registerOutputs_205__7, registerOutputs_205__6, registerOutputs_205__5, 
         registerOutputs_205__4, registerOutputs_205__3, registerOutputs_205__2, 
         registerOutputs_205__1, registerOutputs_205__0, registerOutputs_206__15, 
         registerOutputs_206__14, registerOutputs_206__13, 
         registerOutputs_206__12, registerOutputs_206__11, 
         registerOutputs_206__10, registerOutputs_206__9, registerOutputs_206__8, 
         registerOutputs_206__7, registerOutputs_206__6, registerOutputs_206__5, 
         registerOutputs_206__4, registerOutputs_206__3, registerOutputs_206__2, 
         registerOutputs_206__1, registerOutputs_206__0, registerOutputs_207__15, 
         registerOutputs_207__14, registerOutputs_207__13, 
         registerOutputs_207__12, registerOutputs_207__11, 
         registerOutputs_207__10, registerOutputs_207__9, registerOutputs_207__8, 
         registerOutputs_207__7, registerOutputs_207__6, registerOutputs_207__5, 
         registerOutputs_207__4, registerOutputs_207__3, registerOutputs_207__2, 
         registerOutputs_207__1, registerOutputs_207__0, registerOutputs_208__15, 
         registerOutputs_208__14, registerOutputs_208__13, 
         registerOutputs_208__12, registerOutputs_208__11, 
         registerOutputs_208__10, registerOutputs_208__9, registerOutputs_208__8, 
         registerOutputs_208__7, registerOutputs_208__6, registerOutputs_208__5, 
         registerOutputs_208__4, registerOutputs_208__3, registerOutputs_208__2, 
         registerOutputs_208__1, registerOutputs_208__0, registerOutputs_209__15, 
         registerOutputs_209__14, registerOutputs_209__13, 
         registerOutputs_209__12, registerOutputs_209__11, 
         registerOutputs_209__10, registerOutputs_209__9, registerOutputs_209__8, 
         registerOutputs_209__7, registerOutputs_209__6, registerOutputs_209__5, 
         registerOutputs_209__4, registerOutputs_209__3, registerOutputs_209__2, 
         registerOutputs_209__1, registerOutputs_209__0, registerOutputs_210__15, 
         registerOutputs_210__14, registerOutputs_210__13, 
         registerOutputs_210__12, registerOutputs_210__11, 
         registerOutputs_210__10, registerOutputs_210__9, registerOutputs_210__8, 
         registerOutputs_210__7, registerOutputs_210__6, registerOutputs_210__5, 
         registerOutputs_210__4, registerOutputs_210__3, registerOutputs_210__2, 
         registerOutputs_210__1, registerOutputs_210__0, registerOutputs_211__15, 
         registerOutputs_211__14, registerOutputs_211__13, 
         registerOutputs_211__12, registerOutputs_211__11, 
         registerOutputs_211__10, registerOutputs_211__9, registerOutputs_211__8, 
         registerOutputs_211__7, registerOutputs_211__6, registerOutputs_211__5, 
         registerOutputs_211__4, registerOutputs_211__3, registerOutputs_211__2, 
         registerOutputs_211__1, registerOutputs_211__0, registerOutputs_212__15, 
         registerOutputs_212__14, registerOutputs_212__13, 
         registerOutputs_212__12, registerOutputs_212__11, 
         registerOutputs_212__10, registerOutputs_212__9, registerOutputs_212__8, 
         registerOutputs_212__7, registerOutputs_212__6, registerOutputs_212__5, 
         registerOutputs_212__4, registerOutputs_212__3, registerOutputs_212__2, 
         registerOutputs_212__1, registerOutputs_212__0, registerOutputs_213__15, 
         registerOutputs_213__14, registerOutputs_213__13, 
         registerOutputs_213__12, registerOutputs_213__11, 
         registerOutputs_213__10, registerOutputs_213__9, registerOutputs_213__8, 
         registerOutputs_213__7, registerOutputs_213__6, registerOutputs_213__5, 
         registerOutputs_213__4, registerOutputs_213__3, registerOutputs_213__2, 
         registerOutputs_213__1, registerOutputs_213__0, registerOutputs_214__15, 
         registerOutputs_214__14, registerOutputs_214__13, 
         registerOutputs_214__12, registerOutputs_214__11, 
         registerOutputs_214__10, registerOutputs_214__9, registerOutputs_214__8, 
         registerOutputs_214__7, registerOutputs_214__6, registerOutputs_214__5, 
         registerOutputs_214__4, registerOutputs_214__3, registerOutputs_214__2, 
         registerOutputs_214__1, registerOutputs_214__0, registerOutputs_215__15, 
         registerOutputs_215__14, registerOutputs_215__13, 
         registerOutputs_215__12, registerOutputs_215__11, 
         registerOutputs_215__10, registerOutputs_215__9, registerOutputs_215__8, 
         registerOutputs_215__7, registerOutputs_215__6, registerOutputs_215__5, 
         registerOutputs_215__4, registerOutputs_215__3, registerOutputs_215__2, 
         registerOutputs_215__1, registerOutputs_215__0, registerOutputs_216__15, 
         registerOutputs_216__14, registerOutputs_216__13, 
         registerOutputs_216__12, registerOutputs_216__11, 
         registerOutputs_216__10, registerOutputs_216__9, registerOutputs_216__8, 
         registerOutputs_216__7, registerOutputs_216__6, registerOutputs_216__5, 
         registerOutputs_216__4, registerOutputs_216__3, registerOutputs_216__2, 
         registerOutputs_216__1, registerOutputs_216__0, registerOutputs_217__15, 
         registerOutputs_217__14, registerOutputs_217__13, 
         registerOutputs_217__12, registerOutputs_217__11, 
         registerOutputs_217__10, registerOutputs_217__9, registerOutputs_217__8, 
         registerOutputs_217__7, registerOutputs_217__6, registerOutputs_217__5, 
         registerOutputs_217__4, registerOutputs_217__3, registerOutputs_217__2, 
         registerOutputs_217__1, registerOutputs_217__0, registerOutputs_218__15, 
         registerOutputs_218__14, registerOutputs_218__13, 
         registerOutputs_218__12, registerOutputs_218__11, 
         registerOutputs_218__10, registerOutputs_218__9, registerOutputs_218__8, 
         registerOutputs_218__7, registerOutputs_218__6, registerOutputs_218__5, 
         registerOutputs_218__4, registerOutputs_218__3, registerOutputs_218__2, 
         registerOutputs_218__1, registerOutputs_218__0, registerOutputs_219__15, 
         registerOutputs_219__14, registerOutputs_219__13, 
         registerOutputs_219__12, registerOutputs_219__11, 
         registerOutputs_219__10, registerOutputs_219__9, registerOutputs_219__8, 
         registerOutputs_219__7, registerOutputs_219__6, registerOutputs_219__5, 
         registerOutputs_219__4, registerOutputs_219__3, registerOutputs_219__2, 
         registerOutputs_219__1, registerOutputs_219__0, registerOutputs_220__15, 
         registerOutputs_220__14, registerOutputs_220__13, 
         registerOutputs_220__12, registerOutputs_220__11, 
         registerOutputs_220__10, registerOutputs_220__9, registerOutputs_220__8, 
         registerOutputs_220__7, registerOutputs_220__6, registerOutputs_220__5, 
         registerOutputs_220__4, registerOutputs_220__3, registerOutputs_220__2, 
         registerOutputs_220__1, registerOutputs_220__0, registerOutputs_221__15, 
         registerOutputs_221__14, registerOutputs_221__13, 
         registerOutputs_221__12, registerOutputs_221__11, 
         registerOutputs_221__10, registerOutputs_221__9, registerOutputs_221__8, 
         registerOutputs_221__7, registerOutputs_221__6, registerOutputs_221__5, 
         registerOutputs_221__4, registerOutputs_221__3, registerOutputs_221__2, 
         registerOutputs_221__1, registerOutputs_221__0, registerOutputs_222__15, 
         registerOutputs_222__14, registerOutputs_222__13, 
         registerOutputs_222__12, registerOutputs_222__11, 
         registerOutputs_222__10, registerOutputs_222__9, registerOutputs_222__8, 
         registerOutputs_222__7, registerOutputs_222__6, registerOutputs_222__5, 
         registerOutputs_222__4, registerOutputs_222__3, registerOutputs_222__2, 
         registerOutputs_222__1, registerOutputs_222__0, registerOutputs_223__15, 
         registerOutputs_223__14, registerOutputs_223__13, 
         registerOutputs_223__12, registerOutputs_223__11, 
         registerOutputs_223__10, registerOutputs_223__9, registerOutputs_223__8, 
         registerOutputs_223__7, registerOutputs_223__6, registerOutputs_223__5, 
         registerOutputs_223__4, registerOutputs_223__3, registerOutputs_223__2, 
         registerOutputs_223__1, registerOutputs_223__0, registerOutputs_224__15, 
         registerOutputs_224__14, registerOutputs_224__13, 
         registerOutputs_224__12, registerOutputs_224__11, 
         registerOutputs_224__10, registerOutputs_224__9, registerOutputs_224__8, 
         registerOutputs_224__7, registerOutputs_224__6, registerOutputs_224__5, 
         registerOutputs_224__4, registerOutputs_224__3, registerOutputs_224__2, 
         registerOutputs_224__1, registerOutputs_224__0, registerOutputs_225__15, 
         registerOutputs_225__14, registerOutputs_225__13, 
         registerOutputs_225__12, registerOutputs_225__11, 
         registerOutputs_225__10, registerOutputs_225__9, registerOutputs_225__8, 
         registerOutputs_225__7, registerOutputs_225__6, registerOutputs_225__5, 
         registerOutputs_225__4, registerOutputs_225__3, registerOutputs_225__2, 
         registerOutputs_225__1, registerOutputs_225__0, registerOutputs_226__15, 
         registerOutputs_226__14, registerOutputs_226__13, 
         registerOutputs_226__12, registerOutputs_226__11, 
         registerOutputs_226__10, registerOutputs_226__9, registerOutputs_226__8, 
         registerOutputs_226__7, registerOutputs_226__6, registerOutputs_226__5, 
         registerOutputs_226__4, registerOutputs_226__3, registerOutputs_226__2, 
         registerOutputs_226__1, registerOutputs_226__0, registerOutputs_227__15, 
         registerOutputs_227__14, registerOutputs_227__13, 
         registerOutputs_227__12, registerOutputs_227__11, 
         registerOutputs_227__10, registerOutputs_227__9, registerOutputs_227__8, 
         registerOutputs_227__7, registerOutputs_227__6, registerOutputs_227__5, 
         registerOutputs_227__4, registerOutputs_227__3, registerOutputs_227__2, 
         registerOutputs_227__1, registerOutputs_227__0, registerOutputs_228__15, 
         registerOutputs_228__14, registerOutputs_228__13, 
         registerOutputs_228__12, registerOutputs_228__11, 
         registerOutputs_228__10, registerOutputs_228__9, registerOutputs_228__8, 
         registerOutputs_228__7, registerOutputs_228__6, registerOutputs_228__5, 
         registerOutputs_228__4, registerOutputs_228__3, registerOutputs_228__2, 
         registerOutputs_228__1, registerOutputs_228__0, registerOutputs_229__15, 
         registerOutputs_229__14, registerOutputs_229__13, 
         registerOutputs_229__12, registerOutputs_229__11, 
         registerOutputs_229__10, registerOutputs_229__9, registerOutputs_229__8, 
         registerOutputs_229__7, registerOutputs_229__6, registerOutputs_229__5, 
         registerOutputs_229__4, registerOutputs_229__3, registerOutputs_229__2, 
         registerOutputs_229__1, registerOutputs_229__0, registerOutputs_230__15, 
         registerOutputs_230__14, registerOutputs_230__13, 
         registerOutputs_230__12, registerOutputs_230__11, 
         registerOutputs_230__10, registerOutputs_230__9, registerOutputs_230__8, 
         registerOutputs_230__7, registerOutputs_230__6, registerOutputs_230__5, 
         registerOutputs_230__4, registerOutputs_230__3, registerOutputs_230__2, 
         registerOutputs_230__1, registerOutputs_230__0, registerOutputs_231__15, 
         registerOutputs_231__14, registerOutputs_231__13, 
         registerOutputs_231__12, registerOutputs_231__11, 
         registerOutputs_231__10, registerOutputs_231__9, registerOutputs_231__8, 
         registerOutputs_231__7, registerOutputs_231__6, registerOutputs_231__5, 
         registerOutputs_231__4, registerOutputs_231__3, registerOutputs_231__2, 
         registerOutputs_231__1, registerOutputs_231__0, registerOutputs_232__15, 
         registerOutputs_232__14, registerOutputs_232__13, 
         registerOutputs_232__12, registerOutputs_232__11, 
         registerOutputs_232__10, registerOutputs_232__9, registerOutputs_232__8, 
         registerOutputs_232__7, registerOutputs_232__6, registerOutputs_232__5, 
         registerOutputs_232__4, registerOutputs_232__3, registerOutputs_232__2, 
         registerOutputs_232__1, registerOutputs_232__0, registerOutputs_233__15, 
         registerOutputs_233__14, registerOutputs_233__13, 
         registerOutputs_233__12, registerOutputs_233__11, 
         registerOutputs_233__10, registerOutputs_233__9, registerOutputs_233__8, 
         registerOutputs_233__7, registerOutputs_233__6, registerOutputs_233__5, 
         registerOutputs_233__4, registerOutputs_233__3, registerOutputs_233__2, 
         registerOutputs_233__1, registerOutputs_233__0, registerOutputs_234__15, 
         registerOutputs_234__14, registerOutputs_234__13, 
         registerOutputs_234__12, registerOutputs_234__11, 
         registerOutputs_234__10, registerOutputs_234__9, registerOutputs_234__8, 
         registerOutputs_234__7, registerOutputs_234__6, registerOutputs_234__5, 
         registerOutputs_234__4, registerOutputs_234__3, registerOutputs_234__2, 
         registerOutputs_234__1, registerOutputs_234__0, registerOutputs_235__15, 
         registerOutputs_235__14, registerOutputs_235__13, 
         registerOutputs_235__12, registerOutputs_235__11, 
         registerOutputs_235__10, registerOutputs_235__9, registerOutputs_235__8, 
         registerOutputs_235__7, registerOutputs_235__6, registerOutputs_235__5, 
         registerOutputs_235__4, registerOutputs_235__3, registerOutputs_235__2, 
         registerOutputs_235__1, registerOutputs_235__0, registerOutputs_236__15, 
         registerOutputs_236__14, registerOutputs_236__13, 
         registerOutputs_236__12, registerOutputs_236__11, 
         registerOutputs_236__10, registerOutputs_236__9, registerOutputs_236__8, 
         registerOutputs_236__7, registerOutputs_236__6, registerOutputs_236__5, 
         registerOutputs_236__4, registerOutputs_236__3, registerOutputs_236__2, 
         registerOutputs_236__1, registerOutputs_236__0, registerOutputs_237__15, 
         registerOutputs_237__14, registerOutputs_237__13, 
         registerOutputs_237__12, registerOutputs_237__11, 
         registerOutputs_237__10, registerOutputs_237__9, registerOutputs_237__8, 
         registerOutputs_237__7, registerOutputs_237__6, registerOutputs_237__5, 
         registerOutputs_237__4, registerOutputs_237__3, registerOutputs_237__2, 
         registerOutputs_237__1, registerOutputs_237__0, registerOutputs_238__15, 
         registerOutputs_238__14, registerOutputs_238__13, 
         registerOutputs_238__12, registerOutputs_238__11, 
         registerOutputs_238__10, registerOutputs_238__9, registerOutputs_238__8, 
         registerOutputs_238__7, registerOutputs_238__6, registerOutputs_238__5, 
         registerOutputs_238__4, registerOutputs_238__3, registerOutputs_238__2, 
         registerOutputs_238__1, registerOutputs_238__0, registerOutputs_239__15, 
         registerOutputs_239__14, registerOutputs_239__13, 
         registerOutputs_239__12, registerOutputs_239__11, 
         registerOutputs_239__10, registerOutputs_239__9, registerOutputs_239__8, 
         registerOutputs_239__7, registerOutputs_239__6, registerOutputs_239__5, 
         registerOutputs_239__4, registerOutputs_239__3, registerOutputs_239__2, 
         registerOutputs_239__1, registerOutputs_239__0, registerOutputs_240__15, 
         registerOutputs_240__14, registerOutputs_240__13, 
         registerOutputs_240__12, registerOutputs_240__11, 
         registerOutputs_240__10, registerOutputs_240__9, registerOutputs_240__8, 
         registerOutputs_240__7, registerOutputs_240__6, registerOutputs_240__5, 
         registerOutputs_240__4, registerOutputs_240__3, registerOutputs_240__2, 
         registerOutputs_240__1, registerOutputs_240__0, registerOutputs_241__15, 
         registerOutputs_241__14, registerOutputs_241__13, 
         registerOutputs_241__12, registerOutputs_241__11, 
         registerOutputs_241__10, registerOutputs_241__9, registerOutputs_241__8, 
         registerOutputs_241__7, registerOutputs_241__6, registerOutputs_241__5, 
         registerOutputs_241__4, registerOutputs_241__3, registerOutputs_241__2, 
         registerOutputs_241__1, registerOutputs_241__0, registerOutputs_242__15, 
         registerOutputs_242__14, registerOutputs_242__13, 
         registerOutputs_242__12, registerOutputs_242__11, 
         registerOutputs_242__10, registerOutputs_242__9, registerOutputs_242__8, 
         registerOutputs_242__7, registerOutputs_242__6, registerOutputs_242__5, 
         registerOutputs_242__4, registerOutputs_242__3, registerOutputs_242__2, 
         registerOutputs_242__1, registerOutputs_242__0, registerOutputs_243__15, 
         registerOutputs_243__14, registerOutputs_243__13, 
         registerOutputs_243__12, registerOutputs_243__11, 
         registerOutputs_243__10, registerOutputs_243__9, registerOutputs_243__8, 
         registerOutputs_243__7, registerOutputs_243__6, registerOutputs_243__5, 
         registerOutputs_243__4, registerOutputs_243__3, registerOutputs_243__2, 
         registerOutputs_243__1, registerOutputs_243__0, registerOutputs_244__15, 
         registerOutputs_244__14, registerOutputs_244__13, 
         registerOutputs_244__12, registerOutputs_244__11, 
         registerOutputs_244__10, registerOutputs_244__9, registerOutputs_244__8, 
         registerOutputs_244__7, registerOutputs_244__6, registerOutputs_244__5, 
         registerOutputs_244__4, registerOutputs_244__3, registerOutputs_244__2, 
         registerOutputs_244__1, registerOutputs_244__0, registerOutputs_245__15, 
         registerOutputs_245__14, registerOutputs_245__13, 
         registerOutputs_245__12, registerOutputs_245__11, 
         registerOutputs_245__10, registerOutputs_245__9, registerOutputs_245__8, 
         registerOutputs_245__7, registerOutputs_245__6, registerOutputs_245__5, 
         registerOutputs_245__4, registerOutputs_245__3, registerOutputs_245__2, 
         registerOutputs_245__1, registerOutputs_245__0, registerOutputs_246__15, 
         registerOutputs_246__14, registerOutputs_246__13, 
         registerOutputs_246__12, registerOutputs_246__11, 
         registerOutputs_246__10, registerOutputs_246__9, registerOutputs_246__8, 
         registerOutputs_246__7, registerOutputs_246__6, registerOutputs_246__5, 
         registerOutputs_246__4, registerOutputs_246__3, registerOutputs_246__2, 
         registerOutputs_246__1, registerOutputs_246__0, registerOutputs_247__15, 
         registerOutputs_247__14, registerOutputs_247__13, 
         registerOutputs_247__12, registerOutputs_247__11, 
         registerOutputs_247__10, registerOutputs_247__9, registerOutputs_247__8, 
         registerOutputs_247__7, registerOutputs_247__6, registerOutputs_247__5, 
         registerOutputs_247__4, registerOutputs_247__3, registerOutputs_247__2, 
         registerOutputs_247__1, registerOutputs_247__0, registerOutputs_248__15, 
         registerOutputs_248__14, registerOutputs_248__13, 
         registerOutputs_248__12, registerOutputs_248__11, 
         registerOutputs_248__10, registerOutputs_248__9, registerOutputs_248__8, 
         registerOutputs_248__7, registerOutputs_248__6, registerOutputs_248__5, 
         registerOutputs_248__4, registerOutputs_248__3, registerOutputs_248__2, 
         registerOutputs_248__1, registerOutputs_248__0, registerOutputs_249__15, 
         registerOutputs_249__14, registerOutputs_249__13, 
         registerOutputs_249__12, registerOutputs_249__11, 
         registerOutputs_249__10, registerOutputs_249__9, registerOutputs_249__8, 
         registerOutputs_249__7, registerOutputs_249__6, registerOutputs_249__5, 
         registerOutputs_249__4, registerOutputs_249__3, registerOutputs_249__2, 
         registerOutputs_249__1, registerOutputs_249__0, registerOutputs_250__15, 
         registerOutputs_250__14, registerOutputs_250__13, 
         registerOutputs_250__12, registerOutputs_250__11, 
         registerOutputs_250__10, registerOutputs_250__9, registerOutputs_250__8, 
         registerOutputs_250__7, registerOutputs_250__6, registerOutputs_250__5, 
         registerOutputs_250__4, registerOutputs_250__3, registerOutputs_250__2, 
         registerOutputs_250__1, registerOutputs_250__0, registerOutputs_251__15, 
         registerOutputs_251__14, registerOutputs_251__13, 
         registerOutputs_251__12, registerOutputs_251__11, 
         registerOutputs_251__10, registerOutputs_251__9, registerOutputs_251__8, 
         registerOutputs_251__7, registerOutputs_251__6, registerOutputs_251__5, 
         registerOutputs_251__4, registerOutputs_251__3, registerOutputs_251__2, 
         registerOutputs_251__1, registerOutputs_251__0, registerOutputs_252__15, 
         registerOutputs_252__14, registerOutputs_252__13, 
         registerOutputs_252__12, registerOutputs_252__11, 
         registerOutputs_252__10, registerOutputs_252__9, registerOutputs_252__8, 
         registerOutputs_252__7, registerOutputs_252__6, registerOutputs_252__5, 
         registerOutputs_252__4, registerOutputs_252__3, registerOutputs_252__2, 
         registerOutputs_252__1, registerOutputs_252__0, registerOutputs_253__15, 
         registerOutputs_253__14, registerOutputs_253__13, 
         registerOutputs_253__12, registerOutputs_253__11, 
         registerOutputs_253__10, registerOutputs_253__9, registerOutputs_253__8, 
         registerOutputs_253__7, registerOutputs_253__6, registerOutputs_253__5, 
         registerOutputs_253__4, registerOutputs_253__3, registerOutputs_253__2, 
         registerOutputs_253__1, registerOutputs_253__0, registerOutputs_254__15, 
         registerOutputs_254__14, registerOutputs_254__13, 
         registerOutputs_254__12, registerOutputs_254__11, 
         registerOutputs_254__10, registerOutputs_254__9, registerOutputs_254__8, 
         registerOutputs_254__7, registerOutputs_254__6, registerOutputs_254__5, 
         registerOutputs_254__4, registerOutputs_254__3, registerOutputs_254__2, 
         registerOutputs_254__1, registerOutputs_254__0, registerOutputs_255__15, 
         registerOutputs_255__14, registerOutputs_255__13, 
         registerOutputs_255__12, registerOutputs_255__11, 
         registerOutputs_255__10, registerOutputs_255__9, registerOutputs_255__8, 
         registerOutputs_255__7, registerOutputs_255__6, registerOutputs_255__5, 
         registerOutputs_255__4, registerOutputs_255__3, registerOutputs_255__2, 
         registerOutputs_255__1, registerOutputs_255__0, registerOutputs_256__15, 
         registerOutputs_256__14, registerOutputs_256__13, 
         registerOutputs_256__12, registerOutputs_256__11, 
         registerOutputs_256__10, registerOutputs_256__9, registerOutputs_256__8, 
         registerOutputs_256__7, registerOutputs_256__6, registerOutputs_256__5, 
         registerOutputs_256__4, registerOutputs_256__3, registerOutputs_256__2, 
         registerOutputs_256__1, registerOutputs_256__0, registerOutputs_257__15, 
         registerOutputs_257__14, registerOutputs_257__13, 
         registerOutputs_257__12, registerOutputs_257__11, 
         registerOutputs_257__10, registerOutputs_257__9, registerOutputs_257__8, 
         registerOutputs_257__7, registerOutputs_257__6, registerOutputs_257__5, 
         registerOutputs_257__4, registerOutputs_257__3, registerOutputs_257__2, 
         registerOutputs_257__1, registerOutputs_257__0, registerOutputs_258__15, 
         registerOutputs_258__14, registerOutputs_258__13, 
         registerOutputs_258__12, registerOutputs_258__11, 
         registerOutputs_258__10, registerOutputs_258__9, registerOutputs_258__8, 
         registerOutputs_258__7, registerOutputs_258__6, registerOutputs_258__5, 
         registerOutputs_258__4, registerOutputs_258__3, registerOutputs_258__2, 
         registerOutputs_258__1, registerOutputs_258__0, registerOutputs_259__15, 
         registerOutputs_259__14, registerOutputs_259__13, 
         registerOutputs_259__12, registerOutputs_259__11, 
         registerOutputs_259__10, registerOutputs_259__9, registerOutputs_259__8, 
         registerOutputs_259__7, registerOutputs_259__6, registerOutputs_259__5, 
         registerOutputs_259__4, registerOutputs_259__3, registerOutputs_259__2, 
         registerOutputs_259__1, registerOutputs_259__0, registerOutputs_260__15, 
         registerOutputs_260__14, registerOutputs_260__13, 
         registerOutputs_260__12, registerOutputs_260__11, 
         registerOutputs_260__10, registerOutputs_260__9, registerOutputs_260__8, 
         registerOutputs_260__7, registerOutputs_260__6, registerOutputs_260__5, 
         registerOutputs_260__4, registerOutputs_260__3, registerOutputs_260__2, 
         registerOutputs_260__1, registerOutputs_260__0, registerOutputs_261__15, 
         registerOutputs_261__14, registerOutputs_261__13, 
         registerOutputs_261__12, registerOutputs_261__11, 
         registerOutputs_261__10, registerOutputs_261__9, registerOutputs_261__8, 
         registerOutputs_261__7, registerOutputs_261__6, registerOutputs_261__5, 
         registerOutputs_261__4, registerOutputs_261__3, registerOutputs_261__2, 
         registerOutputs_261__1, registerOutputs_261__0, registerOutputs_262__15, 
         registerOutputs_262__14, registerOutputs_262__13, 
         registerOutputs_262__12, registerOutputs_262__11, 
         registerOutputs_262__10, registerOutputs_262__9, registerOutputs_262__8, 
         registerOutputs_262__7, registerOutputs_262__6, registerOutputs_262__5, 
         registerOutputs_262__4, registerOutputs_262__3, registerOutputs_262__2, 
         registerOutputs_262__1, registerOutputs_262__0, registerOutputs_263__15, 
         registerOutputs_263__14, registerOutputs_263__13, 
         registerOutputs_263__12, registerOutputs_263__11, 
         registerOutputs_263__10, registerOutputs_263__9, registerOutputs_263__8, 
         registerOutputs_263__7, registerOutputs_263__6, registerOutputs_263__5, 
         registerOutputs_263__4, registerOutputs_263__3, registerOutputs_263__2, 
         registerOutputs_263__1, registerOutputs_263__0, registerOutputs_264__15, 
         registerOutputs_264__14, registerOutputs_264__13, 
         registerOutputs_264__12, registerOutputs_264__11, 
         registerOutputs_264__10, registerOutputs_264__9, registerOutputs_264__8, 
         registerOutputs_264__7, registerOutputs_264__6, registerOutputs_264__5, 
         registerOutputs_264__4, registerOutputs_264__3, registerOutputs_264__2, 
         registerOutputs_264__1, registerOutputs_264__0, registerOutputs_265__15, 
         registerOutputs_265__14, registerOutputs_265__13, 
         registerOutputs_265__12, registerOutputs_265__11, 
         registerOutputs_265__10, registerOutputs_265__9, registerOutputs_265__8, 
         registerOutputs_265__7, registerOutputs_265__6, registerOutputs_265__5, 
         registerOutputs_265__4, registerOutputs_265__3, registerOutputs_265__2, 
         registerOutputs_265__1, registerOutputs_265__0, registerOutputs_266__15, 
         registerOutputs_266__14, registerOutputs_266__13, 
         registerOutputs_266__12, registerOutputs_266__11, 
         registerOutputs_266__10, registerOutputs_266__9, registerOutputs_266__8, 
         registerOutputs_266__7, registerOutputs_266__6, registerOutputs_266__5, 
         registerOutputs_266__4, registerOutputs_266__3, registerOutputs_266__2, 
         registerOutputs_266__1, registerOutputs_266__0, registerOutputs_267__15, 
         registerOutputs_267__14, registerOutputs_267__13, 
         registerOutputs_267__12, registerOutputs_267__11, 
         registerOutputs_267__10, registerOutputs_267__9, registerOutputs_267__8, 
         registerOutputs_267__7, registerOutputs_267__6, registerOutputs_267__5, 
         registerOutputs_267__4, registerOutputs_267__3, registerOutputs_267__2, 
         registerOutputs_267__1, registerOutputs_267__0, registerOutputs_268__15, 
         registerOutputs_268__14, registerOutputs_268__13, 
         registerOutputs_268__12, registerOutputs_268__11, 
         registerOutputs_268__10, registerOutputs_268__9, registerOutputs_268__8, 
         registerOutputs_268__7, registerOutputs_268__6, registerOutputs_268__5, 
         registerOutputs_268__4, registerOutputs_268__3, registerOutputs_268__2, 
         registerOutputs_268__1, registerOutputs_268__0, registerOutputs_269__15, 
         registerOutputs_269__14, registerOutputs_269__13, 
         registerOutputs_269__12, registerOutputs_269__11, 
         registerOutputs_269__10, registerOutputs_269__9, registerOutputs_269__8, 
         registerOutputs_269__7, registerOutputs_269__6, registerOutputs_269__5, 
         registerOutputs_269__4, registerOutputs_269__3, registerOutputs_269__2, 
         registerOutputs_269__1, registerOutputs_269__0, registerOutputs_270__15, 
         registerOutputs_270__14, registerOutputs_270__13, 
         registerOutputs_270__12, registerOutputs_270__11, 
         registerOutputs_270__10, registerOutputs_270__9, registerOutputs_270__8, 
         registerOutputs_270__7, registerOutputs_270__6, registerOutputs_270__5, 
         registerOutputs_270__4, registerOutputs_270__3, registerOutputs_270__2, 
         registerOutputs_270__1, registerOutputs_270__0, registerOutputs_271__15, 
         registerOutputs_271__14, registerOutputs_271__13, 
         registerOutputs_271__12, registerOutputs_271__11, 
         registerOutputs_271__10, registerOutputs_271__9, registerOutputs_271__8, 
         registerOutputs_271__7, registerOutputs_271__6, registerOutputs_271__5, 
         registerOutputs_271__4, registerOutputs_271__3, registerOutputs_271__2, 
         registerOutputs_271__1, registerOutputs_271__0, registerOutputs_272__15, 
         registerOutputs_272__14, registerOutputs_272__13, 
         registerOutputs_272__12, registerOutputs_272__11, 
         registerOutputs_272__10, registerOutputs_272__9, registerOutputs_272__8, 
         registerOutputs_272__7, registerOutputs_272__6, registerOutputs_272__5, 
         registerOutputs_272__4, registerOutputs_272__3, registerOutputs_272__2, 
         registerOutputs_272__1, registerOutputs_272__0, registerOutputs_273__15, 
         registerOutputs_273__14, registerOutputs_273__13, 
         registerOutputs_273__12, registerOutputs_273__11, 
         registerOutputs_273__10, registerOutputs_273__9, registerOutputs_273__8, 
         registerOutputs_273__7, registerOutputs_273__6, registerOutputs_273__5, 
         registerOutputs_273__4, registerOutputs_273__3, registerOutputs_273__2, 
         registerOutputs_273__1, registerOutputs_273__0, registerOutputs_274__15, 
         registerOutputs_274__14, registerOutputs_274__13, 
         registerOutputs_274__12, registerOutputs_274__11, 
         registerOutputs_274__10, registerOutputs_274__9, registerOutputs_274__8, 
         registerOutputs_274__7, registerOutputs_274__6, registerOutputs_274__5, 
         registerOutputs_274__4, registerOutputs_274__3, registerOutputs_274__2, 
         registerOutputs_274__1, registerOutputs_274__0, registerOutputs_275__15, 
         registerOutputs_275__14, registerOutputs_275__13, 
         registerOutputs_275__12, registerOutputs_275__11, 
         registerOutputs_275__10, registerOutputs_275__9, registerOutputs_275__8, 
         registerOutputs_275__7, registerOutputs_275__6, registerOutputs_275__5, 
         registerOutputs_275__4, registerOutputs_275__3, registerOutputs_275__2, 
         registerOutputs_275__1, registerOutputs_275__0, registerOutputs_276__15, 
         registerOutputs_276__14, registerOutputs_276__13, 
         registerOutputs_276__12, registerOutputs_276__11, 
         registerOutputs_276__10, registerOutputs_276__9, registerOutputs_276__8, 
         registerOutputs_276__7, registerOutputs_276__6, registerOutputs_276__5, 
         registerOutputs_276__4, registerOutputs_276__3, registerOutputs_276__2, 
         registerOutputs_276__1, registerOutputs_276__0, registerOutputs_277__15, 
         registerOutputs_277__14, registerOutputs_277__13, 
         registerOutputs_277__12, registerOutputs_277__11, 
         registerOutputs_277__10, registerOutputs_277__9, registerOutputs_277__8, 
         registerOutputs_277__7, registerOutputs_277__6, registerOutputs_277__5, 
         registerOutputs_277__4, registerOutputs_277__3, registerOutputs_277__2, 
         registerOutputs_277__1, registerOutputs_277__0, registerOutputs_278__15, 
         registerOutputs_278__14, registerOutputs_278__13, 
         registerOutputs_278__12, registerOutputs_278__11, 
         registerOutputs_278__10, registerOutputs_278__9, registerOutputs_278__8, 
         registerOutputs_278__7, registerOutputs_278__6, registerOutputs_278__5, 
         registerOutputs_278__4, registerOutputs_278__3, registerOutputs_278__2, 
         registerOutputs_278__1, registerOutputs_278__0, registerOutputs_279__15, 
         registerOutputs_279__14, registerOutputs_279__13, 
         registerOutputs_279__12, registerOutputs_279__11, 
         registerOutputs_279__10, registerOutputs_279__9, registerOutputs_279__8, 
         registerOutputs_279__7, registerOutputs_279__6, registerOutputs_279__5, 
         registerOutputs_279__4, registerOutputs_279__3, registerOutputs_279__2, 
         registerOutputs_279__1, registerOutputs_279__0, registerOutputs_280__15, 
         registerOutputs_280__14, registerOutputs_280__13, 
         registerOutputs_280__12, registerOutputs_280__11, 
         registerOutputs_280__10, registerOutputs_280__9, registerOutputs_280__8, 
         registerOutputs_280__7, registerOutputs_280__6, registerOutputs_280__5, 
         registerOutputs_280__4, registerOutputs_280__3, registerOutputs_280__2, 
         registerOutputs_280__1, registerOutputs_280__0, registerOutputs_281__15, 
         registerOutputs_281__14, registerOutputs_281__13, 
         registerOutputs_281__12, registerOutputs_281__11, 
         registerOutputs_281__10, registerOutputs_281__9, registerOutputs_281__8, 
         registerOutputs_281__7, registerOutputs_281__6, registerOutputs_281__5, 
         registerOutputs_281__4, registerOutputs_281__3, registerOutputs_281__2, 
         registerOutputs_281__1, registerOutputs_281__0, registerOutputs_282__15, 
         registerOutputs_282__14, registerOutputs_282__13, 
         registerOutputs_282__12, registerOutputs_282__11, 
         registerOutputs_282__10, registerOutputs_282__9, registerOutputs_282__8, 
         registerOutputs_282__7, registerOutputs_282__6, registerOutputs_282__5, 
         registerOutputs_282__4, registerOutputs_282__3, registerOutputs_282__2, 
         registerOutputs_282__1, registerOutputs_282__0, registerOutputs_283__15, 
         registerOutputs_283__14, registerOutputs_283__13, 
         registerOutputs_283__12, registerOutputs_283__11, 
         registerOutputs_283__10, registerOutputs_283__9, registerOutputs_283__8, 
         registerOutputs_283__7, registerOutputs_283__6, registerOutputs_283__5, 
         registerOutputs_283__4, registerOutputs_283__3, registerOutputs_283__2, 
         registerOutputs_283__1, registerOutputs_283__0, registerOutputs_284__15, 
         registerOutputs_284__14, registerOutputs_284__13, 
         registerOutputs_284__12, registerOutputs_284__11, 
         registerOutputs_284__10, registerOutputs_284__9, registerOutputs_284__8, 
         registerOutputs_284__7, registerOutputs_284__6, registerOutputs_284__5, 
         registerOutputs_284__4, registerOutputs_284__3, registerOutputs_284__2, 
         registerOutputs_284__1, registerOutputs_284__0, registerOutputs_285__15, 
         registerOutputs_285__14, registerOutputs_285__13, 
         registerOutputs_285__12, registerOutputs_285__11, 
         registerOutputs_285__10, registerOutputs_285__9, registerOutputs_285__8, 
         registerOutputs_285__7, registerOutputs_285__6, registerOutputs_285__5, 
         registerOutputs_285__4, registerOutputs_285__3, registerOutputs_285__2, 
         registerOutputs_285__1, registerOutputs_285__0, registerOutputs_286__15, 
         registerOutputs_286__14, registerOutputs_286__13, 
         registerOutputs_286__12, registerOutputs_286__11, 
         registerOutputs_286__10, registerOutputs_286__9, registerOutputs_286__8, 
         registerOutputs_286__7, registerOutputs_286__6, registerOutputs_286__5, 
         registerOutputs_286__4, registerOutputs_286__3, registerOutputs_286__2, 
         registerOutputs_286__1, registerOutputs_286__0, registerOutputs_287__15, 
         registerOutputs_287__14, registerOutputs_287__13, 
         registerOutputs_287__12, registerOutputs_287__11, 
         registerOutputs_287__10, registerOutputs_287__9, registerOutputs_287__8, 
         registerOutputs_287__7, registerOutputs_287__6, registerOutputs_287__5, 
         registerOutputs_287__4, registerOutputs_287__3, registerOutputs_287__2, 
         registerOutputs_287__1, registerOutputs_287__0, registerOutputs_288__15, 
         registerOutputs_288__14, registerOutputs_288__13, 
         registerOutputs_288__12, registerOutputs_288__11, 
         registerOutputs_288__10, registerOutputs_288__9, registerOutputs_288__8, 
         registerOutputs_288__7, registerOutputs_288__6, registerOutputs_288__5, 
         registerOutputs_288__4, registerOutputs_288__3, registerOutputs_288__2, 
         registerOutputs_288__1, registerOutputs_288__0, registerOutputs_289__15, 
         registerOutputs_289__14, registerOutputs_289__13, 
         registerOutputs_289__12, registerOutputs_289__11, 
         registerOutputs_289__10, registerOutputs_289__9, registerOutputs_289__8, 
         registerOutputs_289__7, registerOutputs_289__6, registerOutputs_289__5, 
         registerOutputs_289__4, registerOutputs_289__3, registerOutputs_289__2, 
         registerOutputs_289__1, registerOutputs_289__0, registerOutputs_290__15, 
         registerOutputs_290__14, registerOutputs_290__13, 
         registerOutputs_290__12, registerOutputs_290__11, 
         registerOutputs_290__10, registerOutputs_290__9, registerOutputs_290__8, 
         registerOutputs_290__7, registerOutputs_290__6, registerOutputs_290__5, 
         registerOutputs_290__4, registerOutputs_290__3, registerOutputs_290__2, 
         registerOutputs_290__1, registerOutputs_290__0, registerOutputs_291__15, 
         registerOutputs_291__14, registerOutputs_291__13, 
         registerOutputs_291__12, registerOutputs_291__11, 
         registerOutputs_291__10, registerOutputs_291__9, registerOutputs_291__8, 
         registerOutputs_291__7, registerOutputs_291__6, registerOutputs_291__5, 
         registerOutputs_291__4, registerOutputs_291__3, registerOutputs_291__2, 
         registerOutputs_291__1, registerOutputs_291__0, registerOutputs_292__15, 
         registerOutputs_292__14, registerOutputs_292__13, 
         registerOutputs_292__12, registerOutputs_292__11, 
         registerOutputs_292__10, registerOutputs_292__9, registerOutputs_292__8, 
         registerOutputs_292__7, registerOutputs_292__6, registerOutputs_292__5, 
         registerOutputs_292__4, registerOutputs_292__3, registerOutputs_292__2, 
         registerOutputs_292__1, registerOutputs_292__0, registerOutputs_293__15, 
         registerOutputs_293__14, registerOutputs_293__13, 
         registerOutputs_293__12, registerOutputs_293__11, 
         registerOutputs_293__10, registerOutputs_293__9, registerOutputs_293__8, 
         registerOutputs_293__7, registerOutputs_293__6, registerOutputs_293__5, 
         registerOutputs_293__4, registerOutputs_293__3, registerOutputs_293__2, 
         registerOutputs_293__1, registerOutputs_293__0, registerOutputs_294__15, 
         registerOutputs_294__14, registerOutputs_294__13, 
         registerOutputs_294__12, registerOutputs_294__11, 
         registerOutputs_294__10, registerOutputs_294__9, registerOutputs_294__8, 
         registerOutputs_294__7, registerOutputs_294__6, registerOutputs_294__5, 
         registerOutputs_294__4, registerOutputs_294__3, registerOutputs_294__2, 
         registerOutputs_294__1, registerOutputs_294__0, registerOutputs_295__15, 
         registerOutputs_295__14, registerOutputs_295__13, 
         registerOutputs_295__12, registerOutputs_295__11, 
         registerOutputs_295__10, registerOutputs_295__9, registerOutputs_295__8, 
         registerOutputs_295__7, registerOutputs_295__6, registerOutputs_295__5, 
         registerOutputs_295__4, registerOutputs_295__3, registerOutputs_295__2, 
         registerOutputs_295__1, registerOutputs_295__0, registerOutputs_296__15, 
         registerOutputs_296__14, registerOutputs_296__13, 
         registerOutputs_296__12, registerOutputs_296__11, 
         registerOutputs_296__10, registerOutputs_296__9, registerOutputs_296__8, 
         registerOutputs_296__7, registerOutputs_296__6, registerOutputs_296__5, 
         registerOutputs_296__4, registerOutputs_296__3, registerOutputs_296__2, 
         registerOutputs_296__1, registerOutputs_296__0, registerOutputs_297__15, 
         registerOutputs_297__14, registerOutputs_297__13, 
         registerOutputs_297__12, registerOutputs_297__11, 
         registerOutputs_297__10, registerOutputs_297__9, registerOutputs_297__8, 
         registerOutputs_297__7, registerOutputs_297__6, registerOutputs_297__5, 
         registerOutputs_297__4, registerOutputs_297__3, registerOutputs_297__2, 
         registerOutputs_297__1, registerOutputs_297__0, registerOutputs_298__15, 
         registerOutputs_298__14, registerOutputs_298__13, 
         registerOutputs_298__12, registerOutputs_298__11, 
         registerOutputs_298__10, registerOutputs_298__9, registerOutputs_298__8, 
         registerOutputs_298__7, registerOutputs_298__6, registerOutputs_298__5, 
         registerOutputs_298__4, registerOutputs_298__3, registerOutputs_298__2, 
         registerOutputs_298__1, registerOutputs_298__0, registerOutputs_299__15, 
         registerOutputs_299__14, registerOutputs_299__13, 
         registerOutputs_299__12, registerOutputs_299__11, 
         registerOutputs_299__10, registerOutputs_299__9, registerOutputs_299__8, 
         registerOutputs_299__7, registerOutputs_299__6, registerOutputs_299__5, 
         registerOutputs_299__4, registerOutputs_299__3, registerOutputs_299__2, 
         registerOutputs_299__1, registerOutputs_299__0, registerOutputs_300__15, 
         registerOutputs_300__14, registerOutputs_300__13, 
         registerOutputs_300__12, registerOutputs_300__11, 
         registerOutputs_300__10, registerOutputs_300__9, registerOutputs_300__8, 
         registerOutputs_300__7, registerOutputs_300__6, registerOutputs_300__5, 
         registerOutputs_300__4, registerOutputs_300__3, registerOutputs_300__2, 
         registerOutputs_300__1, registerOutputs_300__0, registerOutputs_301__15, 
         registerOutputs_301__14, registerOutputs_301__13, 
         registerOutputs_301__12, registerOutputs_301__11, 
         registerOutputs_301__10, registerOutputs_301__9, registerOutputs_301__8, 
         registerOutputs_301__7, registerOutputs_301__6, registerOutputs_301__5, 
         registerOutputs_301__4, registerOutputs_301__3, registerOutputs_301__2, 
         registerOutputs_301__1, registerOutputs_301__0, registerOutputs_302__15, 
         registerOutputs_302__14, registerOutputs_302__13, 
         registerOutputs_302__12, registerOutputs_302__11, 
         registerOutputs_302__10, registerOutputs_302__9, registerOutputs_302__8, 
         registerOutputs_302__7, registerOutputs_302__6, registerOutputs_302__5, 
         registerOutputs_302__4, registerOutputs_302__3, registerOutputs_302__2, 
         registerOutputs_302__1, registerOutputs_302__0, registerOutputs_303__15, 
         registerOutputs_303__14, registerOutputs_303__13, 
         registerOutputs_303__12, registerOutputs_303__11, 
         registerOutputs_303__10, registerOutputs_303__9, registerOutputs_303__8, 
         registerOutputs_303__7, registerOutputs_303__6, registerOutputs_303__5, 
         registerOutputs_303__4, registerOutputs_303__3, registerOutputs_303__2, 
         registerOutputs_303__1, registerOutputs_303__0, registerOutputs_304__15, 
         registerOutputs_304__14, registerOutputs_304__13, 
         registerOutputs_304__12, registerOutputs_304__11, 
         registerOutputs_304__10, registerOutputs_304__9, registerOutputs_304__8, 
         registerOutputs_304__7, registerOutputs_304__6, registerOutputs_304__5, 
         registerOutputs_304__4, registerOutputs_304__3, registerOutputs_304__2, 
         registerOutputs_304__1, registerOutputs_304__0, registerOutputs_305__15, 
         registerOutputs_305__14, registerOutputs_305__13, 
         registerOutputs_305__12, registerOutputs_305__11, 
         registerOutputs_305__10, registerOutputs_305__9, registerOutputs_305__8, 
         registerOutputs_305__7, registerOutputs_305__6, registerOutputs_305__5, 
         registerOutputs_305__4, registerOutputs_305__3, registerOutputs_305__2, 
         registerOutputs_305__1, registerOutputs_305__0, registerOutputs_306__15, 
         registerOutputs_306__14, registerOutputs_306__13, 
         registerOutputs_306__12, registerOutputs_306__11, 
         registerOutputs_306__10, registerOutputs_306__9, registerOutputs_306__8, 
         registerOutputs_306__7, registerOutputs_306__6, registerOutputs_306__5, 
         registerOutputs_306__4, registerOutputs_306__3, registerOutputs_306__2, 
         registerOutputs_306__1, registerOutputs_306__0, registerOutputs_307__15, 
         registerOutputs_307__14, registerOutputs_307__13, 
         registerOutputs_307__12, registerOutputs_307__11, 
         registerOutputs_307__10, registerOutputs_307__9, registerOutputs_307__8, 
         registerOutputs_307__7, registerOutputs_307__6, registerOutputs_307__5, 
         registerOutputs_307__4, registerOutputs_307__3, registerOutputs_307__2, 
         registerOutputs_307__1, registerOutputs_307__0, registerOutputs_308__15, 
         registerOutputs_308__14, registerOutputs_308__13, 
         registerOutputs_308__12, registerOutputs_308__11, 
         registerOutputs_308__10, registerOutputs_308__9, registerOutputs_308__8, 
         registerOutputs_308__7, registerOutputs_308__6, registerOutputs_308__5, 
         registerOutputs_308__4, registerOutputs_308__3, registerOutputs_308__2, 
         registerOutputs_308__1, registerOutputs_308__0, registerOutputs_309__15, 
         registerOutputs_309__14, registerOutputs_309__13, 
         registerOutputs_309__12, registerOutputs_309__11, 
         registerOutputs_309__10, registerOutputs_309__9, registerOutputs_309__8, 
         registerOutputs_309__7, registerOutputs_309__6, registerOutputs_309__5, 
         registerOutputs_309__4, registerOutputs_309__3, registerOutputs_309__2, 
         registerOutputs_309__1, registerOutputs_309__0, registerOutputs_310__15, 
         registerOutputs_310__14, registerOutputs_310__13, 
         registerOutputs_310__12, registerOutputs_310__11, 
         registerOutputs_310__10, registerOutputs_310__9, registerOutputs_310__8, 
         registerOutputs_310__7, registerOutputs_310__6, registerOutputs_310__5, 
         registerOutputs_310__4, registerOutputs_310__3, registerOutputs_310__2, 
         registerOutputs_310__1, registerOutputs_310__0, registerOutputs_311__15, 
         registerOutputs_311__14, registerOutputs_311__13, 
         registerOutputs_311__12, registerOutputs_311__11, 
         registerOutputs_311__10, registerOutputs_311__9, registerOutputs_311__8, 
         registerOutputs_311__7, registerOutputs_311__6, registerOutputs_311__5, 
         registerOutputs_311__4, registerOutputs_311__3, registerOutputs_311__2, 
         registerOutputs_311__1, registerOutputs_311__0, registerOutputs_312__15, 
         registerOutputs_312__14, registerOutputs_312__13, 
         registerOutputs_312__12, registerOutputs_312__11, 
         registerOutputs_312__10, registerOutputs_312__9, registerOutputs_312__8, 
         registerOutputs_312__7, registerOutputs_312__6, registerOutputs_312__5, 
         registerOutputs_312__4, registerOutputs_312__3, registerOutputs_312__2, 
         registerOutputs_312__1, registerOutputs_312__0, registerOutputs_313__15, 
         registerOutputs_313__14, registerOutputs_313__13, 
         registerOutputs_313__12, registerOutputs_313__11, 
         registerOutputs_313__10, registerOutputs_313__9, registerOutputs_313__8, 
         registerOutputs_313__7, registerOutputs_313__6, registerOutputs_313__5, 
         registerOutputs_313__4, registerOutputs_313__3, registerOutputs_313__2, 
         registerOutputs_313__1, registerOutputs_313__0, registerOutputs_314__15, 
         registerOutputs_314__14, registerOutputs_314__13, 
         registerOutputs_314__12, registerOutputs_314__11, 
         registerOutputs_314__10, registerOutputs_314__9, registerOutputs_314__8, 
         registerOutputs_314__7, registerOutputs_314__6, registerOutputs_314__5, 
         registerOutputs_314__4, registerOutputs_314__3, registerOutputs_314__2, 
         registerOutputs_314__1, registerOutputs_314__0, registerOutputs_315__15, 
         registerOutputs_315__14, registerOutputs_315__13, 
         registerOutputs_315__12, registerOutputs_315__11, 
         registerOutputs_315__10, registerOutputs_315__9, registerOutputs_315__8, 
         registerOutputs_315__7, registerOutputs_315__6, registerOutputs_315__5, 
         registerOutputs_315__4, registerOutputs_315__3, registerOutputs_315__2, 
         registerOutputs_315__1, registerOutputs_315__0, registerOutputs_316__15, 
         registerOutputs_316__14, registerOutputs_316__13, 
         registerOutputs_316__12, registerOutputs_316__11, 
         registerOutputs_316__10, registerOutputs_316__9, registerOutputs_316__8, 
         registerOutputs_316__7, registerOutputs_316__6, registerOutputs_316__5, 
         registerOutputs_316__4, registerOutputs_316__3, registerOutputs_316__2, 
         registerOutputs_316__1, registerOutputs_316__0, registerOutputs_317__15, 
         registerOutputs_317__14, registerOutputs_317__13, 
         registerOutputs_317__12, registerOutputs_317__11, 
         registerOutputs_317__10, registerOutputs_317__9, registerOutputs_317__8, 
         registerOutputs_317__7, registerOutputs_317__6, registerOutputs_317__5, 
         registerOutputs_317__4, registerOutputs_317__3, registerOutputs_317__2, 
         registerOutputs_317__1, registerOutputs_317__0, registerOutputs_318__15, 
         registerOutputs_318__14, registerOutputs_318__13, 
         registerOutputs_318__12, registerOutputs_318__11, 
         registerOutputs_318__10, registerOutputs_318__9, registerOutputs_318__8, 
         registerOutputs_318__7, registerOutputs_318__6, registerOutputs_318__5, 
         registerOutputs_318__4, registerOutputs_318__3, registerOutputs_318__2, 
         registerOutputs_318__1, registerOutputs_318__0, registerOutputs_319__15, 
         registerOutputs_319__14, registerOutputs_319__13, 
         registerOutputs_319__12, registerOutputs_319__11, 
         registerOutputs_319__10, registerOutputs_319__9, registerOutputs_319__8, 
         registerOutputs_319__7, registerOutputs_319__6, registerOutputs_319__5, 
         registerOutputs_319__4, registerOutputs_319__3, registerOutputs_319__2, 
         registerOutputs_319__1, registerOutputs_319__0, registerOutputs_320__15, 
         registerOutputs_320__14, registerOutputs_320__13, 
         registerOutputs_320__12, registerOutputs_320__11, 
         registerOutputs_320__10, registerOutputs_320__9, registerOutputs_320__8, 
         registerOutputs_320__7, registerOutputs_320__6, registerOutputs_320__5, 
         registerOutputs_320__4, registerOutputs_320__3, registerOutputs_320__2, 
         registerOutputs_320__1, registerOutputs_320__0, registerOutputs_321__15, 
         registerOutputs_321__14, registerOutputs_321__13, 
         registerOutputs_321__12, registerOutputs_321__11, 
         registerOutputs_321__10, registerOutputs_321__9, registerOutputs_321__8, 
         registerOutputs_321__7, registerOutputs_321__6, registerOutputs_321__5, 
         registerOutputs_321__4, registerOutputs_321__3, registerOutputs_321__2, 
         registerOutputs_321__1, registerOutputs_321__0, registerOutputs_322__15, 
         registerOutputs_322__14, registerOutputs_322__13, 
         registerOutputs_322__12, registerOutputs_322__11, 
         registerOutputs_322__10, registerOutputs_322__9, registerOutputs_322__8, 
         registerOutputs_322__7, registerOutputs_322__6, registerOutputs_322__5, 
         registerOutputs_322__4, registerOutputs_322__3, registerOutputs_322__2, 
         registerOutputs_322__1, registerOutputs_322__0, registerOutputs_323__15, 
         registerOutputs_323__14, registerOutputs_323__13, 
         registerOutputs_323__12, registerOutputs_323__11, 
         registerOutputs_323__10, registerOutputs_323__9, registerOutputs_323__8, 
         registerOutputs_323__7, registerOutputs_323__6, registerOutputs_323__5, 
         registerOutputs_323__4, registerOutputs_323__3, registerOutputs_323__2, 
         registerOutputs_323__1, registerOutputs_323__0, registerOutputs_324__15, 
         registerOutputs_324__14, registerOutputs_324__13, 
         registerOutputs_324__12, registerOutputs_324__11, 
         registerOutputs_324__10, registerOutputs_324__9, registerOutputs_324__8, 
         registerOutputs_324__7, registerOutputs_324__6, registerOutputs_324__5, 
         registerOutputs_324__4, registerOutputs_324__3, registerOutputs_324__2, 
         registerOutputs_324__1, registerOutputs_324__0, registerOutputs_325__15, 
         registerOutputs_325__14, registerOutputs_325__13, 
         registerOutputs_325__12, registerOutputs_325__11, 
         registerOutputs_325__10, registerOutputs_325__9, registerOutputs_325__8, 
         registerOutputs_325__7, registerOutputs_325__6, registerOutputs_325__5, 
         registerOutputs_325__4, registerOutputs_325__3, registerOutputs_325__2, 
         registerOutputs_325__1, registerOutputs_325__0, registerOutputs_326__15, 
         registerOutputs_326__14, registerOutputs_326__13, 
         registerOutputs_326__12, registerOutputs_326__11, 
         registerOutputs_326__10, registerOutputs_326__9, registerOutputs_326__8, 
         registerOutputs_326__7, registerOutputs_326__6, registerOutputs_326__5, 
         registerOutputs_326__4, registerOutputs_326__3, registerOutputs_326__2, 
         registerOutputs_326__1, registerOutputs_326__0, registerOutputs_327__15, 
         registerOutputs_327__14, registerOutputs_327__13, 
         registerOutputs_327__12, registerOutputs_327__11, 
         registerOutputs_327__10, registerOutputs_327__9, registerOutputs_327__8, 
         registerOutputs_327__7, registerOutputs_327__6, registerOutputs_327__5, 
         registerOutputs_327__4, registerOutputs_327__3, registerOutputs_327__2, 
         registerOutputs_327__1, registerOutputs_327__0, registerOutputs_328__15, 
         registerOutputs_328__14, registerOutputs_328__13, 
         registerOutputs_328__12, registerOutputs_328__11, 
         registerOutputs_328__10, registerOutputs_328__9, registerOutputs_328__8, 
         registerOutputs_328__7, registerOutputs_328__6, registerOutputs_328__5, 
         registerOutputs_328__4, registerOutputs_328__3, registerOutputs_328__2, 
         registerOutputs_328__1, registerOutputs_328__0, registerOutputs_329__15, 
         registerOutputs_329__14, registerOutputs_329__13, 
         registerOutputs_329__12, registerOutputs_329__11, 
         registerOutputs_329__10, registerOutputs_329__9, registerOutputs_329__8, 
         registerOutputs_329__7, registerOutputs_329__6, registerOutputs_329__5, 
         registerOutputs_329__4, registerOutputs_329__3, registerOutputs_329__2, 
         registerOutputs_329__1, registerOutputs_329__0, registerOutputs_330__15, 
         registerOutputs_330__14, registerOutputs_330__13, 
         registerOutputs_330__12, registerOutputs_330__11, 
         registerOutputs_330__10, registerOutputs_330__9, registerOutputs_330__8, 
         registerOutputs_330__7, registerOutputs_330__6, registerOutputs_330__5, 
         registerOutputs_330__4, registerOutputs_330__3, registerOutputs_330__2, 
         registerOutputs_330__1, registerOutputs_330__0, registerOutputs_331__15, 
         registerOutputs_331__14, registerOutputs_331__13, 
         registerOutputs_331__12, registerOutputs_331__11, 
         registerOutputs_331__10, registerOutputs_331__9, registerOutputs_331__8, 
         registerOutputs_331__7, registerOutputs_331__6, registerOutputs_331__5, 
         registerOutputs_331__4, registerOutputs_331__3, registerOutputs_331__2, 
         registerOutputs_331__1, registerOutputs_331__0, registerOutputs_332__15, 
         registerOutputs_332__14, registerOutputs_332__13, 
         registerOutputs_332__12, registerOutputs_332__11, 
         registerOutputs_332__10, registerOutputs_332__9, registerOutputs_332__8, 
         registerOutputs_332__7, registerOutputs_332__6, registerOutputs_332__5, 
         registerOutputs_332__4, registerOutputs_332__3, registerOutputs_332__2, 
         registerOutputs_332__1, registerOutputs_332__0, registerOutputs_333__15, 
         registerOutputs_333__14, registerOutputs_333__13, 
         registerOutputs_333__12, registerOutputs_333__11, 
         registerOutputs_333__10, registerOutputs_333__9, registerOutputs_333__8, 
         registerOutputs_333__7, registerOutputs_333__6, registerOutputs_333__5, 
         registerOutputs_333__4, registerOutputs_333__3, registerOutputs_333__2, 
         registerOutputs_333__1, registerOutputs_333__0, registerOutputs_334__15, 
         registerOutputs_334__14, registerOutputs_334__13, 
         registerOutputs_334__12, registerOutputs_334__11, 
         registerOutputs_334__10, registerOutputs_334__9, registerOutputs_334__8, 
         registerOutputs_334__7, registerOutputs_334__6, registerOutputs_334__5, 
         registerOutputs_334__4, registerOutputs_334__3, registerOutputs_334__2, 
         registerOutputs_334__1, registerOutputs_334__0, registerOutputs_335__15, 
         registerOutputs_335__14, registerOutputs_335__13, 
         registerOutputs_335__12, registerOutputs_335__11, 
         registerOutputs_335__10, registerOutputs_335__9, registerOutputs_335__8, 
         registerOutputs_335__7, registerOutputs_335__6, registerOutputs_335__5, 
         registerOutputs_335__4, registerOutputs_335__3, registerOutputs_335__2, 
         registerOutputs_335__1, registerOutputs_335__0, registerOutputs_336__15, 
         registerOutputs_336__14, registerOutputs_336__13, 
         registerOutputs_336__12, registerOutputs_336__11, 
         registerOutputs_336__10, registerOutputs_336__9, registerOutputs_336__8, 
         registerOutputs_336__7, registerOutputs_336__6, registerOutputs_336__5, 
         registerOutputs_336__4, registerOutputs_336__3, registerOutputs_336__2, 
         registerOutputs_336__1, registerOutputs_336__0, registerOutputs_337__15, 
         registerOutputs_337__14, registerOutputs_337__13, 
         registerOutputs_337__12, registerOutputs_337__11, 
         registerOutputs_337__10, registerOutputs_337__9, registerOutputs_337__8, 
         registerOutputs_337__7, registerOutputs_337__6, registerOutputs_337__5, 
         registerOutputs_337__4, registerOutputs_337__3, registerOutputs_337__2, 
         registerOutputs_337__1, registerOutputs_337__0, registerOutputs_338__15, 
         registerOutputs_338__14, registerOutputs_338__13, 
         registerOutputs_338__12, registerOutputs_338__11, 
         registerOutputs_338__10, registerOutputs_338__9, registerOutputs_338__8, 
         registerOutputs_338__7, registerOutputs_338__6, registerOutputs_338__5, 
         registerOutputs_338__4, registerOutputs_338__3, registerOutputs_338__2, 
         registerOutputs_338__1, registerOutputs_338__0, registerOutputs_339__15, 
         registerOutputs_339__14, registerOutputs_339__13, 
         registerOutputs_339__12, registerOutputs_339__11, 
         registerOutputs_339__10, registerOutputs_339__9, registerOutputs_339__8, 
         registerOutputs_339__7, registerOutputs_339__6, registerOutputs_339__5, 
         registerOutputs_339__4, registerOutputs_339__3, registerOutputs_339__2, 
         registerOutputs_339__1, registerOutputs_339__0, registerOutputs_340__15, 
         registerOutputs_340__14, registerOutputs_340__13, 
         registerOutputs_340__12, registerOutputs_340__11, 
         registerOutputs_340__10, registerOutputs_340__9, registerOutputs_340__8, 
         registerOutputs_340__7, registerOutputs_340__6, registerOutputs_340__5, 
         registerOutputs_340__4, registerOutputs_340__3, registerOutputs_340__2, 
         registerOutputs_340__1, registerOutputs_340__0, registerOutputs_341__15, 
         registerOutputs_341__14, registerOutputs_341__13, 
         registerOutputs_341__12, registerOutputs_341__11, 
         registerOutputs_341__10, registerOutputs_341__9, registerOutputs_341__8, 
         registerOutputs_341__7, registerOutputs_341__6, registerOutputs_341__5, 
         registerOutputs_341__4, registerOutputs_341__3, registerOutputs_341__2, 
         registerOutputs_341__1, registerOutputs_341__0, registerOutputs_342__15, 
         registerOutputs_342__14, registerOutputs_342__13, 
         registerOutputs_342__12, registerOutputs_342__11, 
         registerOutputs_342__10, registerOutputs_342__9, registerOutputs_342__8, 
         registerOutputs_342__7, registerOutputs_342__6, registerOutputs_342__5, 
         registerOutputs_342__4, registerOutputs_342__3, registerOutputs_342__2, 
         registerOutputs_342__1, registerOutputs_342__0, registerOutputs_343__15, 
         registerOutputs_343__14, registerOutputs_343__13, 
         registerOutputs_343__12, registerOutputs_343__11, 
         registerOutputs_343__10, registerOutputs_343__9, registerOutputs_343__8, 
         registerOutputs_343__7, registerOutputs_343__6, registerOutputs_343__5, 
         registerOutputs_343__4, registerOutputs_343__3, registerOutputs_343__2, 
         registerOutputs_343__1, registerOutputs_343__0, registerOutputs_344__15, 
         registerOutputs_344__14, registerOutputs_344__13, 
         registerOutputs_344__12, registerOutputs_344__11, 
         registerOutputs_344__10, registerOutputs_344__9, registerOutputs_344__8, 
         registerOutputs_344__7, registerOutputs_344__6, registerOutputs_344__5, 
         registerOutputs_344__4, registerOutputs_344__3, registerOutputs_344__2, 
         registerOutputs_344__1, registerOutputs_344__0, registerOutputs_345__15, 
         registerOutputs_345__14, registerOutputs_345__13, 
         registerOutputs_345__12, registerOutputs_345__11, 
         registerOutputs_345__10, registerOutputs_345__9, registerOutputs_345__8, 
         registerOutputs_345__7, registerOutputs_345__6, registerOutputs_345__5, 
         registerOutputs_345__4, registerOutputs_345__3, registerOutputs_345__2, 
         registerOutputs_345__1, registerOutputs_345__0, registerOutputs_346__15, 
         registerOutputs_346__14, registerOutputs_346__13, 
         registerOutputs_346__12, registerOutputs_346__11, 
         registerOutputs_346__10, registerOutputs_346__9, registerOutputs_346__8, 
         registerOutputs_346__7, registerOutputs_346__6, registerOutputs_346__5, 
         registerOutputs_346__4, registerOutputs_346__3, registerOutputs_346__2, 
         registerOutputs_346__1, registerOutputs_346__0, registerOutputs_347__15, 
         registerOutputs_347__14, registerOutputs_347__13, 
         registerOutputs_347__12, registerOutputs_347__11, 
         registerOutputs_347__10, registerOutputs_347__9, registerOutputs_347__8, 
         registerOutputs_347__7, registerOutputs_347__6, registerOutputs_347__5, 
         registerOutputs_347__4, registerOutputs_347__3, registerOutputs_347__2, 
         registerOutputs_347__1, registerOutputs_347__0, registerOutputs_348__15, 
         registerOutputs_348__14, registerOutputs_348__13, 
         registerOutputs_348__12, registerOutputs_348__11, 
         registerOutputs_348__10, registerOutputs_348__9, registerOutputs_348__8, 
         registerOutputs_348__7, registerOutputs_348__6, registerOutputs_348__5, 
         registerOutputs_348__4, registerOutputs_348__3, registerOutputs_348__2, 
         registerOutputs_348__1, registerOutputs_348__0, registerOutputs_349__15, 
         registerOutputs_349__14, registerOutputs_349__13, 
         registerOutputs_349__12, registerOutputs_349__11, 
         registerOutputs_349__10, registerOutputs_349__9, registerOutputs_349__8, 
         registerOutputs_349__7, registerOutputs_349__6, registerOutputs_349__5, 
         registerOutputs_349__4, registerOutputs_349__3, registerOutputs_349__2, 
         registerOutputs_349__1, registerOutputs_349__0, registerOutputs_350__15, 
         registerOutputs_350__14, registerOutputs_350__13, 
         registerOutputs_350__12, registerOutputs_350__11, 
         registerOutputs_350__10, registerOutputs_350__9, registerOutputs_350__8, 
         registerOutputs_350__7, registerOutputs_350__6, registerOutputs_350__5, 
         registerOutputs_350__4, registerOutputs_350__3, registerOutputs_350__2, 
         registerOutputs_350__1, registerOutputs_350__0, registerOutputs_351__15, 
         registerOutputs_351__14, registerOutputs_351__13, 
         registerOutputs_351__12, registerOutputs_351__11, 
         registerOutputs_351__10, registerOutputs_351__9, registerOutputs_351__8, 
         registerOutputs_351__7, registerOutputs_351__6, registerOutputs_351__5, 
         registerOutputs_351__4, registerOutputs_351__3, registerOutputs_351__2, 
         registerOutputs_351__1, registerOutputs_351__0, registerOutputs_352__15, 
         registerOutputs_352__14, registerOutputs_352__13, 
         registerOutputs_352__12, registerOutputs_352__11, 
         registerOutputs_352__10, registerOutputs_352__9, registerOutputs_352__8, 
         registerOutputs_352__7, registerOutputs_352__6, registerOutputs_352__5, 
         registerOutputs_352__4, registerOutputs_352__3, registerOutputs_352__2, 
         registerOutputs_352__1, registerOutputs_352__0, registerOutputs_353__15, 
         registerOutputs_353__14, registerOutputs_353__13, 
         registerOutputs_353__12, registerOutputs_353__11, 
         registerOutputs_353__10, registerOutputs_353__9, registerOutputs_353__8, 
         registerOutputs_353__7, registerOutputs_353__6, registerOutputs_353__5, 
         registerOutputs_353__4, registerOutputs_353__3, registerOutputs_353__2, 
         registerOutputs_353__1, registerOutputs_353__0, registerOutputs_354__15, 
         registerOutputs_354__14, registerOutputs_354__13, 
         registerOutputs_354__12, registerOutputs_354__11, 
         registerOutputs_354__10, registerOutputs_354__9, registerOutputs_354__8, 
         registerOutputs_354__7, registerOutputs_354__6, registerOutputs_354__5, 
         registerOutputs_354__4, registerOutputs_354__3, registerOutputs_354__2, 
         registerOutputs_354__1, registerOutputs_354__0, registerOutputs_355__15, 
         registerOutputs_355__14, registerOutputs_355__13, 
         registerOutputs_355__12, registerOutputs_355__11, 
         registerOutputs_355__10, registerOutputs_355__9, registerOutputs_355__8, 
         registerOutputs_355__7, registerOutputs_355__6, registerOutputs_355__5, 
         registerOutputs_355__4, registerOutputs_355__3, registerOutputs_355__2, 
         registerOutputs_355__1, registerOutputs_355__0, registerOutputs_356__15, 
         registerOutputs_356__14, registerOutputs_356__13, 
         registerOutputs_356__12, registerOutputs_356__11, 
         registerOutputs_356__10, registerOutputs_356__9, registerOutputs_356__8, 
         registerOutputs_356__7, registerOutputs_356__6, registerOutputs_356__5, 
         registerOutputs_356__4, registerOutputs_356__3, registerOutputs_356__2, 
         registerOutputs_356__1, registerOutputs_356__0, registerOutputs_357__15, 
         registerOutputs_357__14, registerOutputs_357__13, 
         registerOutputs_357__12, registerOutputs_357__11, 
         registerOutputs_357__10, registerOutputs_357__9, registerOutputs_357__8, 
         registerOutputs_357__7, registerOutputs_357__6, registerOutputs_357__5, 
         registerOutputs_357__4, registerOutputs_357__3, registerOutputs_357__2, 
         registerOutputs_357__1, registerOutputs_357__0, registerOutputs_358__15, 
         registerOutputs_358__14, registerOutputs_358__13, 
         registerOutputs_358__12, registerOutputs_358__11, 
         registerOutputs_358__10, registerOutputs_358__9, registerOutputs_358__8, 
         registerOutputs_358__7, registerOutputs_358__6, registerOutputs_358__5, 
         registerOutputs_358__4, registerOutputs_358__3, registerOutputs_358__2, 
         registerOutputs_358__1, registerOutputs_358__0, registerOutputs_359__15, 
         registerOutputs_359__14, registerOutputs_359__13, 
         registerOutputs_359__12, registerOutputs_359__11, 
         registerOutputs_359__10, registerOutputs_359__9, registerOutputs_359__8, 
         registerOutputs_359__7, registerOutputs_359__6, registerOutputs_359__5, 
         registerOutputs_359__4, registerOutputs_359__3, registerOutputs_359__2, 
         registerOutputs_359__1, registerOutputs_359__0, registerOutputs_360__15, 
         registerOutputs_360__14, registerOutputs_360__13, 
         registerOutputs_360__12, registerOutputs_360__11, 
         registerOutputs_360__10, registerOutputs_360__9, registerOutputs_360__8, 
         registerOutputs_360__7, registerOutputs_360__6, registerOutputs_360__5, 
         registerOutputs_360__4, registerOutputs_360__3, registerOutputs_360__2, 
         registerOutputs_360__1, registerOutputs_360__0, registerOutputs_361__15, 
         registerOutputs_361__14, registerOutputs_361__13, 
         registerOutputs_361__12, registerOutputs_361__11, 
         registerOutputs_361__10, registerOutputs_361__9, registerOutputs_361__8, 
         registerOutputs_361__7, registerOutputs_361__6, registerOutputs_361__5, 
         registerOutputs_361__4, registerOutputs_361__3, registerOutputs_361__2, 
         registerOutputs_361__1, registerOutputs_361__0, registerOutputs_362__15, 
         registerOutputs_362__14, registerOutputs_362__13, 
         registerOutputs_362__12, registerOutputs_362__11, 
         registerOutputs_362__10, registerOutputs_362__9, registerOutputs_362__8, 
         registerOutputs_362__7, registerOutputs_362__6, registerOutputs_362__5, 
         registerOutputs_362__4, registerOutputs_362__3, registerOutputs_362__2, 
         registerOutputs_362__1, registerOutputs_362__0, registerOutputs_363__15, 
         registerOutputs_363__14, registerOutputs_363__13, 
         registerOutputs_363__12, registerOutputs_363__11, 
         registerOutputs_363__10, registerOutputs_363__9, registerOutputs_363__8, 
         registerOutputs_363__7, registerOutputs_363__6, registerOutputs_363__5, 
         registerOutputs_363__4, registerOutputs_363__3, registerOutputs_363__2, 
         registerOutputs_363__1, registerOutputs_363__0, registerOutputs_364__15, 
         registerOutputs_364__14, registerOutputs_364__13, 
         registerOutputs_364__12, registerOutputs_364__11, 
         registerOutputs_364__10, registerOutputs_364__9, registerOutputs_364__8, 
         registerOutputs_364__7, registerOutputs_364__6, registerOutputs_364__5, 
         registerOutputs_364__4, registerOutputs_364__3, registerOutputs_364__2, 
         registerOutputs_364__1, registerOutputs_364__0, registerOutputs_365__15, 
         registerOutputs_365__14, registerOutputs_365__13, 
         registerOutputs_365__12, registerOutputs_365__11, 
         registerOutputs_365__10, registerOutputs_365__9, registerOutputs_365__8, 
         registerOutputs_365__7, registerOutputs_365__6, registerOutputs_365__5, 
         registerOutputs_365__4, registerOutputs_365__3, registerOutputs_365__2, 
         registerOutputs_365__1, registerOutputs_365__0, registerOutputs_366__15, 
         registerOutputs_366__14, registerOutputs_366__13, 
         registerOutputs_366__12, registerOutputs_366__11, 
         registerOutputs_366__10, registerOutputs_366__9, registerOutputs_366__8, 
         registerOutputs_366__7, registerOutputs_366__6, registerOutputs_366__5, 
         registerOutputs_366__4, registerOutputs_366__3, registerOutputs_366__2, 
         registerOutputs_366__1, registerOutputs_366__0, registerOutputs_367__15, 
         registerOutputs_367__14, registerOutputs_367__13, 
         registerOutputs_367__12, registerOutputs_367__11, 
         registerOutputs_367__10, registerOutputs_367__9, registerOutputs_367__8, 
         registerOutputs_367__7, registerOutputs_367__6, registerOutputs_367__5, 
         registerOutputs_367__4, registerOutputs_367__3, registerOutputs_367__2, 
         registerOutputs_367__1, registerOutputs_367__0, registerOutputs_368__15, 
         registerOutputs_368__14, registerOutputs_368__13, 
         registerOutputs_368__12, registerOutputs_368__11, 
         registerOutputs_368__10, registerOutputs_368__9, registerOutputs_368__8, 
         registerOutputs_368__7, registerOutputs_368__6, registerOutputs_368__5, 
         registerOutputs_368__4, registerOutputs_368__3, registerOutputs_368__2, 
         registerOutputs_368__1, registerOutputs_368__0, registerOutputs_369__15, 
         registerOutputs_369__14, registerOutputs_369__13, 
         registerOutputs_369__12, registerOutputs_369__11, 
         registerOutputs_369__10, registerOutputs_369__9, registerOutputs_369__8, 
         registerOutputs_369__7, registerOutputs_369__6, registerOutputs_369__5, 
         registerOutputs_369__4, registerOutputs_369__3, registerOutputs_369__2, 
         registerOutputs_369__1, registerOutputs_369__0, registerOutputs_370__15, 
         registerOutputs_370__14, registerOutputs_370__13, 
         registerOutputs_370__12, registerOutputs_370__11, 
         registerOutputs_370__10, registerOutputs_370__9, registerOutputs_370__8, 
         registerOutputs_370__7, registerOutputs_370__6, registerOutputs_370__5, 
         registerOutputs_370__4, registerOutputs_370__3, registerOutputs_370__2, 
         registerOutputs_370__1, registerOutputs_370__0, registerOutputs_371__15, 
         registerOutputs_371__14, registerOutputs_371__13, 
         registerOutputs_371__12, registerOutputs_371__11, 
         registerOutputs_371__10, registerOutputs_371__9, registerOutputs_371__8, 
         registerOutputs_371__7, registerOutputs_371__6, registerOutputs_371__5, 
         registerOutputs_371__4, registerOutputs_371__3, registerOutputs_371__2, 
         registerOutputs_371__1, registerOutputs_371__0, registerOutputs_372__15, 
         registerOutputs_372__14, registerOutputs_372__13, 
         registerOutputs_372__12, registerOutputs_372__11, 
         registerOutputs_372__10, registerOutputs_372__9, registerOutputs_372__8, 
         registerOutputs_372__7, registerOutputs_372__6, registerOutputs_372__5, 
         registerOutputs_372__4, registerOutputs_372__3, registerOutputs_372__2, 
         registerOutputs_372__1, registerOutputs_372__0, registerOutputs_373__15, 
         registerOutputs_373__14, registerOutputs_373__13, 
         registerOutputs_373__12, registerOutputs_373__11, 
         registerOutputs_373__10, registerOutputs_373__9, registerOutputs_373__8, 
         registerOutputs_373__7, registerOutputs_373__6, registerOutputs_373__5, 
         registerOutputs_373__4, registerOutputs_373__3, registerOutputs_373__2, 
         registerOutputs_373__1, registerOutputs_373__0, registerOutputs_374__15, 
         registerOutputs_374__14, registerOutputs_374__13, 
         registerOutputs_374__12, registerOutputs_374__11, 
         registerOutputs_374__10, registerOutputs_374__9, registerOutputs_374__8, 
         registerOutputs_374__7, registerOutputs_374__6, registerOutputs_374__5, 
         registerOutputs_374__4, registerOutputs_374__3, registerOutputs_374__2, 
         registerOutputs_374__1, registerOutputs_374__0, registerOutputs_375__15, 
         registerOutputs_375__14, registerOutputs_375__13, 
         registerOutputs_375__12, registerOutputs_375__11, 
         registerOutputs_375__10, registerOutputs_375__9, registerOutputs_375__8, 
         registerOutputs_375__7, registerOutputs_375__6, registerOutputs_375__5, 
         registerOutputs_375__4, registerOutputs_375__3, registerOutputs_375__2, 
         registerOutputs_375__1, registerOutputs_375__0, registerOutputs_376__15, 
         registerOutputs_376__14, registerOutputs_376__13, 
         registerOutputs_376__12, registerOutputs_376__11, 
         registerOutputs_376__10, registerOutputs_376__9, registerOutputs_376__8, 
         registerOutputs_376__7, registerOutputs_376__6, registerOutputs_376__5, 
         registerOutputs_376__4, registerOutputs_376__3, registerOutputs_376__2, 
         registerOutputs_376__1, registerOutputs_376__0, registerOutputs_377__15, 
         registerOutputs_377__14, registerOutputs_377__13, 
         registerOutputs_377__12, registerOutputs_377__11, 
         registerOutputs_377__10, registerOutputs_377__9, registerOutputs_377__8, 
         registerOutputs_377__7, registerOutputs_377__6, registerOutputs_377__5, 
         registerOutputs_377__4, registerOutputs_377__3, registerOutputs_377__2, 
         registerOutputs_377__1, registerOutputs_377__0, registerOutputs_378__15, 
         registerOutputs_378__14, registerOutputs_378__13, 
         registerOutputs_378__12, registerOutputs_378__11, 
         registerOutputs_378__10, registerOutputs_378__9, registerOutputs_378__8, 
         registerOutputs_378__7, registerOutputs_378__6, registerOutputs_378__5, 
         registerOutputs_378__4, registerOutputs_378__3, registerOutputs_378__2, 
         registerOutputs_378__1, registerOutputs_378__0, registerOutputs_379__15, 
         registerOutputs_379__14, registerOutputs_379__13, 
         registerOutputs_379__12, registerOutputs_379__11, 
         registerOutputs_379__10, registerOutputs_379__9, registerOutputs_379__8, 
         registerOutputs_379__7, registerOutputs_379__6, registerOutputs_379__5, 
         registerOutputs_379__4, registerOutputs_379__3, registerOutputs_379__2, 
         registerOutputs_379__1, registerOutputs_379__0, registerOutputs_380__15, 
         registerOutputs_380__14, registerOutputs_380__13, 
         registerOutputs_380__12, registerOutputs_380__11, 
         registerOutputs_380__10, registerOutputs_380__9, registerOutputs_380__8, 
         registerOutputs_380__7, registerOutputs_380__6, registerOutputs_380__5, 
         registerOutputs_380__4, registerOutputs_380__3, registerOutputs_380__2, 
         registerOutputs_380__1, registerOutputs_380__0, registerOutputs_381__15, 
         registerOutputs_381__14, registerOutputs_381__13, 
         registerOutputs_381__12, registerOutputs_381__11, 
         registerOutputs_381__10, registerOutputs_381__9, registerOutputs_381__8, 
         registerOutputs_381__7, registerOutputs_381__6, registerOutputs_381__5, 
         registerOutputs_381__4, registerOutputs_381__3, registerOutputs_381__2, 
         registerOutputs_381__1, registerOutputs_381__0, registerOutputs_382__15, 
         registerOutputs_382__14, registerOutputs_382__13, 
         registerOutputs_382__12, registerOutputs_382__11, 
         registerOutputs_382__10, registerOutputs_382__9, registerOutputs_382__8, 
         registerOutputs_382__7, registerOutputs_382__6, registerOutputs_382__5, 
         registerOutputs_382__4, registerOutputs_382__3, registerOutputs_382__2, 
         registerOutputs_382__1, registerOutputs_382__0, registerOutputs_383__15, 
         registerOutputs_383__14, registerOutputs_383__13, 
         registerOutputs_383__12, registerOutputs_383__11, 
         registerOutputs_383__10, registerOutputs_383__9, registerOutputs_383__8, 
         registerOutputs_383__7, registerOutputs_383__6, registerOutputs_383__5, 
         registerOutputs_383__4, registerOutputs_383__3, registerOutputs_383__2, 
         registerOutputs_383__1, registerOutputs_383__0, registerOutputs_384__15, 
         registerOutputs_384__14, registerOutputs_384__13, 
         registerOutputs_384__12, registerOutputs_384__11, 
         registerOutputs_384__10, registerOutputs_384__9, registerOutputs_384__8, 
         registerOutputs_384__7, registerOutputs_384__6, registerOutputs_384__5, 
         registerOutputs_384__4, registerOutputs_384__3, registerOutputs_384__2, 
         registerOutputs_384__1, registerOutputs_384__0, registerOutputs_385__15, 
         registerOutputs_385__14, registerOutputs_385__13, 
         registerOutputs_385__12, registerOutputs_385__11, 
         registerOutputs_385__10, registerOutputs_385__9, registerOutputs_385__8, 
         registerOutputs_385__7, registerOutputs_385__6, registerOutputs_385__5, 
         registerOutputs_385__4, registerOutputs_385__3, registerOutputs_385__2, 
         registerOutputs_385__1, registerOutputs_385__0, registerOutputs_386__15, 
         registerOutputs_386__14, registerOutputs_386__13, 
         registerOutputs_386__12, registerOutputs_386__11, 
         registerOutputs_386__10, registerOutputs_386__9, registerOutputs_386__8, 
         registerOutputs_386__7, registerOutputs_386__6, registerOutputs_386__5, 
         registerOutputs_386__4, registerOutputs_386__3, registerOutputs_386__2, 
         registerOutputs_386__1, registerOutputs_386__0, registerOutputs_387__15, 
         registerOutputs_387__14, registerOutputs_387__13, 
         registerOutputs_387__12, registerOutputs_387__11, 
         registerOutputs_387__10, registerOutputs_387__9, registerOutputs_387__8, 
         registerOutputs_387__7, registerOutputs_387__6, registerOutputs_387__5, 
         registerOutputs_387__4, registerOutputs_387__3, registerOutputs_387__2, 
         registerOutputs_387__1, registerOutputs_387__0, registerOutputs_388__15, 
         registerOutputs_388__14, registerOutputs_388__13, 
         registerOutputs_388__12, registerOutputs_388__11, 
         registerOutputs_388__10, registerOutputs_388__9, registerOutputs_388__8, 
         registerOutputs_388__7, registerOutputs_388__6, registerOutputs_388__5, 
         registerOutputs_388__4, registerOutputs_388__3, registerOutputs_388__2, 
         registerOutputs_388__1, registerOutputs_388__0, registerOutputs_389__15, 
         registerOutputs_389__14, registerOutputs_389__13, 
         registerOutputs_389__12, registerOutputs_389__11, 
         registerOutputs_389__10, registerOutputs_389__9, registerOutputs_389__8, 
         registerOutputs_389__7, registerOutputs_389__6, registerOutputs_389__5, 
         registerOutputs_389__4, registerOutputs_389__3, registerOutputs_389__2, 
         registerOutputs_389__1, registerOutputs_389__0, registerOutputs_390__15, 
         registerOutputs_390__14, registerOutputs_390__13, 
         registerOutputs_390__12, registerOutputs_390__11, 
         registerOutputs_390__10, registerOutputs_390__9, registerOutputs_390__8, 
         registerOutputs_390__7, registerOutputs_390__6, registerOutputs_390__5, 
         registerOutputs_390__4, registerOutputs_390__3, registerOutputs_390__2, 
         registerOutputs_390__1, registerOutputs_390__0, registerOutputs_391__15, 
         registerOutputs_391__14, registerOutputs_391__13, 
         registerOutputs_391__12, registerOutputs_391__11, 
         registerOutputs_391__10, registerOutputs_391__9, registerOutputs_391__8, 
         registerOutputs_391__7, registerOutputs_391__6, registerOutputs_391__5, 
         registerOutputs_391__4, registerOutputs_391__3, registerOutputs_391__2, 
         registerOutputs_391__1, registerOutputs_391__0, registerOutputs_392__15, 
         registerOutputs_392__14, registerOutputs_392__13, 
         registerOutputs_392__12, registerOutputs_392__11, 
         registerOutputs_392__10, registerOutputs_392__9, registerOutputs_392__8, 
         registerOutputs_392__7, registerOutputs_392__6, registerOutputs_392__5, 
         registerOutputs_392__4, registerOutputs_392__3, registerOutputs_392__2, 
         registerOutputs_392__1, registerOutputs_392__0, registerOutputs_393__15, 
         registerOutputs_393__14, registerOutputs_393__13, 
         registerOutputs_393__12, registerOutputs_393__11, 
         registerOutputs_393__10, registerOutputs_393__9, registerOutputs_393__8, 
         registerOutputs_393__7, registerOutputs_393__6, registerOutputs_393__5, 
         registerOutputs_393__4, registerOutputs_393__3, registerOutputs_393__2, 
         registerOutputs_393__1, registerOutputs_393__0, registerOutputs_394__15, 
         registerOutputs_394__14, registerOutputs_394__13, 
         registerOutputs_394__12, registerOutputs_394__11, 
         registerOutputs_394__10, registerOutputs_394__9, registerOutputs_394__8, 
         registerOutputs_394__7, registerOutputs_394__6, registerOutputs_394__5, 
         registerOutputs_394__4, registerOutputs_394__3, registerOutputs_394__2, 
         registerOutputs_394__1, registerOutputs_394__0, registerOutputs_395__15, 
         registerOutputs_395__14, registerOutputs_395__13, 
         registerOutputs_395__12, registerOutputs_395__11, 
         registerOutputs_395__10, registerOutputs_395__9, registerOutputs_395__8, 
         registerOutputs_395__7, registerOutputs_395__6, registerOutputs_395__5, 
         registerOutputs_395__4, registerOutputs_395__3, registerOutputs_395__2, 
         registerOutputs_395__1, registerOutputs_395__0, registerOutputs_396__15, 
         registerOutputs_396__14, registerOutputs_396__13, 
         registerOutputs_396__12, registerOutputs_396__11, 
         registerOutputs_396__10, registerOutputs_396__9, registerOutputs_396__8, 
         registerOutputs_396__7, registerOutputs_396__6, registerOutputs_396__5, 
         registerOutputs_396__4, registerOutputs_396__3, registerOutputs_396__2, 
         registerOutputs_396__1, registerOutputs_396__0, registerOutputs_397__15, 
         registerOutputs_397__14, registerOutputs_397__13, 
         registerOutputs_397__12, registerOutputs_397__11, 
         registerOutputs_397__10, registerOutputs_397__9, registerOutputs_397__8, 
         registerOutputs_397__7, registerOutputs_397__6, registerOutputs_397__5, 
         registerOutputs_397__4, registerOutputs_397__3, registerOutputs_397__2, 
         registerOutputs_397__1, registerOutputs_397__0, registerOutputs_398__15, 
         registerOutputs_398__14, registerOutputs_398__13, 
         registerOutputs_398__12, registerOutputs_398__11, 
         registerOutputs_398__10, registerOutputs_398__9, registerOutputs_398__8, 
         registerOutputs_398__7, registerOutputs_398__6, registerOutputs_398__5, 
         registerOutputs_398__4, registerOutputs_398__3, registerOutputs_398__2, 
         registerOutputs_398__1, registerOutputs_398__0, registerOutputs_399__15, 
         registerOutputs_399__14, registerOutputs_399__13, 
         registerOutputs_399__12, registerOutputs_399__11, 
         registerOutputs_399__10, registerOutputs_399__9, registerOutputs_399__8, 
         registerOutputs_399__7, registerOutputs_399__6, registerOutputs_399__5, 
         registerOutputs_399__4, registerOutputs_399__3, registerOutputs_399__2, 
         registerOutputs_399__1, registerOutputs_399__0, registerOutputs_400__15, 
         registerOutputs_400__14, registerOutputs_400__13, 
         registerOutputs_400__12, registerOutputs_400__11, 
         registerOutputs_400__10, registerOutputs_400__9, registerOutputs_400__8, 
         registerOutputs_400__7, registerOutputs_400__6, registerOutputs_400__5, 
         registerOutputs_400__4, registerOutputs_400__3, registerOutputs_400__2, 
         registerOutputs_400__1, registerOutputs_400__0, registerOutputs_401__15, 
         registerOutputs_401__14, registerOutputs_401__13, 
         registerOutputs_401__12, registerOutputs_401__11, 
         registerOutputs_401__10, registerOutputs_401__9, registerOutputs_401__8, 
         registerOutputs_401__7, registerOutputs_401__6, registerOutputs_401__5, 
         registerOutputs_401__4, registerOutputs_401__3, registerOutputs_401__2, 
         registerOutputs_401__1, registerOutputs_401__0, registerOutputs_402__15, 
         registerOutputs_402__14, registerOutputs_402__13, 
         registerOutputs_402__12, registerOutputs_402__11, 
         registerOutputs_402__10, registerOutputs_402__9, registerOutputs_402__8, 
         registerOutputs_402__7, registerOutputs_402__6, registerOutputs_402__5, 
         registerOutputs_402__4, registerOutputs_402__3, registerOutputs_402__2, 
         registerOutputs_402__1, registerOutputs_402__0, registerOutputs_403__15, 
         registerOutputs_403__14, registerOutputs_403__13, 
         registerOutputs_403__12, registerOutputs_403__11, 
         registerOutputs_403__10, registerOutputs_403__9, registerOutputs_403__8, 
         registerOutputs_403__7, registerOutputs_403__6, registerOutputs_403__5, 
         registerOutputs_403__4, registerOutputs_403__3, registerOutputs_403__2, 
         registerOutputs_403__1, registerOutputs_403__0, registerOutputs_404__15, 
         registerOutputs_404__14, registerOutputs_404__13, 
         registerOutputs_404__12, registerOutputs_404__11, 
         registerOutputs_404__10, registerOutputs_404__9, registerOutputs_404__8, 
         registerOutputs_404__7, registerOutputs_404__6, registerOutputs_404__5, 
         registerOutputs_404__4, registerOutputs_404__3, registerOutputs_404__2, 
         registerOutputs_404__1, registerOutputs_404__0, registerOutputs_405__15, 
         registerOutputs_405__14, registerOutputs_405__13, 
         registerOutputs_405__12, registerOutputs_405__11, 
         registerOutputs_405__10, registerOutputs_405__9, registerOutputs_405__8, 
         registerOutputs_405__7, registerOutputs_405__6, registerOutputs_405__5, 
         registerOutputs_405__4, registerOutputs_405__3, registerOutputs_405__2, 
         registerOutputs_405__1, registerOutputs_405__0, registerOutputs_406__15, 
         registerOutputs_406__14, registerOutputs_406__13, 
         registerOutputs_406__12, registerOutputs_406__11, 
         registerOutputs_406__10, registerOutputs_406__9, registerOutputs_406__8, 
         registerOutputs_406__7, registerOutputs_406__6, registerOutputs_406__5, 
         registerOutputs_406__4, registerOutputs_406__3, registerOutputs_406__2, 
         registerOutputs_406__1, registerOutputs_406__0, registerOutputs_407__15, 
         registerOutputs_407__14, registerOutputs_407__13, 
         registerOutputs_407__12, registerOutputs_407__11, 
         registerOutputs_407__10, registerOutputs_407__9, registerOutputs_407__8, 
         registerOutputs_407__7, registerOutputs_407__6, registerOutputs_407__5, 
         registerOutputs_407__4, registerOutputs_407__3, registerOutputs_407__2, 
         registerOutputs_407__1, registerOutputs_407__0, registerOutputs_408__15, 
         registerOutputs_408__14, registerOutputs_408__13, 
         registerOutputs_408__12, registerOutputs_408__11, 
         registerOutputs_408__10, registerOutputs_408__9, registerOutputs_408__8, 
         registerOutputs_408__7, registerOutputs_408__6, registerOutputs_408__5, 
         registerOutputs_408__4, registerOutputs_408__3, registerOutputs_408__2, 
         registerOutputs_408__1, registerOutputs_408__0, registerOutputs_409__15, 
         registerOutputs_409__14, registerOutputs_409__13, 
         registerOutputs_409__12, registerOutputs_409__11, 
         registerOutputs_409__10, registerOutputs_409__9, registerOutputs_409__8, 
         registerOutputs_409__7, registerOutputs_409__6, registerOutputs_409__5, 
         registerOutputs_409__4, registerOutputs_409__3, registerOutputs_409__2, 
         registerOutputs_409__1, registerOutputs_409__0, registerOutputs_410__15, 
         registerOutputs_410__14, registerOutputs_410__13, 
         registerOutputs_410__12, registerOutputs_410__11, 
         registerOutputs_410__10, registerOutputs_410__9, registerOutputs_410__8, 
         registerOutputs_410__7, registerOutputs_410__6, registerOutputs_410__5, 
         registerOutputs_410__4, registerOutputs_410__3, registerOutputs_410__2, 
         registerOutputs_410__1, registerOutputs_410__0, registerOutputs_411__15, 
         registerOutputs_411__14, registerOutputs_411__13, 
         registerOutputs_411__12, registerOutputs_411__11, 
         registerOutputs_411__10, registerOutputs_411__9, registerOutputs_411__8, 
         registerOutputs_411__7, registerOutputs_411__6, registerOutputs_411__5, 
         registerOutputs_411__4, registerOutputs_411__3, registerOutputs_411__2, 
         registerOutputs_411__1, registerOutputs_411__0, registerOutputs_412__15, 
         registerOutputs_412__14, registerOutputs_412__13, 
         registerOutputs_412__12, registerOutputs_412__11, 
         registerOutputs_412__10, registerOutputs_412__9, registerOutputs_412__8, 
         registerOutputs_412__7, registerOutputs_412__6, registerOutputs_412__5, 
         registerOutputs_412__4, registerOutputs_412__3, registerOutputs_412__2, 
         registerOutputs_412__1, registerOutputs_412__0, registerOutputs_413__15, 
         registerOutputs_413__14, registerOutputs_413__13, 
         registerOutputs_413__12, registerOutputs_413__11, 
         registerOutputs_413__10, registerOutputs_413__9, registerOutputs_413__8, 
         registerOutputs_413__7, registerOutputs_413__6, registerOutputs_413__5, 
         registerOutputs_413__4, registerOutputs_413__3, registerOutputs_413__2, 
         registerOutputs_413__1, registerOutputs_413__0, registerOutputs_414__15, 
         registerOutputs_414__14, registerOutputs_414__13, 
         registerOutputs_414__12, registerOutputs_414__11, 
         registerOutputs_414__10, registerOutputs_414__9, registerOutputs_414__8, 
         registerOutputs_414__7, registerOutputs_414__6, registerOutputs_414__5, 
         registerOutputs_414__4, registerOutputs_414__3, registerOutputs_414__2, 
         registerOutputs_414__1, registerOutputs_414__0, registerOutputs_415__15, 
         registerOutputs_415__14, registerOutputs_415__13, 
         registerOutputs_415__12, registerOutputs_415__11, 
         registerOutputs_415__10, registerOutputs_415__9, registerOutputs_415__8, 
         registerOutputs_415__7, registerOutputs_415__6, registerOutputs_415__5, 
         registerOutputs_415__4, registerOutputs_415__3, registerOutputs_415__2, 
         registerOutputs_415__1, registerOutputs_415__0, registerOutputs_416__15, 
         registerOutputs_416__14, registerOutputs_416__13, 
         registerOutputs_416__12, registerOutputs_416__11, 
         registerOutputs_416__10, registerOutputs_416__9, registerOutputs_416__8, 
         registerOutputs_416__7, registerOutputs_416__6, registerOutputs_416__5, 
         registerOutputs_416__4, registerOutputs_416__3, registerOutputs_416__2, 
         registerOutputs_416__1, registerOutputs_416__0, registerOutputs_417__15, 
         registerOutputs_417__14, registerOutputs_417__13, 
         registerOutputs_417__12, registerOutputs_417__11, 
         registerOutputs_417__10, registerOutputs_417__9, registerOutputs_417__8, 
         registerOutputs_417__7, registerOutputs_417__6, registerOutputs_417__5, 
         registerOutputs_417__4, registerOutputs_417__3, registerOutputs_417__2, 
         registerOutputs_417__1, registerOutputs_417__0, registerOutputs_418__15, 
         registerOutputs_418__14, registerOutputs_418__13, 
         registerOutputs_418__12, registerOutputs_418__11, 
         registerOutputs_418__10, registerOutputs_418__9, registerOutputs_418__8, 
         registerOutputs_418__7, registerOutputs_418__6, registerOutputs_418__5, 
         registerOutputs_418__4, registerOutputs_418__3, registerOutputs_418__2, 
         registerOutputs_418__1, registerOutputs_418__0, registerOutputs_419__15, 
         registerOutputs_419__14, registerOutputs_419__13, 
         registerOutputs_419__12, registerOutputs_419__11, 
         registerOutputs_419__10, registerOutputs_419__9, registerOutputs_419__8, 
         registerOutputs_419__7, registerOutputs_419__6, registerOutputs_419__5, 
         registerOutputs_419__4, registerOutputs_419__3, registerOutputs_419__2, 
         registerOutputs_419__1, registerOutputs_419__0, registerOutputs_420__15, 
         registerOutputs_420__14, registerOutputs_420__13, 
         registerOutputs_420__12, registerOutputs_420__11, 
         registerOutputs_420__10, registerOutputs_420__9, registerOutputs_420__8, 
         registerOutputs_420__7, registerOutputs_420__6, registerOutputs_420__5, 
         registerOutputs_420__4, registerOutputs_420__3, registerOutputs_420__2, 
         registerOutputs_420__1, registerOutputs_420__0, registerOutputs_421__15, 
         registerOutputs_421__14, registerOutputs_421__13, 
         registerOutputs_421__12, registerOutputs_421__11, 
         registerOutputs_421__10, registerOutputs_421__9, registerOutputs_421__8, 
         registerOutputs_421__7, registerOutputs_421__6, registerOutputs_421__5, 
         registerOutputs_421__4, registerOutputs_421__3, registerOutputs_421__2, 
         registerOutputs_421__1, registerOutputs_421__0, registerOutputs_422__15, 
         registerOutputs_422__14, registerOutputs_422__13, 
         registerOutputs_422__12, registerOutputs_422__11, 
         registerOutputs_422__10, registerOutputs_422__9, registerOutputs_422__8, 
         registerOutputs_422__7, registerOutputs_422__6, registerOutputs_422__5, 
         registerOutputs_422__4, registerOutputs_422__3, registerOutputs_422__2, 
         registerOutputs_422__1, registerOutputs_422__0, registerOutputs_423__15, 
         registerOutputs_423__14, registerOutputs_423__13, 
         registerOutputs_423__12, registerOutputs_423__11, 
         registerOutputs_423__10, registerOutputs_423__9, registerOutputs_423__8, 
         registerOutputs_423__7, registerOutputs_423__6, registerOutputs_423__5, 
         registerOutputs_423__4, registerOutputs_423__3, registerOutputs_423__2, 
         registerOutputs_423__1, registerOutputs_423__0, registerOutputs_424__15, 
         registerOutputs_424__14, registerOutputs_424__13, 
         registerOutputs_424__12, registerOutputs_424__11, 
         registerOutputs_424__10, registerOutputs_424__9, registerOutputs_424__8, 
         registerOutputs_424__7, registerOutputs_424__6, registerOutputs_424__5, 
         registerOutputs_424__4, registerOutputs_424__3, registerOutputs_424__2, 
         registerOutputs_424__1, registerOutputs_424__0, registerOutputs_425__15, 
         registerOutputs_425__14, registerOutputs_425__13, 
         registerOutputs_425__12, registerOutputs_425__11, 
         registerOutputs_425__10, registerOutputs_425__9, registerOutputs_425__8, 
         registerOutputs_425__7, registerOutputs_425__6, registerOutputs_425__5, 
         registerOutputs_425__4, registerOutputs_425__3, registerOutputs_425__2, 
         registerOutputs_425__1, registerOutputs_425__0, registerOutputs_426__15, 
         registerOutputs_426__14, registerOutputs_426__13, 
         registerOutputs_426__12, registerOutputs_426__11, 
         registerOutputs_426__10, registerOutputs_426__9, registerOutputs_426__8, 
         registerOutputs_426__7, registerOutputs_426__6, registerOutputs_426__5, 
         registerOutputs_426__4, registerOutputs_426__3, registerOutputs_426__2, 
         registerOutputs_426__1, registerOutputs_426__0, registerOutputs_427__15, 
         registerOutputs_427__14, registerOutputs_427__13, 
         registerOutputs_427__12, registerOutputs_427__11, 
         registerOutputs_427__10, registerOutputs_427__9, registerOutputs_427__8, 
         registerOutputs_427__7, registerOutputs_427__6, registerOutputs_427__5, 
         registerOutputs_427__4, registerOutputs_427__3, registerOutputs_427__2, 
         registerOutputs_427__1, registerOutputs_427__0, registerOutputs_428__15, 
         registerOutputs_428__14, registerOutputs_428__13, 
         registerOutputs_428__12, registerOutputs_428__11, 
         registerOutputs_428__10, registerOutputs_428__9, registerOutputs_428__8, 
         registerOutputs_428__7, registerOutputs_428__6, registerOutputs_428__5, 
         registerOutputs_428__4, registerOutputs_428__3, registerOutputs_428__2, 
         registerOutputs_428__1, registerOutputs_428__0, registerOutputs_429__15, 
         registerOutputs_429__14, registerOutputs_429__13, 
         registerOutputs_429__12, registerOutputs_429__11, 
         registerOutputs_429__10, registerOutputs_429__9, registerOutputs_429__8, 
         registerOutputs_429__7, registerOutputs_429__6, registerOutputs_429__5, 
         registerOutputs_429__4, registerOutputs_429__3, registerOutputs_429__2, 
         registerOutputs_429__1, registerOutputs_429__0, registerOutputs_430__15, 
         registerOutputs_430__14, registerOutputs_430__13, 
         registerOutputs_430__12, registerOutputs_430__11, 
         registerOutputs_430__10, registerOutputs_430__9, registerOutputs_430__8, 
         registerOutputs_430__7, registerOutputs_430__6, registerOutputs_430__5, 
         registerOutputs_430__4, registerOutputs_430__3, registerOutputs_430__2, 
         registerOutputs_430__1, registerOutputs_430__0, registerOutputs_431__15, 
         registerOutputs_431__14, registerOutputs_431__13, 
         registerOutputs_431__12, registerOutputs_431__11, 
         registerOutputs_431__10, registerOutputs_431__9, registerOutputs_431__8, 
         registerOutputs_431__7, registerOutputs_431__6, registerOutputs_431__5, 
         registerOutputs_431__4, registerOutputs_431__3, registerOutputs_431__2, 
         registerOutputs_431__1, registerOutputs_431__0, registerOutputs_432__15, 
         registerOutputs_432__14, registerOutputs_432__13, 
         registerOutputs_432__12, registerOutputs_432__11, 
         registerOutputs_432__10, registerOutputs_432__9, registerOutputs_432__8, 
         registerOutputs_432__7, registerOutputs_432__6, registerOutputs_432__5, 
         registerOutputs_432__4, registerOutputs_432__3, registerOutputs_432__2, 
         registerOutputs_432__1, registerOutputs_432__0, registerOutputs_433__15, 
         registerOutputs_433__14, registerOutputs_433__13, 
         registerOutputs_433__12, registerOutputs_433__11, 
         registerOutputs_433__10, registerOutputs_433__9, registerOutputs_433__8, 
         registerOutputs_433__7, registerOutputs_433__6, registerOutputs_433__5, 
         registerOutputs_433__4, registerOutputs_433__3, registerOutputs_433__2, 
         registerOutputs_433__1, registerOutputs_433__0, registerOutputs_434__15, 
         registerOutputs_434__14, registerOutputs_434__13, 
         registerOutputs_434__12, registerOutputs_434__11, 
         registerOutputs_434__10, registerOutputs_434__9, registerOutputs_434__8, 
         registerOutputs_434__7, registerOutputs_434__6, registerOutputs_434__5, 
         registerOutputs_434__4, registerOutputs_434__3, registerOutputs_434__2, 
         registerOutputs_434__1, registerOutputs_434__0, registerOutputs_435__15, 
         registerOutputs_435__14, registerOutputs_435__13, 
         registerOutputs_435__12, registerOutputs_435__11, 
         registerOutputs_435__10, registerOutputs_435__9, registerOutputs_435__8, 
         registerOutputs_435__7, registerOutputs_435__6, registerOutputs_435__5, 
         registerOutputs_435__4, registerOutputs_435__3, registerOutputs_435__2, 
         registerOutputs_435__1, registerOutputs_435__0, registerOutputs_436__15, 
         registerOutputs_436__14, registerOutputs_436__13, 
         registerOutputs_436__12, registerOutputs_436__11, 
         registerOutputs_436__10, registerOutputs_436__9, registerOutputs_436__8, 
         registerOutputs_436__7, registerOutputs_436__6, registerOutputs_436__5, 
         registerOutputs_436__4, registerOutputs_436__3, registerOutputs_436__2, 
         registerOutputs_436__1, registerOutputs_436__0, registerOutputs_437__15, 
         registerOutputs_437__14, registerOutputs_437__13, 
         registerOutputs_437__12, registerOutputs_437__11, 
         registerOutputs_437__10, registerOutputs_437__9, registerOutputs_437__8, 
         registerOutputs_437__7, registerOutputs_437__6, registerOutputs_437__5, 
         registerOutputs_437__4, registerOutputs_437__3, registerOutputs_437__2, 
         registerOutputs_437__1, registerOutputs_437__0, registerOutputs_438__15, 
         registerOutputs_438__14, registerOutputs_438__13, 
         registerOutputs_438__12, registerOutputs_438__11, 
         registerOutputs_438__10, registerOutputs_438__9, registerOutputs_438__8, 
         registerOutputs_438__7, registerOutputs_438__6, registerOutputs_438__5, 
         registerOutputs_438__4, registerOutputs_438__3, registerOutputs_438__2, 
         registerOutputs_438__1, registerOutputs_438__0, registerOutputs_439__15, 
         registerOutputs_439__14, registerOutputs_439__13, 
         registerOutputs_439__12, registerOutputs_439__11, 
         registerOutputs_439__10, registerOutputs_439__9, registerOutputs_439__8, 
         registerOutputs_439__7, registerOutputs_439__6, registerOutputs_439__5, 
         registerOutputs_439__4, registerOutputs_439__3, registerOutputs_439__2, 
         registerOutputs_439__1, registerOutputs_439__0, registerOutputs_440__15, 
         registerOutputs_440__14, registerOutputs_440__13, 
         registerOutputs_440__12, registerOutputs_440__11, 
         registerOutputs_440__10, registerOutputs_440__9, registerOutputs_440__8, 
         registerOutputs_440__7, registerOutputs_440__6, registerOutputs_440__5, 
         registerOutputs_440__4, registerOutputs_440__3, registerOutputs_440__2, 
         registerOutputs_440__1, registerOutputs_440__0, registerOutputs_441__15, 
         registerOutputs_441__14, registerOutputs_441__13, 
         registerOutputs_441__12, registerOutputs_441__11, 
         registerOutputs_441__10, registerOutputs_441__9, registerOutputs_441__8, 
         registerOutputs_441__7, registerOutputs_441__6, registerOutputs_441__5, 
         registerOutputs_441__4, registerOutputs_441__3, registerOutputs_441__2, 
         registerOutputs_441__1, registerOutputs_441__0, registerOutputs_442__15, 
         registerOutputs_442__14, registerOutputs_442__13, 
         registerOutputs_442__12, registerOutputs_442__11, 
         registerOutputs_442__10, registerOutputs_442__9, registerOutputs_442__8, 
         registerOutputs_442__7, registerOutputs_442__6, registerOutputs_442__5, 
         registerOutputs_442__4, registerOutputs_442__3, registerOutputs_442__2, 
         registerOutputs_442__1, registerOutputs_442__0, registerOutputs_443__15, 
         registerOutputs_443__14, registerOutputs_443__13, 
         registerOutputs_443__12, registerOutputs_443__11, 
         registerOutputs_443__10, registerOutputs_443__9, registerOutputs_443__8, 
         registerOutputs_443__7, registerOutputs_443__6, registerOutputs_443__5, 
         registerOutputs_443__4, registerOutputs_443__3, registerOutputs_443__2, 
         registerOutputs_443__1, registerOutputs_443__0, registerOutputs_444__15, 
         registerOutputs_444__14, registerOutputs_444__13, 
         registerOutputs_444__12, registerOutputs_444__11, 
         registerOutputs_444__10, registerOutputs_444__9, registerOutputs_444__8, 
         registerOutputs_444__7, registerOutputs_444__6, registerOutputs_444__5, 
         registerOutputs_444__4, registerOutputs_444__3, registerOutputs_444__2, 
         registerOutputs_444__1, registerOutputs_444__0, registerOutputs_445__15, 
         registerOutputs_445__14, registerOutputs_445__13, 
         registerOutputs_445__12, registerOutputs_445__11, 
         registerOutputs_445__10, registerOutputs_445__9, registerOutputs_445__8, 
         registerOutputs_445__7, registerOutputs_445__6, registerOutputs_445__5, 
         registerOutputs_445__4, registerOutputs_445__3, registerOutputs_445__2, 
         registerOutputs_445__1, registerOutputs_445__0, registerOutputs_446__15, 
         registerOutputs_446__14, registerOutputs_446__13, 
         registerOutputs_446__12, registerOutputs_446__11, 
         registerOutputs_446__10, registerOutputs_446__9, registerOutputs_446__8, 
         registerOutputs_446__7, registerOutputs_446__6, registerOutputs_446__5, 
         registerOutputs_446__4, registerOutputs_446__3, registerOutputs_446__2, 
         registerOutputs_446__1, registerOutputs_446__0, registerOutputs_447__15, 
         registerOutputs_447__14, registerOutputs_447__13, 
         registerOutputs_447__12, registerOutputs_447__11, 
         registerOutputs_447__10, registerOutputs_447__9, registerOutputs_447__8, 
         registerOutputs_447__7, registerOutputs_447__6, registerOutputs_447__5, 
         registerOutputs_447__4, registerOutputs_447__3, registerOutputs_447__2, 
         registerOutputs_447__1, registerOutputs_447__0, registerOutputs_448__15, 
         registerOutputs_448__14, registerOutputs_448__13, 
         registerOutputs_448__12, registerOutputs_448__11, 
         registerOutputs_448__10, registerOutputs_448__9, registerOutputs_448__8, 
         registerOutputs_448__7, registerOutputs_448__6, registerOutputs_448__5, 
         registerOutputs_448__4, registerOutputs_448__3, registerOutputs_448__2, 
         registerOutputs_448__1, registerOutputs_448__0, registerOutputs_449__15, 
         registerOutputs_449__14, registerOutputs_449__13, 
         registerOutputs_449__12, registerOutputs_449__11, 
         registerOutputs_449__10, registerOutputs_449__9, registerOutputs_449__8, 
         registerOutputs_449__7, registerOutputs_449__6, registerOutputs_449__5, 
         registerOutputs_449__4, registerOutputs_449__3, registerOutputs_449__2, 
         registerOutputs_449__1, registerOutputs_449__0, registerOutputs_450__15, 
         registerOutputs_450__14, registerOutputs_450__13, 
         registerOutputs_450__12, registerOutputs_450__11, 
         registerOutputs_450__10, registerOutputs_450__9, registerOutputs_450__8, 
         registerOutputs_450__7, registerOutputs_450__6, registerOutputs_450__5, 
         registerOutputs_450__4, registerOutputs_450__3, registerOutputs_450__2, 
         registerOutputs_450__1, registerOutputs_450__0, registerOutputs_451__15, 
         registerOutputs_451__14, registerOutputs_451__13, 
         registerOutputs_451__12, registerOutputs_451__11, 
         registerOutputs_451__10, registerOutputs_451__9, registerOutputs_451__8, 
         registerOutputs_451__7, registerOutputs_451__6, registerOutputs_451__5, 
         registerOutputs_451__4, registerOutputs_451__3, registerOutputs_451__2, 
         registerOutputs_451__1, registerOutputs_451__0, registerOutputs_452__15, 
         registerOutputs_452__14, registerOutputs_452__13, 
         registerOutputs_452__12, registerOutputs_452__11, 
         registerOutputs_452__10, registerOutputs_452__9, registerOutputs_452__8, 
         registerOutputs_452__7, registerOutputs_452__6, registerOutputs_452__5, 
         registerOutputs_452__4, registerOutputs_452__3, registerOutputs_452__2, 
         registerOutputs_452__1, registerOutputs_452__0, registerOutputs_453__15, 
         registerOutputs_453__14, registerOutputs_453__13, 
         registerOutputs_453__12, registerOutputs_453__11, 
         registerOutputs_453__10, registerOutputs_453__9, registerOutputs_453__8, 
         registerOutputs_453__7, registerOutputs_453__6, registerOutputs_453__5, 
         registerOutputs_453__4, registerOutputs_453__3, registerOutputs_453__2, 
         registerOutputs_453__1, registerOutputs_453__0, registerOutputs_454__15, 
         registerOutputs_454__14, registerOutputs_454__13, 
         registerOutputs_454__12, registerOutputs_454__11, 
         registerOutputs_454__10, registerOutputs_454__9, registerOutputs_454__8, 
         registerOutputs_454__7, registerOutputs_454__6, registerOutputs_454__5, 
         registerOutputs_454__4, registerOutputs_454__3, registerOutputs_454__2, 
         registerOutputs_454__1, registerOutputs_454__0, registerOutputs_455__15, 
         registerOutputs_455__14, registerOutputs_455__13, 
         registerOutputs_455__12, registerOutputs_455__11, 
         registerOutputs_455__10, registerOutputs_455__9, registerOutputs_455__8, 
         registerOutputs_455__7, registerOutputs_455__6, registerOutputs_455__5, 
         registerOutputs_455__4, registerOutputs_455__3, registerOutputs_455__2, 
         registerOutputs_455__1, registerOutputs_455__0, registerOutputs_456__15, 
         registerOutputs_456__14, registerOutputs_456__13, 
         registerOutputs_456__12, registerOutputs_456__11, 
         registerOutputs_456__10, registerOutputs_456__9, registerOutputs_456__8, 
         registerOutputs_456__7, registerOutputs_456__6, registerOutputs_456__5, 
         registerOutputs_456__4, registerOutputs_456__3, registerOutputs_456__2, 
         registerOutputs_456__1, registerOutputs_456__0, registerOutputs_457__15, 
         registerOutputs_457__14, registerOutputs_457__13, 
         registerOutputs_457__12, registerOutputs_457__11, 
         registerOutputs_457__10, registerOutputs_457__9, registerOutputs_457__8, 
         registerOutputs_457__7, registerOutputs_457__6, registerOutputs_457__5, 
         registerOutputs_457__4, registerOutputs_457__3, registerOutputs_457__2, 
         registerOutputs_457__1, registerOutputs_457__0, registerOutputs_458__15, 
         registerOutputs_458__14, registerOutputs_458__13, 
         registerOutputs_458__12, registerOutputs_458__11, 
         registerOutputs_458__10, registerOutputs_458__9, registerOutputs_458__8, 
         registerOutputs_458__7, registerOutputs_458__6, registerOutputs_458__5, 
         registerOutputs_458__4, registerOutputs_458__3, registerOutputs_458__2, 
         registerOutputs_458__1, registerOutputs_458__0, registerOutputs_459__15, 
         registerOutputs_459__14, registerOutputs_459__13, 
         registerOutputs_459__12, registerOutputs_459__11, 
         registerOutputs_459__10, registerOutputs_459__9, registerOutputs_459__8, 
         registerOutputs_459__7, registerOutputs_459__6, registerOutputs_459__5, 
         registerOutputs_459__4, registerOutputs_459__3, registerOutputs_459__2, 
         registerOutputs_459__1, registerOutputs_459__0, registerOutputs_460__15, 
         registerOutputs_460__14, registerOutputs_460__13, 
         registerOutputs_460__12, registerOutputs_460__11, 
         registerOutputs_460__10, registerOutputs_460__9, registerOutputs_460__8, 
         registerOutputs_460__7, registerOutputs_460__6, registerOutputs_460__5, 
         registerOutputs_460__4, registerOutputs_460__3, registerOutputs_460__2, 
         registerOutputs_460__1, registerOutputs_460__0, registerOutputs_461__15, 
         registerOutputs_461__14, registerOutputs_461__13, 
         registerOutputs_461__12, registerOutputs_461__11, 
         registerOutputs_461__10, registerOutputs_461__9, registerOutputs_461__8, 
         registerOutputs_461__7, registerOutputs_461__6, registerOutputs_461__5, 
         registerOutputs_461__4, registerOutputs_461__3, registerOutputs_461__2, 
         registerOutputs_461__1, registerOutputs_461__0, registerOutputs_462__15, 
         registerOutputs_462__14, registerOutputs_462__13, 
         registerOutputs_462__12, registerOutputs_462__11, 
         registerOutputs_462__10, registerOutputs_462__9, registerOutputs_462__8, 
         registerOutputs_462__7, registerOutputs_462__6, registerOutputs_462__5, 
         registerOutputs_462__4, registerOutputs_462__3, registerOutputs_462__2, 
         registerOutputs_462__1, registerOutputs_462__0, registerOutputs_463__15, 
         registerOutputs_463__14, registerOutputs_463__13, 
         registerOutputs_463__12, registerOutputs_463__11, 
         registerOutputs_463__10, registerOutputs_463__9, registerOutputs_463__8, 
         registerOutputs_463__7, registerOutputs_463__6, registerOutputs_463__5, 
         registerOutputs_463__4, registerOutputs_463__3, registerOutputs_463__2, 
         registerOutputs_463__1, registerOutputs_463__0, registerOutputs_464__15, 
         registerOutputs_464__14, registerOutputs_464__13, 
         registerOutputs_464__12, registerOutputs_464__11, 
         registerOutputs_464__10, registerOutputs_464__9, registerOutputs_464__8, 
         registerOutputs_464__7, registerOutputs_464__6, registerOutputs_464__5, 
         registerOutputs_464__4, registerOutputs_464__3, registerOutputs_464__2, 
         registerOutputs_464__1, registerOutputs_464__0, registerOutputs_465__15, 
         registerOutputs_465__14, registerOutputs_465__13, 
         registerOutputs_465__12, registerOutputs_465__11, 
         registerOutputs_465__10, registerOutputs_465__9, registerOutputs_465__8, 
         registerOutputs_465__7, registerOutputs_465__6, registerOutputs_465__5, 
         registerOutputs_465__4, registerOutputs_465__3, registerOutputs_465__2, 
         registerOutputs_465__1, registerOutputs_465__0, registerOutputs_466__15, 
         registerOutputs_466__14, registerOutputs_466__13, 
         registerOutputs_466__12, registerOutputs_466__11, 
         registerOutputs_466__10, registerOutputs_466__9, registerOutputs_466__8, 
         registerOutputs_466__7, registerOutputs_466__6, registerOutputs_466__5, 
         registerOutputs_466__4, registerOutputs_466__3, registerOutputs_466__2, 
         registerOutputs_466__1, registerOutputs_466__0, registerOutputs_467__15, 
         registerOutputs_467__14, registerOutputs_467__13, 
         registerOutputs_467__12, registerOutputs_467__11, 
         registerOutputs_467__10, registerOutputs_467__9, registerOutputs_467__8, 
         registerOutputs_467__7, registerOutputs_467__6, registerOutputs_467__5, 
         registerOutputs_467__4, registerOutputs_467__3, registerOutputs_467__2, 
         registerOutputs_467__1, registerOutputs_467__0, registerOutputs_468__15, 
         registerOutputs_468__14, registerOutputs_468__13, 
         registerOutputs_468__12, registerOutputs_468__11, 
         registerOutputs_468__10, registerOutputs_468__9, registerOutputs_468__8, 
         registerOutputs_468__7, registerOutputs_468__6, registerOutputs_468__5, 
         registerOutputs_468__4, registerOutputs_468__3, registerOutputs_468__2, 
         registerOutputs_468__1, registerOutputs_468__0, registerOutputs_469__15, 
         registerOutputs_469__14, registerOutputs_469__13, 
         registerOutputs_469__12, registerOutputs_469__11, 
         registerOutputs_469__10, registerOutputs_469__9, registerOutputs_469__8, 
         registerOutputs_469__7, registerOutputs_469__6, registerOutputs_469__5, 
         registerOutputs_469__4, registerOutputs_469__3, registerOutputs_469__2, 
         registerOutputs_469__1, registerOutputs_469__0, registerOutputs_470__15, 
         registerOutputs_470__14, registerOutputs_470__13, 
         registerOutputs_470__12, registerOutputs_470__11, 
         registerOutputs_470__10, registerOutputs_470__9, registerOutputs_470__8, 
         registerOutputs_470__7, registerOutputs_470__6, registerOutputs_470__5, 
         registerOutputs_470__4, registerOutputs_470__3, registerOutputs_470__2, 
         registerOutputs_470__1, registerOutputs_470__0, registerOutputs_471__15, 
         registerOutputs_471__14, registerOutputs_471__13, 
         registerOutputs_471__12, registerOutputs_471__11, 
         registerOutputs_471__10, registerOutputs_471__9, registerOutputs_471__8, 
         registerOutputs_471__7, registerOutputs_471__6, registerOutputs_471__5, 
         registerOutputs_471__4, registerOutputs_471__3, registerOutputs_471__2, 
         registerOutputs_471__1, registerOutputs_471__0, registerOutputs_472__15, 
         registerOutputs_472__14, registerOutputs_472__13, 
         registerOutputs_472__12, registerOutputs_472__11, 
         registerOutputs_472__10, registerOutputs_472__9, registerOutputs_472__8, 
         registerOutputs_472__7, registerOutputs_472__6, registerOutputs_472__5, 
         registerOutputs_472__4, registerOutputs_472__3, registerOutputs_472__2, 
         registerOutputs_472__1, registerOutputs_472__0, registerOutputs_473__15, 
         registerOutputs_473__14, registerOutputs_473__13, 
         registerOutputs_473__12, registerOutputs_473__11, 
         registerOutputs_473__10, registerOutputs_473__9, registerOutputs_473__8, 
         registerOutputs_473__7, registerOutputs_473__6, registerOutputs_473__5, 
         registerOutputs_473__4, registerOutputs_473__3, registerOutputs_473__2, 
         registerOutputs_473__1, registerOutputs_473__0, registerOutputs_474__15, 
         registerOutputs_474__14, registerOutputs_474__13, 
         registerOutputs_474__12, registerOutputs_474__11, 
         registerOutputs_474__10, registerOutputs_474__9, registerOutputs_474__8, 
         registerOutputs_474__7, registerOutputs_474__6, registerOutputs_474__5, 
         registerOutputs_474__4, registerOutputs_474__3, registerOutputs_474__2, 
         registerOutputs_474__1, registerOutputs_474__0, registerOutputs_475__15, 
         registerOutputs_475__14, registerOutputs_475__13, 
         registerOutputs_475__12, registerOutputs_475__11, 
         registerOutputs_475__10, registerOutputs_475__9, registerOutputs_475__8, 
         registerOutputs_475__7, registerOutputs_475__6, registerOutputs_475__5, 
         registerOutputs_475__4, registerOutputs_475__3, registerOutputs_475__2, 
         registerOutputs_475__1, registerOutputs_475__0, registerOutputs_476__15, 
         registerOutputs_476__14, registerOutputs_476__13, 
         registerOutputs_476__12, registerOutputs_476__11, 
         registerOutputs_476__10, registerOutputs_476__9, registerOutputs_476__8, 
         registerOutputs_476__7, registerOutputs_476__6, registerOutputs_476__5, 
         registerOutputs_476__4, registerOutputs_476__3, registerOutputs_476__2, 
         registerOutputs_476__1, registerOutputs_476__0, registerOutputs_477__15, 
         registerOutputs_477__14, registerOutputs_477__13, 
         registerOutputs_477__12, registerOutputs_477__11, 
         registerOutputs_477__10, registerOutputs_477__9, registerOutputs_477__8, 
         registerOutputs_477__7, registerOutputs_477__6, registerOutputs_477__5, 
         registerOutputs_477__4, registerOutputs_477__3, registerOutputs_477__2, 
         registerOutputs_477__1, registerOutputs_477__0, registerOutputs_478__15, 
         registerOutputs_478__14, registerOutputs_478__13, 
         registerOutputs_478__12, registerOutputs_478__11, 
         registerOutputs_478__10, registerOutputs_478__9, registerOutputs_478__8, 
         registerOutputs_478__7, registerOutputs_478__6, registerOutputs_478__5, 
         registerOutputs_478__4, registerOutputs_478__3, registerOutputs_478__2, 
         registerOutputs_478__1, registerOutputs_478__0, registerOutputs_479__15, 
         registerOutputs_479__14, registerOutputs_479__13, 
         registerOutputs_479__12, registerOutputs_479__11, 
         registerOutputs_479__10, registerOutputs_479__9, registerOutputs_479__8, 
         registerOutputs_479__7, registerOutputs_479__6, registerOutputs_479__5, 
         registerOutputs_479__4, registerOutputs_479__3, registerOutputs_479__2, 
         registerOutputs_479__1, registerOutputs_479__0, registerOutputs_480__15, 
         registerOutputs_480__14, registerOutputs_480__13, 
         registerOutputs_480__12, registerOutputs_480__11, 
         registerOutputs_480__10, registerOutputs_480__9, registerOutputs_480__8, 
         registerOutputs_480__7, registerOutputs_480__6, registerOutputs_480__5, 
         registerOutputs_480__4, registerOutputs_480__3, registerOutputs_480__2, 
         registerOutputs_480__1, registerOutputs_480__0, registerOutputs_481__15, 
         registerOutputs_481__14, registerOutputs_481__13, 
         registerOutputs_481__12, registerOutputs_481__11, 
         registerOutputs_481__10, registerOutputs_481__9, registerOutputs_481__8, 
         registerOutputs_481__7, registerOutputs_481__6, registerOutputs_481__5, 
         registerOutputs_481__4, registerOutputs_481__3, registerOutputs_481__2, 
         registerOutputs_481__1, registerOutputs_481__0, registerOutputs_482__15, 
         registerOutputs_482__14, registerOutputs_482__13, 
         registerOutputs_482__12, registerOutputs_482__11, 
         registerOutputs_482__10, registerOutputs_482__9, registerOutputs_482__8, 
         registerOutputs_482__7, registerOutputs_482__6, registerOutputs_482__5, 
         registerOutputs_482__4, registerOutputs_482__3, registerOutputs_482__2, 
         registerOutputs_482__1, registerOutputs_482__0, registerOutputs_483__15, 
         registerOutputs_483__14, registerOutputs_483__13, 
         registerOutputs_483__12, registerOutputs_483__11, 
         registerOutputs_483__10, registerOutputs_483__9, registerOutputs_483__8, 
         registerOutputs_483__7, registerOutputs_483__6, registerOutputs_483__5, 
         registerOutputs_483__4, registerOutputs_483__3, registerOutputs_483__2, 
         registerOutputs_483__1, registerOutputs_483__0, inputRegisters_0__15, 
         inputRegisters_0__14, inputRegisters_0__13, inputRegisters_0__12, 
         inputRegisters_0__11, inputRegisters_0__10, inputRegisters_0__9, 
         inputRegisters_0__8, inputRegisters_0__7, inputRegisters_0__6, 
         inputRegisters_0__5, inputRegisters_0__4, inputRegisters_0__3, 
         inputRegisters_0__2, inputRegisters_0__1, inputRegisters_0__0, 
         inputRegisters_1__15, inputRegisters_1__14, inputRegisters_1__13, 
         inputRegisters_1__12, inputRegisters_1__11, inputRegisters_1__10, 
         inputRegisters_1__9, inputRegisters_1__8, inputRegisters_1__7, 
         inputRegisters_1__6, inputRegisters_1__5, inputRegisters_1__4, 
         inputRegisters_1__3, inputRegisters_1__2, inputRegisters_1__1, 
         inputRegisters_1__0, inputRegisters_2__15, inputRegisters_2__14, 
         inputRegisters_2__13, inputRegisters_2__12, inputRegisters_2__11, 
         inputRegisters_2__10, inputRegisters_2__9, inputRegisters_2__8, 
         inputRegisters_2__7, inputRegisters_2__6, inputRegisters_2__5, 
         inputRegisters_2__4, inputRegisters_2__3, inputRegisters_2__2, 
         inputRegisters_2__1, inputRegisters_2__0, inputRegisters_3__15, 
         inputRegisters_3__14, inputRegisters_3__13, inputRegisters_3__12, 
         inputRegisters_3__11, inputRegisters_3__10, inputRegisters_3__9, 
         inputRegisters_3__8, inputRegisters_3__7, inputRegisters_3__6, 
         inputRegisters_3__5, inputRegisters_3__4, inputRegisters_3__3, 
         inputRegisters_3__2, inputRegisters_3__1, inputRegisters_3__0, 
         inputRegisters_4__15, inputRegisters_4__14, inputRegisters_4__13, 
         inputRegisters_4__12, inputRegisters_4__11, inputRegisters_4__10, 
         inputRegisters_4__9, inputRegisters_4__8, inputRegisters_4__7, 
         inputRegisters_4__6, inputRegisters_4__5, inputRegisters_4__4, 
         inputRegisters_4__3, inputRegisters_4__2, inputRegisters_4__1, 
         inputRegisters_4__0, inputRegisters_5__15, inputRegisters_5__14, 
         inputRegisters_5__13, inputRegisters_5__12, inputRegisters_5__11, 
         inputRegisters_5__10, inputRegisters_5__9, inputRegisters_5__8, 
         inputRegisters_5__7, inputRegisters_5__6, inputRegisters_5__5, 
         inputRegisters_5__4, inputRegisters_5__3, inputRegisters_5__2, 
         inputRegisters_5__1, inputRegisters_5__0, inputRegisters_6__15, 
         inputRegisters_6__14, inputRegisters_6__13, inputRegisters_6__12, 
         inputRegisters_6__11, inputRegisters_6__10, inputRegisters_6__9, 
         inputRegisters_6__8, inputRegisters_6__7, inputRegisters_6__6, 
         inputRegisters_6__5, inputRegisters_6__4, inputRegisters_6__3, 
         inputRegisters_6__2, inputRegisters_6__1, inputRegisters_6__0, 
         inputRegisters_7__15, inputRegisters_7__14, inputRegisters_7__13, 
         inputRegisters_7__12, inputRegisters_7__11, inputRegisters_7__10, 
         inputRegisters_7__9, inputRegisters_7__8, inputRegisters_7__7, 
         inputRegisters_7__6, inputRegisters_7__5, inputRegisters_7__4, 
         inputRegisters_7__3, inputRegisters_7__2, inputRegisters_7__1, 
         inputRegisters_7__0, inputRegisters_8__15, inputRegisters_8__14, 
         inputRegisters_8__13, inputRegisters_8__12, inputRegisters_8__11, 
         inputRegisters_8__10, inputRegisters_8__9, inputRegisters_8__8, 
         inputRegisters_8__7, inputRegisters_8__6, inputRegisters_8__5, 
         inputRegisters_8__4, inputRegisters_8__3, inputRegisters_8__2, 
         inputRegisters_8__1, inputRegisters_8__0, inputRegisters_9__15, 
         inputRegisters_9__14, inputRegisters_9__13, inputRegisters_9__12, 
         inputRegisters_9__11, inputRegisters_9__10, inputRegisters_9__9, 
         inputRegisters_9__8, inputRegisters_9__7, inputRegisters_9__6, 
         inputRegisters_9__5, inputRegisters_9__4, inputRegisters_9__3, 
         inputRegisters_9__2, inputRegisters_9__1, inputRegisters_9__0, 
         inputRegisters_10__15, inputRegisters_10__14, inputRegisters_10__13, 
         inputRegisters_10__12, inputRegisters_10__11, inputRegisters_10__10, 
         inputRegisters_10__9, inputRegisters_10__8, inputRegisters_10__7, 
         inputRegisters_10__6, inputRegisters_10__5, inputRegisters_10__4, 
         inputRegisters_10__3, inputRegisters_10__2, inputRegisters_10__1, 
         inputRegisters_10__0, inputRegisters_11__15, inputRegisters_11__14, 
         inputRegisters_11__13, inputRegisters_11__12, inputRegisters_11__11, 
         inputRegisters_11__10, inputRegisters_11__9, inputRegisters_11__8, 
         inputRegisters_11__7, inputRegisters_11__6, inputRegisters_11__5, 
         inputRegisters_11__4, inputRegisters_11__3, inputRegisters_11__2, 
         inputRegisters_11__1, inputRegisters_11__0, inputRegisters_12__15, 
         inputRegisters_12__14, inputRegisters_12__13, inputRegisters_12__12, 
         inputRegisters_12__11, inputRegisters_12__10, inputRegisters_12__9, 
         inputRegisters_12__8, inputRegisters_12__7, inputRegisters_12__6, 
         inputRegisters_12__5, inputRegisters_12__4, inputRegisters_12__3, 
         inputRegisters_12__2, inputRegisters_12__1, inputRegisters_12__0, 
         inputRegisters_13__15, inputRegisters_13__14, inputRegisters_13__13, 
         inputRegisters_13__12, inputRegisters_13__11, inputRegisters_13__10, 
         inputRegisters_13__9, inputRegisters_13__8, inputRegisters_13__7, 
         inputRegisters_13__6, inputRegisters_13__5, inputRegisters_13__4, 
         inputRegisters_13__3, inputRegisters_13__2, inputRegisters_13__1, 
         inputRegisters_13__0, inputRegisters_14__15, inputRegisters_14__14, 
         inputRegisters_14__13, inputRegisters_14__12, inputRegisters_14__11, 
         inputRegisters_14__10, inputRegisters_14__9, inputRegisters_14__8, 
         inputRegisters_14__7, inputRegisters_14__6, inputRegisters_14__5, 
         inputRegisters_14__4, inputRegisters_14__3, inputRegisters_14__2, 
         inputRegisters_14__1, inputRegisters_14__0, inputRegisters_15__15, 
         inputRegisters_15__14, inputRegisters_15__13, inputRegisters_15__12, 
         inputRegisters_15__11, inputRegisters_15__10, inputRegisters_15__9, 
         inputRegisters_15__8, inputRegisters_15__7, inputRegisters_15__6, 
         inputRegisters_15__5, inputRegisters_15__4, inputRegisters_15__3, 
         inputRegisters_15__2, inputRegisters_15__1, inputRegisters_15__0, 
         inputRegisters_16__15, inputRegisters_16__14, inputRegisters_16__13, 
         inputRegisters_16__12, inputRegisters_16__11, inputRegisters_16__10, 
         inputRegisters_16__9, inputRegisters_16__8, inputRegisters_16__7, 
         inputRegisters_16__6, inputRegisters_16__5, inputRegisters_16__4, 
         inputRegisters_16__3, inputRegisters_16__2, inputRegisters_16__1, 
         inputRegisters_16__0, inputRegisters_17__15, inputRegisters_17__14, 
         inputRegisters_17__13, inputRegisters_17__12, inputRegisters_17__11, 
         inputRegisters_17__10, inputRegisters_17__9, inputRegisters_17__8, 
         inputRegisters_17__7, inputRegisters_17__6, inputRegisters_17__5, 
         inputRegisters_17__4, inputRegisters_17__3, inputRegisters_17__2, 
         inputRegisters_17__1, inputRegisters_17__0, inputRegisters_18__15, 
         inputRegisters_18__14, inputRegisters_18__13, inputRegisters_18__12, 
         inputRegisters_18__11, inputRegisters_18__10, inputRegisters_18__9, 
         inputRegisters_18__8, inputRegisters_18__7, inputRegisters_18__6, 
         inputRegisters_18__5, inputRegisters_18__4, inputRegisters_18__3, 
         inputRegisters_18__2, inputRegisters_18__1, inputRegisters_18__0, 
         inputRegisters_19__15, inputRegisters_19__14, inputRegisters_19__13, 
         inputRegisters_19__12, inputRegisters_19__11, inputRegisters_19__10, 
         inputRegisters_19__9, inputRegisters_19__8, inputRegisters_19__7, 
         inputRegisters_19__6, inputRegisters_19__5, inputRegisters_19__4, 
         inputRegisters_19__3, inputRegisters_19__2, inputRegisters_19__1, 
         inputRegisters_19__0, inputRegisters_20__15, inputRegisters_20__14, 
         inputRegisters_20__13, inputRegisters_20__12, inputRegisters_20__11, 
         inputRegisters_20__10, inputRegisters_20__9, inputRegisters_20__8, 
         inputRegisters_20__7, inputRegisters_20__6, inputRegisters_20__5, 
         inputRegisters_20__4, inputRegisters_20__3, inputRegisters_20__2, 
         inputRegisters_20__1, inputRegisters_20__0, inputRegisters_21__15, 
         inputRegisters_21__14, inputRegisters_21__13, inputRegisters_21__12, 
         inputRegisters_21__11, inputRegisters_21__10, inputRegisters_21__9, 
         inputRegisters_21__8, inputRegisters_21__7, inputRegisters_21__6, 
         inputRegisters_21__5, inputRegisters_21__4, inputRegisters_21__3, 
         inputRegisters_21__2, inputRegisters_21__1, inputRegisters_21__0, 
         inputRegisters_22__15, inputRegisters_22__14, inputRegisters_22__13, 
         inputRegisters_22__12, inputRegisters_22__11, inputRegisters_22__10, 
         inputRegisters_22__9, inputRegisters_22__8, inputRegisters_22__7, 
         inputRegisters_22__6, inputRegisters_22__5, inputRegisters_22__4, 
         inputRegisters_22__3, inputRegisters_22__2, inputRegisters_22__1, 
         inputRegisters_22__0, inputRegisters_23__15, inputRegisters_23__14, 
         inputRegisters_23__13, inputRegisters_23__12, inputRegisters_23__11, 
         inputRegisters_23__10, inputRegisters_23__9, inputRegisters_23__8, 
         inputRegisters_23__7, inputRegisters_23__6, inputRegisters_23__5, 
         inputRegisters_23__4, inputRegisters_23__3, inputRegisters_23__2, 
         inputRegisters_23__1, inputRegisters_23__0, inputRegisters_24__15, 
         inputRegisters_24__14, inputRegisters_24__13, inputRegisters_24__12, 
         inputRegisters_24__11, inputRegisters_24__10, inputRegisters_24__9, 
         inputRegisters_24__8, inputRegisters_24__7, inputRegisters_24__6, 
         inputRegisters_24__5, inputRegisters_24__4, inputRegisters_24__3, 
         inputRegisters_24__2, inputRegisters_24__1, inputRegisters_24__0, 
         inputRegisters_25__15, inputRegisters_25__14, inputRegisters_25__13, 
         inputRegisters_25__12, inputRegisters_25__11, inputRegisters_25__10, 
         inputRegisters_25__9, inputRegisters_25__8, inputRegisters_25__7, 
         inputRegisters_25__6, inputRegisters_25__5, inputRegisters_25__4, 
         inputRegisters_25__3, inputRegisters_25__2, inputRegisters_25__1, 
         inputRegisters_25__0, inputRegisters_26__15, inputRegisters_26__14, 
         inputRegisters_26__13, inputRegisters_26__12, inputRegisters_26__11, 
         inputRegisters_26__10, inputRegisters_26__9, inputRegisters_26__8, 
         inputRegisters_26__7, inputRegisters_26__6, inputRegisters_26__5, 
         inputRegisters_26__4, inputRegisters_26__3, inputRegisters_26__2, 
         inputRegisters_26__1, inputRegisters_26__0, inputRegisters_27__15, 
         inputRegisters_27__14, inputRegisters_27__13, inputRegisters_27__12, 
         inputRegisters_27__11, inputRegisters_27__10, inputRegisters_27__9, 
         inputRegisters_27__8, inputRegisters_27__7, inputRegisters_27__6, 
         inputRegisters_27__5, inputRegisters_27__4, inputRegisters_27__3, 
         inputRegisters_27__2, inputRegisters_27__1, inputRegisters_27__0, 
         inputRegisters_28__15, inputRegisters_28__14, inputRegisters_28__13, 
         inputRegisters_28__12, inputRegisters_28__11, inputRegisters_28__10, 
         inputRegisters_28__9, inputRegisters_28__8, inputRegisters_28__7, 
         inputRegisters_28__6, inputRegisters_28__5, inputRegisters_28__4, 
         inputRegisters_28__3, inputRegisters_28__2, inputRegisters_28__1, 
         inputRegisters_28__0, inputRegisters_29__15, inputRegisters_29__14, 
         inputRegisters_29__13, inputRegisters_29__12, inputRegisters_29__11, 
         inputRegisters_29__10, inputRegisters_29__9, inputRegisters_29__8, 
         inputRegisters_29__7, inputRegisters_29__6, inputRegisters_29__5, 
         inputRegisters_29__4, inputRegisters_29__3, inputRegisters_29__2, 
         inputRegisters_29__1, inputRegisters_29__0, inputRegisters_30__15, 
         inputRegisters_30__14, inputRegisters_30__13, inputRegisters_30__12, 
         inputRegisters_30__11, inputRegisters_30__10, inputRegisters_30__9, 
         inputRegisters_30__8, inputRegisters_30__7, inputRegisters_30__6, 
         inputRegisters_30__5, inputRegisters_30__4, inputRegisters_30__3, 
         inputRegisters_30__2, inputRegisters_30__1, inputRegisters_30__0, 
         inputRegisters_31__15, inputRegisters_31__14, inputRegisters_31__13, 
         inputRegisters_31__12, inputRegisters_31__11, inputRegisters_31__10, 
         inputRegisters_31__9, inputRegisters_31__8, inputRegisters_31__7, 
         inputRegisters_31__6, inputRegisters_31__5, inputRegisters_31__4, 
         inputRegisters_31__3, inputRegisters_31__2, inputRegisters_31__1, 
         inputRegisters_31__0, inputRegisters_32__15, inputRegisters_32__14, 
         inputRegisters_32__13, inputRegisters_32__12, inputRegisters_32__11, 
         inputRegisters_32__10, inputRegisters_32__9, inputRegisters_32__8, 
         inputRegisters_32__7, inputRegisters_32__6, inputRegisters_32__5, 
         inputRegisters_32__4, inputRegisters_32__3, inputRegisters_32__2, 
         inputRegisters_32__1, inputRegisters_32__0, inputRegisters_33__15, 
         inputRegisters_33__14, inputRegisters_33__13, inputRegisters_33__12, 
         inputRegisters_33__11, inputRegisters_33__10, inputRegisters_33__9, 
         inputRegisters_33__8, inputRegisters_33__7, inputRegisters_33__6, 
         inputRegisters_33__5, inputRegisters_33__4, inputRegisters_33__3, 
         inputRegisters_33__2, inputRegisters_33__1, inputRegisters_33__0, 
         inputRegisters_34__15, inputRegisters_34__14, inputRegisters_34__13, 
         inputRegisters_34__12, inputRegisters_34__11, inputRegisters_34__10, 
         inputRegisters_34__9, inputRegisters_34__8, inputRegisters_34__7, 
         inputRegisters_34__6, inputRegisters_34__5, inputRegisters_34__4, 
         inputRegisters_34__3, inputRegisters_34__2, inputRegisters_34__1, 
         inputRegisters_34__0, inputRegisters_35__15, inputRegisters_35__14, 
         inputRegisters_35__13, inputRegisters_35__12, inputRegisters_35__11, 
         inputRegisters_35__10, inputRegisters_35__9, inputRegisters_35__8, 
         inputRegisters_35__7, inputRegisters_35__6, inputRegisters_35__5, 
         inputRegisters_35__4, inputRegisters_35__3, inputRegisters_35__2, 
         inputRegisters_35__1, inputRegisters_35__0, inputRegisters_36__15, 
         inputRegisters_36__14, inputRegisters_36__13, inputRegisters_36__12, 
         inputRegisters_36__11, inputRegisters_36__10, inputRegisters_36__9, 
         inputRegisters_36__8, inputRegisters_36__7, inputRegisters_36__6, 
         inputRegisters_36__5, inputRegisters_36__4, inputRegisters_36__3, 
         inputRegisters_36__2, inputRegisters_36__1, inputRegisters_36__0, 
         inputRegisters_37__15, inputRegisters_37__14, inputRegisters_37__13, 
         inputRegisters_37__12, inputRegisters_37__11, inputRegisters_37__10, 
         inputRegisters_37__9, inputRegisters_37__8, inputRegisters_37__7, 
         inputRegisters_37__6, inputRegisters_37__5, inputRegisters_37__4, 
         inputRegisters_37__3, inputRegisters_37__2, inputRegisters_37__1, 
         inputRegisters_37__0, inputRegisters_38__15, inputRegisters_38__14, 
         inputRegisters_38__13, inputRegisters_38__12, inputRegisters_38__11, 
         inputRegisters_38__10, inputRegisters_38__9, inputRegisters_38__8, 
         inputRegisters_38__7, inputRegisters_38__6, inputRegisters_38__5, 
         inputRegisters_38__4, inputRegisters_38__3, inputRegisters_38__2, 
         inputRegisters_38__1, inputRegisters_38__0, inputRegisters_39__15, 
         inputRegisters_39__14, inputRegisters_39__13, inputRegisters_39__12, 
         inputRegisters_39__11, inputRegisters_39__10, inputRegisters_39__9, 
         inputRegisters_39__8, inputRegisters_39__7, inputRegisters_39__6, 
         inputRegisters_39__5, inputRegisters_39__4, inputRegisters_39__3, 
         inputRegisters_39__2, inputRegisters_39__1, inputRegisters_39__0, 
         inputRegisters_40__15, inputRegisters_40__14, inputRegisters_40__13, 
         inputRegisters_40__12, inputRegisters_40__11, inputRegisters_40__10, 
         inputRegisters_40__9, inputRegisters_40__8, inputRegisters_40__7, 
         inputRegisters_40__6, inputRegisters_40__5, inputRegisters_40__4, 
         inputRegisters_40__3, inputRegisters_40__2, inputRegisters_40__1, 
         inputRegisters_40__0, inputRegisters_41__15, inputRegisters_41__14, 
         inputRegisters_41__13, inputRegisters_41__12, inputRegisters_41__11, 
         inputRegisters_41__10, inputRegisters_41__9, inputRegisters_41__8, 
         inputRegisters_41__7, inputRegisters_41__6, inputRegisters_41__5, 
         inputRegisters_41__4, inputRegisters_41__3, inputRegisters_41__2, 
         inputRegisters_41__1, inputRegisters_41__0, inputRegisters_42__15, 
         inputRegisters_42__14, inputRegisters_42__13, inputRegisters_42__12, 
         inputRegisters_42__11, inputRegisters_42__10, inputRegisters_42__9, 
         inputRegisters_42__8, inputRegisters_42__7, inputRegisters_42__6, 
         inputRegisters_42__5, inputRegisters_42__4, inputRegisters_42__3, 
         inputRegisters_42__2, inputRegisters_42__1, inputRegisters_42__0, 
         inputRegisters_43__15, inputRegisters_43__14, inputRegisters_43__13, 
         inputRegisters_43__12, inputRegisters_43__11, inputRegisters_43__10, 
         inputRegisters_43__9, inputRegisters_43__8, inputRegisters_43__7, 
         inputRegisters_43__6, inputRegisters_43__5, inputRegisters_43__4, 
         inputRegisters_43__3, inputRegisters_43__2, inputRegisters_43__1, 
         inputRegisters_43__0, inputRegisters_44__15, inputRegisters_44__14, 
         inputRegisters_44__13, inputRegisters_44__12, inputRegisters_44__11, 
         inputRegisters_44__10, inputRegisters_44__9, inputRegisters_44__8, 
         inputRegisters_44__7, inputRegisters_44__6, inputRegisters_44__5, 
         inputRegisters_44__4, inputRegisters_44__3, inputRegisters_44__2, 
         inputRegisters_44__1, inputRegisters_44__0, inputRegisters_45__15, 
         inputRegisters_45__14, inputRegisters_45__13, inputRegisters_45__12, 
         inputRegisters_45__11, inputRegisters_45__10, inputRegisters_45__9, 
         inputRegisters_45__8, inputRegisters_45__7, inputRegisters_45__6, 
         inputRegisters_45__5, inputRegisters_45__4, inputRegisters_45__3, 
         inputRegisters_45__2, inputRegisters_45__1, inputRegisters_45__0, 
         inputRegisters_46__15, inputRegisters_46__14, inputRegisters_46__13, 
         inputRegisters_46__12, inputRegisters_46__11, inputRegisters_46__10, 
         inputRegisters_46__9, inputRegisters_46__8, inputRegisters_46__7, 
         inputRegisters_46__6, inputRegisters_46__5, inputRegisters_46__4, 
         inputRegisters_46__3, inputRegisters_46__2, inputRegisters_46__1, 
         inputRegisters_46__0, inputRegisters_47__15, inputRegisters_47__14, 
         inputRegisters_47__13, inputRegisters_47__12, inputRegisters_47__11, 
         inputRegisters_47__10, inputRegisters_47__9, inputRegisters_47__8, 
         inputRegisters_47__7, inputRegisters_47__6, inputRegisters_47__5, 
         inputRegisters_47__4, inputRegisters_47__3, inputRegisters_47__2, 
         inputRegisters_47__1, inputRegisters_47__0, inputRegisters_48__15, 
         inputRegisters_48__14, inputRegisters_48__13, inputRegisters_48__12, 
         inputRegisters_48__11, inputRegisters_48__10, inputRegisters_48__9, 
         inputRegisters_48__8, inputRegisters_48__7, inputRegisters_48__6, 
         inputRegisters_48__5, inputRegisters_48__4, inputRegisters_48__3, 
         inputRegisters_48__2, inputRegisters_48__1, inputRegisters_48__0, 
         inputRegisters_49__15, inputRegisters_49__14, inputRegisters_49__13, 
         inputRegisters_49__12, inputRegisters_49__11, inputRegisters_49__10, 
         inputRegisters_49__9, inputRegisters_49__8, inputRegisters_49__7, 
         inputRegisters_49__6, inputRegisters_49__5, inputRegisters_49__4, 
         inputRegisters_49__3, inputRegisters_49__2, inputRegisters_49__1, 
         inputRegisters_49__0, inputRegisters_50__15, inputRegisters_50__14, 
         inputRegisters_50__13, inputRegisters_50__12, inputRegisters_50__11, 
         inputRegisters_50__10, inputRegisters_50__9, inputRegisters_50__8, 
         inputRegisters_50__7, inputRegisters_50__6, inputRegisters_50__5, 
         inputRegisters_50__4, inputRegisters_50__3, inputRegisters_50__2, 
         inputRegisters_50__1, inputRegisters_50__0, inputRegisters_51__15, 
         inputRegisters_51__14, inputRegisters_51__13, inputRegisters_51__12, 
         inputRegisters_51__11, inputRegisters_51__10, inputRegisters_51__9, 
         inputRegisters_51__8, inputRegisters_51__7, inputRegisters_51__6, 
         inputRegisters_51__5, inputRegisters_51__4, inputRegisters_51__3, 
         inputRegisters_51__2, inputRegisters_51__1, inputRegisters_51__0, 
         inputRegisters_52__15, inputRegisters_52__14, inputRegisters_52__13, 
         inputRegisters_52__12, inputRegisters_52__11, inputRegisters_52__10, 
         inputRegisters_52__9, inputRegisters_52__8, inputRegisters_52__7, 
         inputRegisters_52__6, inputRegisters_52__5, inputRegisters_52__4, 
         inputRegisters_52__3, inputRegisters_52__2, inputRegisters_52__1, 
         inputRegisters_52__0, inputRegisters_53__15, inputRegisters_53__14, 
         inputRegisters_53__13, inputRegisters_53__12, inputRegisters_53__11, 
         inputRegisters_53__10, inputRegisters_53__9, inputRegisters_53__8, 
         inputRegisters_53__7, inputRegisters_53__6, inputRegisters_53__5, 
         inputRegisters_53__4, inputRegisters_53__3, inputRegisters_53__2, 
         inputRegisters_53__1, inputRegisters_53__0, inputRegisters_54__15, 
         inputRegisters_54__14, inputRegisters_54__13, inputRegisters_54__12, 
         inputRegisters_54__11, inputRegisters_54__10, inputRegisters_54__9, 
         inputRegisters_54__8, inputRegisters_54__7, inputRegisters_54__6, 
         inputRegisters_54__5, inputRegisters_54__4, inputRegisters_54__3, 
         inputRegisters_54__2, inputRegisters_54__1, inputRegisters_54__0, 
         inputRegisters_55__15, inputRegisters_55__14, inputRegisters_55__13, 
         inputRegisters_55__12, inputRegisters_55__11, inputRegisters_55__10, 
         inputRegisters_55__9, inputRegisters_55__8, inputRegisters_55__7, 
         inputRegisters_55__6, inputRegisters_55__5, inputRegisters_55__4, 
         inputRegisters_55__3, inputRegisters_55__2, inputRegisters_55__1, 
         inputRegisters_55__0, inputRegisters_56__15, inputRegisters_56__14, 
         inputRegisters_56__13, inputRegisters_56__12, inputRegisters_56__11, 
         inputRegisters_56__10, inputRegisters_56__9, inputRegisters_56__8, 
         inputRegisters_56__7, inputRegisters_56__6, inputRegisters_56__5, 
         inputRegisters_56__4, inputRegisters_56__3, inputRegisters_56__2, 
         inputRegisters_56__1, inputRegisters_56__0, inputRegisters_57__15, 
         inputRegisters_57__14, inputRegisters_57__13, inputRegisters_57__12, 
         inputRegisters_57__11, inputRegisters_57__10, inputRegisters_57__9, 
         inputRegisters_57__8, inputRegisters_57__7, inputRegisters_57__6, 
         inputRegisters_57__5, inputRegisters_57__4, inputRegisters_57__3, 
         inputRegisters_57__2, inputRegisters_57__1, inputRegisters_57__0, 
         inputRegisters_58__15, inputRegisters_58__14, inputRegisters_58__13, 
         inputRegisters_58__12, inputRegisters_58__11, inputRegisters_58__10, 
         inputRegisters_58__9, inputRegisters_58__8, inputRegisters_58__7, 
         inputRegisters_58__6, inputRegisters_58__5, inputRegisters_58__4, 
         inputRegisters_58__3, inputRegisters_58__2, inputRegisters_58__1, 
         inputRegisters_58__0, inputRegisters_59__15, inputRegisters_59__14, 
         inputRegisters_59__13, inputRegisters_59__12, inputRegisters_59__11, 
         inputRegisters_59__10, inputRegisters_59__9, inputRegisters_59__8, 
         inputRegisters_59__7, inputRegisters_59__6, inputRegisters_59__5, 
         inputRegisters_59__4, inputRegisters_59__3, inputRegisters_59__2, 
         inputRegisters_59__1, inputRegisters_59__0, inputRegisters_60__15, 
         inputRegisters_60__14, inputRegisters_60__13, inputRegisters_60__12, 
         inputRegisters_60__11, inputRegisters_60__10, inputRegisters_60__9, 
         inputRegisters_60__8, inputRegisters_60__7, inputRegisters_60__6, 
         inputRegisters_60__5, inputRegisters_60__4, inputRegisters_60__3, 
         inputRegisters_60__2, inputRegisters_60__1, inputRegisters_60__0, 
         inputRegisters_61__15, inputRegisters_61__14, inputRegisters_61__13, 
         inputRegisters_61__12, inputRegisters_61__11, inputRegisters_61__10, 
         inputRegisters_61__9, inputRegisters_61__8, inputRegisters_61__7, 
         inputRegisters_61__6, inputRegisters_61__5, inputRegisters_61__4, 
         inputRegisters_61__3, inputRegisters_61__2, inputRegisters_61__1, 
         inputRegisters_61__0, inputRegisters_62__15, inputRegisters_62__14, 
         inputRegisters_62__13, inputRegisters_62__12, inputRegisters_62__11, 
         inputRegisters_62__10, inputRegisters_62__9, inputRegisters_62__8, 
         inputRegisters_62__7, inputRegisters_62__6, inputRegisters_62__5, 
         inputRegisters_62__4, inputRegisters_62__3, inputRegisters_62__2, 
         inputRegisters_62__1, inputRegisters_62__0, inputRegisters_63__15, 
         inputRegisters_63__14, inputRegisters_63__13, inputRegisters_63__12, 
         inputRegisters_63__11, inputRegisters_63__10, inputRegisters_63__9, 
         inputRegisters_63__8, inputRegisters_63__7, inputRegisters_63__6, 
         inputRegisters_63__5, inputRegisters_63__4, inputRegisters_63__3, 
         inputRegisters_63__2, inputRegisters_63__1, inputRegisters_63__0, 
         inputRegisters_64__15, inputRegisters_64__14, inputRegisters_64__13, 
         inputRegisters_64__12, inputRegisters_64__11, inputRegisters_64__10, 
         inputRegisters_64__9, inputRegisters_64__8, inputRegisters_64__7, 
         inputRegisters_64__6, inputRegisters_64__5, inputRegisters_64__4, 
         inputRegisters_64__3, inputRegisters_64__2, inputRegisters_64__1, 
         inputRegisters_64__0, inputRegisters_65__15, inputRegisters_65__14, 
         inputRegisters_65__13, inputRegisters_65__12, inputRegisters_65__11, 
         inputRegisters_65__10, inputRegisters_65__9, inputRegisters_65__8, 
         inputRegisters_65__7, inputRegisters_65__6, inputRegisters_65__5, 
         inputRegisters_65__4, inputRegisters_65__3, inputRegisters_65__2, 
         inputRegisters_65__1, inputRegisters_65__0, inputRegisters_66__15, 
         inputRegisters_66__14, inputRegisters_66__13, inputRegisters_66__12, 
         inputRegisters_66__11, inputRegisters_66__10, inputRegisters_66__9, 
         inputRegisters_66__8, inputRegisters_66__7, inputRegisters_66__6, 
         inputRegisters_66__5, inputRegisters_66__4, inputRegisters_66__3, 
         inputRegisters_66__2, inputRegisters_66__1, inputRegisters_66__0, 
         inputRegisters_67__15, inputRegisters_67__14, inputRegisters_67__13, 
         inputRegisters_67__12, inputRegisters_67__11, inputRegisters_67__10, 
         inputRegisters_67__9, inputRegisters_67__8, inputRegisters_67__7, 
         inputRegisters_67__6, inputRegisters_67__5, inputRegisters_67__4, 
         inputRegisters_67__3, inputRegisters_67__2, inputRegisters_67__1, 
         inputRegisters_67__0, inputRegisters_68__15, inputRegisters_68__14, 
         inputRegisters_68__13, inputRegisters_68__12, inputRegisters_68__11, 
         inputRegisters_68__10, inputRegisters_68__9, inputRegisters_68__8, 
         inputRegisters_68__7, inputRegisters_68__6, inputRegisters_68__5, 
         inputRegisters_68__4, inputRegisters_68__3, inputRegisters_68__2, 
         inputRegisters_68__1, inputRegisters_68__0, inputRegisters_69__15, 
         inputRegisters_69__14, inputRegisters_69__13, inputRegisters_69__12, 
         inputRegisters_69__11, inputRegisters_69__10, inputRegisters_69__9, 
         inputRegisters_69__8, inputRegisters_69__7, inputRegisters_69__6, 
         inputRegisters_69__5, inputRegisters_69__4, inputRegisters_69__3, 
         inputRegisters_69__2, inputRegisters_69__1, inputRegisters_69__0, 
         inputRegisters_70__15, inputRegisters_70__14, inputRegisters_70__13, 
         inputRegisters_70__12, inputRegisters_70__11, inputRegisters_70__10, 
         inputRegisters_70__9, inputRegisters_70__8, inputRegisters_70__7, 
         inputRegisters_70__6, inputRegisters_70__5, inputRegisters_70__4, 
         inputRegisters_70__3, inputRegisters_70__2, inputRegisters_70__1, 
         inputRegisters_70__0, inputRegisters_71__15, inputRegisters_71__14, 
         inputRegisters_71__13, inputRegisters_71__12, inputRegisters_71__11, 
         inputRegisters_71__10, inputRegisters_71__9, inputRegisters_71__8, 
         inputRegisters_71__7, inputRegisters_71__6, inputRegisters_71__5, 
         inputRegisters_71__4, inputRegisters_71__3, inputRegisters_71__2, 
         inputRegisters_71__1, inputRegisters_71__0, inputRegisters_72__15, 
         inputRegisters_72__14, inputRegisters_72__13, inputRegisters_72__12, 
         inputRegisters_72__11, inputRegisters_72__10, inputRegisters_72__9, 
         inputRegisters_72__8, inputRegisters_72__7, inputRegisters_72__6, 
         inputRegisters_72__5, inputRegisters_72__4, inputRegisters_72__3, 
         inputRegisters_72__2, inputRegisters_72__1, inputRegisters_72__0, 
         inputRegisters_73__15, inputRegisters_73__14, inputRegisters_73__13, 
         inputRegisters_73__12, inputRegisters_73__11, inputRegisters_73__10, 
         inputRegisters_73__9, inputRegisters_73__8, inputRegisters_73__7, 
         inputRegisters_73__6, inputRegisters_73__5, inputRegisters_73__4, 
         inputRegisters_73__3, inputRegisters_73__2, inputRegisters_73__1, 
         inputRegisters_73__0, inputRegisters_74__15, inputRegisters_74__14, 
         inputRegisters_74__13, inputRegisters_74__12, inputRegisters_74__11, 
         inputRegisters_74__10, inputRegisters_74__9, inputRegisters_74__8, 
         inputRegisters_74__7, inputRegisters_74__6, inputRegisters_74__5, 
         inputRegisters_74__4, inputRegisters_74__3, inputRegisters_74__2, 
         inputRegisters_74__1, inputRegisters_74__0, inputRegisters_75__15, 
         inputRegisters_75__14, inputRegisters_75__13, inputRegisters_75__12, 
         inputRegisters_75__11, inputRegisters_75__10, inputRegisters_75__9, 
         inputRegisters_75__8, inputRegisters_75__7, inputRegisters_75__6, 
         inputRegisters_75__5, inputRegisters_75__4, inputRegisters_75__3, 
         inputRegisters_75__2, inputRegisters_75__1, inputRegisters_75__0, 
         inputRegisters_76__15, inputRegisters_76__14, inputRegisters_76__13, 
         inputRegisters_76__12, inputRegisters_76__11, inputRegisters_76__10, 
         inputRegisters_76__9, inputRegisters_76__8, inputRegisters_76__7, 
         inputRegisters_76__6, inputRegisters_76__5, inputRegisters_76__4, 
         inputRegisters_76__3, inputRegisters_76__2, inputRegisters_76__1, 
         inputRegisters_76__0, inputRegisters_77__15, inputRegisters_77__14, 
         inputRegisters_77__13, inputRegisters_77__12, inputRegisters_77__11, 
         inputRegisters_77__10, inputRegisters_77__9, inputRegisters_77__8, 
         inputRegisters_77__7, inputRegisters_77__6, inputRegisters_77__5, 
         inputRegisters_77__4, inputRegisters_77__3, inputRegisters_77__2, 
         inputRegisters_77__1, inputRegisters_77__0, inputRegisters_78__15, 
         inputRegisters_78__14, inputRegisters_78__13, inputRegisters_78__12, 
         inputRegisters_78__11, inputRegisters_78__10, inputRegisters_78__9, 
         inputRegisters_78__8, inputRegisters_78__7, inputRegisters_78__6, 
         inputRegisters_78__5, inputRegisters_78__4, inputRegisters_78__3, 
         inputRegisters_78__2, inputRegisters_78__1, inputRegisters_78__0, 
         inputRegisters_79__15, inputRegisters_79__14, inputRegisters_79__13, 
         inputRegisters_79__12, inputRegisters_79__11, inputRegisters_79__10, 
         inputRegisters_79__9, inputRegisters_79__8, inputRegisters_79__7, 
         inputRegisters_79__6, inputRegisters_79__5, inputRegisters_79__4, 
         inputRegisters_79__3, inputRegisters_79__2, inputRegisters_79__1, 
         inputRegisters_79__0, inputRegisters_80__15, inputRegisters_80__14, 
         inputRegisters_80__13, inputRegisters_80__12, inputRegisters_80__11, 
         inputRegisters_80__10, inputRegisters_80__9, inputRegisters_80__8, 
         inputRegisters_80__7, inputRegisters_80__6, inputRegisters_80__5, 
         inputRegisters_80__4, inputRegisters_80__3, inputRegisters_80__2, 
         inputRegisters_80__1, inputRegisters_80__0, inputRegisters_81__15, 
         inputRegisters_81__14, inputRegisters_81__13, inputRegisters_81__12, 
         inputRegisters_81__11, inputRegisters_81__10, inputRegisters_81__9, 
         inputRegisters_81__8, inputRegisters_81__7, inputRegisters_81__6, 
         inputRegisters_81__5, inputRegisters_81__4, inputRegisters_81__3, 
         inputRegisters_81__2, inputRegisters_81__1, inputRegisters_81__0, 
         inputRegisters_82__15, inputRegisters_82__14, inputRegisters_82__13, 
         inputRegisters_82__12, inputRegisters_82__11, inputRegisters_82__10, 
         inputRegisters_82__9, inputRegisters_82__8, inputRegisters_82__7, 
         inputRegisters_82__6, inputRegisters_82__5, inputRegisters_82__4, 
         inputRegisters_82__3, inputRegisters_82__2, inputRegisters_82__1, 
         inputRegisters_82__0, inputRegisters_83__15, inputRegisters_83__14, 
         inputRegisters_83__13, inputRegisters_83__12, inputRegisters_83__11, 
         inputRegisters_83__10, inputRegisters_83__9, inputRegisters_83__8, 
         inputRegisters_83__7, inputRegisters_83__6, inputRegisters_83__5, 
         inputRegisters_83__4, inputRegisters_83__3, inputRegisters_83__2, 
         inputRegisters_83__1, inputRegisters_83__0, inputRegisters_84__15, 
         inputRegisters_84__14, inputRegisters_84__13, inputRegisters_84__12, 
         inputRegisters_84__11, inputRegisters_84__10, inputRegisters_84__9, 
         inputRegisters_84__8, inputRegisters_84__7, inputRegisters_84__6, 
         inputRegisters_84__5, inputRegisters_84__4, inputRegisters_84__3, 
         inputRegisters_84__2, inputRegisters_84__1, inputRegisters_84__0, 
         inputRegisters_85__15, inputRegisters_85__14, inputRegisters_85__13, 
         inputRegisters_85__12, inputRegisters_85__11, inputRegisters_85__10, 
         inputRegisters_85__9, inputRegisters_85__8, inputRegisters_85__7, 
         inputRegisters_85__6, inputRegisters_85__5, inputRegisters_85__4, 
         inputRegisters_85__3, inputRegisters_85__2, inputRegisters_85__1, 
         inputRegisters_85__0, inputRegisters_86__15, inputRegisters_86__14, 
         inputRegisters_86__13, inputRegisters_86__12, inputRegisters_86__11, 
         inputRegisters_86__10, inputRegisters_86__9, inputRegisters_86__8, 
         inputRegisters_86__7, inputRegisters_86__6, inputRegisters_86__5, 
         inputRegisters_86__4, inputRegisters_86__3, inputRegisters_86__2, 
         inputRegisters_86__1, inputRegisters_86__0, inputRegisters_87__15, 
         inputRegisters_87__14, inputRegisters_87__13, inputRegisters_87__12, 
         inputRegisters_87__11, inputRegisters_87__10, inputRegisters_87__9, 
         inputRegisters_87__8, inputRegisters_87__7, inputRegisters_87__6, 
         inputRegisters_87__5, inputRegisters_87__4, inputRegisters_87__3, 
         inputRegisters_87__2, inputRegisters_87__1, inputRegisters_87__0, 
         inputRegisters_88__15, inputRegisters_88__14, inputRegisters_88__13, 
         inputRegisters_88__12, inputRegisters_88__11, inputRegisters_88__10, 
         inputRegisters_88__9, inputRegisters_88__8, inputRegisters_88__7, 
         inputRegisters_88__6, inputRegisters_88__5, inputRegisters_88__4, 
         inputRegisters_88__3, inputRegisters_88__2, inputRegisters_88__1, 
         inputRegisters_88__0, inputRegisters_89__15, inputRegisters_89__14, 
         inputRegisters_89__13, inputRegisters_89__12, inputRegisters_89__11, 
         inputRegisters_89__10, inputRegisters_89__9, inputRegisters_89__8, 
         inputRegisters_89__7, inputRegisters_89__6, inputRegisters_89__5, 
         inputRegisters_89__4, inputRegisters_89__3, inputRegisters_89__2, 
         inputRegisters_89__1, inputRegisters_89__0, inputRegisters_90__15, 
         inputRegisters_90__14, inputRegisters_90__13, inputRegisters_90__12, 
         inputRegisters_90__11, inputRegisters_90__10, inputRegisters_90__9, 
         inputRegisters_90__8, inputRegisters_90__7, inputRegisters_90__6, 
         inputRegisters_90__5, inputRegisters_90__4, inputRegisters_90__3, 
         inputRegisters_90__2, inputRegisters_90__1, inputRegisters_90__0, 
         inputRegisters_91__15, inputRegisters_91__14, inputRegisters_91__13, 
         inputRegisters_91__12, inputRegisters_91__11, inputRegisters_91__10, 
         inputRegisters_91__9, inputRegisters_91__8, inputRegisters_91__7, 
         inputRegisters_91__6, inputRegisters_91__5, inputRegisters_91__4, 
         inputRegisters_91__3, inputRegisters_91__2, inputRegisters_91__1, 
         inputRegisters_91__0, inputRegisters_92__15, inputRegisters_92__14, 
         inputRegisters_92__13, inputRegisters_92__12, inputRegisters_92__11, 
         inputRegisters_92__10, inputRegisters_92__9, inputRegisters_92__8, 
         inputRegisters_92__7, inputRegisters_92__6, inputRegisters_92__5, 
         inputRegisters_92__4, inputRegisters_92__3, inputRegisters_92__2, 
         inputRegisters_92__1, inputRegisters_92__0, inputRegisters_93__15, 
         inputRegisters_93__14, inputRegisters_93__13, inputRegisters_93__12, 
         inputRegisters_93__11, inputRegisters_93__10, inputRegisters_93__9, 
         inputRegisters_93__8, inputRegisters_93__7, inputRegisters_93__6, 
         inputRegisters_93__5, inputRegisters_93__4, inputRegisters_93__3, 
         inputRegisters_93__2, inputRegisters_93__1, inputRegisters_93__0, 
         inputRegisters_94__15, inputRegisters_94__14, inputRegisters_94__13, 
         inputRegisters_94__12, inputRegisters_94__11, inputRegisters_94__10, 
         inputRegisters_94__9, inputRegisters_94__8, inputRegisters_94__7, 
         inputRegisters_94__6, inputRegisters_94__5, inputRegisters_94__4, 
         inputRegisters_94__3, inputRegisters_94__2, inputRegisters_94__1, 
         inputRegisters_94__0, inputRegisters_95__15, inputRegisters_95__14, 
         inputRegisters_95__13, inputRegisters_95__12, inputRegisters_95__11, 
         inputRegisters_95__10, inputRegisters_95__9, inputRegisters_95__8, 
         inputRegisters_95__7, inputRegisters_95__6, inputRegisters_95__5, 
         inputRegisters_95__4, inputRegisters_95__3, inputRegisters_95__2, 
         inputRegisters_95__1, inputRegisters_95__0, inputRegisters_96__15, 
         inputRegisters_96__14, inputRegisters_96__13, inputRegisters_96__12, 
         inputRegisters_96__11, inputRegisters_96__10, inputRegisters_96__9, 
         inputRegisters_96__8, inputRegisters_96__7, inputRegisters_96__6, 
         inputRegisters_96__5, inputRegisters_96__4, inputRegisters_96__3, 
         inputRegisters_96__2, inputRegisters_96__1, inputRegisters_96__0, 
         inputRegisters_97__15, inputRegisters_97__14, inputRegisters_97__13, 
         inputRegisters_97__12, inputRegisters_97__11, inputRegisters_97__10, 
         inputRegisters_97__9, inputRegisters_97__8, inputRegisters_97__7, 
         inputRegisters_97__6, inputRegisters_97__5, inputRegisters_97__4, 
         inputRegisters_97__3, inputRegisters_97__2, inputRegisters_97__1, 
         inputRegisters_97__0, inputRegisters_98__15, inputRegisters_98__14, 
         inputRegisters_98__13, inputRegisters_98__12, inputRegisters_98__11, 
         inputRegisters_98__10, inputRegisters_98__9, inputRegisters_98__8, 
         inputRegisters_98__7, inputRegisters_98__6, inputRegisters_98__5, 
         inputRegisters_98__4, inputRegisters_98__3, inputRegisters_98__2, 
         inputRegisters_98__1, inputRegisters_98__0, inputRegisters_99__15, 
         inputRegisters_99__14, inputRegisters_99__13, inputRegisters_99__12, 
         inputRegisters_99__11, inputRegisters_99__10, inputRegisters_99__9, 
         inputRegisters_99__8, inputRegisters_99__7, inputRegisters_99__6, 
         inputRegisters_99__5, inputRegisters_99__4, inputRegisters_99__3, 
         inputRegisters_99__2, inputRegisters_99__1, inputRegisters_99__0, 
         inputRegisters_100__15, inputRegisters_100__14, inputRegisters_100__13, 
         inputRegisters_100__12, inputRegisters_100__11, inputRegisters_100__10, 
         inputRegisters_100__9, inputRegisters_100__8, inputRegisters_100__7, 
         inputRegisters_100__6, inputRegisters_100__5, inputRegisters_100__4, 
         inputRegisters_100__3, inputRegisters_100__2, inputRegisters_100__1, 
         inputRegisters_100__0, inputRegisters_101__15, inputRegisters_101__14, 
         inputRegisters_101__13, inputRegisters_101__12, inputRegisters_101__11, 
         inputRegisters_101__10, inputRegisters_101__9, inputRegisters_101__8, 
         inputRegisters_101__7, inputRegisters_101__6, inputRegisters_101__5, 
         inputRegisters_101__4, inputRegisters_101__3, inputRegisters_101__2, 
         inputRegisters_101__1, inputRegisters_101__0, inputRegisters_102__15, 
         inputRegisters_102__14, inputRegisters_102__13, inputRegisters_102__12, 
         inputRegisters_102__11, inputRegisters_102__10, inputRegisters_102__9, 
         inputRegisters_102__8, inputRegisters_102__7, inputRegisters_102__6, 
         inputRegisters_102__5, inputRegisters_102__4, inputRegisters_102__3, 
         inputRegisters_102__2, inputRegisters_102__1, inputRegisters_102__0, 
         inputRegisters_103__15, inputRegisters_103__14, inputRegisters_103__13, 
         inputRegisters_103__12, inputRegisters_103__11, inputRegisters_103__10, 
         inputRegisters_103__9, inputRegisters_103__8, inputRegisters_103__7, 
         inputRegisters_103__6, inputRegisters_103__5, inputRegisters_103__4, 
         inputRegisters_103__3, inputRegisters_103__2, inputRegisters_103__1, 
         inputRegisters_103__0, inputRegisters_104__15, inputRegisters_104__14, 
         inputRegisters_104__13, inputRegisters_104__12, inputRegisters_104__11, 
         inputRegisters_104__10, inputRegisters_104__9, inputRegisters_104__8, 
         inputRegisters_104__7, inputRegisters_104__6, inputRegisters_104__5, 
         inputRegisters_104__4, inputRegisters_104__3, inputRegisters_104__2, 
         inputRegisters_104__1, inputRegisters_104__0, inputRegisters_105__15, 
         inputRegisters_105__14, inputRegisters_105__13, inputRegisters_105__12, 
         inputRegisters_105__11, inputRegisters_105__10, inputRegisters_105__9, 
         inputRegisters_105__8, inputRegisters_105__7, inputRegisters_105__6, 
         inputRegisters_105__5, inputRegisters_105__4, inputRegisters_105__3, 
         inputRegisters_105__2, inputRegisters_105__1, inputRegisters_105__0, 
         inputRegisters_106__15, inputRegisters_106__14, inputRegisters_106__13, 
         inputRegisters_106__12, inputRegisters_106__11, inputRegisters_106__10, 
         inputRegisters_106__9, inputRegisters_106__8, inputRegisters_106__7, 
         inputRegisters_106__6, inputRegisters_106__5, inputRegisters_106__4, 
         inputRegisters_106__3, inputRegisters_106__2, inputRegisters_106__1, 
         inputRegisters_106__0, inputRegisters_107__15, inputRegisters_107__14, 
         inputRegisters_107__13, inputRegisters_107__12, inputRegisters_107__11, 
         inputRegisters_107__10, inputRegisters_107__9, inputRegisters_107__8, 
         inputRegisters_107__7, inputRegisters_107__6, inputRegisters_107__5, 
         inputRegisters_107__4, inputRegisters_107__3, inputRegisters_107__2, 
         inputRegisters_107__1, inputRegisters_107__0, inputRegisters_108__15, 
         inputRegisters_108__14, inputRegisters_108__13, inputRegisters_108__12, 
         inputRegisters_108__11, inputRegisters_108__10, inputRegisters_108__9, 
         inputRegisters_108__8, inputRegisters_108__7, inputRegisters_108__6, 
         inputRegisters_108__5, inputRegisters_108__4, inputRegisters_108__3, 
         inputRegisters_108__2, inputRegisters_108__1, inputRegisters_108__0, 
         inputRegisters_109__15, inputRegisters_109__14, inputRegisters_109__13, 
         inputRegisters_109__12, inputRegisters_109__11, inputRegisters_109__10, 
         inputRegisters_109__9, inputRegisters_109__8, inputRegisters_109__7, 
         inputRegisters_109__6, inputRegisters_109__5, inputRegisters_109__4, 
         inputRegisters_109__3, inputRegisters_109__2, inputRegisters_109__1, 
         inputRegisters_109__0, inputRegisters_110__15, inputRegisters_110__14, 
         inputRegisters_110__13, inputRegisters_110__12, inputRegisters_110__11, 
         inputRegisters_110__10, inputRegisters_110__9, inputRegisters_110__8, 
         inputRegisters_110__7, inputRegisters_110__6, inputRegisters_110__5, 
         inputRegisters_110__4, inputRegisters_110__3, inputRegisters_110__2, 
         inputRegisters_110__1, inputRegisters_110__0, inputRegisters_111__15, 
         inputRegisters_111__14, inputRegisters_111__13, inputRegisters_111__12, 
         inputRegisters_111__11, inputRegisters_111__10, inputRegisters_111__9, 
         inputRegisters_111__8, inputRegisters_111__7, inputRegisters_111__6, 
         inputRegisters_111__5, inputRegisters_111__4, inputRegisters_111__3, 
         inputRegisters_111__2, inputRegisters_111__1, inputRegisters_111__0, 
         inputRegisters_112__15, inputRegisters_112__14, inputRegisters_112__13, 
         inputRegisters_112__12, inputRegisters_112__11, inputRegisters_112__10, 
         inputRegisters_112__9, inputRegisters_112__8, inputRegisters_112__7, 
         inputRegisters_112__6, inputRegisters_112__5, inputRegisters_112__4, 
         inputRegisters_112__3, inputRegisters_112__2, inputRegisters_112__1, 
         inputRegisters_112__0, inputRegisters_113__15, inputRegisters_113__14, 
         inputRegisters_113__13, inputRegisters_113__12, inputRegisters_113__11, 
         inputRegisters_113__10, inputRegisters_113__9, inputRegisters_113__8, 
         inputRegisters_113__7, inputRegisters_113__6, inputRegisters_113__5, 
         inputRegisters_113__4, inputRegisters_113__3, inputRegisters_113__2, 
         inputRegisters_113__1, inputRegisters_113__0, inputRegisters_114__15, 
         inputRegisters_114__14, inputRegisters_114__13, inputRegisters_114__12, 
         inputRegisters_114__11, inputRegisters_114__10, inputRegisters_114__9, 
         inputRegisters_114__8, inputRegisters_114__7, inputRegisters_114__6, 
         inputRegisters_114__5, inputRegisters_114__4, inputRegisters_114__3, 
         inputRegisters_114__2, inputRegisters_114__1, inputRegisters_114__0, 
         inputRegisters_115__15, inputRegisters_115__14, inputRegisters_115__13, 
         inputRegisters_115__12, inputRegisters_115__11, inputRegisters_115__10, 
         inputRegisters_115__9, inputRegisters_115__8, inputRegisters_115__7, 
         inputRegisters_115__6, inputRegisters_115__5, inputRegisters_115__4, 
         inputRegisters_115__3, inputRegisters_115__2, inputRegisters_115__1, 
         inputRegisters_115__0, inputRegisters_116__15, inputRegisters_116__14, 
         inputRegisters_116__13, inputRegisters_116__12, inputRegisters_116__11, 
         inputRegisters_116__10, inputRegisters_116__9, inputRegisters_116__8, 
         inputRegisters_116__7, inputRegisters_116__6, inputRegisters_116__5, 
         inputRegisters_116__4, inputRegisters_116__3, inputRegisters_116__2, 
         inputRegisters_116__1, inputRegisters_116__0, inputRegisters_117__15, 
         inputRegisters_117__14, inputRegisters_117__13, inputRegisters_117__12, 
         inputRegisters_117__11, inputRegisters_117__10, inputRegisters_117__9, 
         inputRegisters_117__8, inputRegisters_117__7, inputRegisters_117__6, 
         inputRegisters_117__5, inputRegisters_117__4, inputRegisters_117__3, 
         inputRegisters_117__2, inputRegisters_117__1, inputRegisters_117__0, 
         inputRegisters_118__15, inputRegisters_118__14, inputRegisters_118__13, 
         inputRegisters_118__12, inputRegisters_118__11, inputRegisters_118__10, 
         inputRegisters_118__9, inputRegisters_118__8, inputRegisters_118__7, 
         inputRegisters_118__6, inputRegisters_118__5, inputRegisters_118__4, 
         inputRegisters_118__3, inputRegisters_118__2, inputRegisters_118__1, 
         inputRegisters_118__0, inputRegisters_119__15, inputRegisters_119__14, 
         inputRegisters_119__13, inputRegisters_119__12, inputRegisters_119__11, 
         inputRegisters_119__10, inputRegisters_119__9, inputRegisters_119__8, 
         inputRegisters_119__7, inputRegisters_119__6, inputRegisters_119__5, 
         inputRegisters_119__4, inputRegisters_119__3, inputRegisters_119__2, 
         inputRegisters_119__1, inputRegisters_119__0, inputRegisters_120__15, 
         inputRegisters_120__14, inputRegisters_120__13, inputRegisters_120__12, 
         inputRegisters_120__11, inputRegisters_120__10, inputRegisters_120__9, 
         inputRegisters_120__8, inputRegisters_120__7, inputRegisters_120__6, 
         inputRegisters_120__5, inputRegisters_120__4, inputRegisters_120__3, 
         inputRegisters_120__2, inputRegisters_120__1, inputRegisters_120__0, 
         inputRegisters_121__15, inputRegisters_121__14, inputRegisters_121__13, 
         inputRegisters_121__12, inputRegisters_121__11, inputRegisters_121__10, 
         inputRegisters_121__9, inputRegisters_121__8, inputRegisters_121__7, 
         inputRegisters_121__6, inputRegisters_121__5, inputRegisters_121__4, 
         inputRegisters_121__3, inputRegisters_121__2, inputRegisters_121__1, 
         inputRegisters_121__0, inputRegisters_122__15, inputRegisters_122__14, 
         inputRegisters_122__13, inputRegisters_122__12, inputRegisters_122__11, 
         inputRegisters_122__10, inputRegisters_122__9, inputRegisters_122__8, 
         inputRegisters_122__7, inputRegisters_122__6, inputRegisters_122__5, 
         inputRegisters_122__4, inputRegisters_122__3, inputRegisters_122__2, 
         inputRegisters_122__1, inputRegisters_122__0, inputRegisters_123__15, 
         inputRegisters_123__14, inputRegisters_123__13, inputRegisters_123__12, 
         inputRegisters_123__11, inputRegisters_123__10, inputRegisters_123__9, 
         inputRegisters_123__8, inputRegisters_123__7, inputRegisters_123__6, 
         inputRegisters_123__5, inputRegisters_123__4, inputRegisters_123__3, 
         inputRegisters_123__2, inputRegisters_123__1, inputRegisters_123__0, 
         inputRegisters_124__15, inputRegisters_124__14, inputRegisters_124__13, 
         inputRegisters_124__12, inputRegisters_124__11, inputRegisters_124__10, 
         inputRegisters_124__9, inputRegisters_124__8, inputRegisters_124__7, 
         inputRegisters_124__6, inputRegisters_124__5, inputRegisters_124__4, 
         inputRegisters_124__3, inputRegisters_124__2, inputRegisters_124__1, 
         inputRegisters_124__0, inputRegisters_125__15, inputRegisters_125__14, 
         inputRegisters_125__13, inputRegisters_125__12, inputRegisters_125__11, 
         inputRegisters_125__10, inputRegisters_125__9, inputRegisters_125__8, 
         inputRegisters_125__7, inputRegisters_125__6, inputRegisters_125__5, 
         inputRegisters_125__4, inputRegisters_125__3, inputRegisters_125__2, 
         inputRegisters_125__1, inputRegisters_125__0, inputRegisters_126__15, 
         inputRegisters_126__14, inputRegisters_126__13, inputRegisters_126__12, 
         inputRegisters_126__11, inputRegisters_126__10, inputRegisters_126__9, 
         inputRegisters_126__8, inputRegisters_126__7, inputRegisters_126__6, 
         inputRegisters_126__5, inputRegisters_126__4, inputRegisters_126__3, 
         inputRegisters_126__2, inputRegisters_126__1, inputRegisters_126__0, 
         inputRegisters_127__15, inputRegisters_127__14, inputRegisters_127__13, 
         inputRegisters_127__12, inputRegisters_127__11, inputRegisters_127__10, 
         inputRegisters_127__9, inputRegisters_127__8, inputRegisters_127__7, 
         inputRegisters_127__6, inputRegisters_127__5, inputRegisters_127__4, 
         inputRegisters_127__3, inputRegisters_127__2, inputRegisters_127__1, 
         inputRegisters_127__0, inputRegisters_128__15, inputRegisters_128__14, 
         inputRegisters_128__13, inputRegisters_128__12, inputRegisters_128__11, 
         inputRegisters_128__10, inputRegisters_128__9, inputRegisters_128__8, 
         inputRegisters_128__7, inputRegisters_128__6, inputRegisters_128__5, 
         inputRegisters_128__4, inputRegisters_128__3, inputRegisters_128__2, 
         inputRegisters_128__1, inputRegisters_128__0, inputRegisters_129__15, 
         inputRegisters_129__14, inputRegisters_129__13, inputRegisters_129__12, 
         inputRegisters_129__11, inputRegisters_129__10, inputRegisters_129__9, 
         inputRegisters_129__8, inputRegisters_129__7, inputRegisters_129__6, 
         inputRegisters_129__5, inputRegisters_129__4, inputRegisters_129__3, 
         inputRegisters_129__2, inputRegisters_129__1, inputRegisters_129__0, 
         inputRegisters_130__15, inputRegisters_130__14, inputRegisters_130__13, 
         inputRegisters_130__12, inputRegisters_130__11, inputRegisters_130__10, 
         inputRegisters_130__9, inputRegisters_130__8, inputRegisters_130__7, 
         inputRegisters_130__6, inputRegisters_130__5, inputRegisters_130__4, 
         inputRegisters_130__3, inputRegisters_130__2, inputRegisters_130__1, 
         inputRegisters_130__0, inputRegisters_131__15, inputRegisters_131__14, 
         inputRegisters_131__13, inputRegisters_131__12, inputRegisters_131__11, 
         inputRegisters_131__10, inputRegisters_131__9, inputRegisters_131__8, 
         inputRegisters_131__7, inputRegisters_131__6, inputRegisters_131__5, 
         inputRegisters_131__4, inputRegisters_131__3, inputRegisters_131__2, 
         inputRegisters_131__1, inputRegisters_131__0, inputRegisters_132__15, 
         inputRegisters_132__14, inputRegisters_132__13, inputRegisters_132__12, 
         inputRegisters_132__11, inputRegisters_132__10, inputRegisters_132__9, 
         inputRegisters_132__8, inputRegisters_132__7, inputRegisters_132__6, 
         inputRegisters_132__5, inputRegisters_132__4, inputRegisters_132__3, 
         inputRegisters_132__2, inputRegisters_132__1, inputRegisters_132__0, 
         inputRegisters_133__15, inputRegisters_133__14, inputRegisters_133__13, 
         inputRegisters_133__12, inputRegisters_133__11, inputRegisters_133__10, 
         inputRegisters_133__9, inputRegisters_133__8, inputRegisters_133__7, 
         inputRegisters_133__6, inputRegisters_133__5, inputRegisters_133__4, 
         inputRegisters_133__3, inputRegisters_133__2, inputRegisters_133__1, 
         inputRegisters_133__0, inputRegisters_134__15, inputRegisters_134__14, 
         inputRegisters_134__13, inputRegisters_134__12, inputRegisters_134__11, 
         inputRegisters_134__10, inputRegisters_134__9, inputRegisters_134__8, 
         inputRegisters_134__7, inputRegisters_134__6, inputRegisters_134__5, 
         inputRegisters_134__4, inputRegisters_134__3, inputRegisters_134__2, 
         inputRegisters_134__1, inputRegisters_134__0, inputRegisters_135__15, 
         inputRegisters_135__14, inputRegisters_135__13, inputRegisters_135__12, 
         inputRegisters_135__11, inputRegisters_135__10, inputRegisters_135__9, 
         inputRegisters_135__8, inputRegisters_135__7, inputRegisters_135__6, 
         inputRegisters_135__5, inputRegisters_135__4, inputRegisters_135__3, 
         inputRegisters_135__2, inputRegisters_135__1, inputRegisters_135__0, 
         inputRegisters_136__15, inputRegisters_136__14, inputRegisters_136__13, 
         inputRegisters_136__12, inputRegisters_136__11, inputRegisters_136__10, 
         inputRegisters_136__9, inputRegisters_136__8, inputRegisters_136__7, 
         inputRegisters_136__6, inputRegisters_136__5, inputRegisters_136__4, 
         inputRegisters_136__3, inputRegisters_136__2, inputRegisters_136__1, 
         inputRegisters_136__0, inputRegisters_137__15, inputRegisters_137__14, 
         inputRegisters_137__13, inputRegisters_137__12, inputRegisters_137__11, 
         inputRegisters_137__10, inputRegisters_137__9, inputRegisters_137__8, 
         inputRegisters_137__7, inputRegisters_137__6, inputRegisters_137__5, 
         inputRegisters_137__4, inputRegisters_137__3, inputRegisters_137__2, 
         inputRegisters_137__1, inputRegisters_137__0, inputRegisters_138__15, 
         inputRegisters_138__14, inputRegisters_138__13, inputRegisters_138__12, 
         inputRegisters_138__11, inputRegisters_138__10, inputRegisters_138__9, 
         inputRegisters_138__8, inputRegisters_138__7, inputRegisters_138__6, 
         inputRegisters_138__5, inputRegisters_138__4, inputRegisters_138__3, 
         inputRegisters_138__2, inputRegisters_138__1, inputRegisters_138__0, 
         inputRegisters_139__15, inputRegisters_139__14, inputRegisters_139__13, 
         inputRegisters_139__12, inputRegisters_139__11, inputRegisters_139__10, 
         inputRegisters_139__9, inputRegisters_139__8, inputRegisters_139__7, 
         inputRegisters_139__6, inputRegisters_139__5, inputRegisters_139__4, 
         inputRegisters_139__3, inputRegisters_139__2, inputRegisters_139__1, 
         inputRegisters_139__0, inputRegisters_140__15, inputRegisters_140__14, 
         inputRegisters_140__13, inputRegisters_140__12, inputRegisters_140__11, 
         inputRegisters_140__10, inputRegisters_140__9, inputRegisters_140__8, 
         inputRegisters_140__7, inputRegisters_140__6, inputRegisters_140__5, 
         inputRegisters_140__4, inputRegisters_140__3, inputRegisters_140__2, 
         inputRegisters_140__1, inputRegisters_140__0, inputRegisters_141__15, 
         inputRegisters_141__14, inputRegisters_141__13, inputRegisters_141__12, 
         inputRegisters_141__11, inputRegisters_141__10, inputRegisters_141__9, 
         inputRegisters_141__8, inputRegisters_141__7, inputRegisters_141__6, 
         inputRegisters_141__5, inputRegisters_141__4, inputRegisters_141__3, 
         inputRegisters_141__2, inputRegisters_141__1, inputRegisters_141__0, 
         inputRegisters_142__15, inputRegisters_142__14, inputRegisters_142__13, 
         inputRegisters_142__12, inputRegisters_142__11, inputRegisters_142__10, 
         inputRegisters_142__9, inputRegisters_142__8, inputRegisters_142__7, 
         inputRegisters_142__6, inputRegisters_142__5, inputRegisters_142__4, 
         inputRegisters_142__3, inputRegisters_142__2, inputRegisters_142__1, 
         inputRegisters_142__0, inputRegisters_143__15, inputRegisters_143__14, 
         inputRegisters_143__13, inputRegisters_143__12, inputRegisters_143__11, 
         inputRegisters_143__10, inputRegisters_143__9, inputRegisters_143__8, 
         inputRegisters_143__7, inputRegisters_143__6, inputRegisters_143__5, 
         inputRegisters_143__4, inputRegisters_143__3, inputRegisters_143__2, 
         inputRegisters_143__1, inputRegisters_143__0, inputRegisters_144__15, 
         inputRegisters_144__14, inputRegisters_144__13, inputRegisters_144__12, 
         inputRegisters_144__11, inputRegisters_144__10, inputRegisters_144__9, 
         inputRegisters_144__8, inputRegisters_144__7, inputRegisters_144__6, 
         inputRegisters_144__5, inputRegisters_144__4, inputRegisters_144__3, 
         inputRegisters_144__2, inputRegisters_144__1, inputRegisters_144__0, 
         inputRegisters_145__15, inputRegisters_145__14, inputRegisters_145__13, 
         inputRegisters_145__12, inputRegisters_145__11, inputRegisters_145__10, 
         inputRegisters_145__9, inputRegisters_145__8, inputRegisters_145__7, 
         inputRegisters_145__6, inputRegisters_145__5, inputRegisters_145__4, 
         inputRegisters_145__3, inputRegisters_145__2, inputRegisters_145__1, 
         inputRegisters_145__0, inputRegisters_146__15, inputRegisters_146__14, 
         inputRegisters_146__13, inputRegisters_146__12, inputRegisters_146__11, 
         inputRegisters_146__10, inputRegisters_146__9, inputRegisters_146__8, 
         inputRegisters_146__7, inputRegisters_146__6, inputRegisters_146__5, 
         inputRegisters_146__4, inputRegisters_146__3, inputRegisters_146__2, 
         inputRegisters_146__1, inputRegisters_146__0, inputRegisters_147__15, 
         inputRegisters_147__14, inputRegisters_147__13, inputRegisters_147__12, 
         inputRegisters_147__11, inputRegisters_147__10, inputRegisters_147__9, 
         inputRegisters_147__8, inputRegisters_147__7, inputRegisters_147__6, 
         inputRegisters_147__5, inputRegisters_147__4, inputRegisters_147__3, 
         inputRegisters_147__2, inputRegisters_147__1, inputRegisters_147__0, 
         inputRegisters_148__15, inputRegisters_148__14, inputRegisters_148__13, 
         inputRegisters_148__12, inputRegisters_148__11, inputRegisters_148__10, 
         inputRegisters_148__9, inputRegisters_148__8, inputRegisters_148__7, 
         inputRegisters_148__6, inputRegisters_148__5, inputRegisters_148__4, 
         inputRegisters_148__3, inputRegisters_148__2, inputRegisters_148__1, 
         inputRegisters_148__0, inputRegisters_149__15, inputRegisters_149__14, 
         inputRegisters_149__13, inputRegisters_149__12, inputRegisters_149__11, 
         inputRegisters_149__10, inputRegisters_149__9, inputRegisters_149__8, 
         inputRegisters_149__7, inputRegisters_149__6, inputRegisters_149__5, 
         inputRegisters_149__4, inputRegisters_149__3, inputRegisters_149__2, 
         inputRegisters_149__1, inputRegisters_149__0, inputRegisters_150__15, 
         inputRegisters_150__14, inputRegisters_150__13, inputRegisters_150__12, 
         inputRegisters_150__11, inputRegisters_150__10, inputRegisters_150__9, 
         inputRegisters_150__8, inputRegisters_150__7, inputRegisters_150__6, 
         inputRegisters_150__5, inputRegisters_150__4, inputRegisters_150__3, 
         inputRegisters_150__2, inputRegisters_150__1, inputRegisters_150__0, 
         inputRegisters_151__15, inputRegisters_151__14, inputRegisters_151__13, 
         inputRegisters_151__12, inputRegisters_151__11, inputRegisters_151__10, 
         inputRegisters_151__9, inputRegisters_151__8, inputRegisters_151__7, 
         inputRegisters_151__6, inputRegisters_151__5, inputRegisters_151__4, 
         inputRegisters_151__3, inputRegisters_151__2, inputRegisters_151__1, 
         inputRegisters_151__0, inputRegisters_152__15, inputRegisters_152__14, 
         inputRegisters_152__13, inputRegisters_152__12, inputRegisters_152__11, 
         inputRegisters_152__10, inputRegisters_152__9, inputRegisters_152__8, 
         inputRegisters_152__7, inputRegisters_152__6, inputRegisters_152__5, 
         inputRegisters_152__4, inputRegisters_152__3, inputRegisters_152__2, 
         inputRegisters_152__1, inputRegisters_152__0, inputRegisters_153__15, 
         inputRegisters_153__14, inputRegisters_153__13, inputRegisters_153__12, 
         inputRegisters_153__11, inputRegisters_153__10, inputRegisters_153__9, 
         inputRegisters_153__8, inputRegisters_153__7, inputRegisters_153__6, 
         inputRegisters_153__5, inputRegisters_153__4, inputRegisters_153__3, 
         inputRegisters_153__2, inputRegisters_153__1, inputRegisters_153__0, 
         inputRegisters_154__15, inputRegisters_154__14, inputRegisters_154__13, 
         inputRegisters_154__12, inputRegisters_154__11, inputRegisters_154__10, 
         inputRegisters_154__9, inputRegisters_154__8, inputRegisters_154__7, 
         inputRegisters_154__6, inputRegisters_154__5, inputRegisters_154__4, 
         inputRegisters_154__3, inputRegisters_154__2, inputRegisters_154__1, 
         inputRegisters_154__0, inputRegisters_155__15, inputRegisters_155__14, 
         inputRegisters_155__13, inputRegisters_155__12, inputRegisters_155__11, 
         inputRegisters_155__10, inputRegisters_155__9, inputRegisters_155__8, 
         inputRegisters_155__7, inputRegisters_155__6, inputRegisters_155__5, 
         inputRegisters_155__4, inputRegisters_155__3, inputRegisters_155__2, 
         inputRegisters_155__1, inputRegisters_155__0, inputRegisters_156__15, 
         inputRegisters_156__14, inputRegisters_156__13, inputRegisters_156__12, 
         inputRegisters_156__11, inputRegisters_156__10, inputRegisters_156__9, 
         inputRegisters_156__8, inputRegisters_156__7, inputRegisters_156__6, 
         inputRegisters_156__5, inputRegisters_156__4, inputRegisters_156__3, 
         inputRegisters_156__2, inputRegisters_156__1, inputRegisters_156__0, 
         inputRegisters_157__15, inputRegisters_157__14, inputRegisters_157__13, 
         inputRegisters_157__12, inputRegisters_157__11, inputRegisters_157__10, 
         inputRegisters_157__9, inputRegisters_157__8, inputRegisters_157__7, 
         inputRegisters_157__6, inputRegisters_157__5, inputRegisters_157__4, 
         inputRegisters_157__3, inputRegisters_157__2, inputRegisters_157__1, 
         inputRegisters_157__0, inputRegisters_158__15, inputRegisters_158__14, 
         inputRegisters_158__13, inputRegisters_158__12, inputRegisters_158__11, 
         inputRegisters_158__10, inputRegisters_158__9, inputRegisters_158__8, 
         inputRegisters_158__7, inputRegisters_158__6, inputRegisters_158__5, 
         inputRegisters_158__4, inputRegisters_158__3, inputRegisters_158__2, 
         inputRegisters_158__1, inputRegisters_158__0, inputRegisters_159__15, 
         inputRegisters_159__14, inputRegisters_159__13, inputRegisters_159__12, 
         inputRegisters_159__11, inputRegisters_159__10, inputRegisters_159__9, 
         inputRegisters_159__8, inputRegisters_159__7, inputRegisters_159__6, 
         inputRegisters_159__5, inputRegisters_159__4, inputRegisters_159__3, 
         inputRegisters_159__2, inputRegisters_159__1, inputRegisters_159__0, 
         inputRegisters_160__15, inputRegisters_160__14, inputRegisters_160__13, 
         inputRegisters_160__12, inputRegisters_160__11, inputRegisters_160__10, 
         inputRegisters_160__9, inputRegisters_160__8, inputRegisters_160__7, 
         inputRegisters_160__6, inputRegisters_160__5, inputRegisters_160__4, 
         inputRegisters_160__3, inputRegisters_160__2, inputRegisters_160__1, 
         inputRegisters_160__0, inputRegisters_161__15, inputRegisters_161__14, 
         inputRegisters_161__13, inputRegisters_161__12, inputRegisters_161__11, 
         inputRegisters_161__10, inputRegisters_161__9, inputRegisters_161__8, 
         inputRegisters_161__7, inputRegisters_161__6, inputRegisters_161__5, 
         inputRegisters_161__4, inputRegisters_161__3, inputRegisters_161__2, 
         inputRegisters_161__1, inputRegisters_161__0, inputRegisters_162__15, 
         inputRegisters_162__14, inputRegisters_162__13, inputRegisters_162__12, 
         inputRegisters_162__11, inputRegisters_162__10, inputRegisters_162__9, 
         inputRegisters_162__8, inputRegisters_162__7, inputRegisters_162__6, 
         inputRegisters_162__5, inputRegisters_162__4, inputRegisters_162__3, 
         inputRegisters_162__2, inputRegisters_162__1, inputRegisters_162__0, 
         inputRegisters_163__15, inputRegisters_163__14, inputRegisters_163__13, 
         inputRegisters_163__12, inputRegisters_163__11, inputRegisters_163__10, 
         inputRegisters_163__9, inputRegisters_163__8, inputRegisters_163__7, 
         inputRegisters_163__6, inputRegisters_163__5, inputRegisters_163__4, 
         inputRegisters_163__3, inputRegisters_163__2, inputRegisters_163__1, 
         inputRegisters_163__0, inputRegisters_164__15, inputRegisters_164__14, 
         inputRegisters_164__13, inputRegisters_164__12, inputRegisters_164__11, 
         inputRegisters_164__10, inputRegisters_164__9, inputRegisters_164__8, 
         inputRegisters_164__7, inputRegisters_164__6, inputRegisters_164__5, 
         inputRegisters_164__4, inputRegisters_164__3, inputRegisters_164__2, 
         inputRegisters_164__1, inputRegisters_164__0, inputRegisters_165__15, 
         inputRegisters_165__14, inputRegisters_165__13, inputRegisters_165__12, 
         inputRegisters_165__11, inputRegisters_165__10, inputRegisters_165__9, 
         inputRegisters_165__8, inputRegisters_165__7, inputRegisters_165__6, 
         inputRegisters_165__5, inputRegisters_165__4, inputRegisters_165__3, 
         inputRegisters_165__2, inputRegisters_165__1, inputRegisters_165__0, 
         inputRegisters_166__15, inputRegisters_166__14, inputRegisters_166__13, 
         inputRegisters_166__12, inputRegisters_166__11, inputRegisters_166__10, 
         inputRegisters_166__9, inputRegisters_166__8, inputRegisters_166__7, 
         inputRegisters_166__6, inputRegisters_166__5, inputRegisters_166__4, 
         inputRegisters_166__3, inputRegisters_166__2, inputRegisters_166__1, 
         inputRegisters_166__0, inputRegisters_167__15, inputRegisters_167__14, 
         inputRegisters_167__13, inputRegisters_167__12, inputRegisters_167__11, 
         inputRegisters_167__10, inputRegisters_167__9, inputRegisters_167__8, 
         inputRegisters_167__7, inputRegisters_167__6, inputRegisters_167__5, 
         inputRegisters_167__4, inputRegisters_167__3, inputRegisters_167__2, 
         inputRegisters_167__1, inputRegisters_167__0, inputRegisters_168__15, 
         inputRegisters_168__14, inputRegisters_168__13, inputRegisters_168__12, 
         inputRegisters_168__11, inputRegisters_168__10, inputRegisters_168__9, 
         inputRegisters_168__8, inputRegisters_168__7, inputRegisters_168__6, 
         inputRegisters_168__5, inputRegisters_168__4, inputRegisters_168__3, 
         inputRegisters_168__2, inputRegisters_168__1, inputRegisters_168__0, 
         inputRegisters_169__15, inputRegisters_169__14, inputRegisters_169__13, 
         inputRegisters_169__12, inputRegisters_169__11, inputRegisters_169__10, 
         inputRegisters_169__9, inputRegisters_169__8, inputRegisters_169__7, 
         inputRegisters_169__6, inputRegisters_169__5, inputRegisters_169__4, 
         inputRegisters_169__3, inputRegisters_169__2, inputRegisters_169__1, 
         inputRegisters_169__0, inputRegisters_170__15, inputRegisters_170__14, 
         inputRegisters_170__13, inputRegisters_170__12, inputRegisters_170__11, 
         inputRegisters_170__10, inputRegisters_170__9, inputRegisters_170__8, 
         inputRegisters_170__7, inputRegisters_170__6, inputRegisters_170__5, 
         inputRegisters_170__4, inputRegisters_170__3, inputRegisters_170__2, 
         inputRegisters_170__1, inputRegisters_170__0, inputRegisters_171__15, 
         inputRegisters_171__14, inputRegisters_171__13, inputRegisters_171__12, 
         inputRegisters_171__11, inputRegisters_171__10, inputRegisters_171__9, 
         inputRegisters_171__8, inputRegisters_171__7, inputRegisters_171__6, 
         inputRegisters_171__5, inputRegisters_171__4, inputRegisters_171__3, 
         inputRegisters_171__2, inputRegisters_171__1, inputRegisters_171__0, 
         inputRegisters_172__15, inputRegisters_172__14, inputRegisters_172__13, 
         inputRegisters_172__12, inputRegisters_172__11, inputRegisters_172__10, 
         inputRegisters_172__9, inputRegisters_172__8, inputRegisters_172__7, 
         inputRegisters_172__6, inputRegisters_172__5, inputRegisters_172__4, 
         inputRegisters_172__3, inputRegisters_172__2, inputRegisters_172__1, 
         inputRegisters_172__0, inputRegisters_173__15, inputRegisters_173__14, 
         inputRegisters_173__13, inputRegisters_173__12, inputRegisters_173__11, 
         inputRegisters_173__10, inputRegisters_173__9, inputRegisters_173__8, 
         inputRegisters_173__7, inputRegisters_173__6, inputRegisters_173__5, 
         inputRegisters_173__4, inputRegisters_173__3, inputRegisters_173__2, 
         inputRegisters_173__1, inputRegisters_173__0, inputRegisters_174__15, 
         inputRegisters_174__14, inputRegisters_174__13, inputRegisters_174__12, 
         inputRegisters_174__11, inputRegisters_174__10, inputRegisters_174__9, 
         inputRegisters_174__8, inputRegisters_174__7, inputRegisters_174__6, 
         inputRegisters_174__5, inputRegisters_174__4, inputRegisters_174__3, 
         inputRegisters_174__2, inputRegisters_174__1, inputRegisters_174__0, 
         inputRegisters_175__15, inputRegisters_175__14, inputRegisters_175__13, 
         inputRegisters_175__12, inputRegisters_175__11, inputRegisters_175__10, 
         inputRegisters_175__9, inputRegisters_175__8, inputRegisters_175__7, 
         inputRegisters_175__6, inputRegisters_175__5, inputRegisters_175__4, 
         inputRegisters_175__3, inputRegisters_175__2, inputRegisters_175__1, 
         inputRegisters_175__0, inputRegisters_176__15, inputRegisters_176__14, 
         inputRegisters_176__13, inputRegisters_176__12, inputRegisters_176__11, 
         inputRegisters_176__10, inputRegisters_176__9, inputRegisters_176__8, 
         inputRegisters_176__7, inputRegisters_176__6, inputRegisters_176__5, 
         inputRegisters_176__4, inputRegisters_176__3, inputRegisters_176__2, 
         inputRegisters_176__1, inputRegisters_176__0, inputRegisters_177__15, 
         inputRegisters_177__14, inputRegisters_177__13, inputRegisters_177__12, 
         inputRegisters_177__11, inputRegisters_177__10, inputRegisters_177__9, 
         inputRegisters_177__8, inputRegisters_177__7, inputRegisters_177__6, 
         inputRegisters_177__5, inputRegisters_177__4, inputRegisters_177__3, 
         inputRegisters_177__2, inputRegisters_177__1, inputRegisters_177__0, 
         inputRegisters_178__15, inputRegisters_178__14, inputRegisters_178__13, 
         inputRegisters_178__12, inputRegisters_178__11, inputRegisters_178__10, 
         inputRegisters_178__9, inputRegisters_178__8, inputRegisters_178__7, 
         inputRegisters_178__6, inputRegisters_178__5, inputRegisters_178__4, 
         inputRegisters_178__3, inputRegisters_178__2, inputRegisters_178__1, 
         inputRegisters_178__0, inputRegisters_179__15, inputRegisters_179__14, 
         inputRegisters_179__13, inputRegisters_179__12, inputRegisters_179__11, 
         inputRegisters_179__10, inputRegisters_179__9, inputRegisters_179__8, 
         inputRegisters_179__7, inputRegisters_179__6, inputRegisters_179__5, 
         inputRegisters_179__4, inputRegisters_179__3, inputRegisters_179__2, 
         inputRegisters_179__1, inputRegisters_179__0, inputRegisters_180__15, 
         inputRegisters_180__14, inputRegisters_180__13, inputRegisters_180__12, 
         inputRegisters_180__11, inputRegisters_180__10, inputRegisters_180__9, 
         inputRegisters_180__8, inputRegisters_180__7, inputRegisters_180__6, 
         inputRegisters_180__5, inputRegisters_180__4, inputRegisters_180__3, 
         inputRegisters_180__2, inputRegisters_180__1, inputRegisters_180__0, 
         inputRegisters_181__15, inputRegisters_181__14, inputRegisters_181__13, 
         inputRegisters_181__12, inputRegisters_181__11, inputRegisters_181__10, 
         inputRegisters_181__9, inputRegisters_181__8, inputRegisters_181__7, 
         inputRegisters_181__6, inputRegisters_181__5, inputRegisters_181__4, 
         inputRegisters_181__3, inputRegisters_181__2, inputRegisters_181__1, 
         inputRegisters_181__0, inputRegisters_182__15, inputRegisters_182__14, 
         inputRegisters_182__13, inputRegisters_182__12, inputRegisters_182__11, 
         inputRegisters_182__10, inputRegisters_182__9, inputRegisters_182__8, 
         inputRegisters_182__7, inputRegisters_182__6, inputRegisters_182__5, 
         inputRegisters_182__4, inputRegisters_182__3, inputRegisters_182__2, 
         inputRegisters_182__1, inputRegisters_182__0, inputRegisters_183__15, 
         inputRegisters_183__14, inputRegisters_183__13, inputRegisters_183__12, 
         inputRegisters_183__11, inputRegisters_183__10, inputRegisters_183__9, 
         inputRegisters_183__8, inputRegisters_183__7, inputRegisters_183__6, 
         inputRegisters_183__5, inputRegisters_183__4, inputRegisters_183__3, 
         inputRegisters_183__2, inputRegisters_183__1, inputRegisters_183__0, 
         inputRegisters_184__15, inputRegisters_184__14, inputRegisters_184__13, 
         inputRegisters_184__12, inputRegisters_184__11, inputRegisters_184__10, 
         inputRegisters_184__9, inputRegisters_184__8, inputRegisters_184__7, 
         inputRegisters_184__6, inputRegisters_184__5, inputRegisters_184__4, 
         inputRegisters_184__3, inputRegisters_184__2, inputRegisters_184__1, 
         inputRegisters_184__0, inputRegisters_185__15, inputRegisters_185__14, 
         inputRegisters_185__13, inputRegisters_185__12, inputRegisters_185__11, 
         inputRegisters_185__10, inputRegisters_185__9, inputRegisters_185__8, 
         inputRegisters_185__7, inputRegisters_185__6, inputRegisters_185__5, 
         inputRegisters_185__4, inputRegisters_185__3, inputRegisters_185__2, 
         inputRegisters_185__1, inputRegisters_185__0, inputRegisters_186__15, 
         inputRegisters_186__14, inputRegisters_186__13, inputRegisters_186__12, 
         inputRegisters_186__11, inputRegisters_186__10, inputRegisters_186__9, 
         inputRegisters_186__8, inputRegisters_186__7, inputRegisters_186__6, 
         inputRegisters_186__5, inputRegisters_186__4, inputRegisters_186__3, 
         inputRegisters_186__2, inputRegisters_186__1, inputRegisters_186__0, 
         inputRegisters_187__15, inputRegisters_187__14, inputRegisters_187__13, 
         inputRegisters_187__12, inputRegisters_187__11, inputRegisters_187__10, 
         inputRegisters_187__9, inputRegisters_187__8, inputRegisters_187__7, 
         inputRegisters_187__6, inputRegisters_187__5, inputRegisters_187__4, 
         inputRegisters_187__3, inputRegisters_187__2, inputRegisters_187__1, 
         inputRegisters_187__0, inputRegisters_188__15, inputRegisters_188__14, 
         inputRegisters_188__13, inputRegisters_188__12, inputRegisters_188__11, 
         inputRegisters_188__10, inputRegisters_188__9, inputRegisters_188__8, 
         inputRegisters_188__7, inputRegisters_188__6, inputRegisters_188__5, 
         inputRegisters_188__4, inputRegisters_188__3, inputRegisters_188__2, 
         inputRegisters_188__1, inputRegisters_188__0, inputRegisters_189__15, 
         inputRegisters_189__14, inputRegisters_189__13, inputRegisters_189__12, 
         inputRegisters_189__11, inputRegisters_189__10, inputRegisters_189__9, 
         inputRegisters_189__8, inputRegisters_189__7, inputRegisters_189__6, 
         inputRegisters_189__5, inputRegisters_189__4, inputRegisters_189__3, 
         inputRegisters_189__2, inputRegisters_189__1, inputRegisters_189__0, 
         inputRegisters_190__15, inputRegisters_190__14, inputRegisters_190__13, 
         inputRegisters_190__12, inputRegisters_190__11, inputRegisters_190__10, 
         inputRegisters_190__9, inputRegisters_190__8, inputRegisters_190__7, 
         inputRegisters_190__6, inputRegisters_190__5, inputRegisters_190__4, 
         inputRegisters_190__3, inputRegisters_190__2, inputRegisters_190__1, 
         inputRegisters_190__0, inputRegisters_191__15, inputRegisters_191__14, 
         inputRegisters_191__13, inputRegisters_191__12, inputRegisters_191__11, 
         inputRegisters_191__10, inputRegisters_191__9, inputRegisters_191__8, 
         inputRegisters_191__7, inputRegisters_191__6, inputRegisters_191__5, 
         inputRegisters_191__4, inputRegisters_191__3, inputRegisters_191__2, 
         inputRegisters_191__1, inputRegisters_191__0, inputRegisters_192__15, 
         inputRegisters_192__14, inputRegisters_192__13, inputRegisters_192__12, 
         inputRegisters_192__11, inputRegisters_192__10, inputRegisters_192__9, 
         inputRegisters_192__8, inputRegisters_192__7, inputRegisters_192__6, 
         inputRegisters_192__5, inputRegisters_192__4, inputRegisters_192__3, 
         inputRegisters_192__2, inputRegisters_192__1, inputRegisters_192__0, 
         inputRegisters_193__15, inputRegisters_193__14, inputRegisters_193__13, 
         inputRegisters_193__12, inputRegisters_193__11, inputRegisters_193__10, 
         inputRegisters_193__9, inputRegisters_193__8, inputRegisters_193__7, 
         inputRegisters_193__6, inputRegisters_193__5, inputRegisters_193__4, 
         inputRegisters_193__3, inputRegisters_193__2, inputRegisters_193__1, 
         inputRegisters_193__0, inputRegisters_194__15, inputRegisters_194__14, 
         inputRegisters_194__13, inputRegisters_194__12, inputRegisters_194__11, 
         inputRegisters_194__10, inputRegisters_194__9, inputRegisters_194__8, 
         inputRegisters_194__7, inputRegisters_194__6, inputRegisters_194__5, 
         inputRegisters_194__4, inputRegisters_194__3, inputRegisters_194__2, 
         inputRegisters_194__1, inputRegisters_194__0, inputRegisters_195__15, 
         inputRegisters_195__14, inputRegisters_195__13, inputRegisters_195__12, 
         inputRegisters_195__11, inputRegisters_195__10, inputRegisters_195__9, 
         inputRegisters_195__8, inputRegisters_195__7, inputRegisters_195__6, 
         inputRegisters_195__5, inputRegisters_195__4, inputRegisters_195__3, 
         inputRegisters_195__2, inputRegisters_195__1, inputRegisters_195__0, 
         inputRegisters_196__15, inputRegisters_196__14, inputRegisters_196__13, 
         inputRegisters_196__12, inputRegisters_196__11, inputRegisters_196__10, 
         inputRegisters_196__9, inputRegisters_196__8, inputRegisters_196__7, 
         inputRegisters_196__6, inputRegisters_196__5, inputRegisters_196__4, 
         inputRegisters_196__3, inputRegisters_196__2, inputRegisters_196__1, 
         inputRegisters_196__0, inputRegisters_197__15, inputRegisters_197__14, 
         inputRegisters_197__13, inputRegisters_197__12, inputRegisters_197__11, 
         inputRegisters_197__10, inputRegisters_197__9, inputRegisters_197__8, 
         inputRegisters_197__7, inputRegisters_197__6, inputRegisters_197__5, 
         inputRegisters_197__4, inputRegisters_197__3, inputRegisters_197__2, 
         inputRegisters_197__1, inputRegisters_197__0, inputRegisters_198__15, 
         inputRegisters_198__14, inputRegisters_198__13, inputRegisters_198__12, 
         inputRegisters_198__11, inputRegisters_198__10, inputRegisters_198__9, 
         inputRegisters_198__8, inputRegisters_198__7, inputRegisters_198__6, 
         inputRegisters_198__5, inputRegisters_198__4, inputRegisters_198__3, 
         inputRegisters_198__2, inputRegisters_198__1, inputRegisters_198__0, 
         inputRegisters_199__15, inputRegisters_199__14, inputRegisters_199__13, 
         inputRegisters_199__12, inputRegisters_199__11, inputRegisters_199__10, 
         inputRegisters_199__9, inputRegisters_199__8, inputRegisters_199__7, 
         inputRegisters_199__6, inputRegisters_199__5, inputRegisters_199__4, 
         inputRegisters_199__3, inputRegisters_199__2, inputRegisters_199__1, 
         inputRegisters_199__0, inputRegisters_200__15, inputRegisters_200__14, 
         inputRegisters_200__13, inputRegisters_200__12, inputRegisters_200__11, 
         inputRegisters_200__10, inputRegisters_200__9, inputRegisters_200__8, 
         inputRegisters_200__7, inputRegisters_200__6, inputRegisters_200__5, 
         inputRegisters_200__4, inputRegisters_200__3, inputRegisters_200__2, 
         inputRegisters_200__1, inputRegisters_200__0, inputRegisters_201__15, 
         inputRegisters_201__14, inputRegisters_201__13, inputRegisters_201__12, 
         inputRegisters_201__11, inputRegisters_201__10, inputRegisters_201__9, 
         inputRegisters_201__8, inputRegisters_201__7, inputRegisters_201__6, 
         inputRegisters_201__5, inputRegisters_201__4, inputRegisters_201__3, 
         inputRegisters_201__2, inputRegisters_201__1, inputRegisters_201__0, 
         inputRegisters_202__15, inputRegisters_202__14, inputRegisters_202__13, 
         inputRegisters_202__12, inputRegisters_202__11, inputRegisters_202__10, 
         inputRegisters_202__9, inputRegisters_202__8, inputRegisters_202__7, 
         inputRegisters_202__6, inputRegisters_202__5, inputRegisters_202__4, 
         inputRegisters_202__3, inputRegisters_202__2, inputRegisters_202__1, 
         inputRegisters_202__0, inputRegisters_203__15, inputRegisters_203__14, 
         inputRegisters_203__13, inputRegisters_203__12, inputRegisters_203__11, 
         inputRegisters_203__10, inputRegisters_203__9, inputRegisters_203__8, 
         inputRegisters_203__7, inputRegisters_203__6, inputRegisters_203__5, 
         inputRegisters_203__4, inputRegisters_203__3, inputRegisters_203__2, 
         inputRegisters_203__1, inputRegisters_203__0, inputRegisters_204__15, 
         inputRegisters_204__14, inputRegisters_204__13, inputRegisters_204__12, 
         inputRegisters_204__11, inputRegisters_204__10, inputRegisters_204__9, 
         inputRegisters_204__8, inputRegisters_204__7, inputRegisters_204__6, 
         inputRegisters_204__5, inputRegisters_204__4, inputRegisters_204__3, 
         inputRegisters_204__2, inputRegisters_204__1, inputRegisters_204__0, 
         inputRegisters_205__15, inputRegisters_205__14, inputRegisters_205__13, 
         inputRegisters_205__12, inputRegisters_205__11, inputRegisters_205__10, 
         inputRegisters_205__9, inputRegisters_205__8, inputRegisters_205__7, 
         inputRegisters_205__6, inputRegisters_205__5, inputRegisters_205__4, 
         inputRegisters_205__3, inputRegisters_205__2, inputRegisters_205__1, 
         inputRegisters_205__0, inputRegisters_206__15, inputRegisters_206__14, 
         inputRegisters_206__13, inputRegisters_206__12, inputRegisters_206__11, 
         inputRegisters_206__10, inputRegisters_206__9, inputRegisters_206__8, 
         inputRegisters_206__7, inputRegisters_206__6, inputRegisters_206__5, 
         inputRegisters_206__4, inputRegisters_206__3, inputRegisters_206__2, 
         inputRegisters_206__1, inputRegisters_206__0, inputRegisters_207__15, 
         inputRegisters_207__14, inputRegisters_207__13, inputRegisters_207__12, 
         inputRegisters_207__11, inputRegisters_207__10, inputRegisters_207__9, 
         inputRegisters_207__8, inputRegisters_207__7, inputRegisters_207__6, 
         inputRegisters_207__5, inputRegisters_207__4, inputRegisters_207__3, 
         inputRegisters_207__2, inputRegisters_207__1, inputRegisters_207__0, 
         inputRegisters_208__15, inputRegisters_208__14, inputRegisters_208__13, 
         inputRegisters_208__12, inputRegisters_208__11, inputRegisters_208__10, 
         inputRegisters_208__9, inputRegisters_208__8, inputRegisters_208__7, 
         inputRegisters_208__6, inputRegisters_208__5, inputRegisters_208__4, 
         inputRegisters_208__3, inputRegisters_208__2, inputRegisters_208__1, 
         inputRegisters_208__0, inputRegisters_209__15, inputRegisters_209__14, 
         inputRegisters_209__13, inputRegisters_209__12, inputRegisters_209__11, 
         inputRegisters_209__10, inputRegisters_209__9, inputRegisters_209__8, 
         inputRegisters_209__7, inputRegisters_209__6, inputRegisters_209__5, 
         inputRegisters_209__4, inputRegisters_209__3, inputRegisters_209__2, 
         inputRegisters_209__1, inputRegisters_209__0, inputRegisters_210__15, 
         inputRegisters_210__14, inputRegisters_210__13, inputRegisters_210__12, 
         inputRegisters_210__11, inputRegisters_210__10, inputRegisters_210__9, 
         inputRegisters_210__8, inputRegisters_210__7, inputRegisters_210__6, 
         inputRegisters_210__5, inputRegisters_210__4, inputRegisters_210__3, 
         inputRegisters_210__2, inputRegisters_210__1, inputRegisters_210__0, 
         inputRegisters_211__15, inputRegisters_211__14, inputRegisters_211__13, 
         inputRegisters_211__12, inputRegisters_211__11, inputRegisters_211__10, 
         inputRegisters_211__9, inputRegisters_211__8, inputRegisters_211__7, 
         inputRegisters_211__6, inputRegisters_211__5, inputRegisters_211__4, 
         inputRegisters_211__3, inputRegisters_211__2, inputRegisters_211__1, 
         inputRegisters_211__0, inputRegisters_212__15, inputRegisters_212__14, 
         inputRegisters_212__13, inputRegisters_212__12, inputRegisters_212__11, 
         inputRegisters_212__10, inputRegisters_212__9, inputRegisters_212__8, 
         inputRegisters_212__7, inputRegisters_212__6, inputRegisters_212__5, 
         inputRegisters_212__4, inputRegisters_212__3, inputRegisters_212__2, 
         inputRegisters_212__1, inputRegisters_212__0, inputRegisters_213__15, 
         inputRegisters_213__14, inputRegisters_213__13, inputRegisters_213__12, 
         inputRegisters_213__11, inputRegisters_213__10, inputRegisters_213__9, 
         inputRegisters_213__8, inputRegisters_213__7, inputRegisters_213__6, 
         inputRegisters_213__5, inputRegisters_213__4, inputRegisters_213__3, 
         inputRegisters_213__2, inputRegisters_213__1, inputRegisters_213__0, 
         inputRegisters_214__15, inputRegisters_214__14, inputRegisters_214__13, 
         inputRegisters_214__12, inputRegisters_214__11, inputRegisters_214__10, 
         inputRegisters_214__9, inputRegisters_214__8, inputRegisters_214__7, 
         inputRegisters_214__6, inputRegisters_214__5, inputRegisters_214__4, 
         inputRegisters_214__3, inputRegisters_214__2, inputRegisters_214__1, 
         inputRegisters_214__0, inputRegisters_215__15, inputRegisters_215__14, 
         inputRegisters_215__13, inputRegisters_215__12, inputRegisters_215__11, 
         inputRegisters_215__10, inputRegisters_215__9, inputRegisters_215__8, 
         inputRegisters_215__7, inputRegisters_215__6, inputRegisters_215__5, 
         inputRegisters_215__4, inputRegisters_215__3, inputRegisters_215__2, 
         inputRegisters_215__1, inputRegisters_215__0, inputRegisters_216__15, 
         inputRegisters_216__14, inputRegisters_216__13, inputRegisters_216__12, 
         inputRegisters_216__11, inputRegisters_216__10, inputRegisters_216__9, 
         inputRegisters_216__8, inputRegisters_216__7, inputRegisters_216__6, 
         inputRegisters_216__5, inputRegisters_216__4, inputRegisters_216__3, 
         inputRegisters_216__2, inputRegisters_216__1, inputRegisters_216__0, 
         inputRegisters_217__15, inputRegisters_217__14, inputRegisters_217__13, 
         inputRegisters_217__12, inputRegisters_217__11, inputRegisters_217__10, 
         inputRegisters_217__9, inputRegisters_217__8, inputRegisters_217__7, 
         inputRegisters_217__6, inputRegisters_217__5, inputRegisters_217__4, 
         inputRegisters_217__3, inputRegisters_217__2, inputRegisters_217__1, 
         inputRegisters_217__0, inputRegisters_218__15, inputRegisters_218__14, 
         inputRegisters_218__13, inputRegisters_218__12, inputRegisters_218__11, 
         inputRegisters_218__10, inputRegisters_218__9, inputRegisters_218__8, 
         inputRegisters_218__7, inputRegisters_218__6, inputRegisters_218__5, 
         inputRegisters_218__4, inputRegisters_218__3, inputRegisters_218__2, 
         inputRegisters_218__1, inputRegisters_218__0, inputRegisters_219__15, 
         inputRegisters_219__14, inputRegisters_219__13, inputRegisters_219__12, 
         inputRegisters_219__11, inputRegisters_219__10, inputRegisters_219__9, 
         inputRegisters_219__8, inputRegisters_219__7, inputRegisters_219__6, 
         inputRegisters_219__5, inputRegisters_219__4, inputRegisters_219__3, 
         inputRegisters_219__2, inputRegisters_219__1, inputRegisters_219__0, 
         inputRegisters_220__15, inputRegisters_220__14, inputRegisters_220__13, 
         inputRegisters_220__12, inputRegisters_220__11, inputRegisters_220__10, 
         inputRegisters_220__9, inputRegisters_220__8, inputRegisters_220__7, 
         inputRegisters_220__6, inputRegisters_220__5, inputRegisters_220__4, 
         inputRegisters_220__3, inputRegisters_220__2, inputRegisters_220__1, 
         inputRegisters_220__0, inputRegisters_221__15, inputRegisters_221__14, 
         inputRegisters_221__13, inputRegisters_221__12, inputRegisters_221__11, 
         inputRegisters_221__10, inputRegisters_221__9, inputRegisters_221__8, 
         inputRegisters_221__7, inputRegisters_221__6, inputRegisters_221__5, 
         inputRegisters_221__4, inputRegisters_221__3, inputRegisters_221__2, 
         inputRegisters_221__1, inputRegisters_221__0, inputRegisters_222__15, 
         inputRegisters_222__14, inputRegisters_222__13, inputRegisters_222__12, 
         inputRegisters_222__11, inputRegisters_222__10, inputRegisters_222__9, 
         inputRegisters_222__8, inputRegisters_222__7, inputRegisters_222__6, 
         inputRegisters_222__5, inputRegisters_222__4, inputRegisters_222__3, 
         inputRegisters_222__2, inputRegisters_222__1, inputRegisters_222__0, 
         inputRegisters_223__15, inputRegisters_223__14, inputRegisters_223__13, 
         inputRegisters_223__12, inputRegisters_223__11, inputRegisters_223__10, 
         inputRegisters_223__9, inputRegisters_223__8, inputRegisters_223__7, 
         inputRegisters_223__6, inputRegisters_223__5, inputRegisters_223__4, 
         inputRegisters_223__3, inputRegisters_223__2, inputRegisters_223__1, 
         inputRegisters_223__0, inputRegisters_224__15, inputRegisters_224__14, 
         inputRegisters_224__13, inputRegisters_224__12, inputRegisters_224__11, 
         inputRegisters_224__10, inputRegisters_224__9, inputRegisters_224__8, 
         inputRegisters_224__7, inputRegisters_224__6, inputRegisters_224__5, 
         inputRegisters_224__4, inputRegisters_224__3, inputRegisters_224__2, 
         inputRegisters_224__1, inputRegisters_224__0, inputRegisters_225__15, 
         inputRegisters_225__14, inputRegisters_225__13, inputRegisters_225__12, 
         inputRegisters_225__11, inputRegisters_225__10, inputRegisters_225__9, 
         inputRegisters_225__8, inputRegisters_225__7, inputRegisters_225__6, 
         inputRegisters_225__5, inputRegisters_225__4, inputRegisters_225__3, 
         inputRegisters_225__2, inputRegisters_225__1, inputRegisters_225__0, 
         inputRegisters_226__15, inputRegisters_226__14, inputRegisters_226__13, 
         inputRegisters_226__12, inputRegisters_226__11, inputRegisters_226__10, 
         inputRegisters_226__9, inputRegisters_226__8, inputRegisters_226__7, 
         inputRegisters_226__6, inputRegisters_226__5, inputRegisters_226__4, 
         inputRegisters_226__3, inputRegisters_226__2, inputRegisters_226__1, 
         inputRegisters_226__0, inputRegisters_227__15, inputRegisters_227__14, 
         inputRegisters_227__13, inputRegisters_227__12, inputRegisters_227__11, 
         inputRegisters_227__10, inputRegisters_227__9, inputRegisters_227__8, 
         inputRegisters_227__7, inputRegisters_227__6, inputRegisters_227__5, 
         inputRegisters_227__4, inputRegisters_227__3, inputRegisters_227__2, 
         inputRegisters_227__1, inputRegisters_227__0, inputRegisters_228__15, 
         inputRegisters_228__14, inputRegisters_228__13, inputRegisters_228__12, 
         inputRegisters_228__11, inputRegisters_228__10, inputRegisters_228__9, 
         inputRegisters_228__8, inputRegisters_228__7, inputRegisters_228__6, 
         inputRegisters_228__5, inputRegisters_228__4, inputRegisters_228__3, 
         inputRegisters_228__2, inputRegisters_228__1, inputRegisters_228__0, 
         inputRegisters_229__15, inputRegisters_229__14, inputRegisters_229__13, 
         inputRegisters_229__12, inputRegisters_229__11, inputRegisters_229__10, 
         inputRegisters_229__9, inputRegisters_229__8, inputRegisters_229__7, 
         inputRegisters_229__6, inputRegisters_229__5, inputRegisters_229__4, 
         inputRegisters_229__3, inputRegisters_229__2, inputRegisters_229__1, 
         inputRegisters_229__0, inputRegisters_230__15, inputRegisters_230__14, 
         inputRegisters_230__13, inputRegisters_230__12, inputRegisters_230__11, 
         inputRegisters_230__10, inputRegisters_230__9, inputRegisters_230__8, 
         inputRegisters_230__7, inputRegisters_230__6, inputRegisters_230__5, 
         inputRegisters_230__4, inputRegisters_230__3, inputRegisters_230__2, 
         inputRegisters_230__1, inputRegisters_230__0, inputRegisters_231__15, 
         inputRegisters_231__14, inputRegisters_231__13, inputRegisters_231__12, 
         inputRegisters_231__11, inputRegisters_231__10, inputRegisters_231__9, 
         inputRegisters_231__8, inputRegisters_231__7, inputRegisters_231__6, 
         inputRegisters_231__5, inputRegisters_231__4, inputRegisters_231__3, 
         inputRegisters_231__2, inputRegisters_231__1, inputRegisters_231__0, 
         inputRegisters_232__15, inputRegisters_232__14, inputRegisters_232__13, 
         inputRegisters_232__12, inputRegisters_232__11, inputRegisters_232__10, 
         inputRegisters_232__9, inputRegisters_232__8, inputRegisters_232__7, 
         inputRegisters_232__6, inputRegisters_232__5, inputRegisters_232__4, 
         inputRegisters_232__3, inputRegisters_232__2, inputRegisters_232__1, 
         inputRegisters_232__0, inputRegisters_233__15, inputRegisters_233__14, 
         inputRegisters_233__13, inputRegisters_233__12, inputRegisters_233__11, 
         inputRegisters_233__10, inputRegisters_233__9, inputRegisters_233__8, 
         inputRegisters_233__7, inputRegisters_233__6, inputRegisters_233__5, 
         inputRegisters_233__4, inputRegisters_233__3, inputRegisters_233__2, 
         inputRegisters_233__1, inputRegisters_233__0, inputRegisters_234__15, 
         inputRegisters_234__14, inputRegisters_234__13, inputRegisters_234__12, 
         inputRegisters_234__11, inputRegisters_234__10, inputRegisters_234__9, 
         inputRegisters_234__8, inputRegisters_234__7, inputRegisters_234__6, 
         inputRegisters_234__5, inputRegisters_234__4, inputRegisters_234__3, 
         inputRegisters_234__2, inputRegisters_234__1, inputRegisters_234__0, 
         inputRegisters_235__15, inputRegisters_235__14, inputRegisters_235__13, 
         inputRegisters_235__12, inputRegisters_235__11, inputRegisters_235__10, 
         inputRegisters_235__9, inputRegisters_235__8, inputRegisters_235__7, 
         inputRegisters_235__6, inputRegisters_235__5, inputRegisters_235__4, 
         inputRegisters_235__3, inputRegisters_235__2, inputRegisters_235__1, 
         inputRegisters_235__0, inputRegisters_236__15, inputRegisters_236__14, 
         inputRegisters_236__13, inputRegisters_236__12, inputRegisters_236__11, 
         inputRegisters_236__10, inputRegisters_236__9, inputRegisters_236__8, 
         inputRegisters_236__7, inputRegisters_236__6, inputRegisters_236__5, 
         inputRegisters_236__4, inputRegisters_236__3, inputRegisters_236__2, 
         inputRegisters_236__1, inputRegisters_236__0, inputRegisters_237__15, 
         inputRegisters_237__14, inputRegisters_237__13, inputRegisters_237__12, 
         inputRegisters_237__11, inputRegisters_237__10, inputRegisters_237__9, 
         inputRegisters_237__8, inputRegisters_237__7, inputRegisters_237__6, 
         inputRegisters_237__5, inputRegisters_237__4, inputRegisters_237__3, 
         inputRegisters_237__2, inputRegisters_237__1, inputRegisters_237__0, 
         inputRegisters_238__15, inputRegisters_238__14, inputRegisters_238__13, 
         inputRegisters_238__12, inputRegisters_238__11, inputRegisters_238__10, 
         inputRegisters_238__9, inputRegisters_238__8, inputRegisters_238__7, 
         inputRegisters_238__6, inputRegisters_238__5, inputRegisters_238__4, 
         inputRegisters_238__3, inputRegisters_238__2, inputRegisters_238__1, 
         inputRegisters_238__0, inputRegisters_239__15, inputRegisters_239__14, 
         inputRegisters_239__13, inputRegisters_239__12, inputRegisters_239__11, 
         inputRegisters_239__10, inputRegisters_239__9, inputRegisters_239__8, 
         inputRegisters_239__7, inputRegisters_239__6, inputRegisters_239__5, 
         inputRegisters_239__4, inputRegisters_239__3, inputRegisters_239__2, 
         inputRegisters_239__1, inputRegisters_239__0, inputRegisters_240__15, 
         inputRegisters_240__14, inputRegisters_240__13, inputRegisters_240__12, 
         inputRegisters_240__11, inputRegisters_240__10, inputRegisters_240__9, 
         inputRegisters_240__8, inputRegisters_240__7, inputRegisters_240__6, 
         inputRegisters_240__5, inputRegisters_240__4, inputRegisters_240__3, 
         inputRegisters_240__2, inputRegisters_240__1, inputRegisters_240__0, 
         inputRegisters_241__15, inputRegisters_241__14, inputRegisters_241__13, 
         inputRegisters_241__12, inputRegisters_241__11, inputRegisters_241__10, 
         inputRegisters_241__9, inputRegisters_241__8, inputRegisters_241__7, 
         inputRegisters_241__6, inputRegisters_241__5, inputRegisters_241__4, 
         inputRegisters_241__3, inputRegisters_241__2, inputRegisters_241__1, 
         inputRegisters_241__0, inputRegisters_242__15, inputRegisters_242__14, 
         inputRegisters_242__13, inputRegisters_242__12, inputRegisters_242__11, 
         inputRegisters_242__10, inputRegisters_242__9, inputRegisters_242__8, 
         inputRegisters_242__7, inputRegisters_242__6, inputRegisters_242__5, 
         inputRegisters_242__4, inputRegisters_242__3, inputRegisters_242__2, 
         inputRegisters_242__1, inputRegisters_242__0, inputRegisters_243__15, 
         inputRegisters_243__14, inputRegisters_243__13, inputRegisters_243__12, 
         inputRegisters_243__11, inputRegisters_243__10, inputRegisters_243__9, 
         inputRegisters_243__8, inputRegisters_243__7, inputRegisters_243__6, 
         inputRegisters_243__5, inputRegisters_243__4, inputRegisters_243__3, 
         inputRegisters_243__2, inputRegisters_243__1, inputRegisters_243__0, 
         inputRegisters_244__15, inputRegisters_244__14, inputRegisters_244__13, 
         inputRegisters_244__12, inputRegisters_244__11, inputRegisters_244__10, 
         inputRegisters_244__9, inputRegisters_244__8, inputRegisters_244__7, 
         inputRegisters_244__6, inputRegisters_244__5, inputRegisters_244__4, 
         inputRegisters_244__3, inputRegisters_244__2, inputRegisters_244__1, 
         inputRegisters_244__0, inputRegisters_245__15, inputRegisters_245__14, 
         inputRegisters_245__13, inputRegisters_245__12, inputRegisters_245__11, 
         inputRegisters_245__10, inputRegisters_245__9, inputRegisters_245__8, 
         inputRegisters_245__7, inputRegisters_245__6, inputRegisters_245__5, 
         inputRegisters_245__4, inputRegisters_245__3, inputRegisters_245__2, 
         inputRegisters_245__1, inputRegisters_245__0, inputRegisters_246__15, 
         inputRegisters_246__14, inputRegisters_246__13, inputRegisters_246__12, 
         inputRegisters_246__11, inputRegisters_246__10, inputRegisters_246__9, 
         inputRegisters_246__8, inputRegisters_246__7, inputRegisters_246__6, 
         inputRegisters_246__5, inputRegisters_246__4, inputRegisters_246__3, 
         inputRegisters_246__2, inputRegisters_246__1, inputRegisters_246__0, 
         inputRegisters_247__15, inputRegisters_247__14, inputRegisters_247__13, 
         inputRegisters_247__12, inputRegisters_247__11, inputRegisters_247__10, 
         inputRegisters_247__9, inputRegisters_247__8, inputRegisters_247__7, 
         inputRegisters_247__6, inputRegisters_247__5, inputRegisters_247__4, 
         inputRegisters_247__3, inputRegisters_247__2, inputRegisters_247__1, 
         inputRegisters_247__0, inputRegisters_248__15, inputRegisters_248__14, 
         inputRegisters_248__13, inputRegisters_248__12, inputRegisters_248__11, 
         inputRegisters_248__10, inputRegisters_248__9, inputRegisters_248__8, 
         inputRegisters_248__7, inputRegisters_248__6, inputRegisters_248__5, 
         inputRegisters_248__4, inputRegisters_248__3, inputRegisters_248__2, 
         inputRegisters_248__1, inputRegisters_248__0, inputRegisters_249__15, 
         inputRegisters_249__14, inputRegisters_249__13, inputRegisters_249__12, 
         inputRegisters_249__11, inputRegisters_249__10, inputRegisters_249__9, 
         inputRegisters_249__8, inputRegisters_249__7, inputRegisters_249__6, 
         inputRegisters_249__5, inputRegisters_249__4, inputRegisters_249__3, 
         inputRegisters_249__2, inputRegisters_249__1, inputRegisters_249__0, 
         inputRegisters_250__15, inputRegisters_250__14, inputRegisters_250__13, 
         inputRegisters_250__12, inputRegisters_250__11, inputRegisters_250__10, 
         inputRegisters_250__9, inputRegisters_250__8, inputRegisters_250__7, 
         inputRegisters_250__6, inputRegisters_250__5, inputRegisters_250__4, 
         inputRegisters_250__3, inputRegisters_250__2, inputRegisters_250__1, 
         inputRegisters_250__0, inputRegisters_251__15, inputRegisters_251__14, 
         inputRegisters_251__13, inputRegisters_251__12, inputRegisters_251__11, 
         inputRegisters_251__10, inputRegisters_251__9, inputRegisters_251__8, 
         inputRegisters_251__7, inputRegisters_251__6, inputRegisters_251__5, 
         inputRegisters_251__4, inputRegisters_251__3, inputRegisters_251__2, 
         inputRegisters_251__1, inputRegisters_251__0, inputRegisters_252__15, 
         inputRegisters_252__14, inputRegisters_252__13, inputRegisters_252__12, 
         inputRegisters_252__11, inputRegisters_252__10, inputRegisters_252__9, 
         inputRegisters_252__8, inputRegisters_252__7, inputRegisters_252__6, 
         inputRegisters_252__5, inputRegisters_252__4, inputRegisters_252__3, 
         inputRegisters_252__2, inputRegisters_252__1, inputRegisters_252__0, 
         inputRegisters_253__15, inputRegisters_253__14, inputRegisters_253__13, 
         inputRegisters_253__12, inputRegisters_253__11, inputRegisters_253__10, 
         inputRegisters_253__9, inputRegisters_253__8, inputRegisters_253__7, 
         inputRegisters_253__6, inputRegisters_253__5, inputRegisters_253__4, 
         inputRegisters_253__3, inputRegisters_253__2, inputRegisters_253__1, 
         inputRegisters_253__0, inputRegisters_254__15, inputRegisters_254__14, 
         inputRegisters_254__13, inputRegisters_254__12, inputRegisters_254__11, 
         inputRegisters_254__10, inputRegisters_254__9, inputRegisters_254__8, 
         inputRegisters_254__7, inputRegisters_254__6, inputRegisters_254__5, 
         inputRegisters_254__4, inputRegisters_254__3, inputRegisters_254__2, 
         inputRegisters_254__1, inputRegisters_254__0, inputRegisters_255__15, 
         inputRegisters_255__14, inputRegisters_255__13, inputRegisters_255__12, 
         inputRegisters_255__11, inputRegisters_255__10, inputRegisters_255__9, 
         inputRegisters_255__8, inputRegisters_255__7, inputRegisters_255__6, 
         inputRegisters_255__5, inputRegisters_255__4, inputRegisters_255__3, 
         inputRegisters_255__2, inputRegisters_255__1, inputRegisters_255__0, 
         inputRegisters_256__15, inputRegisters_256__14, inputRegisters_256__13, 
         inputRegisters_256__12, inputRegisters_256__11, inputRegisters_256__10, 
         inputRegisters_256__9, inputRegisters_256__8, inputRegisters_256__7, 
         inputRegisters_256__6, inputRegisters_256__5, inputRegisters_256__4, 
         inputRegisters_256__3, inputRegisters_256__2, inputRegisters_256__1, 
         inputRegisters_256__0, inputRegisters_257__15, inputRegisters_257__14, 
         inputRegisters_257__13, inputRegisters_257__12, inputRegisters_257__11, 
         inputRegisters_257__10, inputRegisters_257__9, inputRegisters_257__8, 
         inputRegisters_257__7, inputRegisters_257__6, inputRegisters_257__5, 
         inputRegisters_257__4, inputRegisters_257__3, inputRegisters_257__2, 
         inputRegisters_257__1, inputRegisters_257__0, inputRegisters_258__15, 
         inputRegisters_258__14, inputRegisters_258__13, inputRegisters_258__12, 
         inputRegisters_258__11, inputRegisters_258__10, inputRegisters_258__9, 
         inputRegisters_258__8, inputRegisters_258__7, inputRegisters_258__6, 
         inputRegisters_258__5, inputRegisters_258__4, inputRegisters_258__3, 
         inputRegisters_258__2, inputRegisters_258__1, inputRegisters_258__0, 
         inputRegisters_259__15, inputRegisters_259__14, inputRegisters_259__13, 
         inputRegisters_259__12, inputRegisters_259__11, inputRegisters_259__10, 
         inputRegisters_259__9, inputRegisters_259__8, inputRegisters_259__7, 
         inputRegisters_259__6, inputRegisters_259__5, inputRegisters_259__4, 
         inputRegisters_259__3, inputRegisters_259__2, inputRegisters_259__1, 
         inputRegisters_259__0, inputRegisters_260__15, inputRegisters_260__14, 
         inputRegisters_260__13, inputRegisters_260__12, inputRegisters_260__11, 
         inputRegisters_260__10, inputRegisters_260__9, inputRegisters_260__8, 
         inputRegisters_260__7, inputRegisters_260__6, inputRegisters_260__5, 
         inputRegisters_260__4, inputRegisters_260__3, inputRegisters_260__2, 
         inputRegisters_260__1, inputRegisters_260__0, inputRegisters_261__15, 
         inputRegisters_261__14, inputRegisters_261__13, inputRegisters_261__12, 
         inputRegisters_261__11, inputRegisters_261__10, inputRegisters_261__9, 
         inputRegisters_261__8, inputRegisters_261__7, inputRegisters_261__6, 
         inputRegisters_261__5, inputRegisters_261__4, inputRegisters_261__3, 
         inputRegisters_261__2, inputRegisters_261__1, inputRegisters_261__0, 
         inputRegisters_262__15, inputRegisters_262__14, inputRegisters_262__13, 
         inputRegisters_262__12, inputRegisters_262__11, inputRegisters_262__10, 
         inputRegisters_262__9, inputRegisters_262__8, inputRegisters_262__7, 
         inputRegisters_262__6, inputRegisters_262__5, inputRegisters_262__4, 
         inputRegisters_262__3, inputRegisters_262__2, inputRegisters_262__1, 
         inputRegisters_262__0, inputRegisters_263__15, inputRegisters_263__14, 
         inputRegisters_263__13, inputRegisters_263__12, inputRegisters_263__11, 
         inputRegisters_263__10, inputRegisters_263__9, inputRegisters_263__8, 
         inputRegisters_263__7, inputRegisters_263__6, inputRegisters_263__5, 
         inputRegisters_263__4, inputRegisters_263__3, inputRegisters_263__2, 
         inputRegisters_263__1, inputRegisters_263__0, inputRegisters_264__15, 
         inputRegisters_264__14, inputRegisters_264__13, inputRegisters_264__12, 
         inputRegisters_264__11, inputRegisters_264__10, inputRegisters_264__9, 
         inputRegisters_264__8, inputRegisters_264__7, inputRegisters_264__6, 
         inputRegisters_264__5, inputRegisters_264__4, inputRegisters_264__3, 
         inputRegisters_264__2, inputRegisters_264__1, inputRegisters_264__0, 
         inputRegisters_265__15, inputRegisters_265__14, inputRegisters_265__13, 
         inputRegisters_265__12, inputRegisters_265__11, inputRegisters_265__10, 
         inputRegisters_265__9, inputRegisters_265__8, inputRegisters_265__7, 
         inputRegisters_265__6, inputRegisters_265__5, inputRegisters_265__4, 
         inputRegisters_265__3, inputRegisters_265__2, inputRegisters_265__1, 
         inputRegisters_265__0, inputRegisters_266__15, inputRegisters_266__14, 
         inputRegisters_266__13, inputRegisters_266__12, inputRegisters_266__11, 
         inputRegisters_266__10, inputRegisters_266__9, inputRegisters_266__8, 
         inputRegisters_266__7, inputRegisters_266__6, inputRegisters_266__5, 
         inputRegisters_266__4, inputRegisters_266__3, inputRegisters_266__2, 
         inputRegisters_266__1, inputRegisters_266__0, inputRegisters_267__15, 
         inputRegisters_267__14, inputRegisters_267__13, inputRegisters_267__12, 
         inputRegisters_267__11, inputRegisters_267__10, inputRegisters_267__9, 
         inputRegisters_267__8, inputRegisters_267__7, inputRegisters_267__6, 
         inputRegisters_267__5, inputRegisters_267__4, inputRegisters_267__3, 
         inputRegisters_267__2, inputRegisters_267__1, inputRegisters_267__0, 
         inputRegisters_268__15, inputRegisters_268__14, inputRegisters_268__13, 
         inputRegisters_268__12, inputRegisters_268__11, inputRegisters_268__10, 
         inputRegisters_268__9, inputRegisters_268__8, inputRegisters_268__7, 
         inputRegisters_268__6, inputRegisters_268__5, inputRegisters_268__4, 
         inputRegisters_268__3, inputRegisters_268__2, inputRegisters_268__1, 
         inputRegisters_268__0, inputRegisters_269__15, inputRegisters_269__14, 
         inputRegisters_269__13, inputRegisters_269__12, inputRegisters_269__11, 
         inputRegisters_269__10, inputRegisters_269__9, inputRegisters_269__8, 
         inputRegisters_269__7, inputRegisters_269__6, inputRegisters_269__5, 
         inputRegisters_269__4, inputRegisters_269__3, inputRegisters_269__2, 
         inputRegisters_269__1, inputRegisters_269__0, inputRegisters_270__15, 
         inputRegisters_270__14, inputRegisters_270__13, inputRegisters_270__12, 
         inputRegisters_270__11, inputRegisters_270__10, inputRegisters_270__9, 
         inputRegisters_270__8, inputRegisters_270__7, inputRegisters_270__6, 
         inputRegisters_270__5, inputRegisters_270__4, inputRegisters_270__3, 
         inputRegisters_270__2, inputRegisters_270__1, inputRegisters_270__0, 
         inputRegisters_271__15, inputRegisters_271__14, inputRegisters_271__13, 
         inputRegisters_271__12, inputRegisters_271__11, inputRegisters_271__10, 
         inputRegisters_271__9, inputRegisters_271__8, inputRegisters_271__7, 
         inputRegisters_271__6, inputRegisters_271__5, inputRegisters_271__4, 
         inputRegisters_271__3, inputRegisters_271__2, inputRegisters_271__1, 
         inputRegisters_271__0, inputRegisters_272__15, inputRegisters_272__14, 
         inputRegisters_272__13, inputRegisters_272__12, inputRegisters_272__11, 
         inputRegisters_272__10, inputRegisters_272__9, inputRegisters_272__8, 
         inputRegisters_272__7, inputRegisters_272__6, inputRegisters_272__5, 
         inputRegisters_272__4, inputRegisters_272__3, inputRegisters_272__2, 
         inputRegisters_272__1, inputRegisters_272__0, inputRegisters_273__15, 
         inputRegisters_273__14, inputRegisters_273__13, inputRegisters_273__12, 
         inputRegisters_273__11, inputRegisters_273__10, inputRegisters_273__9, 
         inputRegisters_273__8, inputRegisters_273__7, inputRegisters_273__6, 
         inputRegisters_273__5, inputRegisters_273__4, inputRegisters_273__3, 
         inputRegisters_273__2, inputRegisters_273__1, inputRegisters_273__0, 
         inputRegisters_274__15, inputRegisters_274__14, inputRegisters_274__13, 
         inputRegisters_274__12, inputRegisters_274__11, inputRegisters_274__10, 
         inputRegisters_274__9, inputRegisters_274__8, inputRegisters_274__7, 
         inputRegisters_274__6, inputRegisters_274__5, inputRegisters_274__4, 
         inputRegisters_274__3, inputRegisters_274__2, inputRegisters_274__1, 
         inputRegisters_274__0, inputRegisters_275__15, inputRegisters_275__14, 
         inputRegisters_275__13, inputRegisters_275__12, inputRegisters_275__11, 
         inputRegisters_275__10, inputRegisters_275__9, inputRegisters_275__8, 
         inputRegisters_275__7, inputRegisters_275__6, inputRegisters_275__5, 
         inputRegisters_275__4, inputRegisters_275__3, inputRegisters_275__2, 
         inputRegisters_275__1, inputRegisters_275__0, inputRegisters_276__15, 
         inputRegisters_276__14, inputRegisters_276__13, inputRegisters_276__12, 
         inputRegisters_276__11, inputRegisters_276__10, inputRegisters_276__9, 
         inputRegisters_276__8, inputRegisters_276__7, inputRegisters_276__6, 
         inputRegisters_276__5, inputRegisters_276__4, inputRegisters_276__3, 
         inputRegisters_276__2, inputRegisters_276__1, inputRegisters_276__0, 
         inputRegisters_277__15, inputRegisters_277__14, inputRegisters_277__13, 
         inputRegisters_277__12, inputRegisters_277__11, inputRegisters_277__10, 
         inputRegisters_277__9, inputRegisters_277__8, inputRegisters_277__7, 
         inputRegisters_277__6, inputRegisters_277__5, inputRegisters_277__4, 
         inputRegisters_277__3, inputRegisters_277__2, inputRegisters_277__1, 
         inputRegisters_277__0, inputRegisters_278__15, inputRegisters_278__14, 
         inputRegisters_278__13, inputRegisters_278__12, inputRegisters_278__11, 
         inputRegisters_278__10, inputRegisters_278__9, inputRegisters_278__8, 
         inputRegisters_278__7, inputRegisters_278__6, inputRegisters_278__5, 
         inputRegisters_278__4, inputRegisters_278__3, inputRegisters_278__2, 
         inputRegisters_278__1, inputRegisters_278__0, inputRegisters_279__15, 
         inputRegisters_279__14, inputRegisters_279__13, inputRegisters_279__12, 
         inputRegisters_279__11, inputRegisters_279__10, inputRegisters_279__9, 
         inputRegisters_279__8, inputRegisters_279__7, inputRegisters_279__6, 
         inputRegisters_279__5, inputRegisters_279__4, inputRegisters_279__3, 
         inputRegisters_279__2, inputRegisters_279__1, inputRegisters_279__0, 
         inputRegisters_280__15, inputRegisters_280__14, inputRegisters_280__13, 
         inputRegisters_280__12, inputRegisters_280__11, inputRegisters_280__10, 
         inputRegisters_280__9, inputRegisters_280__8, inputRegisters_280__7, 
         inputRegisters_280__6, inputRegisters_280__5, inputRegisters_280__4, 
         inputRegisters_280__3, inputRegisters_280__2, inputRegisters_280__1, 
         inputRegisters_280__0, inputRegisters_281__15, inputRegisters_281__14, 
         inputRegisters_281__13, inputRegisters_281__12, inputRegisters_281__11, 
         inputRegisters_281__10, inputRegisters_281__9, inputRegisters_281__8, 
         inputRegisters_281__7, inputRegisters_281__6, inputRegisters_281__5, 
         inputRegisters_281__4, inputRegisters_281__3, inputRegisters_281__2, 
         inputRegisters_281__1, inputRegisters_281__0, inputRegisters_282__15, 
         inputRegisters_282__14, inputRegisters_282__13, inputRegisters_282__12, 
         inputRegisters_282__11, inputRegisters_282__10, inputRegisters_282__9, 
         inputRegisters_282__8, inputRegisters_282__7, inputRegisters_282__6, 
         inputRegisters_282__5, inputRegisters_282__4, inputRegisters_282__3, 
         inputRegisters_282__2, inputRegisters_282__1, inputRegisters_282__0, 
         inputRegisters_283__15, inputRegisters_283__14, inputRegisters_283__13, 
         inputRegisters_283__12, inputRegisters_283__11, inputRegisters_283__10, 
         inputRegisters_283__9, inputRegisters_283__8, inputRegisters_283__7, 
         inputRegisters_283__6, inputRegisters_283__5, inputRegisters_283__4, 
         inputRegisters_283__3, inputRegisters_283__2, inputRegisters_283__1, 
         inputRegisters_283__0, inputRegisters_284__15, inputRegisters_284__14, 
         inputRegisters_284__13, inputRegisters_284__12, inputRegisters_284__11, 
         inputRegisters_284__10, inputRegisters_284__9, inputRegisters_284__8, 
         inputRegisters_284__7, inputRegisters_284__6, inputRegisters_284__5, 
         inputRegisters_284__4, inputRegisters_284__3, inputRegisters_284__2, 
         inputRegisters_284__1, inputRegisters_284__0, inputRegisters_285__15, 
         inputRegisters_285__14, inputRegisters_285__13, inputRegisters_285__12, 
         inputRegisters_285__11, inputRegisters_285__10, inputRegisters_285__9, 
         inputRegisters_285__8, inputRegisters_285__7, inputRegisters_285__6, 
         inputRegisters_285__5, inputRegisters_285__4, inputRegisters_285__3, 
         inputRegisters_285__2, inputRegisters_285__1, inputRegisters_285__0, 
         inputRegisters_286__15, inputRegisters_286__14, inputRegisters_286__13, 
         inputRegisters_286__12, inputRegisters_286__11, inputRegisters_286__10, 
         inputRegisters_286__9, inputRegisters_286__8, inputRegisters_286__7, 
         inputRegisters_286__6, inputRegisters_286__5, inputRegisters_286__4, 
         inputRegisters_286__3, inputRegisters_286__2, inputRegisters_286__1, 
         inputRegisters_286__0, inputRegisters_287__15, inputRegisters_287__14, 
         inputRegisters_287__13, inputRegisters_287__12, inputRegisters_287__11, 
         inputRegisters_287__10, inputRegisters_287__9, inputRegisters_287__8, 
         inputRegisters_287__7, inputRegisters_287__6, inputRegisters_287__5, 
         inputRegisters_287__4, inputRegisters_287__3, inputRegisters_287__2, 
         inputRegisters_287__1, inputRegisters_287__0, inputRegisters_288__15, 
         inputRegisters_288__14, inputRegisters_288__13, inputRegisters_288__12, 
         inputRegisters_288__11, inputRegisters_288__10, inputRegisters_288__9, 
         inputRegisters_288__8, inputRegisters_288__7, inputRegisters_288__6, 
         inputRegisters_288__5, inputRegisters_288__4, inputRegisters_288__3, 
         inputRegisters_288__2, inputRegisters_288__1, inputRegisters_288__0, 
         inputRegisters_289__15, inputRegisters_289__14, inputRegisters_289__13, 
         inputRegisters_289__12, inputRegisters_289__11, inputRegisters_289__10, 
         inputRegisters_289__9, inputRegisters_289__8, inputRegisters_289__7, 
         inputRegisters_289__6, inputRegisters_289__5, inputRegisters_289__4, 
         inputRegisters_289__3, inputRegisters_289__2, inputRegisters_289__1, 
         inputRegisters_289__0, inputRegisters_290__15, inputRegisters_290__14, 
         inputRegisters_290__13, inputRegisters_290__12, inputRegisters_290__11, 
         inputRegisters_290__10, inputRegisters_290__9, inputRegisters_290__8, 
         inputRegisters_290__7, inputRegisters_290__6, inputRegisters_290__5, 
         inputRegisters_290__4, inputRegisters_290__3, inputRegisters_290__2, 
         inputRegisters_290__1, inputRegisters_290__0, inputRegisters_291__15, 
         inputRegisters_291__14, inputRegisters_291__13, inputRegisters_291__12, 
         inputRegisters_291__11, inputRegisters_291__10, inputRegisters_291__9, 
         inputRegisters_291__8, inputRegisters_291__7, inputRegisters_291__6, 
         inputRegisters_291__5, inputRegisters_291__4, inputRegisters_291__3, 
         inputRegisters_291__2, inputRegisters_291__1, inputRegisters_291__0, 
         inputRegisters_292__15, inputRegisters_292__14, inputRegisters_292__13, 
         inputRegisters_292__12, inputRegisters_292__11, inputRegisters_292__10, 
         inputRegisters_292__9, inputRegisters_292__8, inputRegisters_292__7, 
         inputRegisters_292__6, inputRegisters_292__5, inputRegisters_292__4, 
         inputRegisters_292__3, inputRegisters_292__2, inputRegisters_292__1, 
         inputRegisters_292__0, inputRegisters_293__15, inputRegisters_293__14, 
         inputRegisters_293__13, inputRegisters_293__12, inputRegisters_293__11, 
         inputRegisters_293__10, inputRegisters_293__9, inputRegisters_293__8, 
         inputRegisters_293__7, inputRegisters_293__6, inputRegisters_293__5, 
         inputRegisters_293__4, inputRegisters_293__3, inputRegisters_293__2, 
         inputRegisters_293__1, inputRegisters_293__0, inputRegisters_294__15, 
         inputRegisters_294__14, inputRegisters_294__13, inputRegisters_294__12, 
         inputRegisters_294__11, inputRegisters_294__10, inputRegisters_294__9, 
         inputRegisters_294__8, inputRegisters_294__7, inputRegisters_294__6, 
         inputRegisters_294__5, inputRegisters_294__4, inputRegisters_294__3, 
         inputRegisters_294__2, inputRegisters_294__1, inputRegisters_294__0, 
         inputRegisters_295__15, inputRegisters_295__14, inputRegisters_295__13, 
         inputRegisters_295__12, inputRegisters_295__11, inputRegisters_295__10, 
         inputRegisters_295__9, inputRegisters_295__8, inputRegisters_295__7, 
         inputRegisters_295__6, inputRegisters_295__5, inputRegisters_295__4, 
         inputRegisters_295__3, inputRegisters_295__2, inputRegisters_295__1, 
         inputRegisters_295__0, inputRegisters_296__15, inputRegisters_296__14, 
         inputRegisters_296__13, inputRegisters_296__12, inputRegisters_296__11, 
         inputRegisters_296__10, inputRegisters_296__9, inputRegisters_296__8, 
         inputRegisters_296__7, inputRegisters_296__6, inputRegisters_296__5, 
         inputRegisters_296__4, inputRegisters_296__3, inputRegisters_296__2, 
         inputRegisters_296__1, inputRegisters_296__0, inputRegisters_297__15, 
         inputRegisters_297__14, inputRegisters_297__13, inputRegisters_297__12, 
         inputRegisters_297__11, inputRegisters_297__10, inputRegisters_297__9, 
         inputRegisters_297__8, inputRegisters_297__7, inputRegisters_297__6, 
         inputRegisters_297__5, inputRegisters_297__4, inputRegisters_297__3, 
         inputRegisters_297__2, inputRegisters_297__1, inputRegisters_297__0, 
         inputRegisters_298__15, inputRegisters_298__14, inputRegisters_298__13, 
         inputRegisters_298__12, inputRegisters_298__11, inputRegisters_298__10, 
         inputRegisters_298__9, inputRegisters_298__8, inputRegisters_298__7, 
         inputRegisters_298__6, inputRegisters_298__5, inputRegisters_298__4, 
         inputRegisters_298__3, inputRegisters_298__2, inputRegisters_298__1, 
         inputRegisters_298__0, inputRegisters_299__15, inputRegisters_299__14, 
         inputRegisters_299__13, inputRegisters_299__12, inputRegisters_299__11, 
         inputRegisters_299__10, inputRegisters_299__9, inputRegisters_299__8, 
         inputRegisters_299__7, inputRegisters_299__6, inputRegisters_299__5, 
         inputRegisters_299__4, inputRegisters_299__3, inputRegisters_299__2, 
         inputRegisters_299__1, inputRegisters_299__0, inputRegisters_300__15, 
         inputRegisters_300__14, inputRegisters_300__13, inputRegisters_300__12, 
         inputRegisters_300__11, inputRegisters_300__10, inputRegisters_300__9, 
         inputRegisters_300__8, inputRegisters_300__7, inputRegisters_300__6, 
         inputRegisters_300__5, inputRegisters_300__4, inputRegisters_300__3, 
         inputRegisters_300__2, inputRegisters_300__1, inputRegisters_300__0, 
         inputRegisters_301__15, inputRegisters_301__14, inputRegisters_301__13, 
         inputRegisters_301__12, inputRegisters_301__11, inputRegisters_301__10, 
         inputRegisters_301__9, inputRegisters_301__8, inputRegisters_301__7, 
         inputRegisters_301__6, inputRegisters_301__5, inputRegisters_301__4, 
         inputRegisters_301__3, inputRegisters_301__2, inputRegisters_301__1, 
         inputRegisters_301__0, inputRegisters_302__15, inputRegisters_302__14, 
         inputRegisters_302__13, inputRegisters_302__12, inputRegisters_302__11, 
         inputRegisters_302__10, inputRegisters_302__9, inputRegisters_302__8, 
         inputRegisters_302__7, inputRegisters_302__6, inputRegisters_302__5, 
         inputRegisters_302__4, inputRegisters_302__3, inputRegisters_302__2, 
         inputRegisters_302__1, inputRegisters_302__0, inputRegisters_303__15, 
         inputRegisters_303__14, inputRegisters_303__13, inputRegisters_303__12, 
         inputRegisters_303__11, inputRegisters_303__10, inputRegisters_303__9, 
         inputRegisters_303__8, inputRegisters_303__7, inputRegisters_303__6, 
         inputRegisters_303__5, inputRegisters_303__4, inputRegisters_303__3, 
         inputRegisters_303__2, inputRegisters_303__1, inputRegisters_303__0, 
         inputRegisters_304__15, inputRegisters_304__14, inputRegisters_304__13, 
         inputRegisters_304__12, inputRegisters_304__11, inputRegisters_304__10, 
         inputRegisters_304__9, inputRegisters_304__8, inputRegisters_304__7, 
         inputRegisters_304__6, inputRegisters_304__5, inputRegisters_304__4, 
         inputRegisters_304__3, inputRegisters_304__2, inputRegisters_304__1, 
         inputRegisters_304__0, inputRegisters_305__15, inputRegisters_305__14, 
         inputRegisters_305__13, inputRegisters_305__12, inputRegisters_305__11, 
         inputRegisters_305__10, inputRegisters_305__9, inputRegisters_305__8, 
         inputRegisters_305__7, inputRegisters_305__6, inputRegisters_305__5, 
         inputRegisters_305__4, inputRegisters_305__3, inputRegisters_305__2, 
         inputRegisters_305__1, inputRegisters_305__0, inputRegisters_306__15, 
         inputRegisters_306__14, inputRegisters_306__13, inputRegisters_306__12, 
         inputRegisters_306__11, inputRegisters_306__10, inputRegisters_306__9, 
         inputRegisters_306__8, inputRegisters_306__7, inputRegisters_306__6, 
         inputRegisters_306__5, inputRegisters_306__4, inputRegisters_306__3, 
         inputRegisters_306__2, inputRegisters_306__1, inputRegisters_306__0, 
         inputRegisters_307__15, inputRegisters_307__14, inputRegisters_307__13, 
         inputRegisters_307__12, inputRegisters_307__11, inputRegisters_307__10, 
         inputRegisters_307__9, inputRegisters_307__8, inputRegisters_307__7, 
         inputRegisters_307__6, inputRegisters_307__5, inputRegisters_307__4, 
         inputRegisters_307__3, inputRegisters_307__2, inputRegisters_307__1, 
         inputRegisters_307__0, inputRegisters_308__15, inputRegisters_308__14, 
         inputRegisters_308__13, inputRegisters_308__12, inputRegisters_308__11, 
         inputRegisters_308__10, inputRegisters_308__9, inputRegisters_308__8, 
         inputRegisters_308__7, inputRegisters_308__6, inputRegisters_308__5, 
         inputRegisters_308__4, inputRegisters_308__3, inputRegisters_308__2, 
         inputRegisters_308__1, inputRegisters_308__0, inputRegisters_309__15, 
         inputRegisters_309__14, inputRegisters_309__13, inputRegisters_309__12, 
         inputRegisters_309__11, inputRegisters_309__10, inputRegisters_309__9, 
         inputRegisters_309__8, inputRegisters_309__7, inputRegisters_309__6, 
         inputRegisters_309__5, inputRegisters_309__4, inputRegisters_309__3, 
         inputRegisters_309__2, inputRegisters_309__1, inputRegisters_309__0, 
         inputRegisters_310__15, inputRegisters_310__14, inputRegisters_310__13, 
         inputRegisters_310__12, inputRegisters_310__11, inputRegisters_310__10, 
         inputRegisters_310__9, inputRegisters_310__8, inputRegisters_310__7, 
         inputRegisters_310__6, inputRegisters_310__5, inputRegisters_310__4, 
         inputRegisters_310__3, inputRegisters_310__2, inputRegisters_310__1, 
         inputRegisters_310__0, inputRegisters_311__15, inputRegisters_311__14, 
         inputRegisters_311__13, inputRegisters_311__12, inputRegisters_311__11, 
         inputRegisters_311__10, inputRegisters_311__9, inputRegisters_311__8, 
         inputRegisters_311__7, inputRegisters_311__6, inputRegisters_311__5, 
         inputRegisters_311__4, inputRegisters_311__3, inputRegisters_311__2, 
         inputRegisters_311__1, inputRegisters_311__0, inputRegisters_312__15, 
         inputRegisters_312__14, inputRegisters_312__13, inputRegisters_312__12, 
         inputRegisters_312__11, inputRegisters_312__10, inputRegisters_312__9, 
         inputRegisters_312__8, inputRegisters_312__7, inputRegisters_312__6, 
         inputRegisters_312__5, inputRegisters_312__4, inputRegisters_312__3, 
         inputRegisters_312__2, inputRegisters_312__1, inputRegisters_312__0, 
         inputRegisters_313__15, inputRegisters_313__14, inputRegisters_313__13, 
         inputRegisters_313__12, inputRegisters_313__11, inputRegisters_313__10, 
         inputRegisters_313__9, inputRegisters_313__8, inputRegisters_313__7, 
         inputRegisters_313__6, inputRegisters_313__5, inputRegisters_313__4, 
         inputRegisters_313__3, inputRegisters_313__2, inputRegisters_313__1, 
         inputRegisters_313__0, inputRegisters_314__15, inputRegisters_314__14, 
         inputRegisters_314__13, inputRegisters_314__12, inputRegisters_314__11, 
         inputRegisters_314__10, inputRegisters_314__9, inputRegisters_314__8, 
         inputRegisters_314__7, inputRegisters_314__6, inputRegisters_314__5, 
         inputRegisters_314__4, inputRegisters_314__3, inputRegisters_314__2, 
         inputRegisters_314__1, inputRegisters_314__0, inputRegisters_315__15, 
         inputRegisters_315__14, inputRegisters_315__13, inputRegisters_315__12, 
         inputRegisters_315__11, inputRegisters_315__10, inputRegisters_315__9, 
         inputRegisters_315__8, inputRegisters_315__7, inputRegisters_315__6, 
         inputRegisters_315__5, inputRegisters_315__4, inputRegisters_315__3, 
         inputRegisters_315__2, inputRegisters_315__1, inputRegisters_315__0, 
         inputRegisters_316__15, inputRegisters_316__14, inputRegisters_316__13, 
         inputRegisters_316__12, inputRegisters_316__11, inputRegisters_316__10, 
         inputRegisters_316__9, inputRegisters_316__8, inputRegisters_316__7, 
         inputRegisters_316__6, inputRegisters_316__5, inputRegisters_316__4, 
         inputRegisters_316__3, inputRegisters_316__2, inputRegisters_316__1, 
         inputRegisters_316__0, inputRegisters_317__15, inputRegisters_317__14, 
         inputRegisters_317__13, inputRegisters_317__12, inputRegisters_317__11, 
         inputRegisters_317__10, inputRegisters_317__9, inputRegisters_317__8, 
         inputRegisters_317__7, inputRegisters_317__6, inputRegisters_317__5, 
         inputRegisters_317__4, inputRegisters_317__3, inputRegisters_317__2, 
         inputRegisters_317__1, inputRegisters_317__0, inputRegisters_318__15, 
         inputRegisters_318__14, inputRegisters_318__13, inputRegisters_318__12, 
         inputRegisters_318__11, inputRegisters_318__10, inputRegisters_318__9, 
         inputRegisters_318__8, inputRegisters_318__7, inputRegisters_318__6, 
         inputRegisters_318__5, inputRegisters_318__4, inputRegisters_318__3, 
         inputRegisters_318__2, inputRegisters_318__1, inputRegisters_318__0, 
         inputRegisters_319__15, inputRegisters_319__14, inputRegisters_319__13, 
         inputRegisters_319__12, inputRegisters_319__11, inputRegisters_319__10, 
         inputRegisters_319__9, inputRegisters_319__8, inputRegisters_319__7, 
         inputRegisters_319__6, inputRegisters_319__5, inputRegisters_319__4, 
         inputRegisters_319__3, inputRegisters_319__2, inputRegisters_319__1, 
         inputRegisters_319__0, inputRegisters_320__15, inputRegisters_320__14, 
         inputRegisters_320__13, inputRegisters_320__12, inputRegisters_320__11, 
         inputRegisters_320__10, inputRegisters_320__9, inputRegisters_320__8, 
         inputRegisters_320__7, inputRegisters_320__6, inputRegisters_320__5, 
         inputRegisters_320__4, inputRegisters_320__3, inputRegisters_320__2, 
         inputRegisters_320__1, inputRegisters_320__0, inputRegisters_321__15, 
         inputRegisters_321__14, inputRegisters_321__13, inputRegisters_321__12, 
         inputRegisters_321__11, inputRegisters_321__10, inputRegisters_321__9, 
         inputRegisters_321__8, inputRegisters_321__7, inputRegisters_321__6, 
         inputRegisters_321__5, inputRegisters_321__4, inputRegisters_321__3, 
         inputRegisters_321__2, inputRegisters_321__1, inputRegisters_321__0, 
         inputRegisters_322__15, inputRegisters_322__14, inputRegisters_322__13, 
         inputRegisters_322__12, inputRegisters_322__11, inputRegisters_322__10, 
         inputRegisters_322__9, inputRegisters_322__8, inputRegisters_322__7, 
         inputRegisters_322__6, inputRegisters_322__5, inputRegisters_322__4, 
         inputRegisters_322__3, inputRegisters_322__2, inputRegisters_322__1, 
         inputRegisters_322__0, inputRegisters_323__15, inputRegisters_323__14, 
         inputRegisters_323__13, inputRegisters_323__12, inputRegisters_323__11, 
         inputRegisters_323__10, inputRegisters_323__9, inputRegisters_323__8, 
         inputRegisters_323__7, inputRegisters_323__6, inputRegisters_323__5, 
         inputRegisters_323__4, inputRegisters_323__3, inputRegisters_323__2, 
         inputRegisters_323__1, inputRegisters_323__0, inputRegisters_324__15, 
         inputRegisters_324__14, inputRegisters_324__13, inputRegisters_324__12, 
         inputRegisters_324__11, inputRegisters_324__10, inputRegisters_324__9, 
         inputRegisters_324__8, inputRegisters_324__7, inputRegisters_324__6, 
         inputRegisters_324__5, inputRegisters_324__4, inputRegisters_324__3, 
         inputRegisters_324__2, inputRegisters_324__1, inputRegisters_324__0, 
         inputRegisters_325__15, inputRegisters_325__14, inputRegisters_325__13, 
         inputRegisters_325__12, inputRegisters_325__11, inputRegisters_325__10, 
         inputRegisters_325__9, inputRegisters_325__8, inputRegisters_325__7, 
         inputRegisters_325__6, inputRegisters_325__5, inputRegisters_325__4, 
         inputRegisters_325__3, inputRegisters_325__2, inputRegisters_325__1, 
         inputRegisters_325__0, inputRegisters_326__15, inputRegisters_326__14, 
         inputRegisters_326__13, inputRegisters_326__12, inputRegisters_326__11, 
         inputRegisters_326__10, inputRegisters_326__9, inputRegisters_326__8, 
         inputRegisters_326__7, inputRegisters_326__6, inputRegisters_326__5, 
         inputRegisters_326__4, inputRegisters_326__3, inputRegisters_326__2, 
         inputRegisters_326__1, inputRegisters_326__0, inputRegisters_327__15, 
         inputRegisters_327__14, inputRegisters_327__13, inputRegisters_327__12, 
         inputRegisters_327__11, inputRegisters_327__10, inputRegisters_327__9, 
         inputRegisters_327__8, inputRegisters_327__7, inputRegisters_327__6, 
         inputRegisters_327__5, inputRegisters_327__4, inputRegisters_327__3, 
         inputRegisters_327__2, inputRegisters_327__1, inputRegisters_327__0, 
         inputRegisters_328__15, inputRegisters_328__14, inputRegisters_328__13, 
         inputRegisters_328__12, inputRegisters_328__11, inputRegisters_328__10, 
         inputRegisters_328__9, inputRegisters_328__8, inputRegisters_328__7, 
         inputRegisters_328__6, inputRegisters_328__5, inputRegisters_328__4, 
         inputRegisters_328__3, inputRegisters_328__2, inputRegisters_328__1, 
         inputRegisters_328__0, inputRegisters_329__15, inputRegisters_329__14, 
         inputRegisters_329__13, inputRegisters_329__12, inputRegisters_329__11, 
         inputRegisters_329__10, inputRegisters_329__9, inputRegisters_329__8, 
         inputRegisters_329__7, inputRegisters_329__6, inputRegisters_329__5, 
         inputRegisters_329__4, inputRegisters_329__3, inputRegisters_329__2, 
         inputRegisters_329__1, inputRegisters_329__0, inputRegisters_330__15, 
         inputRegisters_330__14, inputRegisters_330__13, inputRegisters_330__12, 
         inputRegisters_330__11, inputRegisters_330__10, inputRegisters_330__9, 
         inputRegisters_330__8, inputRegisters_330__7, inputRegisters_330__6, 
         inputRegisters_330__5, inputRegisters_330__4, inputRegisters_330__3, 
         inputRegisters_330__2, inputRegisters_330__1, inputRegisters_330__0, 
         inputRegisters_331__15, inputRegisters_331__14, inputRegisters_331__13, 
         inputRegisters_331__12, inputRegisters_331__11, inputRegisters_331__10, 
         inputRegisters_331__9, inputRegisters_331__8, inputRegisters_331__7, 
         inputRegisters_331__6, inputRegisters_331__5, inputRegisters_331__4, 
         inputRegisters_331__3, inputRegisters_331__2, inputRegisters_331__1, 
         inputRegisters_331__0, inputRegisters_332__15, inputRegisters_332__14, 
         inputRegisters_332__13, inputRegisters_332__12, inputRegisters_332__11, 
         inputRegisters_332__10, inputRegisters_332__9, inputRegisters_332__8, 
         inputRegisters_332__7, inputRegisters_332__6, inputRegisters_332__5, 
         inputRegisters_332__4, inputRegisters_332__3, inputRegisters_332__2, 
         inputRegisters_332__1, inputRegisters_332__0, inputRegisters_333__15, 
         inputRegisters_333__14, inputRegisters_333__13, inputRegisters_333__12, 
         inputRegisters_333__11, inputRegisters_333__10, inputRegisters_333__9, 
         inputRegisters_333__8, inputRegisters_333__7, inputRegisters_333__6, 
         inputRegisters_333__5, inputRegisters_333__4, inputRegisters_333__3, 
         inputRegisters_333__2, inputRegisters_333__1, inputRegisters_333__0, 
         inputRegisters_334__15, inputRegisters_334__14, inputRegisters_334__13, 
         inputRegisters_334__12, inputRegisters_334__11, inputRegisters_334__10, 
         inputRegisters_334__9, inputRegisters_334__8, inputRegisters_334__7, 
         inputRegisters_334__6, inputRegisters_334__5, inputRegisters_334__4, 
         inputRegisters_334__3, inputRegisters_334__2, inputRegisters_334__1, 
         inputRegisters_334__0, inputRegisters_335__15, inputRegisters_335__14, 
         inputRegisters_335__13, inputRegisters_335__12, inputRegisters_335__11, 
         inputRegisters_335__10, inputRegisters_335__9, inputRegisters_335__8, 
         inputRegisters_335__7, inputRegisters_335__6, inputRegisters_335__5, 
         inputRegisters_335__4, inputRegisters_335__3, inputRegisters_335__2, 
         inputRegisters_335__1, inputRegisters_335__0, inputRegisters_336__15, 
         inputRegisters_336__14, inputRegisters_336__13, inputRegisters_336__12, 
         inputRegisters_336__11, inputRegisters_336__10, inputRegisters_336__9, 
         inputRegisters_336__8, inputRegisters_336__7, inputRegisters_336__6, 
         inputRegisters_336__5, inputRegisters_336__4, inputRegisters_336__3, 
         inputRegisters_336__2, inputRegisters_336__1, inputRegisters_336__0, 
         inputRegisters_337__15, inputRegisters_337__14, inputRegisters_337__13, 
         inputRegisters_337__12, inputRegisters_337__11, inputRegisters_337__10, 
         inputRegisters_337__9, inputRegisters_337__8, inputRegisters_337__7, 
         inputRegisters_337__6, inputRegisters_337__5, inputRegisters_337__4, 
         inputRegisters_337__3, inputRegisters_337__2, inputRegisters_337__1, 
         inputRegisters_337__0, inputRegisters_338__15, inputRegisters_338__14, 
         inputRegisters_338__13, inputRegisters_338__12, inputRegisters_338__11, 
         inputRegisters_338__10, inputRegisters_338__9, inputRegisters_338__8, 
         inputRegisters_338__7, inputRegisters_338__6, inputRegisters_338__5, 
         inputRegisters_338__4, inputRegisters_338__3, inputRegisters_338__2, 
         inputRegisters_338__1, inputRegisters_338__0, inputRegisters_339__15, 
         inputRegisters_339__14, inputRegisters_339__13, inputRegisters_339__12, 
         inputRegisters_339__11, inputRegisters_339__10, inputRegisters_339__9, 
         inputRegisters_339__8, inputRegisters_339__7, inputRegisters_339__6, 
         inputRegisters_339__5, inputRegisters_339__4, inputRegisters_339__3, 
         inputRegisters_339__2, inputRegisters_339__1, inputRegisters_339__0, 
         inputRegisters_340__15, inputRegisters_340__14, inputRegisters_340__13, 
         inputRegisters_340__12, inputRegisters_340__11, inputRegisters_340__10, 
         inputRegisters_340__9, inputRegisters_340__8, inputRegisters_340__7, 
         inputRegisters_340__6, inputRegisters_340__5, inputRegisters_340__4, 
         inputRegisters_340__3, inputRegisters_340__2, inputRegisters_340__1, 
         inputRegisters_340__0, inputRegisters_341__15, inputRegisters_341__14, 
         inputRegisters_341__13, inputRegisters_341__12, inputRegisters_341__11, 
         inputRegisters_341__10, inputRegisters_341__9, inputRegisters_341__8, 
         inputRegisters_341__7, inputRegisters_341__6, inputRegisters_341__5, 
         inputRegisters_341__4, inputRegisters_341__3, inputRegisters_341__2, 
         inputRegisters_341__1, inputRegisters_341__0, inputRegisters_342__15, 
         inputRegisters_342__14, inputRegisters_342__13, inputRegisters_342__12, 
         inputRegisters_342__11, inputRegisters_342__10, inputRegisters_342__9, 
         inputRegisters_342__8, inputRegisters_342__7, inputRegisters_342__6, 
         inputRegisters_342__5, inputRegisters_342__4, inputRegisters_342__3, 
         inputRegisters_342__2, inputRegisters_342__1, inputRegisters_342__0, 
         inputRegisters_343__15, inputRegisters_343__14, inputRegisters_343__13, 
         inputRegisters_343__12, inputRegisters_343__11, inputRegisters_343__10, 
         inputRegisters_343__9, inputRegisters_343__8, inputRegisters_343__7, 
         inputRegisters_343__6, inputRegisters_343__5, inputRegisters_343__4, 
         inputRegisters_343__3, inputRegisters_343__2, inputRegisters_343__1, 
         inputRegisters_343__0, inputRegisters_344__15, inputRegisters_344__14, 
         inputRegisters_344__13, inputRegisters_344__12, inputRegisters_344__11, 
         inputRegisters_344__10, inputRegisters_344__9, inputRegisters_344__8, 
         inputRegisters_344__7, inputRegisters_344__6, inputRegisters_344__5, 
         inputRegisters_344__4, inputRegisters_344__3, inputRegisters_344__2, 
         inputRegisters_344__1, inputRegisters_344__0, inputRegisters_345__15, 
         inputRegisters_345__14, inputRegisters_345__13, inputRegisters_345__12, 
         inputRegisters_345__11, inputRegisters_345__10, inputRegisters_345__9, 
         inputRegisters_345__8, inputRegisters_345__7, inputRegisters_345__6, 
         inputRegisters_345__5, inputRegisters_345__4, inputRegisters_345__3, 
         inputRegisters_345__2, inputRegisters_345__1, inputRegisters_345__0, 
         inputRegisters_346__15, inputRegisters_346__14, inputRegisters_346__13, 
         inputRegisters_346__12, inputRegisters_346__11, inputRegisters_346__10, 
         inputRegisters_346__9, inputRegisters_346__8, inputRegisters_346__7, 
         inputRegisters_346__6, inputRegisters_346__5, inputRegisters_346__4, 
         inputRegisters_346__3, inputRegisters_346__2, inputRegisters_346__1, 
         inputRegisters_346__0, inputRegisters_347__15, inputRegisters_347__14, 
         inputRegisters_347__13, inputRegisters_347__12, inputRegisters_347__11, 
         inputRegisters_347__10, inputRegisters_347__9, inputRegisters_347__8, 
         inputRegisters_347__7, inputRegisters_347__6, inputRegisters_347__5, 
         inputRegisters_347__4, inputRegisters_347__3, inputRegisters_347__2, 
         inputRegisters_347__1, inputRegisters_347__0, inputRegisters_348__15, 
         inputRegisters_348__14, inputRegisters_348__13, inputRegisters_348__12, 
         inputRegisters_348__11, inputRegisters_348__10, inputRegisters_348__9, 
         inputRegisters_348__8, inputRegisters_348__7, inputRegisters_348__6, 
         inputRegisters_348__5, inputRegisters_348__4, inputRegisters_348__3, 
         inputRegisters_348__2, inputRegisters_348__1, inputRegisters_348__0, 
         inputRegisters_349__15, inputRegisters_349__14, inputRegisters_349__13, 
         inputRegisters_349__12, inputRegisters_349__11, inputRegisters_349__10, 
         inputRegisters_349__9, inputRegisters_349__8, inputRegisters_349__7, 
         inputRegisters_349__6, inputRegisters_349__5, inputRegisters_349__4, 
         inputRegisters_349__3, inputRegisters_349__2, inputRegisters_349__1, 
         inputRegisters_349__0, inputRegisters_350__15, inputRegisters_350__14, 
         inputRegisters_350__13, inputRegisters_350__12, inputRegisters_350__11, 
         inputRegisters_350__10, inputRegisters_350__9, inputRegisters_350__8, 
         inputRegisters_350__7, inputRegisters_350__6, inputRegisters_350__5, 
         inputRegisters_350__4, inputRegisters_350__3, inputRegisters_350__2, 
         inputRegisters_350__1, inputRegisters_350__0, inputRegisters_351__15, 
         inputRegisters_351__14, inputRegisters_351__13, inputRegisters_351__12, 
         inputRegisters_351__11, inputRegisters_351__10, inputRegisters_351__9, 
         inputRegisters_351__8, inputRegisters_351__7, inputRegisters_351__6, 
         inputRegisters_351__5, inputRegisters_351__4, inputRegisters_351__3, 
         inputRegisters_351__2, inputRegisters_351__1, inputRegisters_351__0, 
         inputRegisters_352__15, inputRegisters_352__14, inputRegisters_352__13, 
         inputRegisters_352__12, inputRegisters_352__11, inputRegisters_352__10, 
         inputRegisters_352__9, inputRegisters_352__8, inputRegisters_352__7, 
         inputRegisters_352__6, inputRegisters_352__5, inputRegisters_352__4, 
         inputRegisters_352__3, inputRegisters_352__2, inputRegisters_352__1, 
         inputRegisters_352__0, inputRegisters_353__15, inputRegisters_353__14, 
         inputRegisters_353__13, inputRegisters_353__12, inputRegisters_353__11, 
         inputRegisters_353__10, inputRegisters_353__9, inputRegisters_353__8, 
         inputRegisters_353__7, inputRegisters_353__6, inputRegisters_353__5, 
         inputRegisters_353__4, inputRegisters_353__3, inputRegisters_353__2, 
         inputRegisters_353__1, inputRegisters_353__0, inputRegisters_354__15, 
         inputRegisters_354__14, inputRegisters_354__13, inputRegisters_354__12, 
         inputRegisters_354__11, inputRegisters_354__10, inputRegisters_354__9, 
         inputRegisters_354__8, inputRegisters_354__7, inputRegisters_354__6, 
         inputRegisters_354__5, inputRegisters_354__4, inputRegisters_354__3, 
         inputRegisters_354__2, inputRegisters_354__1, inputRegisters_354__0, 
         inputRegisters_355__15, inputRegisters_355__14, inputRegisters_355__13, 
         inputRegisters_355__12, inputRegisters_355__11, inputRegisters_355__10, 
         inputRegisters_355__9, inputRegisters_355__8, inputRegisters_355__7, 
         inputRegisters_355__6, inputRegisters_355__5, inputRegisters_355__4, 
         inputRegisters_355__3, inputRegisters_355__2, inputRegisters_355__1, 
         inputRegisters_355__0, inputRegisters_356__15, inputRegisters_356__14, 
         inputRegisters_356__13, inputRegisters_356__12, inputRegisters_356__11, 
         inputRegisters_356__10, inputRegisters_356__9, inputRegisters_356__8, 
         inputRegisters_356__7, inputRegisters_356__6, inputRegisters_356__5, 
         inputRegisters_356__4, inputRegisters_356__3, inputRegisters_356__2, 
         inputRegisters_356__1, inputRegisters_356__0, inputRegisters_357__15, 
         inputRegisters_357__14, inputRegisters_357__13, inputRegisters_357__12, 
         inputRegisters_357__11, inputRegisters_357__10, inputRegisters_357__9, 
         inputRegisters_357__8, inputRegisters_357__7, inputRegisters_357__6, 
         inputRegisters_357__5, inputRegisters_357__4, inputRegisters_357__3, 
         inputRegisters_357__2, inputRegisters_357__1, inputRegisters_357__0, 
         inputRegisters_358__15, inputRegisters_358__14, inputRegisters_358__13, 
         inputRegisters_358__12, inputRegisters_358__11, inputRegisters_358__10, 
         inputRegisters_358__9, inputRegisters_358__8, inputRegisters_358__7, 
         inputRegisters_358__6, inputRegisters_358__5, inputRegisters_358__4, 
         inputRegisters_358__3, inputRegisters_358__2, inputRegisters_358__1, 
         inputRegisters_358__0, inputRegisters_359__15, inputRegisters_359__14, 
         inputRegisters_359__13, inputRegisters_359__12, inputRegisters_359__11, 
         inputRegisters_359__10, inputRegisters_359__9, inputRegisters_359__8, 
         inputRegisters_359__7, inputRegisters_359__6, inputRegisters_359__5, 
         inputRegisters_359__4, inputRegisters_359__3, inputRegisters_359__2, 
         inputRegisters_359__1, inputRegisters_359__0, inputRegisters_360__15, 
         inputRegisters_360__14, inputRegisters_360__13, inputRegisters_360__12, 
         inputRegisters_360__11, inputRegisters_360__10, inputRegisters_360__9, 
         inputRegisters_360__8, inputRegisters_360__7, inputRegisters_360__6, 
         inputRegisters_360__5, inputRegisters_360__4, inputRegisters_360__3, 
         inputRegisters_360__2, inputRegisters_360__1, inputRegisters_360__0, 
         inputRegisters_361__15, inputRegisters_361__14, inputRegisters_361__13, 
         inputRegisters_361__12, inputRegisters_361__11, inputRegisters_361__10, 
         inputRegisters_361__9, inputRegisters_361__8, inputRegisters_361__7, 
         inputRegisters_361__6, inputRegisters_361__5, inputRegisters_361__4, 
         inputRegisters_361__3, inputRegisters_361__2, inputRegisters_361__1, 
         inputRegisters_361__0, inputRegisters_362__15, inputRegisters_362__14, 
         inputRegisters_362__13, inputRegisters_362__12, inputRegisters_362__11, 
         inputRegisters_362__10, inputRegisters_362__9, inputRegisters_362__8, 
         inputRegisters_362__7, inputRegisters_362__6, inputRegisters_362__5, 
         inputRegisters_362__4, inputRegisters_362__3, inputRegisters_362__2, 
         inputRegisters_362__1, inputRegisters_362__0, inputRegisters_363__15, 
         inputRegisters_363__14, inputRegisters_363__13, inputRegisters_363__12, 
         inputRegisters_363__11, inputRegisters_363__10, inputRegisters_363__9, 
         inputRegisters_363__8, inputRegisters_363__7, inputRegisters_363__6, 
         inputRegisters_363__5, inputRegisters_363__4, inputRegisters_363__3, 
         inputRegisters_363__2, inputRegisters_363__1, inputRegisters_363__0, 
         inputRegisters_364__15, inputRegisters_364__14, inputRegisters_364__13, 
         inputRegisters_364__12, inputRegisters_364__11, inputRegisters_364__10, 
         inputRegisters_364__9, inputRegisters_364__8, inputRegisters_364__7, 
         inputRegisters_364__6, inputRegisters_364__5, inputRegisters_364__4, 
         inputRegisters_364__3, inputRegisters_364__2, inputRegisters_364__1, 
         inputRegisters_364__0, inputRegisters_365__15, inputRegisters_365__14, 
         inputRegisters_365__13, inputRegisters_365__12, inputRegisters_365__11, 
         inputRegisters_365__10, inputRegisters_365__9, inputRegisters_365__8, 
         inputRegisters_365__7, inputRegisters_365__6, inputRegisters_365__5, 
         inputRegisters_365__4, inputRegisters_365__3, inputRegisters_365__2, 
         inputRegisters_365__1, inputRegisters_365__0, inputRegisters_366__15, 
         inputRegisters_366__14, inputRegisters_366__13, inputRegisters_366__12, 
         inputRegisters_366__11, inputRegisters_366__10, inputRegisters_366__9, 
         inputRegisters_366__8, inputRegisters_366__7, inputRegisters_366__6, 
         inputRegisters_366__5, inputRegisters_366__4, inputRegisters_366__3, 
         inputRegisters_366__2, inputRegisters_366__1, inputRegisters_366__0, 
         inputRegisters_367__15, inputRegisters_367__14, inputRegisters_367__13, 
         inputRegisters_367__12, inputRegisters_367__11, inputRegisters_367__10, 
         inputRegisters_367__9, inputRegisters_367__8, inputRegisters_367__7, 
         inputRegisters_367__6, inputRegisters_367__5, inputRegisters_367__4, 
         inputRegisters_367__3, inputRegisters_367__2, inputRegisters_367__1, 
         inputRegisters_367__0, inputRegisters_368__15, inputRegisters_368__14, 
         inputRegisters_368__13, inputRegisters_368__12, inputRegisters_368__11, 
         inputRegisters_368__10, inputRegisters_368__9, inputRegisters_368__8, 
         inputRegisters_368__7, inputRegisters_368__6, inputRegisters_368__5, 
         inputRegisters_368__4, inputRegisters_368__3, inputRegisters_368__2, 
         inputRegisters_368__1, inputRegisters_368__0, inputRegisters_369__15, 
         inputRegisters_369__14, inputRegisters_369__13, inputRegisters_369__12, 
         inputRegisters_369__11, inputRegisters_369__10, inputRegisters_369__9, 
         inputRegisters_369__8, inputRegisters_369__7, inputRegisters_369__6, 
         inputRegisters_369__5, inputRegisters_369__4, inputRegisters_369__3, 
         inputRegisters_369__2, inputRegisters_369__1, inputRegisters_369__0, 
         inputRegisters_370__15, inputRegisters_370__14, inputRegisters_370__13, 
         inputRegisters_370__12, inputRegisters_370__11, inputRegisters_370__10, 
         inputRegisters_370__9, inputRegisters_370__8, inputRegisters_370__7, 
         inputRegisters_370__6, inputRegisters_370__5, inputRegisters_370__4, 
         inputRegisters_370__3, inputRegisters_370__2, inputRegisters_370__1, 
         inputRegisters_370__0, inputRegisters_371__15, inputRegisters_371__14, 
         inputRegisters_371__13, inputRegisters_371__12, inputRegisters_371__11, 
         inputRegisters_371__10, inputRegisters_371__9, inputRegisters_371__8, 
         inputRegisters_371__7, inputRegisters_371__6, inputRegisters_371__5, 
         inputRegisters_371__4, inputRegisters_371__3, inputRegisters_371__2, 
         inputRegisters_371__1, inputRegisters_371__0, inputRegisters_372__15, 
         inputRegisters_372__14, inputRegisters_372__13, inputRegisters_372__12, 
         inputRegisters_372__11, inputRegisters_372__10, inputRegisters_372__9, 
         inputRegisters_372__8, inputRegisters_372__7, inputRegisters_372__6, 
         inputRegisters_372__5, inputRegisters_372__4, inputRegisters_372__3, 
         inputRegisters_372__2, inputRegisters_372__1, inputRegisters_372__0, 
         inputRegisters_373__15, inputRegisters_373__14, inputRegisters_373__13, 
         inputRegisters_373__12, inputRegisters_373__11, inputRegisters_373__10, 
         inputRegisters_373__9, inputRegisters_373__8, inputRegisters_373__7, 
         inputRegisters_373__6, inputRegisters_373__5, inputRegisters_373__4, 
         inputRegisters_373__3, inputRegisters_373__2, inputRegisters_373__1, 
         inputRegisters_373__0, inputRegisters_374__15, inputRegisters_374__14, 
         inputRegisters_374__13, inputRegisters_374__12, inputRegisters_374__11, 
         inputRegisters_374__10, inputRegisters_374__9, inputRegisters_374__8, 
         inputRegisters_374__7, inputRegisters_374__6, inputRegisters_374__5, 
         inputRegisters_374__4, inputRegisters_374__3, inputRegisters_374__2, 
         inputRegisters_374__1, inputRegisters_374__0, inputRegisters_375__15, 
         inputRegisters_375__14, inputRegisters_375__13, inputRegisters_375__12, 
         inputRegisters_375__11, inputRegisters_375__10, inputRegisters_375__9, 
         inputRegisters_375__8, inputRegisters_375__7, inputRegisters_375__6, 
         inputRegisters_375__5, inputRegisters_375__4, inputRegisters_375__3, 
         inputRegisters_375__2, inputRegisters_375__1, inputRegisters_375__0, 
         inputRegisters_376__15, inputRegisters_376__14, inputRegisters_376__13, 
         inputRegisters_376__12, inputRegisters_376__11, inputRegisters_376__10, 
         inputRegisters_376__9, inputRegisters_376__8, inputRegisters_376__7, 
         inputRegisters_376__6, inputRegisters_376__5, inputRegisters_376__4, 
         inputRegisters_376__3, inputRegisters_376__2, inputRegisters_376__1, 
         inputRegisters_376__0, inputRegisters_377__15, inputRegisters_377__14, 
         inputRegisters_377__13, inputRegisters_377__12, inputRegisters_377__11, 
         inputRegisters_377__10, inputRegisters_377__9, inputRegisters_377__8, 
         inputRegisters_377__7, inputRegisters_377__6, inputRegisters_377__5, 
         inputRegisters_377__4, inputRegisters_377__3, inputRegisters_377__2, 
         inputRegisters_377__1, inputRegisters_377__0, inputRegisters_378__15, 
         inputRegisters_378__14, inputRegisters_378__13, inputRegisters_378__12, 
         inputRegisters_378__11, inputRegisters_378__10, inputRegisters_378__9, 
         inputRegisters_378__8, inputRegisters_378__7, inputRegisters_378__6, 
         inputRegisters_378__5, inputRegisters_378__4, inputRegisters_378__3, 
         inputRegisters_378__2, inputRegisters_378__1, inputRegisters_378__0, 
         inputRegisters_379__15, inputRegisters_379__14, inputRegisters_379__13, 
         inputRegisters_379__12, inputRegisters_379__11, inputRegisters_379__10, 
         inputRegisters_379__9, inputRegisters_379__8, inputRegisters_379__7, 
         inputRegisters_379__6, inputRegisters_379__5, inputRegisters_379__4, 
         inputRegisters_379__3, inputRegisters_379__2, inputRegisters_379__1, 
         inputRegisters_379__0, inputRegisters_380__15, inputRegisters_380__14, 
         inputRegisters_380__13, inputRegisters_380__12, inputRegisters_380__11, 
         inputRegisters_380__10, inputRegisters_380__9, inputRegisters_380__8, 
         inputRegisters_380__7, inputRegisters_380__6, inputRegisters_380__5, 
         inputRegisters_380__4, inputRegisters_380__3, inputRegisters_380__2, 
         inputRegisters_380__1, inputRegisters_380__0, inputRegisters_381__15, 
         inputRegisters_381__14, inputRegisters_381__13, inputRegisters_381__12, 
         inputRegisters_381__11, inputRegisters_381__10, inputRegisters_381__9, 
         inputRegisters_381__8, inputRegisters_381__7, inputRegisters_381__6, 
         inputRegisters_381__5, inputRegisters_381__4, inputRegisters_381__3, 
         inputRegisters_381__2, inputRegisters_381__1, inputRegisters_381__0, 
         inputRegisters_382__15, inputRegisters_382__14, inputRegisters_382__13, 
         inputRegisters_382__12, inputRegisters_382__11, inputRegisters_382__10, 
         inputRegisters_382__9, inputRegisters_382__8, inputRegisters_382__7, 
         inputRegisters_382__6, inputRegisters_382__5, inputRegisters_382__4, 
         inputRegisters_382__3, inputRegisters_382__2, inputRegisters_382__1, 
         inputRegisters_382__0, inputRegisters_383__15, inputRegisters_383__14, 
         inputRegisters_383__13, inputRegisters_383__12, inputRegisters_383__11, 
         inputRegisters_383__10, inputRegisters_383__9, inputRegisters_383__8, 
         inputRegisters_383__7, inputRegisters_383__6, inputRegisters_383__5, 
         inputRegisters_383__4, inputRegisters_383__3, inputRegisters_383__2, 
         inputRegisters_383__1, inputRegisters_383__0, inputRegisters_384__15, 
         inputRegisters_384__14, inputRegisters_384__13, inputRegisters_384__12, 
         inputRegisters_384__11, inputRegisters_384__10, inputRegisters_384__9, 
         inputRegisters_384__8, inputRegisters_384__7, inputRegisters_384__6, 
         inputRegisters_384__5, inputRegisters_384__4, inputRegisters_384__3, 
         inputRegisters_384__2, inputRegisters_384__1, inputRegisters_384__0, 
         inputRegisters_385__15, inputRegisters_385__14, inputRegisters_385__13, 
         inputRegisters_385__12, inputRegisters_385__11, inputRegisters_385__10, 
         inputRegisters_385__9, inputRegisters_385__8, inputRegisters_385__7, 
         inputRegisters_385__6, inputRegisters_385__5, inputRegisters_385__4, 
         inputRegisters_385__3, inputRegisters_385__2, inputRegisters_385__1, 
         inputRegisters_385__0, inputRegisters_386__15, inputRegisters_386__14, 
         inputRegisters_386__13, inputRegisters_386__12, inputRegisters_386__11, 
         inputRegisters_386__10, inputRegisters_386__9, inputRegisters_386__8, 
         inputRegisters_386__7, inputRegisters_386__6, inputRegisters_386__5, 
         inputRegisters_386__4, inputRegisters_386__3, inputRegisters_386__2, 
         inputRegisters_386__1, inputRegisters_386__0, inputRegisters_387__15, 
         inputRegisters_387__14, inputRegisters_387__13, inputRegisters_387__12, 
         inputRegisters_387__11, inputRegisters_387__10, inputRegisters_387__9, 
         inputRegisters_387__8, inputRegisters_387__7, inputRegisters_387__6, 
         inputRegisters_387__5, inputRegisters_387__4, inputRegisters_387__3, 
         inputRegisters_387__2, inputRegisters_387__1, inputRegisters_387__0, 
         inputRegisters_388__15, inputRegisters_388__14, inputRegisters_388__13, 
         inputRegisters_388__12, inputRegisters_388__11, inputRegisters_388__10, 
         inputRegisters_388__9, inputRegisters_388__8, inputRegisters_388__7, 
         inputRegisters_388__6, inputRegisters_388__5, inputRegisters_388__4, 
         inputRegisters_388__3, inputRegisters_388__2, inputRegisters_388__1, 
         inputRegisters_388__0, inputRegisters_389__15, inputRegisters_389__14, 
         inputRegisters_389__13, inputRegisters_389__12, inputRegisters_389__11, 
         inputRegisters_389__10, inputRegisters_389__9, inputRegisters_389__8, 
         inputRegisters_389__7, inputRegisters_389__6, inputRegisters_389__5, 
         inputRegisters_389__4, inputRegisters_389__3, inputRegisters_389__2, 
         inputRegisters_389__1, inputRegisters_389__0, inputRegisters_390__15, 
         inputRegisters_390__14, inputRegisters_390__13, inputRegisters_390__12, 
         inputRegisters_390__11, inputRegisters_390__10, inputRegisters_390__9, 
         inputRegisters_390__8, inputRegisters_390__7, inputRegisters_390__6, 
         inputRegisters_390__5, inputRegisters_390__4, inputRegisters_390__3, 
         inputRegisters_390__2, inputRegisters_390__1, inputRegisters_390__0, 
         inputRegisters_391__15, inputRegisters_391__14, inputRegisters_391__13, 
         inputRegisters_391__12, inputRegisters_391__11, inputRegisters_391__10, 
         inputRegisters_391__9, inputRegisters_391__8, inputRegisters_391__7, 
         inputRegisters_391__6, inputRegisters_391__5, inputRegisters_391__4, 
         inputRegisters_391__3, inputRegisters_391__2, inputRegisters_391__1, 
         inputRegisters_391__0, inputRegisters_392__15, inputRegisters_392__14, 
         inputRegisters_392__13, inputRegisters_392__12, inputRegisters_392__11, 
         inputRegisters_392__10, inputRegisters_392__9, inputRegisters_392__8, 
         inputRegisters_392__7, inputRegisters_392__6, inputRegisters_392__5, 
         inputRegisters_392__4, inputRegisters_392__3, inputRegisters_392__2, 
         inputRegisters_392__1, inputRegisters_392__0, inputRegisters_393__15, 
         inputRegisters_393__14, inputRegisters_393__13, inputRegisters_393__12, 
         inputRegisters_393__11, inputRegisters_393__10, inputRegisters_393__9, 
         inputRegisters_393__8, inputRegisters_393__7, inputRegisters_393__6, 
         inputRegisters_393__5, inputRegisters_393__4, inputRegisters_393__3, 
         inputRegisters_393__2, inputRegisters_393__1, inputRegisters_393__0, 
         inputRegisters_394__15, inputRegisters_394__14, inputRegisters_394__13, 
         inputRegisters_394__12, inputRegisters_394__11, inputRegisters_394__10, 
         inputRegisters_394__9, inputRegisters_394__8, inputRegisters_394__7, 
         inputRegisters_394__6, inputRegisters_394__5, inputRegisters_394__4, 
         inputRegisters_394__3, inputRegisters_394__2, inputRegisters_394__1, 
         inputRegisters_394__0, inputRegisters_395__15, inputRegisters_395__14, 
         inputRegisters_395__13, inputRegisters_395__12, inputRegisters_395__11, 
         inputRegisters_395__10, inputRegisters_395__9, inputRegisters_395__8, 
         inputRegisters_395__7, inputRegisters_395__6, inputRegisters_395__5, 
         inputRegisters_395__4, inputRegisters_395__3, inputRegisters_395__2, 
         inputRegisters_395__1, inputRegisters_395__0, inputRegisters_396__15, 
         inputRegisters_396__14, inputRegisters_396__13, inputRegisters_396__12, 
         inputRegisters_396__11, inputRegisters_396__10, inputRegisters_396__9, 
         inputRegisters_396__8, inputRegisters_396__7, inputRegisters_396__6, 
         inputRegisters_396__5, inputRegisters_396__4, inputRegisters_396__3, 
         inputRegisters_396__2, inputRegisters_396__1, inputRegisters_396__0, 
         inputRegisters_397__15, inputRegisters_397__14, inputRegisters_397__13, 
         inputRegisters_397__12, inputRegisters_397__11, inputRegisters_397__10, 
         inputRegisters_397__9, inputRegisters_397__8, inputRegisters_397__7, 
         inputRegisters_397__6, inputRegisters_397__5, inputRegisters_397__4, 
         inputRegisters_397__3, inputRegisters_397__2, inputRegisters_397__1, 
         inputRegisters_397__0, inputRegisters_398__15, inputRegisters_398__14, 
         inputRegisters_398__13, inputRegisters_398__12, inputRegisters_398__11, 
         inputRegisters_398__10, inputRegisters_398__9, inputRegisters_398__8, 
         inputRegisters_398__7, inputRegisters_398__6, inputRegisters_398__5, 
         inputRegisters_398__4, inputRegisters_398__3, inputRegisters_398__2, 
         inputRegisters_398__1, inputRegisters_398__0, inputRegisters_399__15, 
         inputRegisters_399__14, inputRegisters_399__13, inputRegisters_399__12, 
         inputRegisters_399__11, inputRegisters_399__10, inputRegisters_399__9, 
         inputRegisters_399__8, inputRegisters_399__7, inputRegisters_399__6, 
         inputRegisters_399__5, inputRegisters_399__4, inputRegisters_399__3, 
         inputRegisters_399__2, inputRegisters_399__1, inputRegisters_399__0, 
         inputRegisters_400__15, inputRegisters_400__14, inputRegisters_400__13, 
         inputRegisters_400__12, inputRegisters_400__11, inputRegisters_400__10, 
         inputRegisters_400__9, inputRegisters_400__8, inputRegisters_400__7, 
         inputRegisters_400__6, inputRegisters_400__5, inputRegisters_400__4, 
         inputRegisters_400__3, inputRegisters_400__2, inputRegisters_400__1, 
         inputRegisters_400__0, inputRegisters_401__15, inputRegisters_401__14, 
         inputRegisters_401__13, inputRegisters_401__12, inputRegisters_401__11, 
         inputRegisters_401__10, inputRegisters_401__9, inputRegisters_401__8, 
         inputRegisters_401__7, inputRegisters_401__6, inputRegisters_401__5, 
         inputRegisters_401__4, inputRegisters_401__3, inputRegisters_401__2, 
         inputRegisters_401__1, inputRegisters_401__0, inputRegisters_402__15, 
         inputRegisters_402__14, inputRegisters_402__13, inputRegisters_402__12, 
         inputRegisters_402__11, inputRegisters_402__10, inputRegisters_402__9, 
         inputRegisters_402__8, inputRegisters_402__7, inputRegisters_402__6, 
         inputRegisters_402__5, inputRegisters_402__4, inputRegisters_402__3, 
         inputRegisters_402__2, inputRegisters_402__1, inputRegisters_402__0, 
         inputRegisters_403__15, inputRegisters_403__14, inputRegisters_403__13, 
         inputRegisters_403__12, inputRegisters_403__11, inputRegisters_403__10, 
         inputRegisters_403__9, inputRegisters_403__8, inputRegisters_403__7, 
         inputRegisters_403__6, inputRegisters_403__5, inputRegisters_403__4, 
         inputRegisters_403__3, inputRegisters_403__2, inputRegisters_403__1, 
         inputRegisters_403__0, inputRegisters_404__15, inputRegisters_404__14, 
         inputRegisters_404__13, inputRegisters_404__12, inputRegisters_404__11, 
         inputRegisters_404__10, inputRegisters_404__9, inputRegisters_404__8, 
         inputRegisters_404__7, inputRegisters_404__6, inputRegisters_404__5, 
         inputRegisters_404__4, inputRegisters_404__3, inputRegisters_404__2, 
         inputRegisters_404__1, inputRegisters_404__0, inputRegisters_405__15, 
         inputRegisters_405__14, inputRegisters_405__13, inputRegisters_405__12, 
         inputRegisters_405__11, inputRegisters_405__10, inputRegisters_405__9, 
         inputRegisters_405__8, inputRegisters_405__7, inputRegisters_405__6, 
         inputRegisters_405__5, inputRegisters_405__4, inputRegisters_405__3, 
         inputRegisters_405__2, inputRegisters_405__1, inputRegisters_405__0, 
         inputRegisters_406__15, inputRegisters_406__14, inputRegisters_406__13, 
         inputRegisters_406__12, inputRegisters_406__11, inputRegisters_406__10, 
         inputRegisters_406__9, inputRegisters_406__8, inputRegisters_406__7, 
         inputRegisters_406__6, inputRegisters_406__5, inputRegisters_406__4, 
         inputRegisters_406__3, inputRegisters_406__2, inputRegisters_406__1, 
         inputRegisters_406__0, inputRegisters_407__15, inputRegisters_407__14, 
         inputRegisters_407__13, inputRegisters_407__12, inputRegisters_407__11, 
         inputRegisters_407__10, inputRegisters_407__9, inputRegisters_407__8, 
         inputRegisters_407__7, inputRegisters_407__6, inputRegisters_407__5, 
         inputRegisters_407__4, inputRegisters_407__3, inputRegisters_407__2, 
         inputRegisters_407__1, inputRegisters_407__0, inputRegisters_408__15, 
         inputRegisters_408__14, inputRegisters_408__13, inputRegisters_408__12, 
         inputRegisters_408__11, inputRegisters_408__10, inputRegisters_408__9, 
         inputRegisters_408__8, inputRegisters_408__7, inputRegisters_408__6, 
         inputRegisters_408__5, inputRegisters_408__4, inputRegisters_408__3, 
         inputRegisters_408__2, inputRegisters_408__1, inputRegisters_408__0, 
         inputRegisters_409__15, inputRegisters_409__14, inputRegisters_409__13, 
         inputRegisters_409__12, inputRegisters_409__11, inputRegisters_409__10, 
         inputRegisters_409__9, inputRegisters_409__8, inputRegisters_409__7, 
         inputRegisters_409__6, inputRegisters_409__5, inputRegisters_409__4, 
         inputRegisters_409__3, inputRegisters_409__2, inputRegisters_409__1, 
         inputRegisters_409__0, inputRegisters_410__15, inputRegisters_410__14, 
         inputRegisters_410__13, inputRegisters_410__12, inputRegisters_410__11, 
         inputRegisters_410__10, inputRegisters_410__9, inputRegisters_410__8, 
         inputRegisters_410__7, inputRegisters_410__6, inputRegisters_410__5, 
         inputRegisters_410__4, inputRegisters_410__3, inputRegisters_410__2, 
         inputRegisters_410__1, inputRegisters_410__0, inputRegisters_411__15, 
         inputRegisters_411__14, inputRegisters_411__13, inputRegisters_411__12, 
         inputRegisters_411__11, inputRegisters_411__10, inputRegisters_411__9, 
         inputRegisters_411__8, inputRegisters_411__7, inputRegisters_411__6, 
         inputRegisters_411__5, inputRegisters_411__4, inputRegisters_411__3, 
         inputRegisters_411__2, inputRegisters_411__1, inputRegisters_411__0, 
         inputRegisters_412__15, inputRegisters_412__14, inputRegisters_412__13, 
         inputRegisters_412__12, inputRegisters_412__11, inputRegisters_412__10, 
         inputRegisters_412__9, inputRegisters_412__8, inputRegisters_412__7, 
         inputRegisters_412__6, inputRegisters_412__5, inputRegisters_412__4, 
         inputRegisters_412__3, inputRegisters_412__2, inputRegisters_412__1, 
         inputRegisters_412__0, inputRegisters_413__15, inputRegisters_413__14, 
         inputRegisters_413__13, inputRegisters_413__12, inputRegisters_413__11, 
         inputRegisters_413__10, inputRegisters_413__9, inputRegisters_413__8, 
         inputRegisters_413__7, inputRegisters_413__6, inputRegisters_413__5, 
         inputRegisters_413__4, inputRegisters_413__3, inputRegisters_413__2, 
         inputRegisters_413__1, inputRegisters_413__0, inputRegisters_414__15, 
         inputRegisters_414__14, inputRegisters_414__13, inputRegisters_414__12, 
         inputRegisters_414__11, inputRegisters_414__10, inputRegisters_414__9, 
         inputRegisters_414__8, inputRegisters_414__7, inputRegisters_414__6, 
         inputRegisters_414__5, inputRegisters_414__4, inputRegisters_414__3, 
         inputRegisters_414__2, inputRegisters_414__1, inputRegisters_414__0, 
         inputRegisters_415__15, inputRegisters_415__14, inputRegisters_415__13, 
         inputRegisters_415__12, inputRegisters_415__11, inputRegisters_415__10, 
         inputRegisters_415__9, inputRegisters_415__8, inputRegisters_415__7, 
         inputRegisters_415__6, inputRegisters_415__5, inputRegisters_415__4, 
         inputRegisters_415__3, inputRegisters_415__2, inputRegisters_415__1, 
         inputRegisters_415__0, inputRegisters_416__15, inputRegisters_416__14, 
         inputRegisters_416__13, inputRegisters_416__12, inputRegisters_416__11, 
         inputRegisters_416__10, inputRegisters_416__9, inputRegisters_416__8, 
         inputRegisters_416__7, inputRegisters_416__6, inputRegisters_416__5, 
         inputRegisters_416__4, inputRegisters_416__3, inputRegisters_416__2, 
         inputRegisters_416__1, inputRegisters_416__0, inputRegisters_417__15, 
         inputRegisters_417__14, inputRegisters_417__13, inputRegisters_417__12, 
         inputRegisters_417__11, inputRegisters_417__10, inputRegisters_417__9, 
         inputRegisters_417__8, inputRegisters_417__7, inputRegisters_417__6, 
         inputRegisters_417__5, inputRegisters_417__4, inputRegisters_417__3, 
         inputRegisters_417__2, inputRegisters_417__1, inputRegisters_417__0, 
         inputRegisters_418__15, inputRegisters_418__14, inputRegisters_418__13, 
         inputRegisters_418__12, inputRegisters_418__11, inputRegisters_418__10, 
         inputRegisters_418__9, inputRegisters_418__8, inputRegisters_418__7, 
         inputRegisters_418__6, inputRegisters_418__5, inputRegisters_418__4, 
         inputRegisters_418__3, inputRegisters_418__2, inputRegisters_418__1, 
         inputRegisters_418__0, inputRegisters_419__15, inputRegisters_419__14, 
         inputRegisters_419__13, inputRegisters_419__12, inputRegisters_419__11, 
         inputRegisters_419__10, inputRegisters_419__9, inputRegisters_419__8, 
         inputRegisters_419__7, inputRegisters_419__6, inputRegisters_419__5, 
         inputRegisters_419__4, inputRegisters_419__3, inputRegisters_419__2, 
         inputRegisters_419__1, inputRegisters_419__0, inputRegisters_420__15, 
         inputRegisters_420__14, inputRegisters_420__13, inputRegisters_420__12, 
         inputRegisters_420__11, inputRegisters_420__10, inputRegisters_420__9, 
         inputRegisters_420__8, inputRegisters_420__7, inputRegisters_420__6, 
         inputRegisters_420__5, inputRegisters_420__4, inputRegisters_420__3, 
         inputRegisters_420__2, inputRegisters_420__1, inputRegisters_420__0, 
         inputRegisters_421__15, inputRegisters_421__14, inputRegisters_421__13, 
         inputRegisters_421__12, inputRegisters_421__11, inputRegisters_421__10, 
         inputRegisters_421__9, inputRegisters_421__8, inputRegisters_421__7, 
         inputRegisters_421__6, inputRegisters_421__5, inputRegisters_421__4, 
         inputRegisters_421__3, inputRegisters_421__2, inputRegisters_421__1, 
         inputRegisters_421__0, inputRegisters_422__15, inputRegisters_422__14, 
         inputRegisters_422__13, inputRegisters_422__12, inputRegisters_422__11, 
         inputRegisters_422__10, inputRegisters_422__9, inputRegisters_422__8, 
         inputRegisters_422__7, inputRegisters_422__6, inputRegisters_422__5, 
         inputRegisters_422__4, inputRegisters_422__3, inputRegisters_422__2, 
         inputRegisters_422__1, inputRegisters_422__0, inputRegisters_423__15, 
         inputRegisters_423__14, inputRegisters_423__13, inputRegisters_423__12, 
         inputRegisters_423__11, inputRegisters_423__10, inputRegisters_423__9, 
         inputRegisters_423__8, inputRegisters_423__7, inputRegisters_423__6, 
         inputRegisters_423__5, inputRegisters_423__4, inputRegisters_423__3, 
         inputRegisters_423__2, inputRegisters_423__1, inputRegisters_423__0, 
         inputRegisters_424__15, inputRegisters_424__14, inputRegisters_424__13, 
         inputRegisters_424__12, inputRegisters_424__11, inputRegisters_424__10, 
         inputRegisters_424__9, inputRegisters_424__8, inputRegisters_424__7, 
         inputRegisters_424__6, inputRegisters_424__5, inputRegisters_424__4, 
         inputRegisters_424__3, inputRegisters_424__2, inputRegisters_424__1, 
         inputRegisters_424__0, inputRegisters_425__15, inputRegisters_425__14, 
         inputRegisters_425__13, inputRegisters_425__12, inputRegisters_425__11, 
         inputRegisters_425__10, inputRegisters_425__9, inputRegisters_425__8, 
         inputRegisters_425__7, inputRegisters_425__6, inputRegisters_425__5, 
         inputRegisters_425__4, inputRegisters_425__3, inputRegisters_425__2, 
         inputRegisters_425__1, inputRegisters_425__0, inputRegisters_426__15, 
         inputRegisters_426__14, inputRegisters_426__13, inputRegisters_426__12, 
         inputRegisters_426__11, inputRegisters_426__10, inputRegisters_426__9, 
         inputRegisters_426__8, inputRegisters_426__7, inputRegisters_426__6, 
         inputRegisters_426__5, inputRegisters_426__4, inputRegisters_426__3, 
         inputRegisters_426__2, inputRegisters_426__1, inputRegisters_426__0, 
         inputRegisters_427__15, inputRegisters_427__14, inputRegisters_427__13, 
         inputRegisters_427__12, inputRegisters_427__11, inputRegisters_427__10, 
         inputRegisters_427__9, inputRegisters_427__8, inputRegisters_427__7, 
         inputRegisters_427__6, inputRegisters_427__5, inputRegisters_427__4, 
         inputRegisters_427__3, inputRegisters_427__2, inputRegisters_427__1, 
         inputRegisters_427__0, inputRegisters_428__15, inputRegisters_428__14, 
         inputRegisters_428__13, inputRegisters_428__12, inputRegisters_428__11, 
         inputRegisters_428__10, inputRegisters_428__9, inputRegisters_428__8, 
         inputRegisters_428__7, inputRegisters_428__6, inputRegisters_428__5, 
         inputRegisters_428__4, inputRegisters_428__3, inputRegisters_428__2, 
         inputRegisters_428__1, inputRegisters_428__0, inputRegisters_429__15, 
         inputRegisters_429__14, inputRegisters_429__13, inputRegisters_429__12, 
         inputRegisters_429__11, inputRegisters_429__10, inputRegisters_429__9, 
         inputRegisters_429__8, inputRegisters_429__7, inputRegisters_429__6, 
         inputRegisters_429__5, inputRegisters_429__4, inputRegisters_429__3, 
         inputRegisters_429__2, inputRegisters_429__1, inputRegisters_429__0, 
         inputRegisters_430__15, inputRegisters_430__14, inputRegisters_430__13, 
         inputRegisters_430__12, inputRegisters_430__11, inputRegisters_430__10, 
         inputRegisters_430__9, inputRegisters_430__8, inputRegisters_430__7, 
         inputRegisters_430__6, inputRegisters_430__5, inputRegisters_430__4, 
         inputRegisters_430__3, inputRegisters_430__2, inputRegisters_430__1, 
         inputRegisters_430__0, inputRegisters_431__15, inputRegisters_431__14, 
         inputRegisters_431__13, inputRegisters_431__12, inputRegisters_431__11, 
         inputRegisters_431__10, inputRegisters_431__9, inputRegisters_431__8, 
         inputRegisters_431__7, inputRegisters_431__6, inputRegisters_431__5, 
         inputRegisters_431__4, inputRegisters_431__3, inputRegisters_431__2, 
         inputRegisters_431__1, inputRegisters_431__0, inputRegisters_432__15, 
         inputRegisters_432__14, inputRegisters_432__13, inputRegisters_432__12, 
         inputRegisters_432__11, inputRegisters_432__10, inputRegisters_432__9, 
         inputRegisters_432__8, inputRegisters_432__7, inputRegisters_432__6, 
         inputRegisters_432__5, inputRegisters_432__4, inputRegisters_432__3, 
         inputRegisters_432__2, inputRegisters_432__1, inputRegisters_432__0, 
         inputRegisters_433__15, inputRegisters_433__14, inputRegisters_433__13, 
         inputRegisters_433__12, inputRegisters_433__11, inputRegisters_433__10, 
         inputRegisters_433__9, inputRegisters_433__8, inputRegisters_433__7, 
         inputRegisters_433__6, inputRegisters_433__5, inputRegisters_433__4, 
         inputRegisters_433__3, inputRegisters_433__2, inputRegisters_433__1, 
         inputRegisters_433__0, inputRegisters_434__15, inputRegisters_434__14, 
         inputRegisters_434__13, inputRegisters_434__12, inputRegisters_434__11, 
         inputRegisters_434__10, inputRegisters_434__9, inputRegisters_434__8, 
         inputRegisters_434__7, inputRegisters_434__6, inputRegisters_434__5, 
         inputRegisters_434__4, inputRegisters_434__3, inputRegisters_434__2, 
         inputRegisters_434__1, inputRegisters_434__0, inputRegisters_435__15, 
         inputRegisters_435__14, inputRegisters_435__13, inputRegisters_435__12, 
         inputRegisters_435__11, inputRegisters_435__10, inputRegisters_435__9, 
         inputRegisters_435__8, inputRegisters_435__7, inputRegisters_435__6, 
         inputRegisters_435__5, inputRegisters_435__4, inputRegisters_435__3, 
         inputRegisters_435__2, inputRegisters_435__1, inputRegisters_435__0, 
         inputRegisters_436__15, inputRegisters_436__14, inputRegisters_436__13, 
         inputRegisters_436__12, inputRegisters_436__11, inputRegisters_436__10, 
         inputRegisters_436__9, inputRegisters_436__8, inputRegisters_436__7, 
         inputRegisters_436__6, inputRegisters_436__5, inputRegisters_436__4, 
         inputRegisters_436__3, inputRegisters_436__2, inputRegisters_436__1, 
         inputRegisters_436__0, inputRegisters_437__15, inputRegisters_437__14, 
         inputRegisters_437__13, inputRegisters_437__12, inputRegisters_437__11, 
         inputRegisters_437__10, inputRegisters_437__9, inputRegisters_437__8, 
         inputRegisters_437__7, inputRegisters_437__6, inputRegisters_437__5, 
         inputRegisters_437__4, inputRegisters_437__3, inputRegisters_437__2, 
         inputRegisters_437__1, inputRegisters_437__0, inputRegisters_438__15, 
         inputRegisters_438__14, inputRegisters_438__13, inputRegisters_438__12, 
         inputRegisters_438__11, inputRegisters_438__10, inputRegisters_438__9, 
         inputRegisters_438__8, inputRegisters_438__7, inputRegisters_438__6, 
         inputRegisters_438__5, inputRegisters_438__4, inputRegisters_438__3, 
         inputRegisters_438__2, inputRegisters_438__1, inputRegisters_438__0, 
         inputRegisters_439__15, inputRegisters_439__14, inputRegisters_439__13, 
         inputRegisters_439__12, inputRegisters_439__11, inputRegisters_439__10, 
         inputRegisters_439__9, inputRegisters_439__8, inputRegisters_439__7, 
         inputRegisters_439__6, inputRegisters_439__5, inputRegisters_439__4, 
         inputRegisters_439__3, inputRegisters_439__2, inputRegisters_439__1, 
         inputRegisters_439__0, inputRegisters_440__15, inputRegisters_440__14, 
         inputRegisters_440__13, inputRegisters_440__12, inputRegisters_440__11, 
         inputRegisters_440__10, inputRegisters_440__9, inputRegisters_440__8, 
         inputRegisters_440__7, inputRegisters_440__6, inputRegisters_440__5, 
         inputRegisters_440__4, inputRegisters_440__3, inputRegisters_440__2, 
         inputRegisters_440__1, inputRegisters_440__0, inputRegisters_441__15, 
         inputRegisters_441__14, inputRegisters_441__13, inputRegisters_441__12, 
         inputRegisters_441__11, inputRegisters_441__10, inputRegisters_441__9, 
         inputRegisters_441__8, inputRegisters_441__7, inputRegisters_441__6, 
         inputRegisters_441__5, inputRegisters_441__4, inputRegisters_441__3, 
         inputRegisters_441__2, inputRegisters_441__1, inputRegisters_441__0, 
         inputRegisters_442__15, inputRegisters_442__14, inputRegisters_442__13, 
         inputRegisters_442__12, inputRegisters_442__11, inputRegisters_442__10, 
         inputRegisters_442__9, inputRegisters_442__8, inputRegisters_442__7, 
         inputRegisters_442__6, inputRegisters_442__5, inputRegisters_442__4, 
         inputRegisters_442__3, inputRegisters_442__2, inputRegisters_442__1, 
         inputRegisters_442__0, inputRegisters_443__15, inputRegisters_443__14, 
         inputRegisters_443__13, inputRegisters_443__12, inputRegisters_443__11, 
         inputRegisters_443__10, inputRegisters_443__9, inputRegisters_443__8, 
         inputRegisters_443__7, inputRegisters_443__6, inputRegisters_443__5, 
         inputRegisters_443__4, inputRegisters_443__3, inputRegisters_443__2, 
         inputRegisters_443__1, inputRegisters_443__0, inputRegisters_444__15, 
         inputRegisters_444__14, inputRegisters_444__13, inputRegisters_444__12, 
         inputRegisters_444__11, inputRegisters_444__10, inputRegisters_444__9, 
         inputRegisters_444__8, inputRegisters_444__7, inputRegisters_444__6, 
         inputRegisters_444__5, inputRegisters_444__4, inputRegisters_444__3, 
         inputRegisters_444__2, inputRegisters_444__1, inputRegisters_444__0, 
         inputRegisters_445__15, inputRegisters_445__14, inputRegisters_445__13, 
         inputRegisters_445__12, inputRegisters_445__11, inputRegisters_445__10, 
         inputRegisters_445__9, inputRegisters_445__8, inputRegisters_445__7, 
         inputRegisters_445__6, inputRegisters_445__5, inputRegisters_445__4, 
         inputRegisters_445__3, inputRegisters_445__2, inputRegisters_445__1, 
         inputRegisters_445__0, inputRegisters_446__15, inputRegisters_446__14, 
         inputRegisters_446__13, inputRegisters_446__12, inputRegisters_446__11, 
         inputRegisters_446__10, inputRegisters_446__9, inputRegisters_446__8, 
         inputRegisters_446__7, inputRegisters_446__6, inputRegisters_446__5, 
         inputRegisters_446__4, inputRegisters_446__3, inputRegisters_446__2, 
         inputRegisters_446__1, inputRegisters_446__0, inputRegisters_447__15, 
         inputRegisters_447__14, inputRegisters_447__13, inputRegisters_447__12, 
         inputRegisters_447__11, inputRegisters_447__10, inputRegisters_447__9, 
         inputRegisters_447__8, inputRegisters_447__7, inputRegisters_447__6, 
         inputRegisters_447__5, inputRegisters_447__4, inputRegisters_447__3, 
         inputRegisters_447__2, inputRegisters_447__1, inputRegisters_447__0, 
         inputRegisters_448__15, inputRegisters_448__14, inputRegisters_448__13, 
         inputRegisters_448__12, inputRegisters_448__11, inputRegisters_448__10, 
         inputRegisters_448__9, inputRegisters_448__8, inputRegisters_448__7, 
         inputRegisters_448__6, inputRegisters_448__5, inputRegisters_448__4, 
         inputRegisters_448__3, inputRegisters_448__2, inputRegisters_448__1, 
         inputRegisters_448__0, inputRegisters_449__15, inputRegisters_449__14, 
         inputRegisters_449__13, inputRegisters_449__12, inputRegisters_449__11, 
         inputRegisters_449__10, inputRegisters_449__9, inputRegisters_449__8, 
         inputRegisters_449__7, inputRegisters_449__6, inputRegisters_449__5, 
         inputRegisters_449__4, inputRegisters_449__3, inputRegisters_449__2, 
         inputRegisters_449__1, inputRegisters_449__0, inputRegisters_450__15, 
         inputRegisters_450__14, inputRegisters_450__13, inputRegisters_450__12, 
         inputRegisters_450__11, inputRegisters_450__10, inputRegisters_450__9, 
         inputRegisters_450__8, inputRegisters_450__7, inputRegisters_450__6, 
         inputRegisters_450__5, inputRegisters_450__4, inputRegisters_450__3, 
         inputRegisters_450__2, inputRegisters_450__1, inputRegisters_450__0, 
         inputRegisters_451__15, inputRegisters_451__14, inputRegisters_451__13, 
         inputRegisters_451__12, inputRegisters_451__11, inputRegisters_451__10, 
         inputRegisters_451__9, inputRegisters_451__8, inputRegisters_451__7, 
         inputRegisters_451__6, inputRegisters_451__5, inputRegisters_451__4, 
         inputRegisters_451__3, inputRegisters_451__2, inputRegisters_451__1, 
         inputRegisters_451__0, inputRegisters_452__15, inputRegisters_452__14, 
         inputRegisters_452__13, inputRegisters_452__12, inputRegisters_452__11, 
         inputRegisters_452__10, inputRegisters_452__9, inputRegisters_452__8, 
         inputRegisters_452__7, inputRegisters_452__6, inputRegisters_452__5, 
         inputRegisters_452__4, inputRegisters_452__3, inputRegisters_452__2, 
         inputRegisters_452__1, inputRegisters_452__0, inputRegisters_453__15, 
         inputRegisters_453__14, inputRegisters_453__13, inputRegisters_453__12, 
         inputRegisters_453__11, inputRegisters_453__10, inputRegisters_453__9, 
         inputRegisters_453__8, inputRegisters_453__7, inputRegisters_453__6, 
         inputRegisters_453__5, inputRegisters_453__4, inputRegisters_453__3, 
         inputRegisters_453__2, inputRegisters_453__1, inputRegisters_453__0, 
         inputRegisters_454__15, inputRegisters_454__14, inputRegisters_454__13, 
         inputRegisters_454__12, inputRegisters_454__11, inputRegisters_454__10, 
         inputRegisters_454__9, inputRegisters_454__8, inputRegisters_454__7, 
         inputRegisters_454__6, inputRegisters_454__5, inputRegisters_454__4, 
         inputRegisters_454__3, inputRegisters_454__2, inputRegisters_454__1, 
         inputRegisters_454__0, inputRegisters_455__15, inputRegisters_455__14, 
         inputRegisters_455__13, inputRegisters_455__12, inputRegisters_455__11, 
         inputRegisters_455__10, inputRegisters_455__9, inputRegisters_455__8, 
         inputRegisters_455__7, inputRegisters_455__6, inputRegisters_455__5, 
         inputRegisters_455__4, inputRegisters_455__3, inputRegisters_455__2, 
         inputRegisters_455__1, inputRegisters_455__0, inputRegisters_456__15, 
         inputRegisters_456__14, inputRegisters_456__13, inputRegisters_456__12, 
         inputRegisters_456__11, inputRegisters_456__10, inputRegisters_456__9, 
         inputRegisters_456__8, inputRegisters_456__7, inputRegisters_456__6, 
         inputRegisters_456__5, inputRegisters_456__4, inputRegisters_456__3, 
         inputRegisters_456__2, inputRegisters_456__1, inputRegisters_456__0, 
         inputRegisters_457__15, inputRegisters_457__14, inputRegisters_457__13, 
         inputRegisters_457__12, inputRegisters_457__11, inputRegisters_457__10, 
         inputRegisters_457__9, inputRegisters_457__8, inputRegisters_457__7, 
         inputRegisters_457__6, inputRegisters_457__5, inputRegisters_457__4, 
         inputRegisters_457__3, inputRegisters_457__2, inputRegisters_457__1, 
         inputRegisters_457__0, inputRegisters_458__15, inputRegisters_458__14, 
         inputRegisters_458__13, inputRegisters_458__12, inputRegisters_458__11, 
         inputRegisters_458__10, inputRegisters_458__9, inputRegisters_458__8, 
         inputRegisters_458__7, inputRegisters_458__6, inputRegisters_458__5, 
         inputRegisters_458__4, inputRegisters_458__3, inputRegisters_458__2, 
         inputRegisters_458__1, inputRegisters_458__0, inputRegisters_459__15, 
         inputRegisters_459__14, inputRegisters_459__13, inputRegisters_459__12, 
         inputRegisters_459__11, inputRegisters_459__10, inputRegisters_459__9, 
         inputRegisters_459__8, inputRegisters_459__7, inputRegisters_459__6, 
         inputRegisters_459__5, inputRegisters_459__4, inputRegisters_459__3, 
         inputRegisters_459__2, inputRegisters_459__1, inputRegisters_459__0, 
         inputRegisters_460__15, inputRegisters_460__14, inputRegisters_460__13, 
         inputRegisters_460__12, inputRegisters_460__11, inputRegisters_460__10, 
         inputRegisters_460__9, inputRegisters_460__8, inputRegisters_460__7, 
         inputRegisters_460__6, inputRegisters_460__5, inputRegisters_460__4, 
         inputRegisters_460__3, inputRegisters_460__2, inputRegisters_460__1, 
         inputRegisters_460__0, inputRegisters_461__15, inputRegisters_461__14, 
         inputRegisters_461__13, inputRegisters_461__12, inputRegisters_461__11, 
         inputRegisters_461__10, inputRegisters_461__9, inputRegisters_461__8, 
         inputRegisters_461__7, inputRegisters_461__6, inputRegisters_461__5, 
         inputRegisters_461__4, inputRegisters_461__3, inputRegisters_461__2, 
         inputRegisters_461__1, inputRegisters_461__0, inputRegisters_462__15, 
         inputRegisters_462__14, inputRegisters_462__13, inputRegisters_462__12, 
         inputRegisters_462__11, inputRegisters_462__10, inputRegisters_462__9, 
         inputRegisters_462__8, inputRegisters_462__7, inputRegisters_462__6, 
         inputRegisters_462__5, inputRegisters_462__4, inputRegisters_462__3, 
         inputRegisters_462__2, inputRegisters_462__1, inputRegisters_462__0, 
         inputRegisters_463__15, inputRegisters_463__14, inputRegisters_463__13, 
         inputRegisters_463__12, inputRegisters_463__11, inputRegisters_463__10, 
         inputRegisters_463__9, inputRegisters_463__8, inputRegisters_463__7, 
         inputRegisters_463__6, inputRegisters_463__5, inputRegisters_463__4, 
         inputRegisters_463__3, inputRegisters_463__2, inputRegisters_463__1, 
         inputRegisters_463__0, inputRegisters_464__15, inputRegisters_464__14, 
         inputRegisters_464__13, inputRegisters_464__12, inputRegisters_464__11, 
         inputRegisters_464__10, inputRegisters_464__9, inputRegisters_464__8, 
         inputRegisters_464__7, inputRegisters_464__6, inputRegisters_464__5, 
         inputRegisters_464__4, inputRegisters_464__3, inputRegisters_464__2, 
         inputRegisters_464__1, inputRegisters_464__0, inputRegisters_465__15, 
         inputRegisters_465__14, inputRegisters_465__13, inputRegisters_465__12, 
         inputRegisters_465__11, inputRegisters_465__10, inputRegisters_465__9, 
         inputRegisters_465__8, inputRegisters_465__7, inputRegisters_465__6, 
         inputRegisters_465__5, inputRegisters_465__4, inputRegisters_465__3, 
         inputRegisters_465__2, inputRegisters_465__1, inputRegisters_465__0, 
         inputRegisters_466__15, inputRegisters_466__14, inputRegisters_466__13, 
         inputRegisters_466__12, inputRegisters_466__11, inputRegisters_466__10, 
         inputRegisters_466__9, inputRegisters_466__8, inputRegisters_466__7, 
         inputRegisters_466__6, inputRegisters_466__5, inputRegisters_466__4, 
         inputRegisters_466__3, inputRegisters_466__2, inputRegisters_466__1, 
         inputRegisters_466__0, inputRegisters_467__15, inputRegisters_467__14, 
         inputRegisters_467__13, inputRegisters_467__12, inputRegisters_467__11, 
         inputRegisters_467__10, inputRegisters_467__9, inputRegisters_467__8, 
         inputRegisters_467__7, inputRegisters_467__6, inputRegisters_467__5, 
         inputRegisters_467__4, inputRegisters_467__3, inputRegisters_467__2, 
         inputRegisters_467__1, inputRegisters_467__0, inputRegisters_468__15, 
         inputRegisters_468__14, inputRegisters_468__13, inputRegisters_468__12, 
         inputRegisters_468__11, inputRegisters_468__10, inputRegisters_468__9, 
         inputRegisters_468__8, inputRegisters_468__7, inputRegisters_468__6, 
         inputRegisters_468__5, inputRegisters_468__4, inputRegisters_468__3, 
         inputRegisters_468__2, inputRegisters_468__1, inputRegisters_468__0, 
         inputRegisters_469__15, inputRegisters_469__14, inputRegisters_469__13, 
         inputRegisters_469__12, inputRegisters_469__11, inputRegisters_469__10, 
         inputRegisters_469__9, inputRegisters_469__8, inputRegisters_469__7, 
         inputRegisters_469__6, inputRegisters_469__5, inputRegisters_469__4, 
         inputRegisters_469__3, inputRegisters_469__2, inputRegisters_469__1, 
         inputRegisters_469__0, inputRegisters_470__15, inputRegisters_470__14, 
         inputRegisters_470__13, inputRegisters_470__12, inputRegisters_470__11, 
         inputRegisters_470__10, inputRegisters_470__9, inputRegisters_470__8, 
         inputRegisters_470__7, inputRegisters_470__6, inputRegisters_470__5, 
         inputRegisters_470__4, inputRegisters_470__3, inputRegisters_470__2, 
         inputRegisters_470__1, inputRegisters_470__0, inputRegisters_471__15, 
         inputRegisters_471__14, inputRegisters_471__13, inputRegisters_471__12, 
         inputRegisters_471__11, inputRegisters_471__10, inputRegisters_471__9, 
         inputRegisters_471__8, inputRegisters_471__7, inputRegisters_471__6, 
         inputRegisters_471__5, inputRegisters_471__4, inputRegisters_471__3, 
         inputRegisters_471__2, inputRegisters_471__1, inputRegisters_471__0, 
         inputRegisters_472__15, inputRegisters_472__14, inputRegisters_472__13, 
         inputRegisters_472__12, inputRegisters_472__11, inputRegisters_472__10, 
         inputRegisters_472__9, inputRegisters_472__8, inputRegisters_472__7, 
         inputRegisters_472__6, inputRegisters_472__5, inputRegisters_472__4, 
         inputRegisters_472__3, inputRegisters_472__2, inputRegisters_472__1, 
         inputRegisters_472__0, inputRegisters_473__15, inputRegisters_473__14, 
         inputRegisters_473__13, inputRegisters_473__12, inputRegisters_473__11, 
         inputRegisters_473__10, inputRegisters_473__9, inputRegisters_473__8, 
         inputRegisters_473__7, inputRegisters_473__6, inputRegisters_473__5, 
         inputRegisters_473__4, inputRegisters_473__3, inputRegisters_473__2, 
         inputRegisters_473__1, inputRegisters_473__0, inputRegisters_474__15, 
         inputRegisters_474__14, inputRegisters_474__13, inputRegisters_474__12, 
         inputRegisters_474__11, inputRegisters_474__10, inputRegisters_474__9, 
         inputRegisters_474__8, inputRegisters_474__7, inputRegisters_474__6, 
         inputRegisters_474__5, inputRegisters_474__4, inputRegisters_474__3, 
         inputRegisters_474__2, inputRegisters_474__1, inputRegisters_474__0, 
         inputRegisters_475__15, inputRegisters_475__14, inputRegisters_475__13, 
         inputRegisters_475__12, inputRegisters_475__11, inputRegisters_475__10, 
         inputRegisters_475__9, inputRegisters_475__8, inputRegisters_475__7, 
         inputRegisters_475__6, inputRegisters_475__5, inputRegisters_475__4, 
         inputRegisters_475__3, inputRegisters_475__2, inputRegisters_475__1, 
         inputRegisters_475__0, inputRegisters_476__15, inputRegisters_476__14, 
         inputRegisters_476__13, inputRegisters_476__12, inputRegisters_476__11, 
         inputRegisters_476__10, inputRegisters_476__9, inputRegisters_476__8, 
         inputRegisters_476__7, inputRegisters_476__6, inputRegisters_476__5, 
         inputRegisters_476__4, inputRegisters_476__3, inputRegisters_476__2, 
         inputRegisters_476__1, inputRegisters_476__0, inputRegisters_477__15, 
         inputRegisters_477__14, inputRegisters_477__13, inputRegisters_477__12, 
         inputRegisters_477__11, inputRegisters_477__10, inputRegisters_477__9, 
         inputRegisters_477__8, inputRegisters_477__7, inputRegisters_477__6, 
         inputRegisters_477__5, inputRegisters_477__4, inputRegisters_477__3, 
         inputRegisters_477__2, inputRegisters_477__1, inputRegisters_477__0, 
         inputRegisters_478__15, inputRegisters_478__14, inputRegisters_478__13, 
         inputRegisters_478__12, inputRegisters_478__11, inputRegisters_478__10, 
         inputRegisters_478__9, inputRegisters_478__8, inputRegisters_478__7, 
         inputRegisters_478__6, inputRegisters_478__5, inputRegisters_478__4, 
         inputRegisters_478__3, inputRegisters_478__2, inputRegisters_478__1, 
         inputRegisters_478__0, inputRegisters_479__15, inputRegisters_479__14, 
         inputRegisters_479__13, inputRegisters_479__12, inputRegisters_479__11, 
         inputRegisters_479__10, inputRegisters_479__9, inputRegisters_479__8, 
         inputRegisters_479__7, inputRegisters_479__6, inputRegisters_479__5, 
         inputRegisters_479__4, inputRegisters_479__3, inputRegisters_479__2, 
         inputRegisters_479__1, inputRegisters_479__0, inputRegisters_480__15, 
         inputRegisters_480__14, inputRegisters_480__13, inputRegisters_480__12, 
         inputRegisters_480__11, inputRegisters_480__10, inputRegisters_480__9, 
         inputRegisters_480__8, inputRegisters_480__7, inputRegisters_480__6, 
         inputRegisters_480__5, inputRegisters_480__4, inputRegisters_480__3, 
         inputRegisters_480__2, inputRegisters_480__1, inputRegisters_480__0, 
         inputRegisters_481__15, inputRegisters_481__14, inputRegisters_481__13, 
         inputRegisters_481__12, inputRegisters_481__11, inputRegisters_481__10, 
         inputRegisters_481__9, inputRegisters_481__8, inputRegisters_481__7, 
         inputRegisters_481__6, inputRegisters_481__5, inputRegisters_481__4, 
         inputRegisters_481__3, inputRegisters_481__2, inputRegisters_481__1, 
         inputRegisters_481__0, inputRegisters_482__15, inputRegisters_482__14, 
         inputRegisters_482__13, inputRegisters_482__12, inputRegisters_482__11, 
         inputRegisters_482__10, inputRegisters_482__9, inputRegisters_482__8, 
         inputRegisters_482__7, inputRegisters_482__6, inputRegisters_482__5, 
         inputRegisters_482__4, inputRegisters_482__3, inputRegisters_482__2, 
         inputRegisters_482__1, inputRegisters_482__0, inputRegisters_483__15, 
         inputRegisters_483__14, inputRegisters_483__13, inputRegisters_483__12, 
         inputRegisters_483__11, inputRegisters_483__10, inputRegisters_483__9, 
         inputRegisters_483__8, inputRegisters_483__7, inputRegisters_483__6, 
         inputRegisters_483__5, inputRegisters_483__4, inputRegisters_483__3, 
         inputRegisters_483__2, inputRegisters_483__1, inputRegisters_483__0, 
         reluMuxOutuput_15, reluMuxOutuput_14, reluMuxOutuput_13, 
         reluMuxOutuput_12, reluMuxOutuput_11, reluMuxOutuput_10, 
         reluMuxOutuput_9, reluMuxOutuput_8, reluMuxOutuput_7, reluMuxOutuput_6, 
         reluMuxOutuput_5, reluMuxOutuput_4, reluMuxOutuput_3, reluMuxOutuput_2, 
         reluMuxOutuput_1, reluMuxOutuput_0, enableRegister_483, 
         enableRegister_482, enableRegister_481, enableRegister_480, 
         enableRegister_479, enableRegister_478, enableRegister_477, 
         enableRegister_476, enableRegister_475, enableRegister_474, 
         enableRegister_473, enableRegister_472, enableRegister_471, 
         enableRegister_470, enableRegister_469, enableRegister_468, 
         enableRegister_467, enableRegister_466, enableRegister_465, 
         enableRegister_464, enableRegister_463, enableRegister_462, 
         enableRegister_461, enableRegister_460, enableRegister_459, 
         enableRegister_458, enableRegister_457, enableRegister_456, 
         enableRegister_455, enableRegister_454, enableRegister_453, 
         enableRegister_452, enableRegister_451, enableRegister_450, 
         enableRegister_449, enableRegister_448, enableRegister_447, 
         enableRegister_446, enableRegister_445, enableRegister_444, 
         enableRegister_443, enableRegister_442, enableRegister_441, 
         enableRegister_440, enableRegister_439, enableRegister_438, 
         enableRegister_437, enableRegister_436, enableRegister_435, 
         enableRegister_434, enableRegister_433, enableRegister_432, 
         enableRegister_431, enableRegister_430, enableRegister_429, 
         enableRegister_428, enableRegister_427, enableRegister_426, 
         enableRegister_425, enableRegister_424, enableRegister_423, 
         enableRegister_422, enableRegister_421, enableRegister_420, 
         enableRegister_419, enableRegister_418, enableRegister_417, 
         enableRegister_416, enableRegister_415, enableRegister_414, 
         enableRegister_413, enableRegister_412, enableRegister_411, 
         enableRegister_410, enableRegister_409, enableRegister_408, 
         enableRegister_407, enableRegister_406, enableRegister_405, 
         enableRegister_404, enableRegister_403, enableRegister_402, 
         enableRegister_401, enableRegister_400, enableRegister_399, 
         enableRegister_398, enableRegister_397, enableRegister_396, 
         enableRegister_395, enableRegister_394, enableRegister_393, 
         enableRegister_392, enableRegister_391, enableRegister_390, 
         enableRegister_389, enableRegister_388, enableRegister_387, 
         enableRegister_386, enableRegister_385, enableRegister_384, 
         enableRegister_383, enableRegister_382, enableRegister_381, 
         enableRegister_380, enableRegister_379, enableRegister_378, 
         enableRegister_377, enableRegister_376, enableRegister_375, 
         enableRegister_374, enableRegister_373, enableRegister_372, 
         enableRegister_371, enableRegister_370, enableRegister_369, 
         enableRegister_368, enableRegister_367, enableRegister_366, 
         enableRegister_365, enableRegister_364, enableRegister_363, 
         enableRegister_362, enableRegister_361, enableRegister_360, 
         enableRegister_359, enableRegister_358, enableRegister_357, 
         enableRegister_356, enableRegister_355, enableRegister_354, 
         enableRegister_353, enableRegister_352, enableRegister_351, 
         enableRegister_350, enableRegister_349, enableRegister_348, 
         enableRegister_347, enableRegister_346, enableRegister_345, 
         enableRegister_344, enableRegister_343, enableRegister_342, 
         enableRegister_341, enableRegister_340, enableRegister_339, 
         enableRegister_338, enableRegister_337, enableRegister_336, 
         enableRegister_335, enableRegister_334, enableRegister_333, 
         enableRegister_332, enableRegister_331, enableRegister_330, 
         enableRegister_329, enableRegister_328, enableRegister_327, 
         enableRegister_326, enableRegister_325, enableRegister_324, 
         enableRegister_323, enableRegister_322, enableRegister_321, 
         enableRegister_320, enableRegister_319, enableRegister_318, 
         enableRegister_317, enableRegister_316, enableRegister_315, 
         enableRegister_314, enableRegister_313, enableRegister_312, 
         enableRegister_311, enableRegister_310, enableRegister_309, 
         enableRegister_308, enableRegister_307, enableRegister_306, 
         enableRegister_305, enableRegister_304, enableRegister_303, 
         enableRegister_302, enableRegister_301, enableRegister_300, 
         enableRegister_299, enableRegister_298, enableRegister_297, 
         enableRegister_296, enableRegister_295, enableRegister_294, 
         enableRegister_293, enableRegister_292, enableRegister_291, 
         enableRegister_290, enableRegister_289, enableRegister_288, 
         enableRegister_287, enableRegister_286, enableRegister_285, 
         enableRegister_284, enableRegister_283, enableRegister_282, 
         enableRegister_281, enableRegister_280, enableRegister_279, 
         enableRegister_278, enableRegister_277, enableRegister_276, 
         enableRegister_275, enableRegister_274, enableRegister_273, 
         enableRegister_272, enableRegister_271, enableRegister_270, 
         enableRegister_269, enableRegister_268, enableRegister_267, 
         enableRegister_266, enableRegister_265, enableRegister_264, 
         enableRegister_263, enableRegister_262, enableRegister_261, 
         enableRegister_260, enableRegister_259, enableRegister_258, 
         enableRegister_257, enableRegister_256, enableRegister_255, 
         enableRegister_254, enableRegister_253, enableRegister_252, 
         enableRegister_251, enableRegister_250, enableRegister_249, 
         enableRegister_248, enableRegister_247, enableRegister_246, 
         enableRegister_245, enableRegister_244, enableRegister_243, 
         enableRegister_242, enableRegister_241, enableRegister_240, 
         enableRegister_239, enableRegister_238, enableRegister_237, 
         enableRegister_236, enableRegister_235, enableRegister_234, 
         enableRegister_233, enableRegister_232, enableRegister_231, 
         enableRegister_230, enableRegister_229, enableRegister_228, 
         enableRegister_227, enableRegister_226, enableRegister_225, 
         enableRegister_224, enableRegister_223, enableRegister_222, 
         enableRegister_221, enableRegister_220, enableRegister_219, 
         enableRegister_218, enableRegister_217, enableRegister_216, 
         enableRegister_215, enableRegister_214, enableRegister_213, 
         enableRegister_212, enableRegister_211, enableRegister_210, 
         enableRegister_209, enableRegister_208, enableRegister_207, 
         enableRegister_206, enableRegister_205, enableRegister_204, 
         enableRegister_203, enableRegister_202, enableRegister_201, 
         enableRegister_200, enableRegister_199, enableRegister_198, 
         enableRegister_197, enableRegister_196, enableRegister_195, 
         enableRegister_194, enableRegister_193, enableRegister_192, 
         enableRegister_191, enableRegister_190, enableRegister_189, 
         enableRegister_188, enableRegister_187, enableRegister_186, 
         enableRegister_185, enableRegister_184, enableRegister_183, 
         enableRegister_182, enableRegister_181, enableRegister_180, 
         enableRegister_179, enableRegister_178, enableRegister_177, 
         enableRegister_176, enableRegister_175, enableRegister_174, 
         enableRegister_173, enableRegister_172, enableRegister_171, 
         enableRegister_170, enableRegister_169, enableRegister_168, 
         enableRegister_167, enableRegister_166, enableRegister_165, 
         enableRegister_164, enableRegister_163, enableRegister_162, 
         enableRegister_161, enableRegister_160, enableRegister_159, 
         enableRegister_158, enableRegister_157, enableRegister_156, 
         enableRegister_155, enableRegister_154, enableRegister_153, 
         enableRegister_152, enableRegister_151, enableRegister_150, 
         enableRegister_149, enableRegister_148, enableRegister_147, 
         enableRegister_146, enableRegister_145, enableRegister_144, 
         enableRegister_143, enableRegister_142, enableRegister_141, 
         enableRegister_140, enableRegister_139, enableRegister_138, 
         enableRegister_137, enableRegister_136, enableRegister_135, 
         enableRegister_134, enableRegister_133, enableRegister_132, 
         enableRegister_131, enableRegister_130, enableRegister_129, 
         enableRegister_128, enableRegister_127, enableRegister_126, 
         enableRegister_125, enableRegister_124, enableRegister_123, 
         enableRegister_122, enableRegister_121, enableRegister_120, 
         enableRegister_119, enableRegister_118, enableRegister_117, 
         enableRegister_116, enableRegister_115, enableRegister_114, 
         enableRegister_113, enableRegister_112, enableRegister_111, 
         enableRegister_110, enableRegister_109, enableRegister_108, 
         enableRegister_107, enableRegister_106, enableRegister_105, 
         enableRegister_104, enableRegister_103, enableRegister_102, 
         enableRegister_101, enableRegister_100, enableRegister_99, 
         enableRegister_98, enableRegister_97, enableRegister_96, 
         enableRegister_95, enableRegister_94, enableRegister_93, 
         enableRegister_92, enableRegister_91, enableRegister_90, 
         enableRegister_89, enableRegister_88, enableRegister_87, 
         enableRegister_86, enableRegister_85, enableRegister_84, 
         enableRegister_83, enableRegister_82, enableRegister_81, 
         enableRegister_80, enableRegister_79, enableRegister_78, 
         enableRegister_77, enableRegister_76, enableRegister_75, 
         enableRegister_74, enableRegister_73, enableRegister_72, 
         enableRegister_71, enableRegister_70, enableRegister_69, 
         enableRegister_68, enableRegister_67, enableRegister_66, 
         enableRegister_65, enableRegister_64, enableRegister_63, 
         enableRegister_62, enableRegister_61, enableRegister_60, 
         enableRegister_59, enableRegister_58, enableRegister_57, 
         enableRegister_56, enableRegister_55, enableRegister_54, 
         enableRegister_53, enableRegister_52, enableRegister_51, 
         enableRegister_50, enableRegister_49, enableRegister_48, 
         enableRegister_47, enableRegister_46, enableRegister_45, 
         enableRegister_44, enableRegister_43, enableRegister_42, 
         enableRegister_41, enableRegister_40, enableRegister_39, 
         enableRegister_38, enableRegister_37, enableRegister_36, 
         enableRegister_35, enableRegister_34, enableRegister_33, 
         enableRegister_32, enableRegister_31, enableRegister_30, 
         enableRegister_29, enableRegister_28, enableRegister_27, 
         enableRegister_26, enableRegister_25, enableRegister_24, 
         enableRegister_23, enableRegister_22, enableRegister_21, 
         enableRegister_20, enableRegister_19, enableRegister_18, 
         enableRegister_17, enableRegister_16, enableRegister_15, 
         enableRegister_14, enableRegister_13, enableRegister_12, 
         enableRegister_11, enableRegister_10, enableRegister_9, 
         enableRegister_8, enableRegister_7, enableRegister_6, enableRegister_5, 
         enableRegister_4, enableRegister_3, enableRegister_2, enableRegister_1, 
         enableRegister_0, registerSelector_8, registerSelector_7, 
         registerSelector_6, registerSelector_5, registerSelector_4, 
         registerSelector_3, registerSelector_2, registerSelector_1, 
         registerSelector_0, notClk, resetCounter, outToRam_15, outToRam_14, 
         outToRam_13, outToRam_12, outToRam_11, outToRam_10, outToRam_9, 
         outToRam_8, outToRam_7, outToRam_6, outToRam_5, outToRam_4, outToRam_3, 
         outToRam_2, outToRam_1, outToRam_0, isRelu, registerOutputs_484__15, 
         nx33625, nx33627, nx33629, nx33631, nx33633, nx33639, nx33641, nx33643, 
         nx33645, nx33647, nx33649, nx33651, nx33653, nx33655, nx33657, nx33659, 
         nx33661, nx33663, nx33665, nx33667, nx33669, nx33671, nx33673, nx33675, 
         nx33677, nx33679, nx33681, nx33683, nx33685, nx33687, nx33689, nx33691, 
         nx33693, nx33695, nx33697, nx33699, nx33701, nx33703, nx33705, nx33707, 
         nx33709, nx33711, nx33713, nx33715, nx33717, nx33719, nx33721, nx33723, 
         nx33725, nx33727, nx33729, nx33731, nx33733, nx33735, nx33737, nx33739, 
         nx33741, nx33743, nx33745, nx33747, nx33749, nx33751, nx33753, nx33755, 
         nx33757, nx33759, nx33761, nx33763, nx33765, nx33767, nx33769, nx33771, 
         nx33773, nx33775, nx33777, nx33779, nx33781, nx33783, nx33785, nx33787, 
         nx33789, nx33791, nx33793, nx33795, nx33797, nx33799, nx33801, nx33803, 
         nx33805, nx33807, nx33809, nx33811, nx33813, nx33815, nx33817, nx33819, 
         nx33821, nx33823, nx33825, nx33827, nx33829, nx33831, nx33833, nx33835, 
         nx33837, nx33839, nx33841, nx33843, nx33845, nx33847, nx33849, nx33851, 
         nx33853, nx33855, nx33857, nx33859, nx33861, nx33863, nx33865, nx33867, 
         nx33869, nx33871, nx33873, nx33875, nx33877, nx33879, nx33881, nx33883, 
         nx33885, nx33887, nx33889, nx33891, nx33893, nx33895, nx33897, nx33899, 
         nx33901, nx33903, nx33905, nx33907, nx33909, nx33911, nx33913, nx33915, 
         nx33917, nx33919, nx33921, nx33923, nx33925, nx33927, nx33929, nx33931, 
         nx33933, nx33935, nx33937, nx33939, nx33941, nx33943, nx33945, nx33947, 
         nx33949, nx33951, nx33953, nx33955, nx33957, nx33959, nx33961, nx33963, 
         nx33965, nx33967, nx33969, nx33971, nx33973, nx33975, nx33977, nx33979, 
         nx33981, nx33983, nx33985, nx33987, nx33989, nx33991, nx33993, nx33995, 
         nx33997, nx33999, nx34001, nx34003, nx34005, nx34007, nx34009, nx34011, 
         nx34013, nx34015, nx34017, nx34019, nx34021, nx34023, nx34025, nx34027, 
         nx34029, nx34031, nx34033, nx34035, nx34037, nx34039, nx34041, nx34043, 
         nx34045, nx34047, nx34049, nx34051, nx34053, nx34055, nx34057, nx34059, 
         nx34061, nx34063, nx34065, nx34067, nx34069, nx34071, nx34073, nx34075, 
         nx34077, nx34079, nx34081, nx34083, nx34085, nx34087, nx34089, nx34091, 
         nx34093, nx34095, nx34097, nx34099, nx34101, nx34103, nx34105, nx34107, 
         nx34109, nx34111, nx34113, nx34115, nx34117, nx34119, nx34121, nx34123, 
         nx34125, nx34127, nx34129, nx34131, nx34133, nx34135, nx34137, nx34139, 
         nx34141, nx34143, nx34145, nx34147, nx34149, nx34151, nx34153, nx34155, 
         nx34157, nx34159, nx34161, nx34163, nx34165, nx34167, nx34169, nx34171, 
         nx34173, nx34175, nx34177, nx34179, nx34181, nx34183, nx34185, nx34187, 
         nx34189, nx34191, nx34193, nx34195, nx34197, nx34199, nx34201, nx34203, 
         nx34205, nx34207, nx34209, nx34211, nx34213, nx34215, nx34217, nx34219, 
         nx34221, nx34223, nx34225, nx34227, nx34229, nx34231, nx34233, nx34235, 
         nx34237, nx34239, nx34241, nx34243, nx34245, nx34247, nx34249, nx34251, 
         nx34253, nx34255, nx34257, nx34259, nx34261, nx34263, nx34265, nx34267, 
         nx34269, nx34271, nx34273, nx34275, nx34277, nx34279, nx34281, nx34283, 
         nx34285, nx34287, nx34289, nx34291, nx34293, nx34295, nx34297, nx34299, 
         nx34301, nx34303, nx34305, nx34307, nx34309, nx34311, nx34313, nx34315, 
         nx34317, nx34319, nx34321, nx34323, nx34325, nx34327, nx34329, nx34331, 
         nx34333, nx34335, nx34337, nx34339, nx34341, nx34343, nx34345, nx34347, 
         nx34349, nx34351, nx34353, nx34355, nx34357, nx34359, nx34361, nx34363, 
         nx34365, nx34367, nx34369, nx34371, nx34373, nx34375, nx34377, nx34379, 
         nx34381, nx34383, nx34385, nx34387, nx34389, nx34391, nx34393, nx34395, 
         nx34397, nx34399, nx34401, nx34403, nx34405, nx34407, nx34409, nx34411, 
         nx34413, nx34415, nx34417, nx34419, nx34421, nx34423, nx34425, nx34427, 
         nx34429, nx34431, nx34433, nx34435, nx34437, nx34439, nx34441, nx34443, 
         nx34445, nx34447, nx34449, nx34451, nx34453, nx34455, nx34457, nx34459, 
         nx34461, nx34463, nx34465, nx34467, nx34469, nx34471, nx34473, nx34475, 
         nx34477, nx34479, nx34481, nx34483, nx34485, nx34487, nx34489, nx34491, 
         nx34493, nx34495, nx34497, nx34499, nx34501, nx34503, nx34505, nx34507, 
         nx34509, nx34511, nx34513, nx34515, nx34517, nx34519, nx34521, nx34523, 
         nx34525, nx34527, nx34529, nx34531, nx34533, nx34535, nx34537, nx34539, 
         nx34541, nx34543, nx34545, nx34547, nx34549, nx34551, nx34553, nx34555, 
         nx34557, nx34559, nx34561, nx34563, nx34565, nx34567, nx34569, nx34571, 
         nx34573, nx34575, nx34577, nx34579, nx34581, nx34583, nx34585, nx34587, 
         nx34589, nx34591, nx34593, nx34595, nx34597, nx34599, nx34601, nx34603, 
         nx34605, nx34607, nx34609, nx34611, nx34613, nx34615, nx34617, nx34619, 
         nx34621, nx34623, nx34625, nx34627, nx34629, nx34631, nx34633, nx34635, 
         nx34637, nx34639, nx34641, nx34643, nx34645, nx34647, nx34649, nx34651, 
         nx34653, nx34655, nx34657, nx34659, nx34661, nx34663, nx34665, nx34667, 
         nx34669, nx34671, nx34673, nx34675, nx34677, nx34679, nx34681, nx34683, 
         nx34685, nx34687, nx34689, nx34691, nx34693, nx34695, nx34697, nx34699, 
         nx34701, nx34703, nx34705, nx34707, nx34709, nx34711, nx34713, nx34715, 
         nx34717, nx34719, nx34721, nx34723, nx34725, nx34727, nx34729, nx34731, 
         nx34733, nx34735, nx34737, nx34739, nx34741, nx34743, nx34745, nx34747, 
         nx34749, nx34751, nx34753, nx34755, nx34757, nx34759, nx34761, nx34763, 
         nx34765, nx34767, nx34769, nx34771, nx34773, nx34775, nx34777, nx34779, 
         nx34781, nx34783, nx34785, nx34787, nx34789, nx34791, nx34793, nx34795, 
         nx34797, nx34799, nx34801, nx34803, nx34805, nx34807, nx34809, nx34811, 
         nx34813, nx34815, nx34817, nx34819, nx34821, nx34823, nx34825, nx34827, 
         nx34829, nx34831, nx34833, nx34835, nx34837, nx34839, nx34841, nx34843, 
         nx34845, nx34847, nx34849, nx34851, nx34853, nx34855, nx34857, nx34859, 
         nx34861, nx34863, nx34865, nx34867, nx34869, nx34871, nx34873, nx34875, 
         nx34877, nx34879, nx34881, nx34883, nx34885, nx34887, nx34889, nx34891, 
         nx34893, nx34895, nx34897, nx34899, nx34901, nx34903, nx34905, nx34907, 
         nx34909, nx34911, nx34913, nx34915, nx34917, nx34919, nx34921, nx34923, 
         nx34925, nx34927, nx34929, nx34931, nx34933, nx34935, nx34937, nx34939, 
         nx34941, nx34943, nx34945, nx34947, nx34949, nx34951, nx34953, nx34955, 
         nx34957, nx34959, nx34961, nx34963, nx34965, nx34967, nx34969, nx34971, 
         nx34973, nx34975, nx34977, nx34979, nx34981, nx34983, nx34985, nx34987, 
         nx34989, nx34991, nx34993, nx34995, nx34997, nx34999, nx35001, nx35003, 
         nx35005, nx35007, nx35009, nx35011, nx35013, nx35015, nx35017, nx35019, 
         nx35021, nx35023, nx35025, nx35027, nx35029, nx35031, nx35033, nx35035, 
         nx35037, nx35039, nx35041, nx35043, nx35045, nx35047, nx35049, nx35051, 
         nx35053, nx35055, nx35057, nx35059, nx35061, nx35063, nx35065, nx35067, 
         nx35069, nx35071, nx35073, nx35075, nx35077, nx35079, nx35081, nx35083, 
         nx35085, nx35087, nx35089, nx35091, nx35093, nx35095, nx35097, nx35099, 
         nx35101, nx35103, nx35105, nx35107, nx35109, nx35111, nx35113, nx35115, 
         nx35117, nx35119, nx35121, nx35123, nx35125, nx35127, nx35129, nx35131, 
         nx35133, nx35135, nx35137, nx35139, nx35141, nx35143, nx35145, nx35147, 
         nx35149, nx35151, nx35153, nx35155, nx35157, nx35159, nx35161, nx35163, 
         nx35165, nx35167, nx35169, nx35171, nx35173, nx35175, nx35177, nx35179, 
         nx35181, nx35183, nx35185, nx35187, nx35189, nx35191, nx35193, nx35195, 
         nx35197, nx35199, nx35201, nx35203, nx35205, nx35207, nx35209, nx35211, 
         nx35213, nx35215, nx35217, nx35219, nx35221, nx35223, nx35225, nx35227, 
         nx35229, nx35231, nx35233, nx35235, nx35237, nx35239, nx35241, nx35243, 
         nx35245, nx35247, nx35249, nx35251, nx35253, nx35255, nx35257, nx35259, 
         nx35261, nx35263, nx35265, nx35267, nx35269, nx35271, nx35273, nx35275, 
         nx35277, nx35279, nx35281, nx35283, nx35285, nx35287, nx35289, nx35291, 
         nx35293, nx35295, nx35297, nx35299, nx35301, nx35303, nx35305, nx35307, 
         nx35309, nx35311, nx35313, nx35315, nx35317, nx35319, nx35321, nx35323, 
         nx35325, nx35327, nx35329, nx35331, nx35333, nx35335, nx35337, nx35339, 
         nx35341, nx35343, nx35345, nx35347, nx35349, nx35351, nx35353, nx35355, 
         nx35357, nx35359, nx35361, nx35363, nx35365, nx35367, nx35369, nx35371, 
         nx35373, nx35375, nx35377, nx35379, nx35381, nx35383, nx35385, nx35387, 
         nx35389, nx35391, nx35393, nx35395, nx35397, nx35399, nx35401, nx35403, 
         nx35405, nx35407, nx35409, nx35411, nx35413, nx35415, nx35417, nx35419, 
         nx35421, nx35423, nx35425, nx35427, nx35429, nx35431, nx35433, nx35435, 
         nx35437, nx35439, nx35441, nx35443, nx35445, nx35447, nx35449, nx35451, 
         nx35453, nx35455, nx35457, nx35459, nx35461, nx35463, nx35465, nx35467, 
         nx35469, nx35471, nx35473, nx35475, nx35477, nx35479, nx35481, nx35483, 
         nx35485, nx35487, nx35489, nx35491, nx35493, nx35495, nx35497, nx35499, 
         nx35501, nx35503, nx35505, nx35507, nx35509, nx35511, nx35513, nx35515, 
         nx35517, nx35519, nx35521, nx35523, nx35525, nx35527, nx35529, nx35531, 
         nx35533, nx35535, nx35537, nx35539, nx35541, nx35543, nx35545, nx35547, 
         nx35549, nx35551, nx35553, nx35555, nx35557, nx35559, nx35561, nx35563, 
         nx35565, nx35567, nx35569, nx35571, nx35573, nx35575, nx35577, nx35579, 
         nx35581, nx35583, nx35585, nx35587, nx35589, nx35591, nx35593, nx35595, 
         nx35597, nx35599, nx35601, nx35603, nx35605, nx35607, nx35609, nx35611, 
         nx35613, nx35615, nx35617, nx35619, nx35621, nx35623, nx35625, nx35627, 
         nx35629, nx35631, nx35633, nx35635, nx35637, nx35639, nx35641, nx35643, 
         nx35645, nx35647, nx35649, nx35651, nx35653, nx35655, nx35657, nx35659, 
         nx35661, nx35663, nx35665, nx35667, nx35669, nx35671, nx35673, nx35675, 
         nx35677, nx35679, nx35681, nx35683, nx35685, nx35687, nx35689, nx35691, 
         nx35693, nx35695, nx35697, nx35699, nx35701, nx35703, nx35705, nx35707, 
         nx35709, nx35711, nx35713, nx35715, nx35717, nx35719, nx35721, nx35723, 
         nx35725, nx35727, nx35729, nx35731, nx35733, nx35735, nx35737, nx35739, 
         nx35741, nx35743, nx35745, nx35747, nx35749, nx35751, nx35753, nx35755, 
         nx35757, nx35759, nx35761, nx35763, nx35765, nx35767, nx35769, nx35771, 
         nx35773, nx35775, nx35777, nx35779, nx35781, nx35783, nx35785, nx35787, 
         nx35789, nx35791, nx35793, nx35795, nx35797, nx35799, nx35801, nx35803, 
         nx35805, nx35807, nx35809, nx35811, nx35813, nx35815, nx35817, nx35819, 
         nx35821, nx35823, nx35825, nx35827, nx35829, nx35831, nx35833, nx35835, 
         nx35837, nx35839, nx35841, nx35843, nx35845, nx35847, nx35849, nx35851, 
         nx35853, nx35855, nx35857, nx35859, nx35861, nx35863, nx35865, nx35867, 
         nx35869, nx35871, nx35873, nx35875, nx35877, nx35879, nx35881, nx35885, 
         nx35887, nx35889, nx35891, nx35893, nx35895, nx35897, nx35899, nx35901, 
         nx35903, nx35905, nx35907, nx35909, nx35911, nx35913, nx35915, nx35917, 
         nx35919, nx35921, nx35923, nx35925, nx35927, nx35929, nx35931, nx35933, 
         nx35935, nx35937, nx35939, nx35941, nx35943, nx35945, nx35947, nx35949, 
         nx35951, nx35953, nx35955, nx35957, nx35959, nx35961, nx35963, nx35965, 
         nx35967, nx35969, nx35971, nx35973, nx35975, nx35977, nx35979, nx35981, 
         nx35983, nx35985, nx35987, nx35989, nx35991, nx35993, nx35995, nx35997, 
         nx35999, nx36001, nx36003, nx36005, nx36007, nx36009, nx36011, nx36013, 
         nx36015, nx36017, nx36019, nx36021, nx36023, nx36027, nx36029, nx36031, 
         nx36033, nx36035, nx36037, nx36039, nx36041, nx36043, nx36045, nx36047, 
         nx36049, nx36051, nx36053, nx36055, nx36057, nx36059, nx36061, nx36063, 
         nx36065, nx36067, nx36069, nx36071, nx36073, nx36075, nx36077, nx36079, 
         nx36081, nx36083, nx36085, nx36087, nx36089, nx36091, nx36093, nx36095, 
         nx36097, nx36099, nx36101, nx36103, nx36105, nx36107, nx36109, nx36111, 
         nx36113, nx36115, nx36117, nx36119, nx36121, nx36123, nx36125, nx36127, 
         nx36129, nx36131, nx36133, nx36135, nx36137, nx36139, nx36141, nx36143, 
         nx36145, nx36147, nx36149, nx36151, nx36153, nx36155, nx36157, nx36159, 
         nx36161, nx36163, nx36165, nx36169, nx36171, nx36173, nx36175, nx36177, 
         nx36179, nx36181, nx36183, nx36185, nx36187, nx36189, nx36191, nx36193, 
         nx36195, nx36197, nx36199, nx36201, nx36203, nx36205, nx36207, nx36209, 
         nx36211, nx36213, nx36215, nx36217, nx36219, nx36221, nx36223, nx36225, 
         nx36227, nx36229, nx36231, nx36233, nx36235, nx36237, nx36239, nx36241, 
         nx36243, nx36245, nx36247, nx36249, nx36251, nx36253, nx36255, nx36257, 
         nx36259, nx36261, nx36263, nx36265, nx36267, nx36269, nx36271, nx36273, 
         nx36275, nx36277, nx36279, nx36281, nx36283, nx36285, nx36287, nx36289, 
         nx36291, nx36293, nx36295, nx36297, nx36299, nx36301, nx36303, nx36305, 
         nx36307, nx36311, nx36313, nx36315, nx36317, nx36319, nx36321, nx36323, 
         nx36325, nx36327, nx36329, nx36331, nx36333, nx36335, nx36337, nx36339, 
         nx36341, nx36343, nx36345, nx36347, nx36349, nx36351, nx36353, nx36355, 
         nx36357, nx36359, nx36361, nx36363, nx36365, nx36367, nx36369, nx36371, 
         nx36373, nx36375, nx36377, nx36379, nx36381, nx36383, nx36385, nx36387, 
         nx36389, nx36391, nx36393, nx36395, nx36397, nx36399, nx36401, nx36403, 
         nx36405, nx36407, nx36409, nx36411, nx36413, nx36415, nx36417, nx36419, 
         nx36421, nx36423, nx36425, nx36427, nx36429, nx36431, nx36433, nx36435, 
         nx36437, nx36439, nx36441, nx36443, nx36445, nx36447, nx36449, nx36453, 
         nx36455, nx36457, nx36459, nx36461, nx36463, nx36465, nx36467, nx36469, 
         nx36471, nx36473, nx36475, nx36477, nx36479, nx36481, nx36483, nx36485, 
         nx36487, nx36489, nx36491, nx36493, nx36495, nx36497, nx36499, nx36501, 
         nx36503, nx36505, nx36507, nx36509, nx36511, nx36513, nx36515, nx36517, 
         nx36519, nx36521, nx36523, nx36525, nx36527, nx36529, nx36531, nx36533, 
         nx36535, nx36537, nx36539, nx36541, nx36543, nx36545, nx36547, nx36549, 
         nx36551, nx36553, nx36555, nx36557, nx36559, nx36561, nx36563, nx36565, 
         nx36567, nx36569, nx36571, nx36573, nx36575, nx36577, nx36579, nx36581, 
         nx36583, nx36585, nx36587, nx36589, nx36591, nx36595, nx36597, nx36599, 
         nx36601, nx36603, nx36605, nx36607, nx36609, nx36611, nx36613, nx36615, 
         nx36617, nx36619, nx36621, nx36623, nx36625, nx36627, nx36629, nx36631, 
         nx36633, nx36635, nx36637, nx36639, nx36641, nx36643, nx36645, nx36647, 
         nx36649, nx36651, nx36653, nx36655, nx36657, nx36659, nx36661, nx36663, 
         nx36665, nx36667, nx36669, nx36671, nx36673, nx36675, nx36677, nx36679, 
         nx36681, nx36683, nx36685, nx36687, nx36689, nx36691, nx36693, nx36695, 
         nx36697, nx36699, nx36701, nx36703, nx36705, nx36707, nx36709, nx36711, 
         nx36713, nx36715, nx36717, nx36719, nx36721, nx36723, nx36725, nx36727, 
         nx36729, nx36731, nx36733, nx36737, nx36739, nx36741, nx36743, nx36745, 
         nx36747, nx36749, nx36751, nx36753, nx36755, nx36757, nx36759, nx36761, 
         nx36763, nx36765, nx36767, nx36769, nx36771, nx36773, nx36775, nx36777, 
         nx36779, nx36781, nx36783, nx36785, nx36787, nx36789, nx36791, nx36793, 
         nx36795, nx36797, nx36799, nx36801, nx36803, nx36805, nx36807, nx36809, 
         nx36811, nx36813, nx36815, nx36817, nx36819, nx36821, nx36823, nx36825, 
         nx36827, nx36829, nx36831, nx36833, nx36835, nx36837, nx36839, nx36841, 
         nx36843, nx36845, nx36847, nx36849, nx36851, nx36853, nx36855, nx36857, 
         nx36859, nx36861, nx36863, nx36865, nx36867, nx36869, nx36871, nx36873, 
         nx36875, nx36879, nx36881, nx36883, nx36885, nx36887, nx36889, nx36891, 
         nx36893, nx36895, nx36897, nx36899, nx36901, nx36903, nx36905, nx36907, 
         nx36909, nx36911, nx36913, nx36915, nx36917, nx36919, nx36921, nx36923, 
         nx36925, nx36927, nx36929, nx36931, nx36933, nx36935, nx36937, nx36939, 
         nx36941, nx36943, nx36945, nx36947, nx36949, nx36951, nx36953, nx36955, 
         nx36957, nx36959, nx36961, nx36963, nx36965, nx36967, nx36969, nx36971, 
         nx36973, nx36975, nx36977, nx36979, nx36981, nx36983, nx36985, nx36987, 
         nx36989, nx36991, nx36993, nx36995, nx36997, nx36999, nx37001, nx37003, 
         nx37005, nx37007, nx37009, nx37011, nx37013, nx37015, nx37017, nx37021, 
         nx37023, nx37025, nx37027, nx37029, nx37031, nx37033, nx37035, nx37037, 
         nx37039, nx37041, nx37043, nx37045, nx37047, nx37049, nx37051, nx37053, 
         nx37055, nx37057, nx37059, nx37061, nx37063, nx37065, nx37067, nx37069, 
         nx37071, nx37073, nx37075, nx37077, nx37079, nx37081, nx37083, nx37085, 
         nx37087, nx37089, nx37091, nx37093, nx37095, nx37097, nx37099, nx37101, 
         nx37103, nx37105, nx37107, nx37109, nx37111, nx37113, nx37115, nx37117, 
         nx37119, nx37121, nx37123, nx37125, nx37127, nx37129, nx37131, nx37133, 
         nx37135, nx37137, nx37139, nx37141, nx37143, nx37145, nx37147, nx37149, 
         nx37151, nx37153, nx37155, nx37157, nx37159, nx37163, nx37165, nx37167, 
         nx37169, nx37171, nx37173, nx37175, nx37177, nx37179, nx37181, nx37183, 
         nx37185, nx37187, nx37189, nx37191, nx37193, nx37195, nx37197, nx37199, 
         nx37201, nx37203, nx37205, nx37207, nx37209, nx37211, nx37213, nx37215, 
         nx37217, nx37219, nx37221, nx37223, nx37225, nx37227, nx37229, nx37231, 
         nx37233, nx37235, nx37237, nx37239, nx37241, nx37243, nx37245, nx37247, 
         nx37249, nx37251, nx37253, nx37255, nx37257, nx37259, nx37261, nx37263, 
         nx37265, nx37267, nx37269, nx37271, nx37273, nx37275, nx37277, nx37279, 
         nx37281, nx37283, nx37285, nx37287, nx37289, nx37291, nx37293, nx37295, 
         nx37297, nx37299, nx37301, nx37305, nx37307, nx37309, nx37311, nx37313, 
         nx37315, nx37317, nx37319, nx37321, nx37323, nx37325, nx37327, nx37329, 
         nx37331, nx37333, nx37335, nx37337, nx37339, nx37341, nx37343, nx37345, 
         nx37347, nx37349, nx37351, nx37353, nx37355, nx37357, nx37359, nx37361, 
         nx37363, nx37365, nx37367, nx37369, nx37371, nx37373, nx37375, nx37377, 
         nx37379, nx37381, nx37383, nx37385, nx37387, nx37389, nx37391, nx37393, 
         nx37395, nx37397, nx37399, nx37401, nx37403, nx37405, nx37407, nx37409, 
         nx37411, nx37413, nx37415, nx37417, nx37419, nx37421, nx37423, nx37425, 
         nx37427, nx37429, nx37431, nx37433, nx37435, nx37437, nx37439, nx37441, 
         nx37443, nx37447, nx37449, nx37451, nx37453, nx37455, nx37457, nx37459, 
         nx37461, nx37463, nx37465, nx37467, nx37469, nx37471, nx37473, nx37475, 
         nx37477, nx37479, nx37481, nx37483, nx37485, nx37487, nx37489, nx37491, 
         nx37493, nx37495, nx37497, nx37499, nx37501, nx37503, nx37505, nx37507, 
         nx37509, nx37511, nx37513, nx37515, nx37517, nx37519, nx37521, nx37523, 
         nx37525, nx37527, nx37529, nx37531, nx37533, nx37535, nx37537, nx37539, 
         nx37541, nx37543, nx37545, nx37547, nx37549, nx37551, nx37553, nx37555, 
         nx37557, nx37559, nx37561, nx37563, nx37565, nx37567, nx37569, nx37571, 
         nx37573, nx37575, nx37577, nx37579, nx37581, nx37583, nx37585, nx37589, 
         nx37591, nx37593, nx37595, nx37597, nx37599, nx37601, nx37603, nx37605, 
         nx37607, nx37609, nx37611, nx37613, nx37615, nx37617, nx37619, nx37621, 
         nx37623, nx37625, nx37627, nx37629, nx37631, nx37633, nx37635, nx37637, 
         nx37639, nx37641, nx37643, nx37645, nx37647, nx37649, nx37651, nx37653, 
         nx37655, nx37657, nx37659, nx37661, nx37663, nx37665, nx37667, nx37669, 
         nx37671, nx37673, nx37675, nx37677, nx37679, nx37681, nx37683, nx37685, 
         nx37687, nx37689, nx37691, nx37693, nx37695, nx37697, nx37699, nx37701, 
         nx37703, nx37705, nx37707, nx37709, nx37711, nx37713, nx37715, nx37717, 
         nx37719, nx37721, nx37723, nx37725, nx37727, nx37731, nx37733, nx37735, 
         nx37737, nx37739, nx37741, nx37743, nx37745, nx37747, nx37749, nx37751, 
         nx37753, nx37755, nx37757, nx37759, nx37761, nx37763, nx37765, nx37767, 
         nx37769, nx37771, nx37773, nx37775, nx37777, nx37779, nx37781, nx37783, 
         nx37785, nx37787, nx37789, nx37791, nx37793, nx37795, nx37797, nx37799, 
         nx37801, nx37803, nx37805, nx37807, nx37809, nx37811, nx37813, nx37815, 
         nx37817, nx37819, nx37821, nx37823, nx37825, nx37827, nx37829, nx37831, 
         nx37833, nx37835, nx37837, nx37839, nx37841, nx37843, nx37845, nx37847, 
         nx37849, nx37851, nx37853, nx37855, nx37857, nx37859, nx37861, nx37863, 
         nx37865, nx37867, nx37869, nx37873, nx37875, nx37877, nx37879, nx37881, 
         nx37883, nx37885, nx37887, nx37889, nx37891, nx37893, nx37895, nx37897, 
         nx37899, nx37901, nx37903, nx37905, nx37907, nx37909, nx37911, nx37913, 
         nx37915, nx37917, nx37919, nx37921, nx37923, nx37925, nx37927, nx37929, 
         nx37931, nx37933, nx37935, nx37937, nx37939, nx37941, nx37943, nx37945, 
         nx37947, nx37949, nx37951, nx37953, nx37955, nx37957, nx37959, nx37961, 
         nx37963, nx37965, nx37967, nx37969, nx37971, nx37973, nx37975, nx37977, 
         nx37979, nx37981, nx37983, nx37985, nx37987, nx37989, nx37991, nx37993, 
         nx37995, nx37997, nx37999, nx38001, nx38003, nx38005, nx38007, nx38009, 
         nx38011, nx38015, nx38017, nx38019, nx38021, nx38023, nx38025, nx38027, 
         nx38029, nx38031, nx38033, nx38035, nx38037, nx38039, nx38041, nx38043, 
         nx38045, nx38047, nx38049, nx38051, nx38053, nx38055, nx38057, nx38059, 
         nx38061, nx38063, nx38065, nx38067, nx38069, nx38071, nx38073, nx38075, 
         nx38077, nx38079, nx38081, nx38083, nx38085, nx38087, nx38089, nx38091, 
         nx38093, nx38095, nx38097, nx38099, nx38101, nx38103, nx38105, nx38107, 
         nx38109, nx38111, nx38113, nx38115, nx38117, nx38119, nx38121, nx38123, 
         nx38125, nx38127, nx38129, nx38131, nx38133, nx38135, nx38137, nx38139, 
         nx38141, nx38143, nx38145, nx38147, nx38149, nx38151, nx38153, nx38155, 
         nx38157, nx38159, nx38161, nx38163, nx38165, nx38167, nx38169, nx38171, 
         nx38173, nx38175, nx38177, nx38179, nx38181, nx38183, nx38185, nx38187, 
         nx38189, nx38191, nx38193, nx38195, nx38197, nx38199, nx38201, nx38203, 
         nx38205, nx38207, nx38209, nx38211, nx38213, nx38215, nx38217, nx38219, 
         nx38221, nx38223, nx38225, nx38227, nx38229, nx38231, nx38233, nx38235, 
         nx38237, nx38239, nx38241, nx38243, nx38245, nx38247, nx38249, nx38251, 
         nx38253, nx38255, nx38257, nx38259, nx38261, nx38263, nx38265, nx38267, 
         nx38269, nx38271, nx38273, nx38275, nx38277, nx38279, nx38281, nx38283, 
         nx38285, nx38287, nx38289, nx38291, nx38293, nx38295, nx38297, nx38299, 
         nx38301, nx38303, nx38305, nx38307, nx38309, nx38311, nx38313, nx38315, 
         nx38317, nx38319, nx38321, nx38323, nx38325, nx38327, nx38329, nx38331, 
         nx38333, nx38335, nx38337, nx38339, nx38341, nx38343, nx38345, nx38347, 
         nx38349, nx38351, nx38353, nx38355, nx38357, nx38359, nx38361, nx38363, 
         nx38365, nx38367, nx38369, nx38371, nx38373, nx38375, nx38377, nx38379, 
         nx38381, nx38383, nx38385, nx38387, nx38389, nx38391, nx38393, nx38395, 
         nx38397, nx38399, nx38401, nx38403, nx38405, nx38407, nx38409, nx38411, 
         nx38413, nx38415, nx38417, nx38419, nx38421, nx38423, nx38425, nx38427, 
         nx38429, nx38431, nx38433, nx38435, nx38437, nx38439, nx38441, nx38443, 
         nx38445, nx38447, nx38449, nx38451, nx38453, nx38455, nx38457, nx38459, 
         nx38461, nx38463, nx38465, nx38467, nx38469, nx38471, nx38473, nx38475, 
         nx38477, nx38479, nx38481, nx38483, nx38485, nx38487, nx38489, nx38491, 
         nx38493, nx38495, nx38497, nx38499, nx38501, nx38503, nx38505, nx38507, 
         nx38509, nx38511, nx38513, nx38515, nx38517, nx38519, nx38521, nx38523, 
         nx38525, nx38527, nx38529, nx38531, nx38533, nx38535, nx38537, nx38539, 
         nx38541, nx38543, nx38545, nx38547, nx38549, nx38551, nx38553, nx38555, 
         nx38557, nx38559, nx38561, nx38563, nx38565, nx38567, nx38569, nx38571, 
         nx38573, nx38575, nx38577, nx38579, nx38581, nx38583, nx38585, nx38587, 
         nx38589, nx38591, nx38593, nx38595, nx38597, nx38599, nx38601, nx38603, 
         nx38605, nx38607, nx38609, nx38611, nx38613, nx38615, nx38617, nx38619, 
         nx38621, nx38623, nx38625, nx38627, nx38629, nx38631, nx38633, nx38635, 
         nx38637, nx38639, nx38641, nx38643, nx38645, nx38647, nx38649, nx38651, 
         nx38653, nx38655, nx38657, nx38659, nx38661, nx38663, nx38665, nx38667, 
         nx38669, nx38671, nx38673, nx38675, nx38677, nx38679, nx38681, nx38683, 
         nx38685, nx38687, nx38689, nx38691, nx38693, nx38695, nx38697, nx38699, 
         nx38701, nx38703, nx38705, nx38707, nx38709, nx38711, nx38713, nx38715, 
         nx38717, nx38719, nx38721, nx38723, nx38725, nx38727, nx38729, nx38731, 
         nx38733, nx38735, nx38737, nx38739, nx38741, nx38743, nx38745, nx38747, 
         nx38749, nx38751, nx38753, nx38755, nx38757, nx38759, nx38761, nx38763, 
         nx38765, nx38767, nx38769, nx38771, nx38773, nx38775, nx38777, nx38779, 
         nx38785, nx38787, nx38789, nx38791, nx38793, nx38795, nx38797, nx38799, 
         nx38801, nx38803, nx38805, nx38807, nx38809, nx38811, nx38813, nx38815, 
         nx38817, nx38819, nx38821, nx38823, nx38825, nx38827, nx38829, nx38831, 
         nx38833, nx38835, nx38837, nx38839, nx38841, nx38843, nx38845, nx38847, 
         nx38849, nx38851, nx38853, nx38855, nx38857, nx38859, nx38861, nx38863, 
         nx38865, nx38867, nx38869, nx38871, nx38873, nx38875, nx38877, nx38879, 
         nx38881, nx38883, nx38885, nx38887, nx38889, nx38891, nx38893, nx38895, 
         nx38897, nx38899, nx38901;
    wire [27:0] \$dummy ;




    Decoder_9 decoderLabel (.T ({nx33625,registerSelector_7,nx38155,
              registerSelector_5,registerSelector_4,nx38157,nx33627,
              registerSelector_1,nx33631}), .en (enableDecoder), .decoded ({
              \$dummy [0],\$dummy [1],\$dummy [2],\$dummy [3],\$dummy [4],
              \$dummy [5],\$dummy [6],\$dummy [7],\$dummy [8],\$dummy [9],
              \$dummy [10],\$dummy [11],\$dummy [12],\$dummy [13],\$dummy [14],
              \$dummy [15],\$dummy [16],\$dummy [17],\$dummy [18],\$dummy [19],
              \$dummy [20],\$dummy [21],\$dummy [22],\$dummy [23],\$dummy [24],
              \$dummy [25],\$dummy [26],\$dummy [27],decoderOutput_483,
              decoderOutput_482,decoderOutput_481,decoderOutput_480,
              decoderOutput_479,decoderOutput_478,decoderOutput_477,
              decoderOutput_476,decoderOutput_475,decoderOutput_474,
              decoderOutput_473,decoderOutput_472,decoderOutput_471,
              decoderOutput_470,decoderOutput_469,decoderOutput_468,
              decoderOutput_467,decoderOutput_466,decoderOutput_465,
              decoderOutput_464,decoderOutput_463,decoderOutput_462,
              decoderOutput_461,decoderOutput_460,decoderOutput_459,
              decoderOutput_458,decoderOutput_457,decoderOutput_456,
              decoderOutput_455,decoderOutput_454,decoderOutput_453,
              decoderOutput_452,decoderOutput_451,decoderOutput_450,
              decoderOutput_449,decoderOutput_448,decoderOutput_447,
              decoderOutput_446,decoderOutput_445,decoderOutput_444,
              decoderOutput_443,decoderOutput_442,decoderOutput_441,
              decoderOutput_440,decoderOutput_439,decoderOutput_438,
              decoderOutput_437,decoderOutput_436,decoderOutput_435,
              decoderOutput_434,decoderOutput_433,decoderOutput_432,
              decoderOutput_431,decoderOutput_430,decoderOutput_429,
              decoderOutput_428,decoderOutput_427,decoderOutput_426,
              decoderOutput_425,decoderOutput_424,decoderOutput_423,
              decoderOutput_422,decoderOutput_421,decoderOutput_420,
              decoderOutput_419,decoderOutput_418,decoderOutput_417,
              decoderOutput_416,decoderOutput_415,decoderOutput_414,
              decoderOutput_413,decoderOutput_412,decoderOutput_411,
              decoderOutput_410,decoderOutput_409,decoderOutput_408,
              decoderOutput_407,decoderOutput_406,decoderOutput_405,
              decoderOutput_404,decoderOutput_403,decoderOutput_402,
              decoderOutput_401,decoderOutput_400,decoderOutput_399,
              decoderOutput_398,decoderOutput_397,decoderOutput_396,
              decoderOutput_395,decoderOutput_394,decoderOutput_393,
              decoderOutput_392,decoderOutput_391,decoderOutput_390,
              decoderOutput_389,decoderOutput_388,decoderOutput_387,
              decoderOutput_386,decoderOutput_385,decoderOutput_384,
              decoderOutput_383,decoderOutput_382,decoderOutput_381,
              decoderOutput_380,decoderOutput_379,decoderOutput_378,
              decoderOutput_377,decoderOutput_376,decoderOutput_375,
              decoderOutput_374,decoderOutput_373,decoderOutput_372,
              decoderOutput_371,decoderOutput_370,decoderOutput_369,
              decoderOutput_368,decoderOutput_367,decoderOutput_366,
              decoderOutput_365,decoderOutput_364,decoderOutput_363,
              decoderOutput_362,decoderOutput_361,decoderOutput_360,
              decoderOutput_359,decoderOutput_358,decoderOutput_357,
              decoderOutput_356,decoderOutput_355,decoderOutput_354,
              decoderOutput_353,decoderOutput_352,decoderOutput_351,
              decoderOutput_350,decoderOutput_349,decoderOutput_348,
              decoderOutput_347,decoderOutput_346,decoderOutput_345,
              decoderOutput_344,decoderOutput_343,decoderOutput_342,
              decoderOutput_341,decoderOutput_340,decoderOutput_339,
              decoderOutput_338,decoderOutput_337,decoderOutput_336,
              decoderOutput_335,decoderOutput_334,decoderOutput_333,
              decoderOutput_332,decoderOutput_331,decoderOutput_330,
              decoderOutput_329,decoderOutput_328,decoderOutput_327,
              decoderOutput_326,decoderOutput_325,decoderOutput_324,
              decoderOutput_323,decoderOutput_322,decoderOutput_321,
              decoderOutput_320,decoderOutput_319,decoderOutput_318,
              decoderOutput_317,decoderOutput_316,decoderOutput_315,
              decoderOutput_314,decoderOutput_313,decoderOutput_312,
              decoderOutput_311,decoderOutput_310,decoderOutput_309,
              decoderOutput_308,decoderOutput_307,decoderOutput_306,
              decoderOutput_305,decoderOutput_304,decoderOutput_303,
              decoderOutput_302,decoderOutput_301,decoderOutput_300,
              decoderOutput_299,decoderOutput_298,decoderOutput_297,
              decoderOutput_296,decoderOutput_295,decoderOutput_294,
              decoderOutput_293,decoderOutput_292,decoderOutput_291,
              decoderOutput_290,decoderOutput_289,decoderOutput_288,
              decoderOutput_287,decoderOutput_286,decoderOutput_285,
              decoderOutput_284,decoderOutput_283,decoderOutput_282,
              decoderOutput_281,decoderOutput_280,decoderOutput_279,
              decoderOutput_278,decoderOutput_277,decoderOutput_276,
              decoderOutput_275,decoderOutput_274,decoderOutput_273,
              decoderOutput_272,decoderOutput_271,decoderOutput_270,
              decoderOutput_269,decoderOutput_268,decoderOutput_267,
              decoderOutput_266,decoderOutput_265,decoderOutput_264,
              decoderOutput_263,decoderOutput_262,decoderOutput_261,
              decoderOutput_260,decoderOutput_259,decoderOutput_258,
              decoderOutput_257,decoderOutput_256,decoderOutput_255,
              decoderOutput_254,decoderOutput_253,decoderOutput_252,
              decoderOutput_251,decoderOutput_250,decoderOutput_249,
              decoderOutput_248,decoderOutput_247,decoderOutput_246,
              decoderOutput_245,decoderOutput_244,decoderOutput_243,
              decoderOutput_242,decoderOutput_241,decoderOutput_240,
              decoderOutput_239,decoderOutput_238,decoderOutput_237,
              decoderOutput_236,decoderOutput_235,decoderOutput_234,
              decoderOutput_233,decoderOutput_232,decoderOutput_231,
              decoderOutput_230,decoderOutput_229,decoderOutput_228,
              decoderOutput_227,decoderOutput_226,decoderOutput_225,
              decoderOutput_224,decoderOutput_223,decoderOutput_222,
              decoderOutput_221,decoderOutput_220,decoderOutput_219,
              decoderOutput_218,decoderOutput_217,decoderOutput_216,
              decoderOutput_215,decoderOutput_214,decoderOutput_213,
              decoderOutput_212,decoderOutput_211,decoderOutput_210,
              decoderOutput_209,decoderOutput_208,decoderOutput_207,
              decoderOutput_206,decoderOutput_205,decoderOutput_204,
              decoderOutput_203,decoderOutput_202,decoderOutput_201,
              decoderOutput_200,decoderOutput_199,decoderOutput_198,
              decoderOutput_197,decoderOutput_196,decoderOutput_195,
              decoderOutput_194,decoderOutput_193,decoderOutput_192,
              decoderOutput_191,decoderOutput_190,decoderOutput_189,
              decoderOutput_188,decoderOutput_187,decoderOutput_186,
              decoderOutput_185,decoderOutput_184,decoderOutput_183,
              decoderOutput_182,decoderOutput_181,decoderOutput_180,
              decoderOutput_179,decoderOutput_178,decoderOutput_177,
              decoderOutput_176,decoderOutput_175,decoderOutput_174,
              decoderOutput_173,decoderOutput_172,decoderOutput_171,
              decoderOutput_170,decoderOutput_169,decoderOutput_168,
              decoderOutput_167,decoderOutput_166,decoderOutput_165,
              decoderOutput_164,decoderOutput_163,decoderOutput_162,
              decoderOutput_161,decoderOutput_160,decoderOutput_159,
              decoderOutput_158,decoderOutput_157,decoderOutput_156,
              decoderOutput_155,decoderOutput_154,decoderOutput_153,
              decoderOutput_152,decoderOutput_151,decoderOutput_150,
              decoderOutput_149,decoderOutput_148,decoderOutput_147,
              decoderOutput_146,decoderOutput_145,decoderOutput_144,
              decoderOutput_143,decoderOutput_142,decoderOutput_141,
              decoderOutput_140,decoderOutput_139,decoderOutput_138,
              decoderOutput_137,decoderOutput_136,decoderOutput_135,
              decoderOutput_134,decoderOutput_133,decoderOutput_132,
              decoderOutput_131,decoderOutput_130,decoderOutput_129,
              decoderOutput_128,decoderOutput_127,decoderOutput_126,
              decoderOutput_125,decoderOutput_124,decoderOutput_123,
              decoderOutput_122,decoderOutput_121,decoderOutput_120,
              decoderOutput_119,decoderOutput_118,decoderOutput_117,
              decoderOutput_116,decoderOutput_115,decoderOutput_114,
              decoderOutput_113,decoderOutput_112,decoderOutput_111,
              decoderOutput_110,decoderOutput_109,decoderOutput_108,
              decoderOutput_107,decoderOutput_106,decoderOutput_105,
              decoderOutput_104,decoderOutput_103,decoderOutput_102,
              decoderOutput_101,decoderOutput_100,decoderOutput_99,
              decoderOutput_98,decoderOutput_97,decoderOutput_96,
              decoderOutput_95,decoderOutput_94,decoderOutput_93,
              decoderOutput_92,decoderOutput_91,decoderOutput_90,
              decoderOutput_89,decoderOutput_88,decoderOutput_87,
              decoderOutput_86,decoderOutput_85,decoderOutput_84,
              decoderOutput_83,decoderOutput_82,decoderOutput_81,
              decoderOutput_80,decoderOutput_79,decoderOutput_78,
              decoderOutput_77,decoderOutput_76,decoderOutput_75,
              decoderOutput_74,decoderOutput_73,decoderOutput_72,
              decoderOutput_71,decoderOutput_70,decoderOutput_69,
              decoderOutput_68,decoderOutput_67,decoderOutput_66,
              decoderOutput_65,decoderOutput_64,decoderOutput_63,
              decoderOutput_62,decoderOutput_61,decoderOutput_60,
              decoderOutput_59,decoderOutput_58,decoderOutput_57,
              decoderOutput_56,decoderOutput_55,decoderOutput_54,
              decoderOutput_53,decoderOutput_52,decoderOutput_51,
              decoderOutput_50,decoderOutput_49,decoderOutput_48,
              decoderOutput_47,decoderOutput_46,decoderOutput_45,
              decoderOutput_44,decoderOutput_43,decoderOutput_42,
              decoderOutput_41,decoderOutput_40,decoderOutput_39,
              decoderOutput_38,decoderOutput_37,decoderOutput_36,
              decoderOutput_35,decoderOutput_34,decoderOutput_33,
              decoderOutput_32,decoderOutput_31,decoderOutput_30,
              decoderOutput_29,decoderOutput_28,decoderOutput_27,
              decoderOutput_26,decoderOutput_25,decoderOutput_24,
              decoderOutput_23,decoderOutput_22,decoderOutput_21,
              decoderOutput_20,decoderOutput_19,decoderOutput_18,
              decoderOutput_17,decoderOutput_16,decoderOutput_15,
              decoderOutput_14,decoderOutput_13,decoderOutput_12,
              decoderOutput_11,decoderOutput_10,decoderOutput_9,decoderOutput_8,
              decoderOutput_7,decoderOutput_6,decoderOutput_5,decoderOutput_4,
              decoderOutput_3,decoderOutput_2,decoderOutput_1,decoderOutput_0})
              ) ;
    Mux2_16 loop1_0_y (.A ({nx35885,nx36027,nx36169,nx36311,nx36453,nx36595,
            nx36737,nx36879,nx37021,nx37163,nx37305,nx37447,nx37589,nx37731,
            nx37873,nx38015}), .B ({nx33641,nx33779,nx33917,nx34055,nx34193,
            nx34331,nx34469,nx34611,nx34753,nx34895,nx35037,nx35179,nx35321,
            nx35463,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35605), .C ({inputRegisters_0__15,inputRegisters_0__14,
            inputRegisters_0__13,inputRegisters_0__12,inputRegisters_0__11,
            inputRegisters_0__10,inputRegisters_0__9,inputRegisters_0__8,
            inputRegisters_0__7,inputRegisters_0__6,inputRegisters_0__5,
            inputRegisters_0__4,inputRegisters_0__3,inputRegisters_0__2,
            inputRegisters_0__1,inputRegisters_0__0})) ;
    Reg_16 loop1_0_x (.D ({inputRegisters_0__15,inputRegisters_0__14,
           inputRegisters_0__13,inputRegisters_0__12,inputRegisters_0__11,
           inputRegisters_0__10,inputRegisters_0__9,inputRegisters_0__8,
           inputRegisters_0__7,inputRegisters_0__6,inputRegisters_0__5,
           inputRegisters_0__4,inputRegisters_0__3,inputRegisters_0__2,
           inputRegisters_0__1,inputRegisters_0__0}), .en (enableRegister_0), .clk (
           clk), .rst (resetRegisters), .Q ({registerOutputs_0__15,
           registerOutputs_0__14,registerOutputs_0__13,registerOutputs_0__12,
           registerOutputs_0__11,registerOutputs_0__10,registerOutputs_0__9,
           registerOutputs_0__8,registerOutputs_0__7,registerOutputs_0__6,
           registerOutputs_0__5,registerOutputs_0__4,registerOutputs_0__3,
           registerOutputs_0__2,registerOutputs_0__1,registerOutputs_0__0})) ;
    Mux2_16 loop1_1_y (.A ({nx35885,nx36027,nx36169,nx36311,nx36453,nx36595,
            nx36737,nx36879,nx37021,nx37163,nx37305,nx37447,nx37589,nx37731,
            nx37873,nx38015}), .B ({nx33641,nx33779,nx33917,nx34055,nx34193,
            nx34331,nx34471,nx34611,nx34753,nx34895,nx35037,nx35179,nx35321,
            nx35463,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35605), .C ({inputRegisters_1__15,inputRegisters_1__14,
            inputRegisters_1__13,inputRegisters_1__12,inputRegisters_1__11,
            inputRegisters_1__10,inputRegisters_1__9,inputRegisters_1__8,
            inputRegisters_1__7,inputRegisters_1__6,inputRegisters_1__5,
            inputRegisters_1__4,inputRegisters_1__3,inputRegisters_1__2,
            inputRegisters_1__1,inputRegisters_1__0})) ;
    Reg_16 loop1_1_x (.D ({inputRegisters_1__15,inputRegisters_1__14,
           inputRegisters_1__13,inputRegisters_1__12,inputRegisters_1__11,
           inputRegisters_1__10,inputRegisters_1__9,inputRegisters_1__8,
           inputRegisters_1__7,inputRegisters_1__6,inputRegisters_1__5,
           inputRegisters_1__4,inputRegisters_1__3,inputRegisters_1__2,
           inputRegisters_1__1,inputRegisters_1__0}), .en (enableRegister_1), .clk (
           clk), .rst (resetRegisters), .Q ({registerOutputs_1__15,
           registerOutputs_1__14,registerOutputs_1__13,registerOutputs_1__12,
           registerOutputs_1__11,registerOutputs_1__10,registerOutputs_1__9,
           registerOutputs_1__8,registerOutputs_1__7,registerOutputs_1__6,
           registerOutputs_1__5,registerOutputs_1__4,registerOutputs_1__3,
           registerOutputs_1__2,registerOutputs_1__1,registerOutputs_1__0})) ;
    Mux2_16 loop1_2_y (.A ({nx35885,nx36027,nx36169,nx36311,nx36453,nx36595,
            nx36737,nx36879,nx37021,nx37163,nx37305,nx37447,nx37589,nx37731,
            nx37873,nx38015}), .B ({nx33641,nx33779,nx33917,nx34055,nx34193,
            nx34333,nx34471,nx34611,nx34753,nx34895,nx35037,nx35179,nx35321,
            nx35463,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35605), .C ({inputRegisters_2__15,inputRegisters_2__14,
            inputRegisters_2__13,inputRegisters_2__12,inputRegisters_2__11,
            inputRegisters_2__10,inputRegisters_2__9,inputRegisters_2__8,
            inputRegisters_2__7,inputRegisters_2__6,inputRegisters_2__5,
            inputRegisters_2__4,inputRegisters_2__3,inputRegisters_2__2,
            inputRegisters_2__1,inputRegisters_2__0})) ;
    Reg_16 loop1_2_x (.D ({inputRegisters_2__15,inputRegisters_2__14,
           inputRegisters_2__13,inputRegisters_2__12,inputRegisters_2__11,
           inputRegisters_2__10,inputRegisters_2__9,inputRegisters_2__8,
           inputRegisters_2__7,inputRegisters_2__6,inputRegisters_2__5,
           inputRegisters_2__4,inputRegisters_2__3,inputRegisters_2__2,
           inputRegisters_2__1,inputRegisters_2__0}), .en (enableRegister_2), .clk (
           clk), .rst (resetRegisters), .Q ({registerOutputs_2__15,
           registerOutputs_2__14,registerOutputs_2__13,registerOutputs_2__12,
           registerOutputs_2__11,registerOutputs_2__10,registerOutputs_2__9,
           registerOutputs_2__8,registerOutputs_2__7,registerOutputs_2__6,
           registerOutputs_2__5,registerOutputs_2__4,registerOutputs_2__3,
           registerOutputs_2__2,registerOutputs_2__1,registerOutputs_2__0})) ;
    Mux2_16 loop1_3_y (.A ({nx35885,nx36027,nx36169,nx36311,nx36453,nx36595,
            nx36737,nx36879,nx37021,nx37163,nx37305,nx37447,nx37589,nx37731,
            nx37873,nx38015}), .B ({nx33641,nx33779,nx33917,nx34055,nx34195,
            nx34333,nx34471,nx34611,nx34753,nx34895,nx35037,nx35179,nx35321,
            nx35463,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35605), .C ({inputRegisters_3__15,inputRegisters_3__14,
            inputRegisters_3__13,inputRegisters_3__12,inputRegisters_3__11,
            inputRegisters_3__10,inputRegisters_3__9,inputRegisters_3__8,
            inputRegisters_3__7,inputRegisters_3__6,inputRegisters_3__5,
            inputRegisters_3__4,inputRegisters_3__3,inputRegisters_3__2,
            inputRegisters_3__1,inputRegisters_3__0})) ;
    Reg_16 loop1_3_x (.D ({inputRegisters_3__15,inputRegisters_3__14,
           inputRegisters_3__13,inputRegisters_3__12,inputRegisters_3__11,
           inputRegisters_3__10,inputRegisters_3__9,inputRegisters_3__8,
           inputRegisters_3__7,inputRegisters_3__6,inputRegisters_3__5,
           inputRegisters_3__4,inputRegisters_3__3,inputRegisters_3__2,
           inputRegisters_3__1,inputRegisters_3__0}), .en (enableRegister_3), .clk (
           clk), .rst (resetRegisters), .Q ({registerOutputs_3__15,
           registerOutputs_3__14,registerOutputs_3__13,registerOutputs_3__12,
           registerOutputs_3__11,registerOutputs_3__10,registerOutputs_3__9,
           registerOutputs_3__8,registerOutputs_3__7,registerOutputs_3__6,
           registerOutputs_3__5,registerOutputs_3__4,registerOutputs_3__3,
           registerOutputs_3__2,registerOutputs_3__1,registerOutputs_3__0})) ;
    Mux2_16 loop1_4_y (.A ({nx35885,nx36027,nx36169,nx36311,nx36453,nx36595,
            nx36737,nx36879,nx37021,nx37163,nx37305,nx37447,nx37589,nx37731,
            nx37873,nx38015}), .B ({nx33641,nx33779,nx33917,nx34057,nx34195,
            nx34333,nx34471,nx34611,nx34753,nx34895,nx35037,nx35179,nx35321,
            nx35463,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35605), .C ({inputRegisters_4__15,inputRegisters_4__14,
            inputRegisters_4__13,inputRegisters_4__12,inputRegisters_4__11,
            inputRegisters_4__10,inputRegisters_4__9,inputRegisters_4__8,
            inputRegisters_4__7,inputRegisters_4__6,inputRegisters_4__5,
            inputRegisters_4__4,inputRegisters_4__3,inputRegisters_4__2,
            inputRegisters_4__1,inputRegisters_4__0})) ;
    Reg_16 loop1_4_x (.D ({inputRegisters_4__15,inputRegisters_4__14,
           inputRegisters_4__13,inputRegisters_4__12,inputRegisters_4__11,
           inputRegisters_4__10,inputRegisters_4__9,inputRegisters_4__8,
           inputRegisters_4__7,inputRegisters_4__6,inputRegisters_4__5,
           inputRegisters_4__4,inputRegisters_4__3,inputRegisters_4__2,
           inputRegisters_4__1,inputRegisters_4__0}), .en (enableRegister_4), .clk (
           clk), .rst (resetRegisters), .Q ({registerOutputs_4__15,
           registerOutputs_4__14,registerOutputs_4__13,registerOutputs_4__12,
           registerOutputs_4__11,registerOutputs_4__10,registerOutputs_4__9,
           registerOutputs_4__8,registerOutputs_4__7,registerOutputs_4__6,
           registerOutputs_4__5,registerOutputs_4__4,registerOutputs_4__3,
           registerOutputs_4__2,registerOutputs_4__1,registerOutputs_4__0})) ;
    Mux2_16 loop1_5_y (.A ({nx35885,nx36027,nx36169,nx36311,nx36453,nx36595,
            nx36737,nx36879,nx37021,nx37163,nx37305,nx37447,nx37589,nx37731,
            nx37873,nx38015}), .B ({nx33641,nx33779,nx33919,nx34057,nx34195,
            nx34333,nx34471,nx34611,nx34753,nx34895,nx35037,nx35179,nx35321,
            nx35463,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35605), .C ({inputRegisters_5__15,inputRegisters_5__14,
            inputRegisters_5__13,inputRegisters_5__12,inputRegisters_5__11,
            inputRegisters_5__10,inputRegisters_5__9,inputRegisters_5__8,
            inputRegisters_5__7,inputRegisters_5__6,inputRegisters_5__5,
            inputRegisters_5__4,inputRegisters_5__3,inputRegisters_5__2,
            inputRegisters_5__1,inputRegisters_5__0})) ;
    Reg_16 loop1_5_x (.D ({inputRegisters_5__15,inputRegisters_5__14,
           inputRegisters_5__13,inputRegisters_5__12,inputRegisters_5__11,
           inputRegisters_5__10,inputRegisters_5__9,inputRegisters_5__8,
           inputRegisters_5__7,inputRegisters_5__6,inputRegisters_5__5,
           inputRegisters_5__4,inputRegisters_5__3,inputRegisters_5__2,
           inputRegisters_5__1,inputRegisters_5__0}), .en (enableRegister_5), .clk (
           clk), .rst (resetRegisters), .Q ({registerOutputs_5__15,
           registerOutputs_5__14,registerOutputs_5__13,registerOutputs_5__12,
           registerOutputs_5__11,registerOutputs_5__10,registerOutputs_5__9,
           registerOutputs_5__8,registerOutputs_5__7,registerOutputs_5__6,
           registerOutputs_5__5,registerOutputs_5__4,registerOutputs_5__3,
           registerOutputs_5__2,registerOutputs_5__1,registerOutputs_5__0})) ;
    Mux2_16 loop1_6_y (.A ({nx35885,nx36027,nx36169,nx36311,nx36453,nx36595,
            nx36737,nx36879,nx37021,nx37163,nx37305,nx37447,nx37589,nx37731,
            nx37873,nx38015}), .B ({nx33641,nx33781,nx33919,nx34057,nx34195,
            nx34333,nx34471,nx34611,nx34753,nx34895,nx35037,nx35179,nx35321,
            nx35463,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35605), .C ({inputRegisters_6__15,inputRegisters_6__14,
            inputRegisters_6__13,inputRegisters_6__12,inputRegisters_6__11,
            inputRegisters_6__10,inputRegisters_6__9,inputRegisters_6__8,
            inputRegisters_6__7,inputRegisters_6__6,inputRegisters_6__5,
            inputRegisters_6__4,inputRegisters_6__3,inputRegisters_6__2,
            inputRegisters_6__1,inputRegisters_6__0})) ;
    Reg_16 loop1_6_x (.D ({inputRegisters_6__15,inputRegisters_6__14,
           inputRegisters_6__13,inputRegisters_6__12,inputRegisters_6__11,
           inputRegisters_6__10,inputRegisters_6__9,inputRegisters_6__8,
           inputRegisters_6__7,inputRegisters_6__6,inputRegisters_6__5,
           inputRegisters_6__4,inputRegisters_6__3,inputRegisters_6__2,
           inputRegisters_6__1,inputRegisters_6__0}), .en (enableRegister_6), .clk (
           clk), .rst (resetRegisters), .Q ({registerOutputs_6__15,
           registerOutputs_6__14,registerOutputs_6__13,registerOutputs_6__12,
           registerOutputs_6__11,registerOutputs_6__10,registerOutputs_6__9,
           registerOutputs_6__8,registerOutputs_6__7,registerOutputs_6__6,
           registerOutputs_6__5,registerOutputs_6__4,registerOutputs_6__3,
           registerOutputs_6__2,registerOutputs_6__1,registerOutputs_6__0})) ;
    Mux2_16 loop1_7_y (.A ({nx35887,nx36029,nx36171,nx36313,nx36455,nx36597,
            nx36739,nx36881,nx37023,nx37165,nx37307,nx37449,nx37591,nx37733,
            nx37875,nx38017}), .B ({nx33643,nx33781,nx33919,nx34057,nx34195,
            nx34333,nx34471,nx34613,nx34755,nx34897,nx35039,nx35181,nx35323,
            nx35465,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35607), .C ({inputRegisters_7__15,inputRegisters_7__14,
            inputRegisters_7__13,inputRegisters_7__12,inputRegisters_7__11,
            inputRegisters_7__10,inputRegisters_7__9,inputRegisters_7__8,
            inputRegisters_7__7,inputRegisters_7__6,inputRegisters_7__5,
            inputRegisters_7__4,inputRegisters_7__3,inputRegisters_7__2,
            inputRegisters_7__1,inputRegisters_7__0})) ;
    Reg_16 loop1_7_x (.D ({inputRegisters_7__15,inputRegisters_7__14,
           inputRegisters_7__13,inputRegisters_7__12,inputRegisters_7__11,
           inputRegisters_7__10,inputRegisters_7__9,inputRegisters_7__8,
           inputRegisters_7__7,inputRegisters_7__6,inputRegisters_7__5,
           inputRegisters_7__4,inputRegisters_7__3,inputRegisters_7__2,
           inputRegisters_7__1,inputRegisters_7__0}), .en (enableRegister_7), .clk (
           clk), .rst (resetRegisters), .Q ({registerOutputs_7__15,
           registerOutputs_7__14,registerOutputs_7__13,registerOutputs_7__12,
           registerOutputs_7__11,registerOutputs_7__10,registerOutputs_7__9,
           registerOutputs_7__8,registerOutputs_7__7,registerOutputs_7__6,
           registerOutputs_7__5,registerOutputs_7__4,registerOutputs_7__3,
           registerOutputs_7__2,registerOutputs_7__1,registerOutputs_7__0})) ;
    Mux2_16 loop1_8_y (.A ({nx35887,nx36029,nx36171,nx36313,nx36455,nx36597,
            nx36739,nx36881,nx37023,nx37165,nx37307,nx37449,nx37591,nx37733,
            nx37875,nx38017}), .B ({nx33643,nx33781,nx33919,nx34057,nx34195,
            nx34333,nx34473,nx34613,nx34755,nx34897,nx35039,nx35181,nx35323,
            nx35465,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35607), .C ({inputRegisters_8__15,inputRegisters_8__14,
            inputRegisters_8__13,inputRegisters_8__12,inputRegisters_8__11,
            inputRegisters_8__10,inputRegisters_8__9,inputRegisters_8__8,
            inputRegisters_8__7,inputRegisters_8__6,inputRegisters_8__5,
            inputRegisters_8__4,inputRegisters_8__3,inputRegisters_8__2,
            inputRegisters_8__1,inputRegisters_8__0})) ;
    Reg_16 loop1_8_x (.D ({inputRegisters_8__15,inputRegisters_8__14,
           inputRegisters_8__13,inputRegisters_8__12,inputRegisters_8__11,
           inputRegisters_8__10,inputRegisters_8__9,inputRegisters_8__8,
           inputRegisters_8__7,inputRegisters_8__6,inputRegisters_8__5,
           inputRegisters_8__4,inputRegisters_8__3,inputRegisters_8__2,
           inputRegisters_8__1,inputRegisters_8__0}), .en (enableRegister_8), .clk (
           clk), .rst (resetRegisters), .Q ({registerOutputs_8__15,
           registerOutputs_8__14,registerOutputs_8__13,registerOutputs_8__12,
           registerOutputs_8__11,registerOutputs_8__10,registerOutputs_8__9,
           registerOutputs_8__8,registerOutputs_8__7,registerOutputs_8__6,
           registerOutputs_8__5,registerOutputs_8__4,registerOutputs_8__3,
           registerOutputs_8__2,registerOutputs_8__1,registerOutputs_8__0})) ;
    Mux2_16 loop1_9_y (.A ({nx35887,nx36029,nx36171,nx36313,nx36455,nx36597,
            nx36739,nx36881,nx37023,nx37165,nx37307,nx37449,nx37591,nx37733,
            nx37875,nx38017}), .B ({nx33643,nx33781,nx33919,nx34057,nx34195,
            nx34335,nx34473,nx34613,nx34755,nx34897,nx35039,nx35181,nx35323,
            nx35465,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35607), .C ({inputRegisters_9__15,inputRegisters_9__14,
            inputRegisters_9__13,inputRegisters_9__12,inputRegisters_9__11,
            inputRegisters_9__10,inputRegisters_9__9,inputRegisters_9__8,
            inputRegisters_9__7,inputRegisters_9__6,inputRegisters_9__5,
            inputRegisters_9__4,inputRegisters_9__3,inputRegisters_9__2,
            inputRegisters_9__1,inputRegisters_9__0})) ;
    Reg_16 loop1_9_x (.D ({inputRegisters_9__15,inputRegisters_9__14,
           inputRegisters_9__13,inputRegisters_9__12,inputRegisters_9__11,
           inputRegisters_9__10,inputRegisters_9__9,inputRegisters_9__8,
           inputRegisters_9__7,inputRegisters_9__6,inputRegisters_9__5,
           inputRegisters_9__4,inputRegisters_9__3,inputRegisters_9__2,
           inputRegisters_9__1,inputRegisters_9__0}), .en (enableRegister_9), .clk (
           clk), .rst (resetRegisters), .Q ({registerOutputs_9__15,
           registerOutputs_9__14,registerOutputs_9__13,registerOutputs_9__12,
           registerOutputs_9__11,registerOutputs_9__10,registerOutputs_9__9,
           registerOutputs_9__8,registerOutputs_9__7,registerOutputs_9__6,
           registerOutputs_9__5,registerOutputs_9__4,registerOutputs_9__3,
           registerOutputs_9__2,registerOutputs_9__1,registerOutputs_9__0})) ;
    Mux2_16 loop1_10_y (.A ({nx35887,nx36029,nx36171,nx36313,nx36455,nx36597,
            nx36739,nx36881,nx37023,nx37165,nx37307,nx37449,nx37591,nx37733,
            nx37875,nx38017}), .B ({nx33643,nx33781,nx33919,nx34057,nx34197,
            nx34335,nx34473,nx34613,nx34755,nx34897,nx35039,nx35181,nx35323,
            nx35465,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35607), .C ({inputRegisters_10__15,inputRegisters_10__14,
            inputRegisters_10__13,inputRegisters_10__12,inputRegisters_10__11,
            inputRegisters_10__10,inputRegisters_10__9,inputRegisters_10__8,
            inputRegisters_10__7,inputRegisters_10__6,inputRegisters_10__5,
            inputRegisters_10__4,inputRegisters_10__3,inputRegisters_10__2,
            inputRegisters_10__1,inputRegisters_10__0})) ;
    Reg_16 loop1_10_x (.D ({inputRegisters_10__15,inputRegisters_10__14,
           inputRegisters_10__13,inputRegisters_10__12,inputRegisters_10__11,
           inputRegisters_10__10,inputRegisters_10__9,inputRegisters_10__8,
           inputRegisters_10__7,inputRegisters_10__6,inputRegisters_10__5,
           inputRegisters_10__4,inputRegisters_10__3,inputRegisters_10__2,
           inputRegisters_10__1,inputRegisters_10__0}), .en (enableRegister_10)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_10__15,
           registerOutputs_10__14,registerOutputs_10__13,registerOutputs_10__12,
           registerOutputs_10__11,registerOutputs_10__10,registerOutputs_10__9,
           registerOutputs_10__8,registerOutputs_10__7,registerOutputs_10__6,
           registerOutputs_10__5,registerOutputs_10__4,registerOutputs_10__3,
           registerOutputs_10__2,registerOutputs_10__1,registerOutputs_10__0})
           ) ;
    Mux2_16 loop1_11_y (.A ({nx35887,nx36029,nx36171,nx36313,nx36455,nx36597,
            nx36739,nx36881,nx37023,nx37165,nx37307,nx37449,nx37591,nx37733,
            nx37875,nx38017}), .B ({nx33643,nx33781,nx33919,nx34059,nx34197,
            nx34335,nx34473,nx34613,nx34755,nx34897,nx35039,nx35181,nx35323,
            nx35465,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35607), .C ({inputRegisters_11__15,inputRegisters_11__14,
            inputRegisters_11__13,inputRegisters_11__12,inputRegisters_11__11,
            inputRegisters_11__10,inputRegisters_11__9,inputRegisters_11__8,
            inputRegisters_11__7,inputRegisters_11__6,inputRegisters_11__5,
            inputRegisters_11__4,inputRegisters_11__3,inputRegisters_11__2,
            inputRegisters_11__1,inputRegisters_11__0})) ;
    Reg_16 loop1_11_x (.D ({inputRegisters_11__15,inputRegisters_11__14,
           inputRegisters_11__13,inputRegisters_11__12,inputRegisters_11__11,
           inputRegisters_11__10,inputRegisters_11__9,inputRegisters_11__8,
           inputRegisters_11__7,inputRegisters_11__6,inputRegisters_11__5,
           inputRegisters_11__4,inputRegisters_11__3,inputRegisters_11__2,
           inputRegisters_11__1,inputRegisters_11__0}), .en (enableRegister_11)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_11__15,
           registerOutputs_11__14,registerOutputs_11__13,registerOutputs_11__12,
           registerOutputs_11__11,registerOutputs_11__10,registerOutputs_11__9,
           registerOutputs_11__8,registerOutputs_11__7,registerOutputs_11__6,
           registerOutputs_11__5,registerOutputs_11__4,registerOutputs_11__3,
           registerOutputs_11__2,registerOutputs_11__1,registerOutputs_11__0})
           ) ;
    Mux2_16 loop1_12_y (.A ({nx35887,nx36029,nx36171,nx36313,nx36455,nx36597,
            nx36739,nx36881,nx37023,nx37165,nx37307,nx37449,nx37591,nx37733,
            nx37875,nx38017}), .B ({nx33643,nx33781,nx33921,nx34059,nx34197,
            nx34335,nx34473,nx34613,nx34755,nx34897,nx35039,nx35181,nx35323,
            nx35465,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35607), .C ({inputRegisters_12__15,inputRegisters_12__14,
            inputRegisters_12__13,inputRegisters_12__12,inputRegisters_12__11,
            inputRegisters_12__10,inputRegisters_12__9,inputRegisters_12__8,
            inputRegisters_12__7,inputRegisters_12__6,inputRegisters_12__5,
            inputRegisters_12__4,inputRegisters_12__3,inputRegisters_12__2,
            inputRegisters_12__1,inputRegisters_12__0})) ;
    Reg_16 loop1_12_x (.D ({inputRegisters_12__15,inputRegisters_12__14,
           inputRegisters_12__13,inputRegisters_12__12,inputRegisters_12__11,
           inputRegisters_12__10,inputRegisters_12__9,inputRegisters_12__8,
           inputRegisters_12__7,inputRegisters_12__6,inputRegisters_12__5,
           inputRegisters_12__4,inputRegisters_12__3,inputRegisters_12__2,
           inputRegisters_12__1,inputRegisters_12__0}), .en (enableRegister_12)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_12__15,
           registerOutputs_12__14,registerOutputs_12__13,registerOutputs_12__12,
           registerOutputs_12__11,registerOutputs_12__10,registerOutputs_12__9,
           registerOutputs_12__8,registerOutputs_12__7,registerOutputs_12__6,
           registerOutputs_12__5,registerOutputs_12__4,registerOutputs_12__3,
           registerOutputs_12__2,registerOutputs_12__1,registerOutputs_12__0})
           ) ;
    Mux2_16 loop1_13_y (.A ({nx35887,nx36029,nx36171,nx36313,nx36455,nx36597,
            nx36739,nx36881,nx37023,nx37165,nx37307,nx37449,nx37591,nx37733,
            nx37875,nx38017}), .B ({nx33643,nx33783,nx33921,nx34059,nx34197,
            nx34335,nx34473,nx34613,nx34755,nx34897,nx35039,nx35181,nx35323,
            nx35465,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35607), .C ({inputRegisters_13__15,inputRegisters_13__14,
            inputRegisters_13__13,inputRegisters_13__12,inputRegisters_13__11,
            inputRegisters_13__10,inputRegisters_13__9,inputRegisters_13__8,
            inputRegisters_13__7,inputRegisters_13__6,inputRegisters_13__5,
            inputRegisters_13__4,inputRegisters_13__3,inputRegisters_13__2,
            inputRegisters_13__1,inputRegisters_13__0})) ;
    Reg_16 loop1_13_x (.D ({inputRegisters_13__15,inputRegisters_13__14,
           inputRegisters_13__13,inputRegisters_13__12,inputRegisters_13__11,
           inputRegisters_13__10,inputRegisters_13__9,inputRegisters_13__8,
           inputRegisters_13__7,inputRegisters_13__6,inputRegisters_13__5,
           inputRegisters_13__4,inputRegisters_13__3,inputRegisters_13__2,
           inputRegisters_13__1,inputRegisters_13__0}), .en (enableRegister_13)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_13__15,
           registerOutputs_13__14,registerOutputs_13__13,registerOutputs_13__12,
           registerOutputs_13__11,registerOutputs_13__10,registerOutputs_13__9,
           registerOutputs_13__8,registerOutputs_13__7,registerOutputs_13__6,
           registerOutputs_13__5,registerOutputs_13__4,registerOutputs_13__3,
           registerOutputs_13__2,registerOutputs_13__1,registerOutputs_13__0})
           ) ;
    Mux2_16 loop1_14_y (.A ({nx35889,nx36031,nx36173,nx36315,nx36457,nx36599,
            nx36741,nx36883,nx37025,nx37167,nx37309,nx37451,nx37593,nx37735,
            nx37877,nx38019}), .B ({nx33645,nx33783,nx33921,nx34059,nx34197,
            nx34335,nx34473,nx34615,nx34757,nx34899,nx35041,nx35183,nx35325,
            nx35467,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35609), .C ({inputRegisters_14__15,inputRegisters_14__14,
            inputRegisters_14__13,inputRegisters_14__12,inputRegisters_14__11,
            inputRegisters_14__10,inputRegisters_14__9,inputRegisters_14__8,
            inputRegisters_14__7,inputRegisters_14__6,inputRegisters_14__5,
            inputRegisters_14__4,inputRegisters_14__3,inputRegisters_14__2,
            inputRegisters_14__1,inputRegisters_14__0})) ;
    Reg_16 loop1_14_x (.D ({inputRegisters_14__15,inputRegisters_14__14,
           inputRegisters_14__13,inputRegisters_14__12,inputRegisters_14__11,
           inputRegisters_14__10,inputRegisters_14__9,inputRegisters_14__8,
           inputRegisters_14__7,inputRegisters_14__6,inputRegisters_14__5,
           inputRegisters_14__4,inputRegisters_14__3,inputRegisters_14__2,
           inputRegisters_14__1,inputRegisters_14__0}), .en (enableRegister_14)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_14__15,
           registerOutputs_14__14,registerOutputs_14__13,registerOutputs_14__12,
           registerOutputs_14__11,registerOutputs_14__10,registerOutputs_14__9,
           registerOutputs_14__8,registerOutputs_14__7,registerOutputs_14__6,
           registerOutputs_14__5,registerOutputs_14__4,registerOutputs_14__3,
           registerOutputs_14__2,registerOutputs_14__1,registerOutputs_14__0})
           ) ;
    Mux2_16 loop1_15_y (.A ({nx35889,nx36031,nx36173,nx36315,nx36457,nx36599,
            nx36741,nx36883,nx37025,nx37167,nx37309,nx37451,nx37593,nx37735,
            nx37877,nx38019}), .B ({nx33645,nx33783,nx33921,nx34059,nx34197,
            nx34335,nx34475,nx34615,nx34757,nx34899,nx35041,nx35183,nx35325,
            nx35467,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35609), .C ({inputRegisters_15__15,inputRegisters_15__14,
            inputRegisters_15__13,inputRegisters_15__12,inputRegisters_15__11,
            inputRegisters_15__10,inputRegisters_15__9,inputRegisters_15__8,
            inputRegisters_15__7,inputRegisters_15__6,inputRegisters_15__5,
            inputRegisters_15__4,inputRegisters_15__3,inputRegisters_15__2,
            inputRegisters_15__1,inputRegisters_15__0})) ;
    Reg_16 loop1_15_x (.D ({inputRegisters_15__15,inputRegisters_15__14,
           inputRegisters_15__13,inputRegisters_15__12,inputRegisters_15__11,
           inputRegisters_15__10,inputRegisters_15__9,inputRegisters_15__8,
           inputRegisters_15__7,inputRegisters_15__6,inputRegisters_15__5,
           inputRegisters_15__4,inputRegisters_15__3,inputRegisters_15__2,
           inputRegisters_15__1,inputRegisters_15__0}), .en (enableRegister_15)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_15__15,
           registerOutputs_15__14,registerOutputs_15__13,registerOutputs_15__12,
           registerOutputs_15__11,registerOutputs_15__10,registerOutputs_15__9,
           registerOutputs_15__8,registerOutputs_15__7,registerOutputs_15__6,
           registerOutputs_15__5,registerOutputs_15__4,registerOutputs_15__3,
           registerOutputs_15__2,registerOutputs_15__1,registerOutputs_15__0})
           ) ;
    Mux2_16 loop1_16_y (.A ({nx35889,nx36031,nx36173,nx36315,nx36457,nx36599,
            nx36741,nx36883,nx37025,nx37167,nx37309,nx37451,nx37593,nx37735,
            nx37877,nx38019}), .B ({nx33645,nx33783,nx33921,nx34059,nx34197,
            nx34337,nx34475,nx34615,nx34757,nx34899,nx35041,nx35183,nx35325,
            nx35467,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35609), .C ({inputRegisters_16__15,inputRegisters_16__14,
            inputRegisters_16__13,inputRegisters_16__12,inputRegisters_16__11,
            inputRegisters_16__10,inputRegisters_16__9,inputRegisters_16__8,
            inputRegisters_16__7,inputRegisters_16__6,inputRegisters_16__5,
            inputRegisters_16__4,inputRegisters_16__3,inputRegisters_16__2,
            inputRegisters_16__1,inputRegisters_16__0})) ;
    Reg_16 loop1_16_x (.D ({inputRegisters_16__15,inputRegisters_16__14,
           inputRegisters_16__13,inputRegisters_16__12,inputRegisters_16__11,
           inputRegisters_16__10,inputRegisters_16__9,inputRegisters_16__8,
           inputRegisters_16__7,inputRegisters_16__6,inputRegisters_16__5,
           inputRegisters_16__4,inputRegisters_16__3,inputRegisters_16__2,
           inputRegisters_16__1,inputRegisters_16__0}), .en (enableRegister_16)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_16__15,
           registerOutputs_16__14,registerOutputs_16__13,registerOutputs_16__12,
           registerOutputs_16__11,registerOutputs_16__10,registerOutputs_16__9,
           registerOutputs_16__8,registerOutputs_16__7,registerOutputs_16__6,
           registerOutputs_16__5,registerOutputs_16__4,registerOutputs_16__3,
           registerOutputs_16__2,registerOutputs_16__1,registerOutputs_16__0})
           ) ;
    Mux2_16 loop1_17_y (.A ({nx35889,nx36031,nx36173,nx36315,nx36457,nx36599,
            nx36741,nx36883,nx37025,nx37167,nx37309,nx37451,nx37593,nx37735,
            nx37877,nx38019}), .B ({nx33645,nx33783,nx33921,nx34059,nx34199,
            nx34337,nx34475,nx34615,nx34757,nx34899,nx35041,nx35183,nx35325,
            nx35467,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35609), .C ({inputRegisters_17__15,inputRegisters_17__14,
            inputRegisters_17__13,inputRegisters_17__12,inputRegisters_17__11,
            inputRegisters_17__10,inputRegisters_17__9,inputRegisters_17__8,
            inputRegisters_17__7,inputRegisters_17__6,inputRegisters_17__5,
            inputRegisters_17__4,inputRegisters_17__3,inputRegisters_17__2,
            inputRegisters_17__1,inputRegisters_17__0})) ;
    Reg_16 loop1_17_x (.D ({inputRegisters_17__15,inputRegisters_17__14,
           inputRegisters_17__13,inputRegisters_17__12,inputRegisters_17__11,
           inputRegisters_17__10,inputRegisters_17__9,inputRegisters_17__8,
           inputRegisters_17__7,inputRegisters_17__6,inputRegisters_17__5,
           inputRegisters_17__4,inputRegisters_17__3,inputRegisters_17__2,
           inputRegisters_17__1,inputRegisters_17__0}), .en (enableRegister_17)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_17__15,
           registerOutputs_17__14,registerOutputs_17__13,registerOutputs_17__12,
           registerOutputs_17__11,registerOutputs_17__10,registerOutputs_17__9,
           registerOutputs_17__8,registerOutputs_17__7,registerOutputs_17__6,
           registerOutputs_17__5,registerOutputs_17__4,registerOutputs_17__3,
           registerOutputs_17__2,registerOutputs_17__1,registerOutputs_17__0})
           ) ;
    Mux2_16 loop1_18_y (.A ({nx35889,nx36031,nx36173,nx36315,nx36457,nx36599,
            nx36741,nx36883,nx37025,nx37167,nx37309,nx37451,nx37593,nx37735,
            nx37877,nx38019}), .B ({nx33645,nx33783,nx33921,nx34061,nx34199,
            nx34337,nx34475,nx34615,nx34757,nx34899,nx35041,nx35183,nx35325,
            nx35467,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35609), .C ({inputRegisters_18__15,inputRegisters_18__14,
            inputRegisters_18__13,inputRegisters_18__12,inputRegisters_18__11,
            inputRegisters_18__10,inputRegisters_18__9,inputRegisters_18__8,
            inputRegisters_18__7,inputRegisters_18__6,inputRegisters_18__5,
            inputRegisters_18__4,inputRegisters_18__3,inputRegisters_18__2,
            inputRegisters_18__1,inputRegisters_18__0})) ;
    Reg_16 loop1_18_x (.D ({inputRegisters_18__15,inputRegisters_18__14,
           inputRegisters_18__13,inputRegisters_18__12,inputRegisters_18__11,
           inputRegisters_18__10,inputRegisters_18__9,inputRegisters_18__8,
           inputRegisters_18__7,inputRegisters_18__6,inputRegisters_18__5,
           inputRegisters_18__4,inputRegisters_18__3,inputRegisters_18__2,
           inputRegisters_18__1,inputRegisters_18__0}), .en (enableRegister_18)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_18__15,
           registerOutputs_18__14,registerOutputs_18__13,registerOutputs_18__12,
           registerOutputs_18__11,registerOutputs_18__10,registerOutputs_18__9,
           registerOutputs_18__8,registerOutputs_18__7,registerOutputs_18__6,
           registerOutputs_18__5,registerOutputs_18__4,registerOutputs_18__3,
           registerOutputs_18__2,registerOutputs_18__1,registerOutputs_18__0})
           ) ;
    Mux2_16 loop1_19_y (.A ({nx35889,nx36031,nx36173,nx36315,nx36457,nx36599,
            nx36741,nx36883,nx37025,nx37167,nx37309,nx37451,nx37593,nx37735,
            nx37877,nx38019}), .B ({nx33645,nx33783,nx33923,nx34061,nx34199,
            nx34337,nx34475,nx34615,nx34757,nx34899,nx35041,nx35183,nx35325,
            nx35467,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35609), .C ({inputRegisters_19__15,inputRegisters_19__14,
            inputRegisters_19__13,inputRegisters_19__12,inputRegisters_19__11,
            inputRegisters_19__10,inputRegisters_19__9,inputRegisters_19__8,
            inputRegisters_19__7,inputRegisters_19__6,inputRegisters_19__5,
            inputRegisters_19__4,inputRegisters_19__3,inputRegisters_19__2,
            inputRegisters_19__1,inputRegisters_19__0})) ;
    Reg_16 loop1_19_x (.D ({inputRegisters_19__15,inputRegisters_19__14,
           inputRegisters_19__13,inputRegisters_19__12,inputRegisters_19__11,
           inputRegisters_19__10,inputRegisters_19__9,inputRegisters_19__8,
           inputRegisters_19__7,inputRegisters_19__6,inputRegisters_19__5,
           inputRegisters_19__4,inputRegisters_19__3,inputRegisters_19__2,
           inputRegisters_19__1,inputRegisters_19__0}), .en (enableRegister_19)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_19__15,
           registerOutputs_19__14,registerOutputs_19__13,registerOutputs_19__12,
           registerOutputs_19__11,registerOutputs_19__10,registerOutputs_19__9,
           registerOutputs_19__8,registerOutputs_19__7,registerOutputs_19__6,
           registerOutputs_19__5,registerOutputs_19__4,registerOutputs_19__3,
           registerOutputs_19__2,registerOutputs_19__1,registerOutputs_19__0})
           ) ;
    Mux2_16 loop1_20_y (.A ({nx35889,nx36031,nx36173,nx36315,nx36457,nx36599,
            nx36741,nx36883,nx37025,nx37167,nx37309,nx37451,nx37593,nx37735,
            nx37877,nx38019}), .B ({nx33645,nx33785,nx33923,nx34061,nx34199,
            nx34337,nx34475,nx34615,nx34757,nx34899,nx35041,nx35183,nx35325,
            nx35467,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35609), .C ({inputRegisters_20__15,inputRegisters_20__14,
            inputRegisters_20__13,inputRegisters_20__12,inputRegisters_20__11,
            inputRegisters_20__10,inputRegisters_20__9,inputRegisters_20__8,
            inputRegisters_20__7,inputRegisters_20__6,inputRegisters_20__5,
            inputRegisters_20__4,inputRegisters_20__3,inputRegisters_20__2,
            inputRegisters_20__1,inputRegisters_20__0})) ;
    Reg_16 loop1_20_x (.D ({inputRegisters_20__15,inputRegisters_20__14,
           inputRegisters_20__13,inputRegisters_20__12,inputRegisters_20__11,
           inputRegisters_20__10,inputRegisters_20__9,inputRegisters_20__8,
           inputRegisters_20__7,inputRegisters_20__6,inputRegisters_20__5,
           inputRegisters_20__4,inputRegisters_20__3,inputRegisters_20__2,
           inputRegisters_20__1,inputRegisters_20__0}), .en (enableRegister_20)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_20__15,
           registerOutputs_20__14,registerOutputs_20__13,registerOutputs_20__12,
           registerOutputs_20__11,registerOutputs_20__10,registerOutputs_20__9,
           registerOutputs_20__8,registerOutputs_20__7,registerOutputs_20__6,
           registerOutputs_20__5,registerOutputs_20__4,registerOutputs_20__3,
           registerOutputs_20__2,registerOutputs_20__1,registerOutputs_20__0})
           ) ;
    Mux2_16 loop1_21_y (.A ({nx35891,nx36033,nx36175,nx36317,nx36459,nx36601,
            nx36743,nx36885,nx37027,nx37169,nx37311,nx37453,nx37595,nx37737,
            nx37879,nx38021}), .B ({nx33647,nx33785,nx33923,nx34061,nx34199,
            nx34337,nx34475,nx34617,nx34759,nx34901,nx35043,nx35185,nx35327,
            nx35469,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35611), .C ({inputRegisters_21__15,inputRegisters_21__14,
            inputRegisters_21__13,inputRegisters_21__12,inputRegisters_21__11,
            inputRegisters_21__10,inputRegisters_21__9,inputRegisters_21__8,
            inputRegisters_21__7,inputRegisters_21__6,inputRegisters_21__5,
            inputRegisters_21__4,inputRegisters_21__3,inputRegisters_21__2,
            inputRegisters_21__1,inputRegisters_21__0})) ;
    Reg_16 loop1_21_x (.D ({inputRegisters_21__15,inputRegisters_21__14,
           inputRegisters_21__13,inputRegisters_21__12,inputRegisters_21__11,
           inputRegisters_21__10,inputRegisters_21__9,inputRegisters_21__8,
           inputRegisters_21__7,inputRegisters_21__6,inputRegisters_21__5,
           inputRegisters_21__4,inputRegisters_21__3,inputRegisters_21__2,
           inputRegisters_21__1,inputRegisters_21__0}), .en (enableRegister_21)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_21__15,
           registerOutputs_21__14,registerOutputs_21__13,registerOutputs_21__12,
           registerOutputs_21__11,registerOutputs_21__10,registerOutputs_21__9,
           registerOutputs_21__8,registerOutputs_21__7,registerOutputs_21__6,
           registerOutputs_21__5,registerOutputs_21__4,registerOutputs_21__3,
           registerOutputs_21__2,registerOutputs_21__1,registerOutputs_21__0})
           ) ;
    Mux2_16 loop1_22_y (.A ({nx35891,nx36033,nx36175,nx36317,nx36459,nx36601,
            nx36743,nx36885,nx37027,nx37169,nx37311,nx37453,nx37595,nx37737,
            nx37879,nx38021}), .B ({nx33647,nx33785,nx33923,nx34061,nx34199,
            nx34337,nx34477,nx34617,nx34759,nx34901,nx35043,nx35185,nx35327,
            nx35469,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35611), .C ({inputRegisters_22__15,inputRegisters_22__14,
            inputRegisters_22__13,inputRegisters_22__12,inputRegisters_22__11,
            inputRegisters_22__10,inputRegisters_22__9,inputRegisters_22__8,
            inputRegisters_22__7,inputRegisters_22__6,inputRegisters_22__5,
            inputRegisters_22__4,inputRegisters_22__3,inputRegisters_22__2,
            inputRegisters_22__1,inputRegisters_22__0})) ;
    Reg_16 loop1_22_x (.D ({inputRegisters_22__15,inputRegisters_22__14,
           inputRegisters_22__13,inputRegisters_22__12,inputRegisters_22__11,
           inputRegisters_22__10,inputRegisters_22__9,inputRegisters_22__8,
           inputRegisters_22__7,inputRegisters_22__6,inputRegisters_22__5,
           inputRegisters_22__4,inputRegisters_22__3,inputRegisters_22__2,
           inputRegisters_22__1,inputRegisters_22__0}), .en (enableRegister_22)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_22__15,
           registerOutputs_22__14,registerOutputs_22__13,registerOutputs_22__12,
           registerOutputs_22__11,registerOutputs_22__10,registerOutputs_22__9,
           registerOutputs_22__8,registerOutputs_22__7,registerOutputs_22__6,
           registerOutputs_22__5,registerOutputs_22__4,registerOutputs_22__3,
           registerOutputs_22__2,registerOutputs_22__1,registerOutputs_22__0})
           ) ;
    Mux2_16 loop1_23_y (.A ({nx35891,nx36033,nx36175,nx36317,nx36459,nx36601,
            nx36743,nx36885,nx37027,nx37169,nx37311,nx37453,nx37595,nx37737,
            nx37879,nx38021}), .B ({nx33647,nx33785,nx33923,nx34061,nx34199,
            nx34339,nx34477,nx34617,nx34759,nx34901,nx35043,nx35185,nx35327,
            nx35469,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35611), .C ({inputRegisters_23__15,inputRegisters_23__14,
            inputRegisters_23__13,inputRegisters_23__12,inputRegisters_23__11,
            inputRegisters_23__10,inputRegisters_23__9,inputRegisters_23__8,
            inputRegisters_23__7,inputRegisters_23__6,inputRegisters_23__5,
            inputRegisters_23__4,inputRegisters_23__3,inputRegisters_23__2,
            inputRegisters_23__1,inputRegisters_23__0})) ;
    Reg_16 loop1_23_x (.D ({inputRegisters_23__15,inputRegisters_23__14,
           inputRegisters_23__13,inputRegisters_23__12,inputRegisters_23__11,
           inputRegisters_23__10,inputRegisters_23__9,inputRegisters_23__8,
           inputRegisters_23__7,inputRegisters_23__6,inputRegisters_23__5,
           inputRegisters_23__4,inputRegisters_23__3,inputRegisters_23__2,
           inputRegisters_23__1,inputRegisters_23__0}), .en (enableRegister_23)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_23__15,
           registerOutputs_23__14,registerOutputs_23__13,registerOutputs_23__12,
           registerOutputs_23__11,registerOutputs_23__10,registerOutputs_23__9,
           registerOutputs_23__8,registerOutputs_23__7,registerOutputs_23__6,
           registerOutputs_23__5,registerOutputs_23__4,registerOutputs_23__3,
           registerOutputs_23__2,registerOutputs_23__1,registerOutputs_23__0})
           ) ;
    Mux2_16 loop1_24_y (.A ({nx35891,nx36033,nx36175,nx36317,nx36459,nx36601,
            nx36743,nx36885,nx37027,nx37169,nx37311,nx37453,nx37595,nx37737,
            nx37879,nx38021}), .B ({nx33647,nx33785,nx33923,nx34061,nx34201,
            nx34339,nx34477,nx34617,nx34759,nx34901,nx35043,nx35185,nx35327,
            nx35469,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35611), .C ({inputRegisters_24__15,inputRegisters_24__14,
            inputRegisters_24__13,inputRegisters_24__12,inputRegisters_24__11,
            inputRegisters_24__10,inputRegisters_24__9,inputRegisters_24__8,
            inputRegisters_24__7,inputRegisters_24__6,inputRegisters_24__5,
            inputRegisters_24__4,inputRegisters_24__3,inputRegisters_24__2,
            inputRegisters_24__1,inputRegisters_24__0})) ;
    Reg_16 loop1_24_x (.D ({inputRegisters_24__15,inputRegisters_24__14,
           inputRegisters_24__13,inputRegisters_24__12,inputRegisters_24__11,
           inputRegisters_24__10,inputRegisters_24__9,inputRegisters_24__8,
           inputRegisters_24__7,inputRegisters_24__6,inputRegisters_24__5,
           inputRegisters_24__4,inputRegisters_24__3,inputRegisters_24__2,
           inputRegisters_24__1,inputRegisters_24__0}), .en (enableRegister_24)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_24__15,
           registerOutputs_24__14,registerOutputs_24__13,registerOutputs_24__12,
           registerOutputs_24__11,registerOutputs_24__10,registerOutputs_24__9,
           registerOutputs_24__8,registerOutputs_24__7,registerOutputs_24__6,
           registerOutputs_24__5,registerOutputs_24__4,registerOutputs_24__3,
           registerOutputs_24__2,registerOutputs_24__1,registerOutputs_24__0})
           ) ;
    Mux2_16 loop1_25_y (.A ({nx35891,nx36033,nx36175,nx36317,nx36459,nx36601,
            nx36743,nx36885,nx37027,nx37169,nx37311,nx37453,nx37595,nx37737,
            nx37879,nx38021}), .B ({nx33647,nx33785,nx33923,nx34063,nx34201,
            nx34339,nx34477,nx34617,nx34759,nx34901,nx35043,nx35185,nx35327,
            nx35469,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35611), .C ({inputRegisters_25__15,inputRegisters_25__14,
            inputRegisters_25__13,inputRegisters_25__12,inputRegisters_25__11,
            inputRegisters_25__10,inputRegisters_25__9,inputRegisters_25__8,
            inputRegisters_25__7,inputRegisters_25__6,inputRegisters_25__5,
            inputRegisters_25__4,inputRegisters_25__3,inputRegisters_25__2,
            inputRegisters_25__1,inputRegisters_25__0})) ;
    Reg_16 loop1_25_x (.D ({inputRegisters_25__15,inputRegisters_25__14,
           inputRegisters_25__13,inputRegisters_25__12,inputRegisters_25__11,
           inputRegisters_25__10,inputRegisters_25__9,inputRegisters_25__8,
           inputRegisters_25__7,inputRegisters_25__6,inputRegisters_25__5,
           inputRegisters_25__4,inputRegisters_25__3,inputRegisters_25__2,
           inputRegisters_25__1,inputRegisters_25__0}), .en (enableRegister_25)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_25__15,
           registerOutputs_25__14,registerOutputs_25__13,registerOutputs_25__12,
           registerOutputs_25__11,registerOutputs_25__10,registerOutputs_25__9,
           registerOutputs_25__8,registerOutputs_25__7,registerOutputs_25__6,
           registerOutputs_25__5,registerOutputs_25__4,registerOutputs_25__3,
           registerOutputs_25__2,registerOutputs_25__1,registerOutputs_25__0})
           ) ;
    Mux2_16 loop1_26_y (.A ({nx35891,nx36033,nx36175,nx36317,nx36459,nx36601,
            nx36743,nx36885,nx37027,nx37169,nx37311,nx37453,nx37595,nx37737,
            nx37879,nx38021}), .B ({nx33647,nx33785,nx33925,nx34063,nx34201,
            nx34339,nx34477,nx34617,nx34759,nx34901,nx35043,nx35185,nx35327,
            nx35469,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35611), .C ({inputRegisters_26__15,inputRegisters_26__14,
            inputRegisters_26__13,inputRegisters_26__12,inputRegisters_26__11,
            inputRegisters_26__10,inputRegisters_26__9,inputRegisters_26__8,
            inputRegisters_26__7,inputRegisters_26__6,inputRegisters_26__5,
            inputRegisters_26__4,inputRegisters_26__3,inputRegisters_26__2,
            inputRegisters_26__1,inputRegisters_26__0})) ;
    Reg_16 loop1_26_x (.D ({inputRegisters_26__15,inputRegisters_26__14,
           inputRegisters_26__13,inputRegisters_26__12,inputRegisters_26__11,
           inputRegisters_26__10,inputRegisters_26__9,inputRegisters_26__8,
           inputRegisters_26__7,inputRegisters_26__6,inputRegisters_26__5,
           inputRegisters_26__4,inputRegisters_26__3,inputRegisters_26__2,
           inputRegisters_26__1,inputRegisters_26__0}), .en (enableRegister_26)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_26__15,
           registerOutputs_26__14,registerOutputs_26__13,registerOutputs_26__12,
           registerOutputs_26__11,registerOutputs_26__10,registerOutputs_26__9,
           registerOutputs_26__8,registerOutputs_26__7,registerOutputs_26__6,
           registerOutputs_26__5,registerOutputs_26__4,registerOutputs_26__3,
           registerOutputs_26__2,registerOutputs_26__1,registerOutputs_26__0})
           ) ;
    Mux2_16 loop1_27_y (.A ({nx35891,nx36033,nx36175,nx36317,nx36459,nx36601,
            nx36743,nx36885,nx37027,nx37169,nx37311,nx37453,nx37595,nx37737,
            nx37879,nx38021}), .B ({nx33647,nx33787,nx33925,nx34063,nx34201,
            nx34339,nx34477,nx34617,nx34759,nx34901,nx35043,nx35185,nx35327,
            nx35469,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35611), .C ({inputRegisters_27__15,inputRegisters_27__14,
            inputRegisters_27__13,inputRegisters_27__12,inputRegisters_27__11,
            inputRegisters_27__10,inputRegisters_27__9,inputRegisters_27__8,
            inputRegisters_27__7,inputRegisters_27__6,inputRegisters_27__5,
            inputRegisters_27__4,inputRegisters_27__3,inputRegisters_27__2,
            inputRegisters_27__1,inputRegisters_27__0})) ;
    Reg_16 loop1_27_x (.D ({inputRegisters_27__15,inputRegisters_27__14,
           inputRegisters_27__13,inputRegisters_27__12,inputRegisters_27__11,
           inputRegisters_27__10,inputRegisters_27__9,inputRegisters_27__8,
           inputRegisters_27__7,inputRegisters_27__6,inputRegisters_27__5,
           inputRegisters_27__4,inputRegisters_27__3,inputRegisters_27__2,
           inputRegisters_27__1,inputRegisters_27__0}), .en (enableRegister_27)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_27__15,
           registerOutputs_27__14,registerOutputs_27__13,registerOutputs_27__12,
           registerOutputs_27__11,registerOutputs_27__10,registerOutputs_27__9,
           registerOutputs_27__8,registerOutputs_27__7,registerOutputs_27__6,
           registerOutputs_27__5,registerOutputs_27__4,registerOutputs_27__3,
           registerOutputs_27__2,registerOutputs_27__1,registerOutputs_27__0})
           ) ;
    Mux2_16 loop1_28_y (.A ({nx35893,nx36035,nx36177,nx36319,nx36461,nx36603,
            nx36745,nx36887,nx37029,nx37171,nx37313,nx37455,nx37597,nx37739,
            nx37881,nx38023}), .B ({nx33649,nx33787,nx33925,nx34063,nx34201,
            nx34339,nx34477,nx34619,nx34761,nx34903,nx35045,nx35187,nx35329,
            nx35471,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35613), .C ({inputRegisters_28__15,inputRegisters_28__14,
            inputRegisters_28__13,inputRegisters_28__12,inputRegisters_28__11,
            inputRegisters_28__10,inputRegisters_28__9,inputRegisters_28__8,
            inputRegisters_28__7,inputRegisters_28__6,inputRegisters_28__5,
            inputRegisters_28__4,inputRegisters_28__3,inputRegisters_28__2,
            inputRegisters_28__1,inputRegisters_28__0})) ;
    Reg_16 loop1_28_x (.D ({inputRegisters_28__15,inputRegisters_28__14,
           inputRegisters_28__13,inputRegisters_28__12,inputRegisters_28__11,
           inputRegisters_28__10,inputRegisters_28__9,inputRegisters_28__8,
           inputRegisters_28__7,inputRegisters_28__6,inputRegisters_28__5,
           inputRegisters_28__4,inputRegisters_28__3,inputRegisters_28__2,
           inputRegisters_28__1,inputRegisters_28__0}), .en (enableRegister_28)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_28__15,
           registerOutputs_28__14,registerOutputs_28__13,registerOutputs_28__12,
           registerOutputs_28__11,registerOutputs_28__10,registerOutputs_28__9,
           registerOutputs_28__8,registerOutputs_28__7,registerOutputs_28__6,
           registerOutputs_28__5,registerOutputs_28__4,registerOutputs_28__3,
           registerOutputs_28__2,registerOutputs_28__1,registerOutputs_28__0})
           ) ;
    Mux2_16 loop1_29_y (.A ({nx35893,nx36035,nx36177,nx36319,nx36461,nx36603,
            nx36745,nx36887,nx37029,nx37171,nx37313,nx37455,nx37597,nx37739,
            nx37881,nx38023}), .B ({nx33649,nx33787,nx33925,nx34063,nx34201,
            nx34339,nx34479,nx34619,nx34761,nx34903,nx35045,nx35187,nx35329,
            nx35471,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35613), .C ({inputRegisters_29__15,inputRegisters_29__14,
            inputRegisters_29__13,inputRegisters_29__12,inputRegisters_29__11,
            inputRegisters_29__10,inputRegisters_29__9,inputRegisters_29__8,
            inputRegisters_29__7,inputRegisters_29__6,inputRegisters_29__5,
            inputRegisters_29__4,inputRegisters_29__3,inputRegisters_29__2,
            inputRegisters_29__1,inputRegisters_29__0})) ;
    Reg_16 loop1_29_x (.D ({inputRegisters_29__15,inputRegisters_29__14,
           inputRegisters_29__13,inputRegisters_29__12,inputRegisters_29__11,
           inputRegisters_29__10,inputRegisters_29__9,inputRegisters_29__8,
           inputRegisters_29__7,inputRegisters_29__6,inputRegisters_29__5,
           inputRegisters_29__4,inputRegisters_29__3,inputRegisters_29__2,
           inputRegisters_29__1,inputRegisters_29__0}), .en (enableRegister_29)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_29__15,
           registerOutputs_29__14,registerOutputs_29__13,registerOutputs_29__12,
           registerOutputs_29__11,registerOutputs_29__10,registerOutputs_29__9,
           registerOutputs_29__8,registerOutputs_29__7,registerOutputs_29__6,
           registerOutputs_29__5,registerOutputs_29__4,registerOutputs_29__3,
           registerOutputs_29__2,registerOutputs_29__1,registerOutputs_29__0})
           ) ;
    Mux2_16 loop1_30_y (.A ({nx35893,nx36035,nx36177,nx36319,nx36461,nx36603,
            nx36745,nx36887,nx37029,nx37171,nx37313,nx37455,nx37597,nx37739,
            nx37881,nx38023}), .B ({nx33649,nx33787,nx33925,nx34063,nx34201,
            nx34341,nx34479,nx34619,nx34761,nx34903,nx35045,nx35187,nx35329,
            nx35471,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35613), .C ({inputRegisters_30__15,inputRegisters_30__14,
            inputRegisters_30__13,inputRegisters_30__12,inputRegisters_30__11,
            inputRegisters_30__10,inputRegisters_30__9,inputRegisters_30__8,
            inputRegisters_30__7,inputRegisters_30__6,inputRegisters_30__5,
            inputRegisters_30__4,inputRegisters_30__3,inputRegisters_30__2,
            inputRegisters_30__1,inputRegisters_30__0})) ;
    Reg_16 loop1_30_x (.D ({inputRegisters_30__15,inputRegisters_30__14,
           inputRegisters_30__13,inputRegisters_30__12,inputRegisters_30__11,
           inputRegisters_30__10,inputRegisters_30__9,inputRegisters_30__8,
           inputRegisters_30__7,inputRegisters_30__6,inputRegisters_30__5,
           inputRegisters_30__4,inputRegisters_30__3,inputRegisters_30__2,
           inputRegisters_30__1,inputRegisters_30__0}), .en (enableRegister_30)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_30__15,
           registerOutputs_30__14,registerOutputs_30__13,registerOutputs_30__12,
           registerOutputs_30__11,registerOutputs_30__10,registerOutputs_30__9,
           registerOutputs_30__8,registerOutputs_30__7,registerOutputs_30__6,
           registerOutputs_30__5,registerOutputs_30__4,registerOutputs_30__3,
           registerOutputs_30__2,registerOutputs_30__1,registerOutputs_30__0})
           ) ;
    Mux2_16 loop1_31_y (.A ({nx35893,nx36035,nx36177,nx36319,nx36461,nx36603,
            nx36745,nx36887,nx37029,nx37171,nx37313,nx37455,nx37597,nx37739,
            nx37881,nx38023}), .B ({nx33649,nx33787,nx33925,nx34063,nx34203,
            nx34341,nx34479,nx34619,nx34761,nx34903,nx35045,nx35187,nx35329,
            nx35471,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35613), .C ({inputRegisters_31__15,inputRegisters_31__14,
            inputRegisters_31__13,inputRegisters_31__12,inputRegisters_31__11,
            inputRegisters_31__10,inputRegisters_31__9,inputRegisters_31__8,
            inputRegisters_31__7,inputRegisters_31__6,inputRegisters_31__5,
            inputRegisters_31__4,inputRegisters_31__3,inputRegisters_31__2,
            inputRegisters_31__1,inputRegisters_31__0})) ;
    Reg_16 loop1_31_x (.D ({inputRegisters_31__15,inputRegisters_31__14,
           inputRegisters_31__13,inputRegisters_31__12,inputRegisters_31__11,
           inputRegisters_31__10,inputRegisters_31__9,inputRegisters_31__8,
           inputRegisters_31__7,inputRegisters_31__6,inputRegisters_31__5,
           inputRegisters_31__4,inputRegisters_31__3,inputRegisters_31__2,
           inputRegisters_31__1,inputRegisters_31__0}), .en (enableRegister_31)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_31__15,
           registerOutputs_31__14,registerOutputs_31__13,registerOutputs_31__12,
           registerOutputs_31__11,registerOutputs_31__10,registerOutputs_31__9,
           registerOutputs_31__8,registerOutputs_31__7,registerOutputs_31__6,
           registerOutputs_31__5,registerOutputs_31__4,registerOutputs_31__3,
           registerOutputs_31__2,registerOutputs_31__1,registerOutputs_31__0})
           ) ;
    Mux2_16 loop1_32_y (.A ({nx35893,nx36035,nx36177,nx36319,nx36461,nx36603,
            nx36745,nx36887,nx37029,nx37171,nx37313,nx37455,nx37597,nx37739,
            nx37881,nx38023}), .B ({nx33649,nx33787,nx33925,nx34065,nx34203,
            nx34341,nx34479,nx34619,nx34761,nx34903,nx35045,nx35187,nx35329,
            nx35471,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35613), .C ({inputRegisters_32__15,inputRegisters_32__14,
            inputRegisters_32__13,inputRegisters_32__12,inputRegisters_32__11,
            inputRegisters_32__10,inputRegisters_32__9,inputRegisters_32__8,
            inputRegisters_32__7,inputRegisters_32__6,inputRegisters_32__5,
            inputRegisters_32__4,inputRegisters_32__3,inputRegisters_32__2,
            inputRegisters_32__1,inputRegisters_32__0})) ;
    Reg_16 loop1_32_x (.D ({inputRegisters_32__15,inputRegisters_32__14,
           inputRegisters_32__13,inputRegisters_32__12,inputRegisters_32__11,
           inputRegisters_32__10,inputRegisters_32__9,inputRegisters_32__8,
           inputRegisters_32__7,inputRegisters_32__6,inputRegisters_32__5,
           inputRegisters_32__4,inputRegisters_32__3,inputRegisters_32__2,
           inputRegisters_32__1,inputRegisters_32__0}), .en (enableRegister_32)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_32__15,
           registerOutputs_32__14,registerOutputs_32__13,registerOutputs_32__12,
           registerOutputs_32__11,registerOutputs_32__10,registerOutputs_32__9,
           registerOutputs_32__8,registerOutputs_32__7,registerOutputs_32__6,
           registerOutputs_32__5,registerOutputs_32__4,registerOutputs_32__3,
           registerOutputs_32__2,registerOutputs_32__1,registerOutputs_32__0})
           ) ;
    Mux2_16 loop1_33_y (.A ({nx35893,nx36035,nx36177,nx36319,nx36461,nx36603,
            nx36745,nx36887,nx37029,nx37171,nx37313,nx37455,nx37597,nx37739,
            nx37881,nx38023}), .B ({nx33649,nx33787,nx33927,nx34065,nx34203,
            nx34341,nx34479,nx34619,nx34761,nx34903,nx35045,nx35187,nx35329,
            nx35471,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35613), .C ({inputRegisters_33__15,inputRegisters_33__14,
            inputRegisters_33__13,inputRegisters_33__12,inputRegisters_33__11,
            inputRegisters_33__10,inputRegisters_33__9,inputRegisters_33__8,
            inputRegisters_33__7,inputRegisters_33__6,inputRegisters_33__5,
            inputRegisters_33__4,inputRegisters_33__3,inputRegisters_33__2,
            inputRegisters_33__1,inputRegisters_33__0})) ;
    Reg_16 loop1_33_x (.D ({inputRegisters_33__15,inputRegisters_33__14,
           inputRegisters_33__13,inputRegisters_33__12,inputRegisters_33__11,
           inputRegisters_33__10,inputRegisters_33__9,inputRegisters_33__8,
           inputRegisters_33__7,inputRegisters_33__6,inputRegisters_33__5,
           inputRegisters_33__4,inputRegisters_33__3,inputRegisters_33__2,
           inputRegisters_33__1,inputRegisters_33__0}), .en (enableRegister_33)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_33__15,
           registerOutputs_33__14,registerOutputs_33__13,registerOutputs_33__12,
           registerOutputs_33__11,registerOutputs_33__10,registerOutputs_33__9,
           registerOutputs_33__8,registerOutputs_33__7,registerOutputs_33__6,
           registerOutputs_33__5,registerOutputs_33__4,registerOutputs_33__3,
           registerOutputs_33__2,registerOutputs_33__1,registerOutputs_33__0})
           ) ;
    Mux2_16 loop1_34_y (.A ({nx35893,nx36035,nx36177,nx36319,nx36461,nx36603,
            nx36745,nx36887,nx37029,nx37171,nx37313,nx37455,nx37597,nx37739,
            nx37881,nx38023}), .B ({nx33649,nx33789,nx33927,nx34065,nx34203,
            nx34341,nx34479,nx34619,nx34761,nx34903,nx35045,nx35187,nx35329,
            nx35471,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35613), .C ({inputRegisters_34__15,inputRegisters_34__14,
            inputRegisters_34__13,inputRegisters_34__12,inputRegisters_34__11,
            inputRegisters_34__10,inputRegisters_34__9,inputRegisters_34__8,
            inputRegisters_34__7,inputRegisters_34__6,inputRegisters_34__5,
            inputRegisters_34__4,inputRegisters_34__3,inputRegisters_34__2,
            inputRegisters_34__1,inputRegisters_34__0})) ;
    Reg_16 loop1_34_x (.D ({inputRegisters_34__15,inputRegisters_34__14,
           inputRegisters_34__13,inputRegisters_34__12,inputRegisters_34__11,
           inputRegisters_34__10,inputRegisters_34__9,inputRegisters_34__8,
           inputRegisters_34__7,inputRegisters_34__6,inputRegisters_34__5,
           inputRegisters_34__4,inputRegisters_34__3,inputRegisters_34__2,
           inputRegisters_34__1,inputRegisters_34__0}), .en (enableRegister_34)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_34__15,
           registerOutputs_34__14,registerOutputs_34__13,registerOutputs_34__12,
           registerOutputs_34__11,registerOutputs_34__10,registerOutputs_34__9,
           registerOutputs_34__8,registerOutputs_34__7,registerOutputs_34__6,
           registerOutputs_34__5,registerOutputs_34__4,registerOutputs_34__3,
           registerOutputs_34__2,registerOutputs_34__1,registerOutputs_34__0})
           ) ;
    Mux2_16 loop1_35_y (.A ({nx35895,nx36037,nx36179,nx36321,nx36463,nx36605,
            nx36747,nx36889,nx37031,nx37173,nx37315,nx37457,nx37599,nx37741,
            nx37883,nx38025}), .B ({nx33651,nx33789,nx33927,nx34065,nx34203,
            nx34341,nx34479,nx34621,nx34763,nx34905,nx35047,nx35189,nx35331,
            nx35473,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35615), .C ({inputRegisters_35__15,inputRegisters_35__14,
            inputRegisters_35__13,inputRegisters_35__12,inputRegisters_35__11,
            inputRegisters_35__10,inputRegisters_35__9,inputRegisters_35__8,
            inputRegisters_35__7,inputRegisters_35__6,inputRegisters_35__5,
            inputRegisters_35__4,inputRegisters_35__3,inputRegisters_35__2,
            inputRegisters_35__1,inputRegisters_35__0})) ;
    Reg_16 loop1_35_x (.D ({inputRegisters_35__15,inputRegisters_35__14,
           inputRegisters_35__13,inputRegisters_35__12,inputRegisters_35__11,
           inputRegisters_35__10,inputRegisters_35__9,inputRegisters_35__8,
           inputRegisters_35__7,inputRegisters_35__6,inputRegisters_35__5,
           inputRegisters_35__4,inputRegisters_35__3,inputRegisters_35__2,
           inputRegisters_35__1,inputRegisters_35__0}), .en (enableRegister_35)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_35__15,
           registerOutputs_35__14,registerOutputs_35__13,registerOutputs_35__12,
           registerOutputs_35__11,registerOutputs_35__10,registerOutputs_35__9,
           registerOutputs_35__8,registerOutputs_35__7,registerOutputs_35__6,
           registerOutputs_35__5,registerOutputs_35__4,registerOutputs_35__3,
           registerOutputs_35__2,registerOutputs_35__1,registerOutputs_35__0})
           ) ;
    Mux2_16 loop1_36_y (.A ({nx35895,nx36037,nx36179,nx36321,nx36463,nx36605,
            nx36747,nx36889,nx37031,nx37173,nx37315,nx37457,nx37599,nx37741,
            nx37883,nx38025}), .B ({nx33651,nx33789,nx33927,nx34065,nx34203,
            nx34341,nx34481,nx34621,nx34763,nx34905,nx35047,nx35189,nx35331,
            nx35473,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35615), .C ({inputRegisters_36__15,inputRegisters_36__14,
            inputRegisters_36__13,inputRegisters_36__12,inputRegisters_36__11,
            inputRegisters_36__10,inputRegisters_36__9,inputRegisters_36__8,
            inputRegisters_36__7,inputRegisters_36__6,inputRegisters_36__5,
            inputRegisters_36__4,inputRegisters_36__3,inputRegisters_36__2,
            inputRegisters_36__1,inputRegisters_36__0})) ;
    Reg_16 loop1_36_x (.D ({inputRegisters_36__15,inputRegisters_36__14,
           inputRegisters_36__13,inputRegisters_36__12,inputRegisters_36__11,
           inputRegisters_36__10,inputRegisters_36__9,inputRegisters_36__8,
           inputRegisters_36__7,inputRegisters_36__6,inputRegisters_36__5,
           inputRegisters_36__4,inputRegisters_36__3,inputRegisters_36__2,
           inputRegisters_36__1,inputRegisters_36__0}), .en (enableRegister_36)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_36__15,
           registerOutputs_36__14,registerOutputs_36__13,registerOutputs_36__12,
           registerOutputs_36__11,registerOutputs_36__10,registerOutputs_36__9,
           registerOutputs_36__8,registerOutputs_36__7,registerOutputs_36__6,
           registerOutputs_36__5,registerOutputs_36__4,registerOutputs_36__3,
           registerOutputs_36__2,registerOutputs_36__1,registerOutputs_36__0})
           ) ;
    Mux2_16 loop1_37_y (.A ({nx35895,nx36037,nx36179,nx36321,nx36463,nx36605,
            nx36747,nx36889,nx37031,nx37173,nx37315,nx37457,nx37599,nx37741,
            nx37883,nx38025}), .B ({nx33651,nx33789,nx33927,nx34065,nx34203,
            nx34343,nx34481,nx34621,nx34763,nx34905,nx35047,nx35189,nx35331,
            nx35473,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35615), .C ({inputRegisters_37__15,inputRegisters_37__14,
            inputRegisters_37__13,inputRegisters_37__12,inputRegisters_37__11,
            inputRegisters_37__10,inputRegisters_37__9,inputRegisters_37__8,
            inputRegisters_37__7,inputRegisters_37__6,inputRegisters_37__5,
            inputRegisters_37__4,inputRegisters_37__3,inputRegisters_37__2,
            inputRegisters_37__1,inputRegisters_37__0})) ;
    Reg_16 loop1_37_x (.D ({inputRegisters_37__15,inputRegisters_37__14,
           inputRegisters_37__13,inputRegisters_37__12,inputRegisters_37__11,
           inputRegisters_37__10,inputRegisters_37__9,inputRegisters_37__8,
           inputRegisters_37__7,inputRegisters_37__6,inputRegisters_37__5,
           inputRegisters_37__4,inputRegisters_37__3,inputRegisters_37__2,
           inputRegisters_37__1,inputRegisters_37__0}), .en (enableRegister_37)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_37__15,
           registerOutputs_37__14,registerOutputs_37__13,registerOutputs_37__12,
           registerOutputs_37__11,registerOutputs_37__10,registerOutputs_37__9,
           registerOutputs_37__8,registerOutputs_37__7,registerOutputs_37__6,
           registerOutputs_37__5,registerOutputs_37__4,registerOutputs_37__3,
           registerOutputs_37__2,registerOutputs_37__1,registerOutputs_37__0})
           ) ;
    Mux2_16 loop1_38_y (.A ({nx35895,nx36037,nx36179,nx36321,nx36463,nx36605,
            nx36747,nx36889,nx37031,nx37173,nx37315,nx37457,nx37599,nx37741,
            nx37883,nx38025}), .B ({nx33651,nx33789,nx33927,nx34065,nx34205,
            nx34343,nx34481,nx34621,nx34763,nx34905,nx35047,nx35189,nx35331,
            nx35473,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35615), .C ({inputRegisters_38__15,inputRegisters_38__14,
            inputRegisters_38__13,inputRegisters_38__12,inputRegisters_38__11,
            inputRegisters_38__10,inputRegisters_38__9,inputRegisters_38__8,
            inputRegisters_38__7,inputRegisters_38__6,inputRegisters_38__5,
            inputRegisters_38__4,inputRegisters_38__3,inputRegisters_38__2,
            inputRegisters_38__1,inputRegisters_38__0})) ;
    Reg_16 loop1_38_x (.D ({inputRegisters_38__15,inputRegisters_38__14,
           inputRegisters_38__13,inputRegisters_38__12,inputRegisters_38__11,
           inputRegisters_38__10,inputRegisters_38__9,inputRegisters_38__8,
           inputRegisters_38__7,inputRegisters_38__6,inputRegisters_38__5,
           inputRegisters_38__4,inputRegisters_38__3,inputRegisters_38__2,
           inputRegisters_38__1,inputRegisters_38__0}), .en (enableRegister_38)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_38__15,
           registerOutputs_38__14,registerOutputs_38__13,registerOutputs_38__12,
           registerOutputs_38__11,registerOutputs_38__10,registerOutputs_38__9,
           registerOutputs_38__8,registerOutputs_38__7,registerOutputs_38__6,
           registerOutputs_38__5,registerOutputs_38__4,registerOutputs_38__3,
           registerOutputs_38__2,registerOutputs_38__1,registerOutputs_38__0})
           ) ;
    Mux2_16 loop1_39_y (.A ({nx35895,nx36037,nx36179,nx36321,nx36463,nx36605,
            nx36747,nx36889,nx37031,nx37173,nx37315,nx37457,nx37599,nx37741,
            nx37883,nx38025}), .B ({nx33651,nx33789,nx33927,nx34067,nx34205,
            nx34343,nx34481,nx34621,nx34763,nx34905,nx35047,nx35189,nx35331,
            nx35473,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35615), .C ({inputRegisters_39__15,inputRegisters_39__14,
            inputRegisters_39__13,inputRegisters_39__12,inputRegisters_39__11,
            inputRegisters_39__10,inputRegisters_39__9,inputRegisters_39__8,
            inputRegisters_39__7,inputRegisters_39__6,inputRegisters_39__5,
            inputRegisters_39__4,inputRegisters_39__3,inputRegisters_39__2,
            inputRegisters_39__1,inputRegisters_39__0})) ;
    Reg_16 loop1_39_x (.D ({inputRegisters_39__15,inputRegisters_39__14,
           inputRegisters_39__13,inputRegisters_39__12,inputRegisters_39__11,
           inputRegisters_39__10,inputRegisters_39__9,inputRegisters_39__8,
           inputRegisters_39__7,inputRegisters_39__6,inputRegisters_39__5,
           inputRegisters_39__4,inputRegisters_39__3,inputRegisters_39__2,
           inputRegisters_39__1,inputRegisters_39__0}), .en (enableRegister_39)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_39__15,
           registerOutputs_39__14,registerOutputs_39__13,registerOutputs_39__12,
           registerOutputs_39__11,registerOutputs_39__10,registerOutputs_39__9,
           registerOutputs_39__8,registerOutputs_39__7,registerOutputs_39__6,
           registerOutputs_39__5,registerOutputs_39__4,registerOutputs_39__3,
           registerOutputs_39__2,registerOutputs_39__1,registerOutputs_39__0})
           ) ;
    Mux2_16 loop1_40_y (.A ({nx35895,nx36037,nx36179,nx36321,nx36463,nx36605,
            nx36747,nx36889,nx37031,nx37173,nx37315,nx37457,nx37599,nx37741,
            nx37883,nx38025}), .B ({nx33651,nx33789,nx33929,nx34067,nx34205,
            nx34343,nx34481,nx34621,nx34763,nx34905,nx35047,nx35189,nx35331,
            nx35473,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35615), .C ({inputRegisters_40__15,inputRegisters_40__14,
            inputRegisters_40__13,inputRegisters_40__12,inputRegisters_40__11,
            inputRegisters_40__10,inputRegisters_40__9,inputRegisters_40__8,
            inputRegisters_40__7,inputRegisters_40__6,inputRegisters_40__5,
            inputRegisters_40__4,inputRegisters_40__3,inputRegisters_40__2,
            inputRegisters_40__1,inputRegisters_40__0})) ;
    Reg_16 loop1_40_x (.D ({inputRegisters_40__15,inputRegisters_40__14,
           inputRegisters_40__13,inputRegisters_40__12,inputRegisters_40__11,
           inputRegisters_40__10,inputRegisters_40__9,inputRegisters_40__8,
           inputRegisters_40__7,inputRegisters_40__6,inputRegisters_40__5,
           inputRegisters_40__4,inputRegisters_40__3,inputRegisters_40__2,
           inputRegisters_40__1,inputRegisters_40__0}), .en (enableRegister_40)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_40__15,
           registerOutputs_40__14,registerOutputs_40__13,registerOutputs_40__12,
           registerOutputs_40__11,registerOutputs_40__10,registerOutputs_40__9,
           registerOutputs_40__8,registerOutputs_40__7,registerOutputs_40__6,
           registerOutputs_40__5,registerOutputs_40__4,registerOutputs_40__3,
           registerOutputs_40__2,registerOutputs_40__1,registerOutputs_40__0})
           ) ;
    Mux2_16 loop1_41_y (.A ({nx35895,nx36037,nx36179,nx36321,nx36463,nx36605,
            nx36747,nx36889,nx37031,nx37173,nx37315,nx37457,nx37599,nx37741,
            nx37883,nx38025}), .B ({nx33651,nx33791,nx33929,nx34067,nx34205,
            nx34343,nx34481,nx34621,nx34763,nx34905,nx35047,nx35189,nx35331,
            nx35473,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35615), .C ({inputRegisters_41__15,inputRegisters_41__14,
            inputRegisters_41__13,inputRegisters_41__12,inputRegisters_41__11,
            inputRegisters_41__10,inputRegisters_41__9,inputRegisters_41__8,
            inputRegisters_41__7,inputRegisters_41__6,inputRegisters_41__5,
            inputRegisters_41__4,inputRegisters_41__3,inputRegisters_41__2,
            inputRegisters_41__1,inputRegisters_41__0})) ;
    Reg_16 loop1_41_x (.D ({inputRegisters_41__15,inputRegisters_41__14,
           inputRegisters_41__13,inputRegisters_41__12,inputRegisters_41__11,
           inputRegisters_41__10,inputRegisters_41__9,inputRegisters_41__8,
           inputRegisters_41__7,inputRegisters_41__6,inputRegisters_41__5,
           inputRegisters_41__4,inputRegisters_41__3,inputRegisters_41__2,
           inputRegisters_41__1,inputRegisters_41__0}), .en (enableRegister_41)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_41__15,
           registerOutputs_41__14,registerOutputs_41__13,registerOutputs_41__12,
           registerOutputs_41__11,registerOutputs_41__10,registerOutputs_41__9,
           registerOutputs_41__8,registerOutputs_41__7,registerOutputs_41__6,
           registerOutputs_41__5,registerOutputs_41__4,registerOutputs_41__3,
           registerOutputs_41__2,registerOutputs_41__1,registerOutputs_41__0})
           ) ;
    Mux2_16 loop1_42_y (.A ({nx35897,nx36039,nx36181,nx36323,nx36465,nx36607,
            nx36749,nx36891,nx37033,nx37175,nx37317,nx37459,nx37601,nx37743,
            nx37885,nx38027}), .B ({nx33653,nx33791,nx33929,nx34067,nx34205,
            nx34343,nx34481,nx34623,nx34765,nx34907,nx35049,nx35191,nx35333,
            nx35475,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35617), .C ({inputRegisters_42__15,inputRegisters_42__14,
            inputRegisters_42__13,inputRegisters_42__12,inputRegisters_42__11,
            inputRegisters_42__10,inputRegisters_42__9,inputRegisters_42__8,
            inputRegisters_42__7,inputRegisters_42__6,inputRegisters_42__5,
            inputRegisters_42__4,inputRegisters_42__3,inputRegisters_42__2,
            inputRegisters_42__1,inputRegisters_42__0})) ;
    Reg_16 loop1_42_x (.D ({inputRegisters_42__15,inputRegisters_42__14,
           inputRegisters_42__13,inputRegisters_42__12,inputRegisters_42__11,
           inputRegisters_42__10,inputRegisters_42__9,inputRegisters_42__8,
           inputRegisters_42__7,inputRegisters_42__6,inputRegisters_42__5,
           inputRegisters_42__4,inputRegisters_42__3,inputRegisters_42__2,
           inputRegisters_42__1,inputRegisters_42__0}), .en (enableRegister_42)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_42__15,
           registerOutputs_42__14,registerOutputs_42__13,registerOutputs_42__12,
           registerOutputs_42__11,registerOutputs_42__10,registerOutputs_42__9,
           registerOutputs_42__8,registerOutputs_42__7,registerOutputs_42__6,
           registerOutputs_42__5,registerOutputs_42__4,registerOutputs_42__3,
           registerOutputs_42__2,registerOutputs_42__1,registerOutputs_42__0})
           ) ;
    Mux2_16 loop1_43_y (.A ({nx35897,nx36039,nx36181,nx36323,nx36465,nx36607,
            nx36749,nx36891,nx37033,nx37175,nx37317,nx37459,nx37601,nx37743,
            nx37885,nx38027}), .B ({nx33653,nx33791,nx33929,nx34067,nx34205,
            nx34343,nx34483,nx34623,nx34765,nx34907,nx35049,nx35191,nx35333,
            nx35475,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35617), .C ({inputRegisters_43__15,inputRegisters_43__14,
            inputRegisters_43__13,inputRegisters_43__12,inputRegisters_43__11,
            inputRegisters_43__10,inputRegisters_43__9,inputRegisters_43__8,
            inputRegisters_43__7,inputRegisters_43__6,inputRegisters_43__5,
            inputRegisters_43__4,inputRegisters_43__3,inputRegisters_43__2,
            inputRegisters_43__1,inputRegisters_43__0})) ;
    Reg_16 loop1_43_x (.D ({inputRegisters_43__15,inputRegisters_43__14,
           inputRegisters_43__13,inputRegisters_43__12,inputRegisters_43__11,
           inputRegisters_43__10,inputRegisters_43__9,inputRegisters_43__8,
           inputRegisters_43__7,inputRegisters_43__6,inputRegisters_43__5,
           inputRegisters_43__4,inputRegisters_43__3,inputRegisters_43__2,
           inputRegisters_43__1,inputRegisters_43__0}), .en (enableRegister_43)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_43__15,
           registerOutputs_43__14,registerOutputs_43__13,registerOutputs_43__12,
           registerOutputs_43__11,registerOutputs_43__10,registerOutputs_43__9,
           registerOutputs_43__8,registerOutputs_43__7,registerOutputs_43__6,
           registerOutputs_43__5,registerOutputs_43__4,registerOutputs_43__3,
           registerOutputs_43__2,registerOutputs_43__1,registerOutputs_43__0})
           ) ;
    Mux2_16 loop1_44_y (.A ({nx35897,nx36039,nx36181,nx36323,nx36465,nx36607,
            nx36749,nx36891,nx37033,nx37175,nx37317,nx37459,nx37601,nx37743,
            nx37885,nx38027}), .B ({nx33653,nx33791,nx33929,nx34067,nx34205,
            nx34345,nx34483,nx34623,nx34765,nx34907,nx35049,nx35191,nx35333,
            nx35475,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35617), .C ({inputRegisters_44__15,inputRegisters_44__14,
            inputRegisters_44__13,inputRegisters_44__12,inputRegisters_44__11,
            inputRegisters_44__10,inputRegisters_44__9,inputRegisters_44__8,
            inputRegisters_44__7,inputRegisters_44__6,inputRegisters_44__5,
            inputRegisters_44__4,inputRegisters_44__3,inputRegisters_44__2,
            inputRegisters_44__1,inputRegisters_44__0})) ;
    Reg_16 loop1_44_x (.D ({inputRegisters_44__15,inputRegisters_44__14,
           inputRegisters_44__13,inputRegisters_44__12,inputRegisters_44__11,
           inputRegisters_44__10,inputRegisters_44__9,inputRegisters_44__8,
           inputRegisters_44__7,inputRegisters_44__6,inputRegisters_44__5,
           inputRegisters_44__4,inputRegisters_44__3,inputRegisters_44__2,
           inputRegisters_44__1,inputRegisters_44__0}), .en (enableRegister_44)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_44__15,
           registerOutputs_44__14,registerOutputs_44__13,registerOutputs_44__12,
           registerOutputs_44__11,registerOutputs_44__10,registerOutputs_44__9,
           registerOutputs_44__8,registerOutputs_44__7,registerOutputs_44__6,
           registerOutputs_44__5,registerOutputs_44__4,registerOutputs_44__3,
           registerOutputs_44__2,registerOutputs_44__1,registerOutputs_44__0})
           ) ;
    Mux2_16 loop1_45_y (.A ({nx35897,nx36039,nx36181,nx36323,nx36465,nx36607,
            nx36749,nx36891,nx37033,nx37175,nx37317,nx37459,nx37601,nx37743,
            nx37885,nx38027}), .B ({nx33653,nx33791,nx33929,nx34067,nx34207,
            nx34345,nx34483,nx34623,nx34765,nx34907,nx35049,nx35191,nx35333,
            nx35475,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35617), .C ({inputRegisters_45__15,inputRegisters_45__14,
            inputRegisters_45__13,inputRegisters_45__12,inputRegisters_45__11,
            inputRegisters_45__10,inputRegisters_45__9,inputRegisters_45__8,
            inputRegisters_45__7,inputRegisters_45__6,inputRegisters_45__5,
            inputRegisters_45__4,inputRegisters_45__3,inputRegisters_45__2,
            inputRegisters_45__1,inputRegisters_45__0})) ;
    Reg_16 loop1_45_x (.D ({inputRegisters_45__15,inputRegisters_45__14,
           inputRegisters_45__13,inputRegisters_45__12,inputRegisters_45__11,
           inputRegisters_45__10,inputRegisters_45__9,inputRegisters_45__8,
           inputRegisters_45__7,inputRegisters_45__6,inputRegisters_45__5,
           inputRegisters_45__4,inputRegisters_45__3,inputRegisters_45__2,
           inputRegisters_45__1,inputRegisters_45__0}), .en (enableRegister_45)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_45__15,
           registerOutputs_45__14,registerOutputs_45__13,registerOutputs_45__12,
           registerOutputs_45__11,registerOutputs_45__10,registerOutputs_45__9,
           registerOutputs_45__8,registerOutputs_45__7,registerOutputs_45__6,
           registerOutputs_45__5,registerOutputs_45__4,registerOutputs_45__3,
           registerOutputs_45__2,registerOutputs_45__1,registerOutputs_45__0})
           ) ;
    Mux2_16 loop1_46_y (.A ({nx35897,nx36039,nx36181,nx36323,nx36465,nx36607,
            nx36749,nx36891,nx37033,nx37175,nx37317,nx37459,nx37601,nx37743,
            nx37885,nx38027}), .B ({nx33653,nx33791,nx33929,nx34069,nx34207,
            nx34345,nx34483,nx34623,nx34765,nx34907,nx35049,nx35191,nx35333,
            nx35475,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35617), .C ({inputRegisters_46__15,inputRegisters_46__14,
            inputRegisters_46__13,inputRegisters_46__12,inputRegisters_46__11,
            inputRegisters_46__10,inputRegisters_46__9,inputRegisters_46__8,
            inputRegisters_46__7,inputRegisters_46__6,inputRegisters_46__5,
            inputRegisters_46__4,inputRegisters_46__3,inputRegisters_46__2,
            inputRegisters_46__1,inputRegisters_46__0})) ;
    Reg_16 loop1_46_x (.D ({inputRegisters_46__15,inputRegisters_46__14,
           inputRegisters_46__13,inputRegisters_46__12,inputRegisters_46__11,
           inputRegisters_46__10,inputRegisters_46__9,inputRegisters_46__8,
           inputRegisters_46__7,inputRegisters_46__6,inputRegisters_46__5,
           inputRegisters_46__4,inputRegisters_46__3,inputRegisters_46__2,
           inputRegisters_46__1,inputRegisters_46__0}), .en (enableRegister_46)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_46__15,
           registerOutputs_46__14,registerOutputs_46__13,registerOutputs_46__12,
           registerOutputs_46__11,registerOutputs_46__10,registerOutputs_46__9,
           registerOutputs_46__8,registerOutputs_46__7,registerOutputs_46__6,
           registerOutputs_46__5,registerOutputs_46__4,registerOutputs_46__3,
           registerOutputs_46__2,registerOutputs_46__1,registerOutputs_46__0})
           ) ;
    Mux2_16 loop1_47_y (.A ({nx35897,nx36039,nx36181,nx36323,nx36465,nx36607,
            nx36749,nx36891,nx37033,nx37175,nx37317,nx37459,nx37601,nx37743,
            nx37885,nx38027}), .B ({nx33653,nx33791,nx33931,nx34069,nx34207,
            nx34345,nx34483,nx34623,nx34765,nx34907,nx35049,nx35191,nx35333,
            nx35475,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35617), .C ({inputRegisters_47__15,inputRegisters_47__14,
            inputRegisters_47__13,inputRegisters_47__12,inputRegisters_47__11,
            inputRegisters_47__10,inputRegisters_47__9,inputRegisters_47__8,
            inputRegisters_47__7,inputRegisters_47__6,inputRegisters_47__5,
            inputRegisters_47__4,inputRegisters_47__3,inputRegisters_47__2,
            inputRegisters_47__1,inputRegisters_47__0})) ;
    Reg_16 loop1_47_x (.D ({inputRegisters_47__15,inputRegisters_47__14,
           inputRegisters_47__13,inputRegisters_47__12,inputRegisters_47__11,
           inputRegisters_47__10,inputRegisters_47__9,inputRegisters_47__8,
           inputRegisters_47__7,inputRegisters_47__6,inputRegisters_47__5,
           inputRegisters_47__4,inputRegisters_47__3,inputRegisters_47__2,
           inputRegisters_47__1,inputRegisters_47__0}), .en (enableRegister_47)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_47__15,
           registerOutputs_47__14,registerOutputs_47__13,registerOutputs_47__12,
           registerOutputs_47__11,registerOutputs_47__10,registerOutputs_47__9,
           registerOutputs_47__8,registerOutputs_47__7,registerOutputs_47__6,
           registerOutputs_47__5,registerOutputs_47__4,registerOutputs_47__3,
           registerOutputs_47__2,registerOutputs_47__1,registerOutputs_47__0})
           ) ;
    Mux2_16 loop1_48_y (.A ({nx35897,nx36039,nx36181,nx36323,nx36465,nx36607,
            nx36749,nx36891,nx37033,nx37175,nx37317,nx37459,nx37601,nx37743,
            nx37885,nx38027}), .B ({nx33653,nx33793,nx33931,nx34069,nx34207,
            nx34345,nx34483,nx34623,nx34765,nx34907,nx35049,nx35191,nx35333,
            nx35475,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35617), .C ({inputRegisters_48__15,inputRegisters_48__14,
            inputRegisters_48__13,inputRegisters_48__12,inputRegisters_48__11,
            inputRegisters_48__10,inputRegisters_48__9,inputRegisters_48__8,
            inputRegisters_48__7,inputRegisters_48__6,inputRegisters_48__5,
            inputRegisters_48__4,inputRegisters_48__3,inputRegisters_48__2,
            inputRegisters_48__1,inputRegisters_48__0})) ;
    Reg_16 loop1_48_x (.D ({inputRegisters_48__15,inputRegisters_48__14,
           inputRegisters_48__13,inputRegisters_48__12,inputRegisters_48__11,
           inputRegisters_48__10,inputRegisters_48__9,inputRegisters_48__8,
           inputRegisters_48__7,inputRegisters_48__6,inputRegisters_48__5,
           inputRegisters_48__4,inputRegisters_48__3,inputRegisters_48__2,
           inputRegisters_48__1,inputRegisters_48__0}), .en (enableRegister_48)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_48__15,
           registerOutputs_48__14,registerOutputs_48__13,registerOutputs_48__12,
           registerOutputs_48__11,registerOutputs_48__10,registerOutputs_48__9,
           registerOutputs_48__8,registerOutputs_48__7,registerOutputs_48__6,
           registerOutputs_48__5,registerOutputs_48__4,registerOutputs_48__3,
           registerOutputs_48__2,registerOutputs_48__1,registerOutputs_48__0})
           ) ;
    Mux2_16 loop1_49_y (.A ({nx35899,nx36041,nx36183,nx36325,nx36467,nx36609,
            nx36751,nx36893,nx37035,nx37177,nx37319,nx37461,nx37603,nx37745,
            nx37887,nx38029}), .B ({nx33655,nx33793,nx33931,nx34069,nx34207,
            nx34345,nx34483,nx34625,nx34767,nx34909,nx35051,nx35193,nx35335,
            nx35477,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35619), .C ({inputRegisters_49__15,inputRegisters_49__14,
            inputRegisters_49__13,inputRegisters_49__12,inputRegisters_49__11,
            inputRegisters_49__10,inputRegisters_49__9,inputRegisters_49__8,
            inputRegisters_49__7,inputRegisters_49__6,inputRegisters_49__5,
            inputRegisters_49__4,inputRegisters_49__3,inputRegisters_49__2,
            inputRegisters_49__1,inputRegisters_49__0})) ;
    Reg_16 loop1_49_x (.D ({inputRegisters_49__15,inputRegisters_49__14,
           inputRegisters_49__13,inputRegisters_49__12,inputRegisters_49__11,
           inputRegisters_49__10,inputRegisters_49__9,inputRegisters_49__8,
           inputRegisters_49__7,inputRegisters_49__6,inputRegisters_49__5,
           inputRegisters_49__4,inputRegisters_49__3,inputRegisters_49__2,
           inputRegisters_49__1,inputRegisters_49__0}), .en (enableRegister_49)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_49__15,
           registerOutputs_49__14,registerOutputs_49__13,registerOutputs_49__12,
           registerOutputs_49__11,registerOutputs_49__10,registerOutputs_49__9,
           registerOutputs_49__8,registerOutputs_49__7,registerOutputs_49__6,
           registerOutputs_49__5,registerOutputs_49__4,registerOutputs_49__3,
           registerOutputs_49__2,registerOutputs_49__1,registerOutputs_49__0})
           ) ;
    Mux2_16 loop1_50_y (.A ({nx35899,nx36041,nx36183,nx36325,nx36467,nx36609,
            nx36751,nx36893,nx37035,nx37177,nx37319,nx37461,nx37603,nx37745,
            nx37887,nx38029}), .B ({nx33655,nx33793,nx33931,nx34069,nx34207,
            nx34345,nx34485,nx34625,nx34767,nx34909,nx35051,nx35193,nx35335,
            nx35477,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35619), .C ({inputRegisters_50__15,inputRegisters_50__14,
            inputRegisters_50__13,inputRegisters_50__12,inputRegisters_50__11,
            inputRegisters_50__10,inputRegisters_50__9,inputRegisters_50__8,
            inputRegisters_50__7,inputRegisters_50__6,inputRegisters_50__5,
            inputRegisters_50__4,inputRegisters_50__3,inputRegisters_50__2,
            inputRegisters_50__1,inputRegisters_50__0})) ;
    Reg_16 loop1_50_x (.D ({inputRegisters_50__15,inputRegisters_50__14,
           inputRegisters_50__13,inputRegisters_50__12,inputRegisters_50__11,
           inputRegisters_50__10,inputRegisters_50__9,inputRegisters_50__8,
           inputRegisters_50__7,inputRegisters_50__6,inputRegisters_50__5,
           inputRegisters_50__4,inputRegisters_50__3,inputRegisters_50__2,
           inputRegisters_50__1,inputRegisters_50__0}), .en (enableRegister_50)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_50__15,
           registerOutputs_50__14,registerOutputs_50__13,registerOutputs_50__12,
           registerOutputs_50__11,registerOutputs_50__10,registerOutputs_50__9,
           registerOutputs_50__8,registerOutputs_50__7,registerOutputs_50__6,
           registerOutputs_50__5,registerOutputs_50__4,registerOutputs_50__3,
           registerOutputs_50__2,registerOutputs_50__1,registerOutputs_50__0})
           ) ;
    Mux2_16 loop1_51_y (.A ({nx35899,nx36041,nx36183,nx36325,nx36467,nx36609,
            nx36751,nx36893,nx37035,nx37177,nx37319,nx37461,nx37603,nx37745,
            nx37887,nx38029}), .B ({nx33655,nx33793,nx33931,nx34069,nx34207,
            nx34347,nx34485,nx34625,nx34767,nx34909,nx35051,nx35193,nx35335,
            nx35477,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35619), .C ({inputRegisters_51__15,inputRegisters_51__14,
            inputRegisters_51__13,inputRegisters_51__12,inputRegisters_51__11,
            inputRegisters_51__10,inputRegisters_51__9,inputRegisters_51__8,
            inputRegisters_51__7,inputRegisters_51__6,inputRegisters_51__5,
            inputRegisters_51__4,inputRegisters_51__3,inputRegisters_51__2,
            inputRegisters_51__1,inputRegisters_51__0})) ;
    Reg_16 loop1_51_x (.D ({inputRegisters_51__15,inputRegisters_51__14,
           inputRegisters_51__13,inputRegisters_51__12,inputRegisters_51__11,
           inputRegisters_51__10,inputRegisters_51__9,inputRegisters_51__8,
           inputRegisters_51__7,inputRegisters_51__6,inputRegisters_51__5,
           inputRegisters_51__4,inputRegisters_51__3,inputRegisters_51__2,
           inputRegisters_51__1,inputRegisters_51__0}), .en (enableRegister_51)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_51__15,
           registerOutputs_51__14,registerOutputs_51__13,registerOutputs_51__12,
           registerOutputs_51__11,registerOutputs_51__10,registerOutputs_51__9,
           registerOutputs_51__8,registerOutputs_51__7,registerOutputs_51__6,
           registerOutputs_51__5,registerOutputs_51__4,registerOutputs_51__3,
           registerOutputs_51__2,registerOutputs_51__1,registerOutputs_51__0})
           ) ;
    Mux2_16 loop1_52_y (.A ({nx35899,nx36041,nx36183,nx36325,nx36467,nx36609,
            nx36751,nx36893,nx37035,nx37177,nx37319,nx37461,nx37603,nx37745,
            nx37887,nx38029}), .B ({nx33655,nx33793,nx33931,nx34069,nx34209,
            nx34347,nx34485,nx34625,nx34767,nx34909,nx35051,nx35193,nx35335,
            nx35477,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35619), .C ({inputRegisters_52__15,inputRegisters_52__14,
            inputRegisters_52__13,inputRegisters_52__12,inputRegisters_52__11,
            inputRegisters_52__10,inputRegisters_52__9,inputRegisters_52__8,
            inputRegisters_52__7,inputRegisters_52__6,inputRegisters_52__5,
            inputRegisters_52__4,inputRegisters_52__3,inputRegisters_52__2,
            inputRegisters_52__1,inputRegisters_52__0})) ;
    Reg_16 loop1_52_x (.D ({inputRegisters_52__15,inputRegisters_52__14,
           inputRegisters_52__13,inputRegisters_52__12,inputRegisters_52__11,
           inputRegisters_52__10,inputRegisters_52__9,inputRegisters_52__8,
           inputRegisters_52__7,inputRegisters_52__6,inputRegisters_52__5,
           inputRegisters_52__4,inputRegisters_52__3,inputRegisters_52__2,
           inputRegisters_52__1,inputRegisters_52__0}), .en (enableRegister_52)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_52__15,
           registerOutputs_52__14,registerOutputs_52__13,registerOutputs_52__12,
           registerOutputs_52__11,registerOutputs_52__10,registerOutputs_52__9,
           registerOutputs_52__8,registerOutputs_52__7,registerOutputs_52__6,
           registerOutputs_52__5,registerOutputs_52__4,registerOutputs_52__3,
           registerOutputs_52__2,registerOutputs_52__1,registerOutputs_52__0})
           ) ;
    Mux2_16 loop1_53_y (.A ({nx35899,nx36041,nx36183,nx36325,nx36467,nx36609,
            nx36751,nx36893,nx37035,nx37177,nx37319,nx37461,nx37603,nx37745,
            nx37887,nx38029}), .B ({nx33655,nx33793,nx33931,nx34071,nx34209,
            nx34347,nx34485,nx34625,nx34767,nx34909,nx35051,nx35193,nx35335,
            nx35477,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35619), .C ({inputRegisters_53__15,inputRegisters_53__14,
            inputRegisters_53__13,inputRegisters_53__12,inputRegisters_53__11,
            inputRegisters_53__10,inputRegisters_53__9,inputRegisters_53__8,
            inputRegisters_53__7,inputRegisters_53__6,inputRegisters_53__5,
            inputRegisters_53__4,inputRegisters_53__3,inputRegisters_53__2,
            inputRegisters_53__1,inputRegisters_53__0})) ;
    Reg_16 loop1_53_x (.D ({inputRegisters_53__15,inputRegisters_53__14,
           inputRegisters_53__13,inputRegisters_53__12,inputRegisters_53__11,
           inputRegisters_53__10,inputRegisters_53__9,inputRegisters_53__8,
           inputRegisters_53__7,inputRegisters_53__6,inputRegisters_53__5,
           inputRegisters_53__4,inputRegisters_53__3,inputRegisters_53__2,
           inputRegisters_53__1,inputRegisters_53__0}), .en (enableRegister_53)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_53__15,
           registerOutputs_53__14,registerOutputs_53__13,registerOutputs_53__12,
           registerOutputs_53__11,registerOutputs_53__10,registerOutputs_53__9,
           registerOutputs_53__8,registerOutputs_53__7,registerOutputs_53__6,
           registerOutputs_53__5,registerOutputs_53__4,registerOutputs_53__3,
           registerOutputs_53__2,registerOutputs_53__1,registerOutputs_53__0})
           ) ;
    Mux2_16 loop1_54_y (.A ({nx35899,nx36041,nx36183,nx36325,nx36467,nx36609,
            nx36751,nx36893,nx37035,nx37177,nx37319,nx37461,nx37603,nx37745,
            nx37887,nx38029}), .B ({nx33655,nx33793,nx33933,nx34071,nx34209,
            nx34347,nx34485,nx34625,nx34767,nx34909,nx35051,nx35193,nx35335,
            nx35477,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35619), .C ({inputRegisters_54__15,inputRegisters_54__14,
            inputRegisters_54__13,inputRegisters_54__12,inputRegisters_54__11,
            inputRegisters_54__10,inputRegisters_54__9,inputRegisters_54__8,
            inputRegisters_54__7,inputRegisters_54__6,inputRegisters_54__5,
            inputRegisters_54__4,inputRegisters_54__3,inputRegisters_54__2,
            inputRegisters_54__1,inputRegisters_54__0})) ;
    Reg_16 loop1_54_x (.D ({inputRegisters_54__15,inputRegisters_54__14,
           inputRegisters_54__13,inputRegisters_54__12,inputRegisters_54__11,
           inputRegisters_54__10,inputRegisters_54__9,inputRegisters_54__8,
           inputRegisters_54__7,inputRegisters_54__6,inputRegisters_54__5,
           inputRegisters_54__4,inputRegisters_54__3,inputRegisters_54__2,
           inputRegisters_54__1,inputRegisters_54__0}), .en (enableRegister_54)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_54__15,
           registerOutputs_54__14,registerOutputs_54__13,registerOutputs_54__12,
           registerOutputs_54__11,registerOutputs_54__10,registerOutputs_54__9,
           registerOutputs_54__8,registerOutputs_54__7,registerOutputs_54__6,
           registerOutputs_54__5,registerOutputs_54__4,registerOutputs_54__3,
           registerOutputs_54__2,registerOutputs_54__1,registerOutputs_54__0})
           ) ;
    Mux2_16 loop1_55_y (.A ({nx35899,nx36041,nx36183,nx36325,nx36467,nx36609,
            nx36751,nx36893,nx37035,nx37177,nx37319,nx37461,nx37603,nx37745,
            nx37887,nx38029}), .B ({nx33655,nx33795,nx33933,nx34071,nx34209,
            nx34347,nx34485,nx34625,nx34767,nx34909,nx35051,nx35193,nx35335,
            nx35477,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35619), .C ({inputRegisters_55__15,inputRegisters_55__14,
            inputRegisters_55__13,inputRegisters_55__12,inputRegisters_55__11,
            inputRegisters_55__10,inputRegisters_55__9,inputRegisters_55__8,
            inputRegisters_55__7,inputRegisters_55__6,inputRegisters_55__5,
            inputRegisters_55__4,inputRegisters_55__3,inputRegisters_55__2,
            inputRegisters_55__1,inputRegisters_55__0})) ;
    Reg_16 loop1_55_x (.D ({inputRegisters_55__15,inputRegisters_55__14,
           inputRegisters_55__13,inputRegisters_55__12,inputRegisters_55__11,
           inputRegisters_55__10,inputRegisters_55__9,inputRegisters_55__8,
           inputRegisters_55__7,inputRegisters_55__6,inputRegisters_55__5,
           inputRegisters_55__4,inputRegisters_55__3,inputRegisters_55__2,
           inputRegisters_55__1,inputRegisters_55__0}), .en (enableRegister_55)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_55__15,
           registerOutputs_55__14,registerOutputs_55__13,registerOutputs_55__12,
           registerOutputs_55__11,registerOutputs_55__10,registerOutputs_55__9,
           registerOutputs_55__8,registerOutputs_55__7,registerOutputs_55__6,
           registerOutputs_55__5,registerOutputs_55__4,registerOutputs_55__3,
           registerOutputs_55__2,registerOutputs_55__1,registerOutputs_55__0})
           ) ;
    Mux2_16 loop1_56_y (.A ({nx35901,nx36043,nx36185,nx36327,nx36469,nx36611,
            nx36753,nx36895,nx37037,nx37179,nx37321,nx37463,nx37605,nx37747,
            nx37889,nx38031}), .B ({nx33657,nx33795,nx33933,nx34071,nx34209,
            nx34347,nx34485,nx34627,nx34769,nx34911,nx35053,nx35195,nx35337,
            nx35479,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35621), .C ({inputRegisters_56__15,inputRegisters_56__14,
            inputRegisters_56__13,inputRegisters_56__12,inputRegisters_56__11,
            inputRegisters_56__10,inputRegisters_56__9,inputRegisters_56__8,
            inputRegisters_56__7,inputRegisters_56__6,inputRegisters_56__5,
            inputRegisters_56__4,inputRegisters_56__3,inputRegisters_56__2,
            inputRegisters_56__1,inputRegisters_56__0})) ;
    Reg_16 loop1_56_x (.D ({inputRegisters_56__15,inputRegisters_56__14,
           inputRegisters_56__13,inputRegisters_56__12,inputRegisters_56__11,
           inputRegisters_56__10,inputRegisters_56__9,inputRegisters_56__8,
           inputRegisters_56__7,inputRegisters_56__6,inputRegisters_56__5,
           inputRegisters_56__4,inputRegisters_56__3,inputRegisters_56__2,
           inputRegisters_56__1,inputRegisters_56__0}), .en (enableRegister_56)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_56__15,
           registerOutputs_56__14,registerOutputs_56__13,registerOutputs_56__12,
           registerOutputs_56__11,registerOutputs_56__10,registerOutputs_56__9,
           registerOutputs_56__8,registerOutputs_56__7,registerOutputs_56__6,
           registerOutputs_56__5,registerOutputs_56__4,registerOutputs_56__3,
           registerOutputs_56__2,registerOutputs_56__1,registerOutputs_56__0})
           ) ;
    Mux2_16 loop1_57_y (.A ({nx35901,nx36043,nx36185,nx36327,nx36469,nx36611,
            nx36753,nx36895,nx37037,nx37179,nx37321,nx37463,nx37605,nx37747,
            nx37889,nx38031}), .B ({nx33657,nx33795,nx33933,nx34071,nx34209,
            nx34347,nx34487,nx34627,nx34769,nx34911,nx35053,nx35195,nx35337,
            nx35479,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35621), .C ({inputRegisters_57__15,inputRegisters_57__14,
            inputRegisters_57__13,inputRegisters_57__12,inputRegisters_57__11,
            inputRegisters_57__10,inputRegisters_57__9,inputRegisters_57__8,
            inputRegisters_57__7,inputRegisters_57__6,inputRegisters_57__5,
            inputRegisters_57__4,inputRegisters_57__3,inputRegisters_57__2,
            inputRegisters_57__1,inputRegisters_57__0})) ;
    Reg_16 loop1_57_x (.D ({inputRegisters_57__15,inputRegisters_57__14,
           inputRegisters_57__13,inputRegisters_57__12,inputRegisters_57__11,
           inputRegisters_57__10,inputRegisters_57__9,inputRegisters_57__8,
           inputRegisters_57__7,inputRegisters_57__6,inputRegisters_57__5,
           inputRegisters_57__4,inputRegisters_57__3,inputRegisters_57__2,
           inputRegisters_57__1,inputRegisters_57__0}), .en (enableRegister_57)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_57__15,
           registerOutputs_57__14,registerOutputs_57__13,registerOutputs_57__12,
           registerOutputs_57__11,registerOutputs_57__10,registerOutputs_57__9,
           registerOutputs_57__8,registerOutputs_57__7,registerOutputs_57__6,
           registerOutputs_57__5,registerOutputs_57__4,registerOutputs_57__3,
           registerOutputs_57__2,registerOutputs_57__1,registerOutputs_57__0})
           ) ;
    Mux2_16 loop1_58_y (.A ({nx35901,nx36043,nx36185,nx36327,nx36469,nx36611,
            nx36753,nx36895,nx37037,nx37179,nx37321,nx37463,nx37605,nx37747,
            nx37889,nx38031}), .B ({nx33657,nx33795,nx33933,nx34071,nx34209,
            nx34349,nx34487,nx34627,nx34769,nx34911,nx35053,nx35195,nx35337,
            nx35479,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35621), .C ({inputRegisters_58__15,inputRegisters_58__14,
            inputRegisters_58__13,inputRegisters_58__12,inputRegisters_58__11,
            inputRegisters_58__10,inputRegisters_58__9,inputRegisters_58__8,
            inputRegisters_58__7,inputRegisters_58__6,inputRegisters_58__5,
            inputRegisters_58__4,inputRegisters_58__3,inputRegisters_58__2,
            inputRegisters_58__1,inputRegisters_58__0})) ;
    Reg_16 loop1_58_x (.D ({inputRegisters_58__15,inputRegisters_58__14,
           inputRegisters_58__13,inputRegisters_58__12,inputRegisters_58__11,
           inputRegisters_58__10,inputRegisters_58__9,inputRegisters_58__8,
           inputRegisters_58__7,inputRegisters_58__6,inputRegisters_58__5,
           inputRegisters_58__4,inputRegisters_58__3,inputRegisters_58__2,
           inputRegisters_58__1,inputRegisters_58__0}), .en (enableRegister_58)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_58__15,
           registerOutputs_58__14,registerOutputs_58__13,registerOutputs_58__12,
           registerOutputs_58__11,registerOutputs_58__10,registerOutputs_58__9,
           registerOutputs_58__8,registerOutputs_58__7,registerOutputs_58__6,
           registerOutputs_58__5,registerOutputs_58__4,registerOutputs_58__3,
           registerOutputs_58__2,registerOutputs_58__1,registerOutputs_58__0})
           ) ;
    Mux2_16 loop1_59_y (.A ({nx35901,nx36043,nx36185,nx36327,nx36469,nx36611,
            nx36753,nx36895,nx37037,nx37179,nx37321,nx37463,nx37605,nx37747,
            nx37889,nx38031}), .B ({nx33657,nx33795,nx33933,nx34071,nx34211,
            nx34349,nx34487,nx34627,nx34769,nx34911,nx35053,nx35195,nx35337,
            nx35479,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35621), .C ({inputRegisters_59__15,inputRegisters_59__14,
            inputRegisters_59__13,inputRegisters_59__12,inputRegisters_59__11,
            inputRegisters_59__10,inputRegisters_59__9,inputRegisters_59__8,
            inputRegisters_59__7,inputRegisters_59__6,inputRegisters_59__5,
            inputRegisters_59__4,inputRegisters_59__3,inputRegisters_59__2,
            inputRegisters_59__1,inputRegisters_59__0})) ;
    Reg_16 loop1_59_x (.D ({inputRegisters_59__15,inputRegisters_59__14,
           inputRegisters_59__13,inputRegisters_59__12,inputRegisters_59__11,
           inputRegisters_59__10,inputRegisters_59__9,inputRegisters_59__8,
           inputRegisters_59__7,inputRegisters_59__6,inputRegisters_59__5,
           inputRegisters_59__4,inputRegisters_59__3,inputRegisters_59__2,
           inputRegisters_59__1,inputRegisters_59__0}), .en (enableRegister_59)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_59__15,
           registerOutputs_59__14,registerOutputs_59__13,registerOutputs_59__12,
           registerOutputs_59__11,registerOutputs_59__10,registerOutputs_59__9,
           registerOutputs_59__8,registerOutputs_59__7,registerOutputs_59__6,
           registerOutputs_59__5,registerOutputs_59__4,registerOutputs_59__3,
           registerOutputs_59__2,registerOutputs_59__1,registerOutputs_59__0})
           ) ;
    Mux2_16 loop1_60_y (.A ({nx35901,nx36043,nx36185,nx36327,nx36469,nx36611,
            nx36753,nx36895,nx37037,nx37179,nx37321,nx37463,nx37605,nx37747,
            nx37889,nx38031}), .B ({nx33657,nx33795,nx33933,nx34073,nx34211,
            nx34349,nx34487,nx34627,nx34769,nx34911,nx35053,nx35195,nx35337,
            nx35479,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35621), .C ({inputRegisters_60__15,inputRegisters_60__14,
            inputRegisters_60__13,inputRegisters_60__12,inputRegisters_60__11,
            inputRegisters_60__10,inputRegisters_60__9,inputRegisters_60__8,
            inputRegisters_60__7,inputRegisters_60__6,inputRegisters_60__5,
            inputRegisters_60__4,inputRegisters_60__3,inputRegisters_60__2,
            inputRegisters_60__1,inputRegisters_60__0})) ;
    Reg_16 loop1_60_x (.D ({inputRegisters_60__15,inputRegisters_60__14,
           inputRegisters_60__13,inputRegisters_60__12,inputRegisters_60__11,
           inputRegisters_60__10,inputRegisters_60__9,inputRegisters_60__8,
           inputRegisters_60__7,inputRegisters_60__6,inputRegisters_60__5,
           inputRegisters_60__4,inputRegisters_60__3,inputRegisters_60__2,
           inputRegisters_60__1,inputRegisters_60__0}), .en (enableRegister_60)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_60__15,
           registerOutputs_60__14,registerOutputs_60__13,registerOutputs_60__12,
           registerOutputs_60__11,registerOutputs_60__10,registerOutputs_60__9,
           registerOutputs_60__8,registerOutputs_60__7,registerOutputs_60__6,
           registerOutputs_60__5,registerOutputs_60__4,registerOutputs_60__3,
           registerOutputs_60__2,registerOutputs_60__1,registerOutputs_60__0})
           ) ;
    Mux2_16 loop1_61_y (.A ({nx35901,nx36043,nx36185,nx36327,nx36469,nx36611,
            nx36753,nx36895,nx37037,nx37179,nx37321,nx37463,nx37605,nx37747,
            nx37889,nx38031}), .B ({nx33657,nx33795,nx33935,nx34073,nx34211,
            nx34349,nx34487,nx34627,nx34769,nx34911,nx35053,nx35195,nx35337,
            nx35479,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35621), .C ({inputRegisters_61__15,inputRegisters_61__14,
            inputRegisters_61__13,inputRegisters_61__12,inputRegisters_61__11,
            inputRegisters_61__10,inputRegisters_61__9,inputRegisters_61__8,
            inputRegisters_61__7,inputRegisters_61__6,inputRegisters_61__5,
            inputRegisters_61__4,inputRegisters_61__3,inputRegisters_61__2,
            inputRegisters_61__1,inputRegisters_61__0})) ;
    Reg_16 loop1_61_x (.D ({inputRegisters_61__15,inputRegisters_61__14,
           inputRegisters_61__13,inputRegisters_61__12,inputRegisters_61__11,
           inputRegisters_61__10,inputRegisters_61__9,inputRegisters_61__8,
           inputRegisters_61__7,inputRegisters_61__6,inputRegisters_61__5,
           inputRegisters_61__4,inputRegisters_61__3,inputRegisters_61__2,
           inputRegisters_61__1,inputRegisters_61__0}), .en (enableRegister_61)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_61__15,
           registerOutputs_61__14,registerOutputs_61__13,registerOutputs_61__12,
           registerOutputs_61__11,registerOutputs_61__10,registerOutputs_61__9,
           registerOutputs_61__8,registerOutputs_61__7,registerOutputs_61__6,
           registerOutputs_61__5,registerOutputs_61__4,registerOutputs_61__3,
           registerOutputs_61__2,registerOutputs_61__1,registerOutputs_61__0})
           ) ;
    Mux2_16 loop1_62_y (.A ({nx35901,nx36043,nx36185,nx36327,nx36469,nx36611,
            nx36753,nx36895,nx37037,nx37179,nx37321,nx37463,nx37605,nx37747,
            nx37889,nx38031}), .B ({nx33657,nx33797,nx33935,nx34073,nx34211,
            nx34349,nx34487,nx34627,nx34769,nx34911,nx35053,nx35195,nx35337,
            nx35479,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35621), .C ({inputRegisters_62__15,inputRegisters_62__14,
            inputRegisters_62__13,inputRegisters_62__12,inputRegisters_62__11,
            inputRegisters_62__10,inputRegisters_62__9,inputRegisters_62__8,
            inputRegisters_62__7,inputRegisters_62__6,inputRegisters_62__5,
            inputRegisters_62__4,inputRegisters_62__3,inputRegisters_62__2,
            inputRegisters_62__1,inputRegisters_62__0})) ;
    Reg_16 loop1_62_x (.D ({inputRegisters_62__15,inputRegisters_62__14,
           inputRegisters_62__13,inputRegisters_62__12,inputRegisters_62__11,
           inputRegisters_62__10,inputRegisters_62__9,inputRegisters_62__8,
           inputRegisters_62__7,inputRegisters_62__6,inputRegisters_62__5,
           inputRegisters_62__4,inputRegisters_62__3,inputRegisters_62__2,
           inputRegisters_62__1,inputRegisters_62__0}), .en (enableRegister_62)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_62__15,
           registerOutputs_62__14,registerOutputs_62__13,registerOutputs_62__12,
           registerOutputs_62__11,registerOutputs_62__10,registerOutputs_62__9,
           registerOutputs_62__8,registerOutputs_62__7,registerOutputs_62__6,
           registerOutputs_62__5,registerOutputs_62__4,registerOutputs_62__3,
           registerOutputs_62__2,registerOutputs_62__1,registerOutputs_62__0})
           ) ;
    Mux2_16 loop1_63_y (.A ({nx35903,nx36045,nx36187,nx36329,nx36471,nx36613,
            nx36755,nx36897,nx37039,nx37181,nx37323,nx37465,nx37607,nx37749,
            nx37891,nx38033}), .B ({nx33659,nx33797,nx33935,nx34073,nx34211,
            nx34349,nx34487,nx34629,nx34771,nx34913,nx35055,nx35197,nx35339,
            nx35481,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35623), .C ({inputRegisters_63__15,inputRegisters_63__14,
            inputRegisters_63__13,inputRegisters_63__12,inputRegisters_63__11,
            inputRegisters_63__10,inputRegisters_63__9,inputRegisters_63__8,
            inputRegisters_63__7,inputRegisters_63__6,inputRegisters_63__5,
            inputRegisters_63__4,inputRegisters_63__3,inputRegisters_63__2,
            inputRegisters_63__1,inputRegisters_63__0})) ;
    Reg_16 loop1_63_x (.D ({inputRegisters_63__15,inputRegisters_63__14,
           inputRegisters_63__13,inputRegisters_63__12,inputRegisters_63__11,
           inputRegisters_63__10,inputRegisters_63__9,inputRegisters_63__8,
           inputRegisters_63__7,inputRegisters_63__6,inputRegisters_63__5,
           inputRegisters_63__4,inputRegisters_63__3,inputRegisters_63__2,
           inputRegisters_63__1,inputRegisters_63__0}), .en (enableRegister_63)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_63__15,
           registerOutputs_63__14,registerOutputs_63__13,registerOutputs_63__12,
           registerOutputs_63__11,registerOutputs_63__10,registerOutputs_63__9,
           registerOutputs_63__8,registerOutputs_63__7,registerOutputs_63__6,
           registerOutputs_63__5,registerOutputs_63__4,registerOutputs_63__3,
           registerOutputs_63__2,registerOutputs_63__1,registerOutputs_63__0})
           ) ;
    Mux2_16 loop1_64_y (.A ({nx35903,nx36045,nx36187,nx36329,nx36471,nx36613,
            nx36755,nx36897,nx37039,nx37181,nx37323,nx37465,nx37607,nx37749,
            nx37891,nx38033}), .B ({nx33659,nx33797,nx33935,nx34073,nx34211,
            nx34349,nx34489,nx34629,nx34771,nx34913,nx35055,nx35197,nx35339,
            nx35481,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35623), .C ({inputRegisters_64__15,inputRegisters_64__14,
            inputRegisters_64__13,inputRegisters_64__12,inputRegisters_64__11,
            inputRegisters_64__10,inputRegisters_64__9,inputRegisters_64__8,
            inputRegisters_64__7,inputRegisters_64__6,inputRegisters_64__5,
            inputRegisters_64__4,inputRegisters_64__3,inputRegisters_64__2,
            inputRegisters_64__1,inputRegisters_64__0})) ;
    Reg_16 loop1_64_x (.D ({inputRegisters_64__15,inputRegisters_64__14,
           inputRegisters_64__13,inputRegisters_64__12,inputRegisters_64__11,
           inputRegisters_64__10,inputRegisters_64__9,inputRegisters_64__8,
           inputRegisters_64__7,inputRegisters_64__6,inputRegisters_64__5,
           inputRegisters_64__4,inputRegisters_64__3,inputRegisters_64__2,
           inputRegisters_64__1,inputRegisters_64__0}), .en (enableRegister_64)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_64__15,
           registerOutputs_64__14,registerOutputs_64__13,registerOutputs_64__12,
           registerOutputs_64__11,registerOutputs_64__10,registerOutputs_64__9,
           registerOutputs_64__8,registerOutputs_64__7,registerOutputs_64__6,
           registerOutputs_64__5,registerOutputs_64__4,registerOutputs_64__3,
           registerOutputs_64__2,registerOutputs_64__1,registerOutputs_64__0})
           ) ;
    Mux2_16 loop1_65_y (.A ({nx35903,nx36045,nx36187,nx36329,nx36471,nx36613,
            nx36755,nx36897,nx37039,nx37181,nx37323,nx37465,nx37607,nx37749,
            nx37891,nx38033}), .B ({nx33659,nx33797,nx33935,nx34073,nx34211,
            nx34351,nx34489,nx34629,nx34771,nx34913,nx35055,nx35197,nx35339,
            nx35481,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35623), .C ({inputRegisters_65__15,inputRegisters_65__14,
            inputRegisters_65__13,inputRegisters_65__12,inputRegisters_65__11,
            inputRegisters_65__10,inputRegisters_65__9,inputRegisters_65__8,
            inputRegisters_65__7,inputRegisters_65__6,inputRegisters_65__5,
            inputRegisters_65__4,inputRegisters_65__3,inputRegisters_65__2,
            inputRegisters_65__1,inputRegisters_65__0})) ;
    Reg_16 loop1_65_x (.D ({inputRegisters_65__15,inputRegisters_65__14,
           inputRegisters_65__13,inputRegisters_65__12,inputRegisters_65__11,
           inputRegisters_65__10,inputRegisters_65__9,inputRegisters_65__8,
           inputRegisters_65__7,inputRegisters_65__6,inputRegisters_65__5,
           inputRegisters_65__4,inputRegisters_65__3,inputRegisters_65__2,
           inputRegisters_65__1,inputRegisters_65__0}), .en (enableRegister_65)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_65__15,
           registerOutputs_65__14,registerOutputs_65__13,registerOutputs_65__12,
           registerOutputs_65__11,registerOutputs_65__10,registerOutputs_65__9,
           registerOutputs_65__8,registerOutputs_65__7,registerOutputs_65__6,
           registerOutputs_65__5,registerOutputs_65__4,registerOutputs_65__3,
           registerOutputs_65__2,registerOutputs_65__1,registerOutputs_65__0})
           ) ;
    Mux2_16 loop1_66_y (.A ({nx35903,nx36045,nx36187,nx36329,nx36471,nx36613,
            nx36755,nx36897,nx37039,nx37181,nx37323,nx37465,nx37607,nx37749,
            nx37891,nx38033}), .B ({nx33659,nx33797,nx33935,nx34073,nx34213,
            nx34351,nx34489,nx34629,nx34771,nx34913,nx35055,nx35197,nx35339,
            nx35481,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35623), .C ({inputRegisters_66__15,inputRegisters_66__14,
            inputRegisters_66__13,inputRegisters_66__12,inputRegisters_66__11,
            inputRegisters_66__10,inputRegisters_66__9,inputRegisters_66__8,
            inputRegisters_66__7,inputRegisters_66__6,inputRegisters_66__5,
            inputRegisters_66__4,inputRegisters_66__3,inputRegisters_66__2,
            inputRegisters_66__1,inputRegisters_66__0})) ;
    Reg_16 loop1_66_x (.D ({inputRegisters_66__15,inputRegisters_66__14,
           inputRegisters_66__13,inputRegisters_66__12,inputRegisters_66__11,
           inputRegisters_66__10,inputRegisters_66__9,inputRegisters_66__8,
           inputRegisters_66__7,inputRegisters_66__6,inputRegisters_66__5,
           inputRegisters_66__4,inputRegisters_66__3,inputRegisters_66__2,
           inputRegisters_66__1,inputRegisters_66__0}), .en (enableRegister_66)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_66__15,
           registerOutputs_66__14,registerOutputs_66__13,registerOutputs_66__12,
           registerOutputs_66__11,registerOutputs_66__10,registerOutputs_66__9,
           registerOutputs_66__8,registerOutputs_66__7,registerOutputs_66__6,
           registerOutputs_66__5,registerOutputs_66__4,registerOutputs_66__3,
           registerOutputs_66__2,registerOutputs_66__1,registerOutputs_66__0})
           ) ;
    Mux2_16 loop1_67_y (.A ({nx35903,nx36045,nx36187,nx36329,nx36471,nx36613,
            nx36755,nx36897,nx37039,nx37181,nx37323,nx37465,nx37607,nx37749,
            nx37891,nx38033}), .B ({nx33659,nx33797,nx33935,nx34075,nx34213,
            nx34351,nx34489,nx34629,nx34771,nx34913,nx35055,nx35197,nx35339,
            nx35481,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35623), .C ({inputRegisters_67__15,inputRegisters_67__14,
            inputRegisters_67__13,inputRegisters_67__12,inputRegisters_67__11,
            inputRegisters_67__10,inputRegisters_67__9,inputRegisters_67__8,
            inputRegisters_67__7,inputRegisters_67__6,inputRegisters_67__5,
            inputRegisters_67__4,inputRegisters_67__3,inputRegisters_67__2,
            inputRegisters_67__1,inputRegisters_67__0})) ;
    Reg_16 loop1_67_x (.D ({inputRegisters_67__15,inputRegisters_67__14,
           inputRegisters_67__13,inputRegisters_67__12,inputRegisters_67__11,
           inputRegisters_67__10,inputRegisters_67__9,inputRegisters_67__8,
           inputRegisters_67__7,inputRegisters_67__6,inputRegisters_67__5,
           inputRegisters_67__4,inputRegisters_67__3,inputRegisters_67__2,
           inputRegisters_67__1,inputRegisters_67__0}), .en (enableRegister_67)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_67__15,
           registerOutputs_67__14,registerOutputs_67__13,registerOutputs_67__12,
           registerOutputs_67__11,registerOutputs_67__10,registerOutputs_67__9,
           registerOutputs_67__8,registerOutputs_67__7,registerOutputs_67__6,
           registerOutputs_67__5,registerOutputs_67__4,registerOutputs_67__3,
           registerOutputs_67__2,registerOutputs_67__1,registerOutputs_67__0})
           ) ;
    Mux2_16 loop1_68_y (.A ({nx35903,nx36045,nx36187,nx36329,nx36471,nx36613,
            nx36755,nx36897,nx37039,nx37181,nx37323,nx37465,nx37607,nx37749,
            nx37891,nx38033}), .B ({nx33659,nx33797,nx33937,nx34075,nx34213,
            nx34351,nx34489,nx34629,nx34771,nx34913,nx35055,nx35197,nx35339,
            nx35481,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35623), .C ({inputRegisters_68__15,inputRegisters_68__14,
            inputRegisters_68__13,inputRegisters_68__12,inputRegisters_68__11,
            inputRegisters_68__10,inputRegisters_68__9,inputRegisters_68__8,
            inputRegisters_68__7,inputRegisters_68__6,inputRegisters_68__5,
            inputRegisters_68__4,inputRegisters_68__3,inputRegisters_68__2,
            inputRegisters_68__1,inputRegisters_68__0})) ;
    Reg_16 loop1_68_x (.D ({inputRegisters_68__15,inputRegisters_68__14,
           inputRegisters_68__13,inputRegisters_68__12,inputRegisters_68__11,
           inputRegisters_68__10,inputRegisters_68__9,inputRegisters_68__8,
           inputRegisters_68__7,inputRegisters_68__6,inputRegisters_68__5,
           inputRegisters_68__4,inputRegisters_68__3,inputRegisters_68__2,
           inputRegisters_68__1,inputRegisters_68__0}), .en (enableRegister_68)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_68__15,
           registerOutputs_68__14,registerOutputs_68__13,registerOutputs_68__12,
           registerOutputs_68__11,registerOutputs_68__10,registerOutputs_68__9,
           registerOutputs_68__8,registerOutputs_68__7,registerOutputs_68__6,
           registerOutputs_68__5,registerOutputs_68__4,registerOutputs_68__3,
           registerOutputs_68__2,registerOutputs_68__1,registerOutputs_68__0})
           ) ;
    Mux2_16 loop1_69_y (.A ({nx35903,nx36045,nx36187,nx36329,nx36471,nx36613,
            nx36755,nx36897,nx37039,nx37181,nx37323,nx37465,nx37607,nx37749,
            nx37891,nx38033}), .B ({nx33659,nx33799,nx33937,nx34075,nx34213,
            nx34351,nx34489,nx34629,nx34771,nx34913,nx35055,nx35197,nx35339,
            nx35481,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35623), .C ({inputRegisters_69__15,inputRegisters_69__14,
            inputRegisters_69__13,inputRegisters_69__12,inputRegisters_69__11,
            inputRegisters_69__10,inputRegisters_69__9,inputRegisters_69__8,
            inputRegisters_69__7,inputRegisters_69__6,inputRegisters_69__5,
            inputRegisters_69__4,inputRegisters_69__3,inputRegisters_69__2,
            inputRegisters_69__1,inputRegisters_69__0})) ;
    Reg_16 loop1_69_x (.D ({inputRegisters_69__15,inputRegisters_69__14,
           inputRegisters_69__13,inputRegisters_69__12,inputRegisters_69__11,
           inputRegisters_69__10,inputRegisters_69__9,inputRegisters_69__8,
           inputRegisters_69__7,inputRegisters_69__6,inputRegisters_69__5,
           inputRegisters_69__4,inputRegisters_69__3,inputRegisters_69__2,
           inputRegisters_69__1,inputRegisters_69__0}), .en (enableRegister_69)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_69__15,
           registerOutputs_69__14,registerOutputs_69__13,registerOutputs_69__12,
           registerOutputs_69__11,registerOutputs_69__10,registerOutputs_69__9,
           registerOutputs_69__8,registerOutputs_69__7,registerOutputs_69__6,
           registerOutputs_69__5,registerOutputs_69__4,registerOutputs_69__3,
           registerOutputs_69__2,registerOutputs_69__1,registerOutputs_69__0})
           ) ;
    Mux2_16 loop1_70_y (.A ({nx35905,nx36047,nx36189,nx36331,nx36473,nx36615,
            nx36757,nx36899,nx37041,nx37183,nx37325,nx37467,nx37609,nx37751,
            nx37893,nx38035}), .B ({nx33661,nx33799,nx33937,nx34075,nx34213,
            nx34351,nx34489,nx34631,nx34773,nx34915,nx35057,nx35199,nx35341,
            nx35483,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35625), .C ({inputRegisters_70__15,inputRegisters_70__14,
            inputRegisters_70__13,inputRegisters_70__12,inputRegisters_70__11,
            inputRegisters_70__10,inputRegisters_70__9,inputRegisters_70__8,
            inputRegisters_70__7,inputRegisters_70__6,inputRegisters_70__5,
            inputRegisters_70__4,inputRegisters_70__3,inputRegisters_70__2,
            inputRegisters_70__1,inputRegisters_70__0})) ;
    Reg_16 loop1_70_x (.D ({inputRegisters_70__15,inputRegisters_70__14,
           inputRegisters_70__13,inputRegisters_70__12,inputRegisters_70__11,
           inputRegisters_70__10,inputRegisters_70__9,inputRegisters_70__8,
           inputRegisters_70__7,inputRegisters_70__6,inputRegisters_70__5,
           inputRegisters_70__4,inputRegisters_70__3,inputRegisters_70__2,
           inputRegisters_70__1,inputRegisters_70__0}), .en (enableRegister_70)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_70__15,
           registerOutputs_70__14,registerOutputs_70__13,registerOutputs_70__12,
           registerOutputs_70__11,registerOutputs_70__10,registerOutputs_70__9,
           registerOutputs_70__8,registerOutputs_70__7,registerOutputs_70__6,
           registerOutputs_70__5,registerOutputs_70__4,registerOutputs_70__3,
           registerOutputs_70__2,registerOutputs_70__1,registerOutputs_70__0})
           ) ;
    Mux2_16 loop1_71_y (.A ({nx35905,nx36047,nx36189,nx36331,nx36473,nx36615,
            nx36757,nx36899,nx37041,nx37183,nx37325,nx37467,nx37609,nx37751,
            nx37893,nx38035}), .B ({nx33661,nx33799,nx33937,nx34075,nx34213,
            nx34351,nx34491,nx34631,nx34773,nx34915,nx35057,nx35199,nx35341,
            nx35483,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35625), .C ({inputRegisters_71__15,inputRegisters_71__14,
            inputRegisters_71__13,inputRegisters_71__12,inputRegisters_71__11,
            inputRegisters_71__10,inputRegisters_71__9,inputRegisters_71__8,
            inputRegisters_71__7,inputRegisters_71__6,inputRegisters_71__5,
            inputRegisters_71__4,inputRegisters_71__3,inputRegisters_71__2,
            inputRegisters_71__1,inputRegisters_71__0})) ;
    Reg_16 loop1_71_x (.D ({inputRegisters_71__15,inputRegisters_71__14,
           inputRegisters_71__13,inputRegisters_71__12,inputRegisters_71__11,
           inputRegisters_71__10,inputRegisters_71__9,inputRegisters_71__8,
           inputRegisters_71__7,inputRegisters_71__6,inputRegisters_71__5,
           inputRegisters_71__4,inputRegisters_71__3,inputRegisters_71__2,
           inputRegisters_71__1,inputRegisters_71__0}), .en (enableRegister_71)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_71__15,
           registerOutputs_71__14,registerOutputs_71__13,registerOutputs_71__12,
           registerOutputs_71__11,registerOutputs_71__10,registerOutputs_71__9,
           registerOutputs_71__8,registerOutputs_71__7,registerOutputs_71__6,
           registerOutputs_71__5,registerOutputs_71__4,registerOutputs_71__3,
           registerOutputs_71__2,registerOutputs_71__1,registerOutputs_71__0})
           ) ;
    Mux2_16 loop1_72_y (.A ({nx35905,nx36047,nx36189,nx36331,nx36473,nx36615,
            nx36757,nx36899,nx37041,nx37183,nx37325,nx37467,nx37609,nx37751,
            nx37893,nx38035}), .B ({nx33661,nx33799,nx33937,nx34075,nx34213,
            nx34353,nx34491,nx34631,nx34773,nx34915,nx35057,nx35199,nx35341,
            nx35483,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35625), .C ({inputRegisters_72__15,inputRegisters_72__14,
            inputRegisters_72__13,inputRegisters_72__12,inputRegisters_72__11,
            inputRegisters_72__10,inputRegisters_72__9,inputRegisters_72__8,
            inputRegisters_72__7,inputRegisters_72__6,inputRegisters_72__5,
            inputRegisters_72__4,inputRegisters_72__3,inputRegisters_72__2,
            inputRegisters_72__1,inputRegisters_72__0})) ;
    Reg_16 loop1_72_x (.D ({inputRegisters_72__15,inputRegisters_72__14,
           inputRegisters_72__13,inputRegisters_72__12,inputRegisters_72__11,
           inputRegisters_72__10,inputRegisters_72__9,inputRegisters_72__8,
           inputRegisters_72__7,inputRegisters_72__6,inputRegisters_72__5,
           inputRegisters_72__4,inputRegisters_72__3,inputRegisters_72__2,
           inputRegisters_72__1,inputRegisters_72__0}), .en (enableRegister_72)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_72__15,
           registerOutputs_72__14,registerOutputs_72__13,registerOutputs_72__12,
           registerOutputs_72__11,registerOutputs_72__10,registerOutputs_72__9,
           registerOutputs_72__8,registerOutputs_72__7,registerOutputs_72__6,
           registerOutputs_72__5,registerOutputs_72__4,registerOutputs_72__3,
           registerOutputs_72__2,registerOutputs_72__1,registerOutputs_72__0})
           ) ;
    Mux2_16 loop1_73_y (.A ({nx35905,nx36047,nx36189,nx36331,nx36473,nx36615,
            nx36757,nx36899,nx37041,nx37183,nx37325,nx37467,nx37609,nx37751,
            nx37893,nx38035}), .B ({nx33661,nx33799,nx33937,nx34075,nx34215,
            nx34353,nx34491,nx34631,nx34773,nx34915,nx35057,nx35199,nx35341,
            nx35483,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35625), .C ({inputRegisters_73__15,inputRegisters_73__14,
            inputRegisters_73__13,inputRegisters_73__12,inputRegisters_73__11,
            inputRegisters_73__10,inputRegisters_73__9,inputRegisters_73__8,
            inputRegisters_73__7,inputRegisters_73__6,inputRegisters_73__5,
            inputRegisters_73__4,inputRegisters_73__3,inputRegisters_73__2,
            inputRegisters_73__1,inputRegisters_73__0})) ;
    Reg_16 loop1_73_x (.D ({inputRegisters_73__15,inputRegisters_73__14,
           inputRegisters_73__13,inputRegisters_73__12,inputRegisters_73__11,
           inputRegisters_73__10,inputRegisters_73__9,inputRegisters_73__8,
           inputRegisters_73__7,inputRegisters_73__6,inputRegisters_73__5,
           inputRegisters_73__4,inputRegisters_73__3,inputRegisters_73__2,
           inputRegisters_73__1,inputRegisters_73__0}), .en (enableRegister_73)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_73__15,
           registerOutputs_73__14,registerOutputs_73__13,registerOutputs_73__12,
           registerOutputs_73__11,registerOutputs_73__10,registerOutputs_73__9,
           registerOutputs_73__8,registerOutputs_73__7,registerOutputs_73__6,
           registerOutputs_73__5,registerOutputs_73__4,registerOutputs_73__3,
           registerOutputs_73__2,registerOutputs_73__1,registerOutputs_73__0})
           ) ;
    Mux2_16 loop1_74_y (.A ({nx35905,nx36047,nx36189,nx36331,nx36473,nx36615,
            nx36757,nx36899,nx37041,nx37183,nx37325,nx37467,nx37609,nx37751,
            nx37893,nx38035}), .B ({nx33661,nx33799,nx33937,nx34077,nx34215,
            nx34353,nx34491,nx34631,nx34773,nx34915,nx35057,nx35199,nx35341,
            nx35483,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35625), .C ({inputRegisters_74__15,inputRegisters_74__14,
            inputRegisters_74__13,inputRegisters_74__12,inputRegisters_74__11,
            inputRegisters_74__10,inputRegisters_74__9,inputRegisters_74__8,
            inputRegisters_74__7,inputRegisters_74__6,inputRegisters_74__5,
            inputRegisters_74__4,inputRegisters_74__3,inputRegisters_74__2,
            inputRegisters_74__1,inputRegisters_74__0})) ;
    Reg_16 loop1_74_x (.D ({inputRegisters_74__15,inputRegisters_74__14,
           inputRegisters_74__13,inputRegisters_74__12,inputRegisters_74__11,
           inputRegisters_74__10,inputRegisters_74__9,inputRegisters_74__8,
           inputRegisters_74__7,inputRegisters_74__6,inputRegisters_74__5,
           inputRegisters_74__4,inputRegisters_74__3,inputRegisters_74__2,
           inputRegisters_74__1,inputRegisters_74__0}), .en (enableRegister_74)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_74__15,
           registerOutputs_74__14,registerOutputs_74__13,registerOutputs_74__12,
           registerOutputs_74__11,registerOutputs_74__10,registerOutputs_74__9,
           registerOutputs_74__8,registerOutputs_74__7,registerOutputs_74__6,
           registerOutputs_74__5,registerOutputs_74__4,registerOutputs_74__3,
           registerOutputs_74__2,registerOutputs_74__1,registerOutputs_74__0})
           ) ;
    Mux2_16 loop1_75_y (.A ({nx35905,nx36047,nx36189,nx36331,nx36473,nx36615,
            nx36757,nx36899,nx37041,nx37183,nx37325,nx37467,nx37609,nx37751,
            nx37893,nx38035}), .B ({nx33661,nx33799,nx33939,nx34077,nx34215,
            nx34353,nx34491,nx34631,nx34773,nx34915,nx35057,nx35199,nx35341,
            nx35483,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35625), .C ({inputRegisters_75__15,inputRegisters_75__14,
            inputRegisters_75__13,inputRegisters_75__12,inputRegisters_75__11,
            inputRegisters_75__10,inputRegisters_75__9,inputRegisters_75__8,
            inputRegisters_75__7,inputRegisters_75__6,inputRegisters_75__5,
            inputRegisters_75__4,inputRegisters_75__3,inputRegisters_75__2,
            inputRegisters_75__1,inputRegisters_75__0})) ;
    Reg_16 loop1_75_x (.D ({inputRegisters_75__15,inputRegisters_75__14,
           inputRegisters_75__13,inputRegisters_75__12,inputRegisters_75__11,
           inputRegisters_75__10,inputRegisters_75__9,inputRegisters_75__8,
           inputRegisters_75__7,inputRegisters_75__6,inputRegisters_75__5,
           inputRegisters_75__4,inputRegisters_75__3,inputRegisters_75__2,
           inputRegisters_75__1,inputRegisters_75__0}), .en (enableRegister_75)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_75__15,
           registerOutputs_75__14,registerOutputs_75__13,registerOutputs_75__12,
           registerOutputs_75__11,registerOutputs_75__10,registerOutputs_75__9,
           registerOutputs_75__8,registerOutputs_75__7,registerOutputs_75__6,
           registerOutputs_75__5,registerOutputs_75__4,registerOutputs_75__3,
           registerOutputs_75__2,registerOutputs_75__1,registerOutputs_75__0})
           ) ;
    Mux2_16 loop1_76_y (.A ({nx35905,nx36047,nx36189,nx36331,nx36473,nx36615,
            nx36757,nx36899,nx37041,nx37183,nx37325,nx37467,nx37609,nx37751,
            nx37893,nx38035}), .B ({nx33661,nx33801,nx33939,nx34077,nx34215,
            nx34353,nx34491,nx34631,nx34773,nx34915,nx35057,nx35199,nx35341,
            nx35483,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35625), .C ({inputRegisters_76__15,inputRegisters_76__14,
            inputRegisters_76__13,inputRegisters_76__12,inputRegisters_76__11,
            inputRegisters_76__10,inputRegisters_76__9,inputRegisters_76__8,
            inputRegisters_76__7,inputRegisters_76__6,inputRegisters_76__5,
            inputRegisters_76__4,inputRegisters_76__3,inputRegisters_76__2,
            inputRegisters_76__1,inputRegisters_76__0})) ;
    Reg_16 loop1_76_x (.D ({inputRegisters_76__15,inputRegisters_76__14,
           inputRegisters_76__13,inputRegisters_76__12,inputRegisters_76__11,
           inputRegisters_76__10,inputRegisters_76__9,inputRegisters_76__8,
           inputRegisters_76__7,inputRegisters_76__6,inputRegisters_76__5,
           inputRegisters_76__4,inputRegisters_76__3,inputRegisters_76__2,
           inputRegisters_76__1,inputRegisters_76__0}), .en (enableRegister_76)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_76__15,
           registerOutputs_76__14,registerOutputs_76__13,registerOutputs_76__12,
           registerOutputs_76__11,registerOutputs_76__10,registerOutputs_76__9,
           registerOutputs_76__8,registerOutputs_76__7,registerOutputs_76__6,
           registerOutputs_76__5,registerOutputs_76__4,registerOutputs_76__3,
           registerOutputs_76__2,registerOutputs_76__1,registerOutputs_76__0})
           ) ;
    Mux2_16 loop1_77_y (.A ({nx35907,nx36049,nx36191,nx36333,nx36475,nx36617,
            nx36759,nx36901,nx37043,nx37185,nx37327,nx37469,nx37611,nx37753,
            nx37895,nx38037}), .B ({nx33663,nx33801,nx33939,nx34077,nx34215,
            nx34353,nx34491,nx34633,nx34775,nx34917,nx35059,nx35201,nx35343,
            nx35485,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35627), .C ({inputRegisters_77__15,inputRegisters_77__14,
            inputRegisters_77__13,inputRegisters_77__12,inputRegisters_77__11,
            inputRegisters_77__10,inputRegisters_77__9,inputRegisters_77__8,
            inputRegisters_77__7,inputRegisters_77__6,inputRegisters_77__5,
            inputRegisters_77__4,inputRegisters_77__3,inputRegisters_77__2,
            inputRegisters_77__1,inputRegisters_77__0})) ;
    Reg_16 loop1_77_x (.D ({inputRegisters_77__15,inputRegisters_77__14,
           inputRegisters_77__13,inputRegisters_77__12,inputRegisters_77__11,
           inputRegisters_77__10,inputRegisters_77__9,inputRegisters_77__8,
           inputRegisters_77__7,inputRegisters_77__6,inputRegisters_77__5,
           inputRegisters_77__4,inputRegisters_77__3,inputRegisters_77__2,
           inputRegisters_77__1,inputRegisters_77__0}), .en (enableRegister_77)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_77__15,
           registerOutputs_77__14,registerOutputs_77__13,registerOutputs_77__12,
           registerOutputs_77__11,registerOutputs_77__10,registerOutputs_77__9,
           registerOutputs_77__8,registerOutputs_77__7,registerOutputs_77__6,
           registerOutputs_77__5,registerOutputs_77__4,registerOutputs_77__3,
           registerOutputs_77__2,registerOutputs_77__1,registerOutputs_77__0})
           ) ;
    Mux2_16 loop1_78_y (.A ({nx35907,nx36049,nx36191,nx36333,nx36475,nx36617,
            nx36759,nx36901,nx37043,nx37185,nx37327,nx37469,nx37611,nx37753,
            nx37895,nx38037}), .B ({nx33663,nx33801,nx33939,nx34077,nx34215,
            nx34353,nx34493,nx34633,nx34775,nx34917,nx35059,nx35201,nx35343,
            nx35485,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35627), .C ({inputRegisters_78__15,inputRegisters_78__14,
            inputRegisters_78__13,inputRegisters_78__12,inputRegisters_78__11,
            inputRegisters_78__10,inputRegisters_78__9,inputRegisters_78__8,
            inputRegisters_78__7,inputRegisters_78__6,inputRegisters_78__5,
            inputRegisters_78__4,inputRegisters_78__3,inputRegisters_78__2,
            inputRegisters_78__1,inputRegisters_78__0})) ;
    Reg_16 loop1_78_x (.D ({inputRegisters_78__15,inputRegisters_78__14,
           inputRegisters_78__13,inputRegisters_78__12,inputRegisters_78__11,
           inputRegisters_78__10,inputRegisters_78__9,inputRegisters_78__8,
           inputRegisters_78__7,inputRegisters_78__6,inputRegisters_78__5,
           inputRegisters_78__4,inputRegisters_78__3,inputRegisters_78__2,
           inputRegisters_78__1,inputRegisters_78__0}), .en (enableRegister_78)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_78__15,
           registerOutputs_78__14,registerOutputs_78__13,registerOutputs_78__12,
           registerOutputs_78__11,registerOutputs_78__10,registerOutputs_78__9,
           registerOutputs_78__8,registerOutputs_78__7,registerOutputs_78__6,
           registerOutputs_78__5,registerOutputs_78__4,registerOutputs_78__3,
           registerOutputs_78__2,registerOutputs_78__1,registerOutputs_78__0})
           ) ;
    Mux2_16 loop1_79_y (.A ({nx35907,nx36049,nx36191,nx36333,nx36475,nx36617,
            nx36759,nx36901,nx37043,nx37185,nx37327,nx37469,nx37611,nx37753,
            nx37895,nx38037}), .B ({nx33663,nx33801,nx33939,nx34077,nx34215,
            nx34355,nx34493,nx34633,nx34775,nx34917,nx35059,nx35201,nx35343,
            nx35485,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35627), .C ({inputRegisters_79__15,inputRegisters_79__14,
            inputRegisters_79__13,inputRegisters_79__12,inputRegisters_79__11,
            inputRegisters_79__10,inputRegisters_79__9,inputRegisters_79__8,
            inputRegisters_79__7,inputRegisters_79__6,inputRegisters_79__5,
            inputRegisters_79__4,inputRegisters_79__3,inputRegisters_79__2,
            inputRegisters_79__1,inputRegisters_79__0})) ;
    Reg_16 loop1_79_x (.D ({inputRegisters_79__15,inputRegisters_79__14,
           inputRegisters_79__13,inputRegisters_79__12,inputRegisters_79__11,
           inputRegisters_79__10,inputRegisters_79__9,inputRegisters_79__8,
           inputRegisters_79__7,inputRegisters_79__6,inputRegisters_79__5,
           inputRegisters_79__4,inputRegisters_79__3,inputRegisters_79__2,
           inputRegisters_79__1,inputRegisters_79__0}), .en (enableRegister_79)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_79__15,
           registerOutputs_79__14,registerOutputs_79__13,registerOutputs_79__12,
           registerOutputs_79__11,registerOutputs_79__10,registerOutputs_79__9,
           registerOutputs_79__8,registerOutputs_79__7,registerOutputs_79__6,
           registerOutputs_79__5,registerOutputs_79__4,registerOutputs_79__3,
           registerOutputs_79__2,registerOutputs_79__1,registerOutputs_79__0})
           ) ;
    Mux2_16 loop1_80_y (.A ({nx35907,nx36049,nx36191,nx36333,nx36475,nx36617,
            nx36759,nx36901,nx37043,nx37185,nx37327,nx37469,nx37611,nx37753,
            nx37895,nx38037}), .B ({nx33663,nx33801,nx33939,nx34077,nx34217,
            nx34355,nx34493,nx34633,nx34775,nx34917,nx35059,nx35201,nx35343,
            nx35485,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35627), .C ({inputRegisters_80__15,inputRegisters_80__14,
            inputRegisters_80__13,inputRegisters_80__12,inputRegisters_80__11,
            inputRegisters_80__10,inputRegisters_80__9,inputRegisters_80__8,
            inputRegisters_80__7,inputRegisters_80__6,inputRegisters_80__5,
            inputRegisters_80__4,inputRegisters_80__3,inputRegisters_80__2,
            inputRegisters_80__1,inputRegisters_80__0})) ;
    Reg_16 loop1_80_x (.D ({inputRegisters_80__15,inputRegisters_80__14,
           inputRegisters_80__13,inputRegisters_80__12,inputRegisters_80__11,
           inputRegisters_80__10,inputRegisters_80__9,inputRegisters_80__8,
           inputRegisters_80__7,inputRegisters_80__6,inputRegisters_80__5,
           inputRegisters_80__4,inputRegisters_80__3,inputRegisters_80__2,
           inputRegisters_80__1,inputRegisters_80__0}), .en (enableRegister_80)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_80__15,
           registerOutputs_80__14,registerOutputs_80__13,registerOutputs_80__12,
           registerOutputs_80__11,registerOutputs_80__10,registerOutputs_80__9,
           registerOutputs_80__8,registerOutputs_80__7,registerOutputs_80__6,
           registerOutputs_80__5,registerOutputs_80__4,registerOutputs_80__3,
           registerOutputs_80__2,registerOutputs_80__1,registerOutputs_80__0})
           ) ;
    Mux2_16 loop1_81_y (.A ({nx35907,nx36049,nx36191,nx36333,nx36475,nx36617,
            nx36759,nx36901,nx37043,nx37185,nx37327,nx37469,nx37611,nx37753,
            nx37895,nx38037}), .B ({nx33663,nx33801,nx33939,nx34079,nx34217,
            nx34355,nx34493,nx34633,nx34775,nx34917,nx35059,nx35201,nx35343,
            nx35485,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35627), .C ({inputRegisters_81__15,inputRegisters_81__14,
            inputRegisters_81__13,inputRegisters_81__12,inputRegisters_81__11,
            inputRegisters_81__10,inputRegisters_81__9,inputRegisters_81__8,
            inputRegisters_81__7,inputRegisters_81__6,inputRegisters_81__5,
            inputRegisters_81__4,inputRegisters_81__3,inputRegisters_81__2,
            inputRegisters_81__1,inputRegisters_81__0})) ;
    Reg_16 loop1_81_x (.D ({inputRegisters_81__15,inputRegisters_81__14,
           inputRegisters_81__13,inputRegisters_81__12,inputRegisters_81__11,
           inputRegisters_81__10,inputRegisters_81__9,inputRegisters_81__8,
           inputRegisters_81__7,inputRegisters_81__6,inputRegisters_81__5,
           inputRegisters_81__4,inputRegisters_81__3,inputRegisters_81__2,
           inputRegisters_81__1,inputRegisters_81__0}), .en (enableRegister_81)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_81__15,
           registerOutputs_81__14,registerOutputs_81__13,registerOutputs_81__12,
           registerOutputs_81__11,registerOutputs_81__10,registerOutputs_81__9,
           registerOutputs_81__8,registerOutputs_81__7,registerOutputs_81__6,
           registerOutputs_81__5,registerOutputs_81__4,registerOutputs_81__3,
           registerOutputs_81__2,registerOutputs_81__1,registerOutputs_81__0})
           ) ;
    Mux2_16 loop1_82_y (.A ({nx35907,nx36049,nx36191,nx36333,nx36475,nx36617,
            nx36759,nx36901,nx37043,nx37185,nx37327,nx37469,nx37611,nx37753,
            nx37895,nx38037}), .B ({nx33663,nx33801,nx33941,nx34079,nx34217,
            nx34355,nx34493,nx34633,nx34775,nx34917,nx35059,nx35201,nx35343,
            nx35485,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35627), .C ({inputRegisters_82__15,inputRegisters_82__14,
            inputRegisters_82__13,inputRegisters_82__12,inputRegisters_82__11,
            inputRegisters_82__10,inputRegisters_82__9,inputRegisters_82__8,
            inputRegisters_82__7,inputRegisters_82__6,inputRegisters_82__5,
            inputRegisters_82__4,inputRegisters_82__3,inputRegisters_82__2,
            inputRegisters_82__1,inputRegisters_82__0})) ;
    Reg_16 loop1_82_x (.D ({inputRegisters_82__15,inputRegisters_82__14,
           inputRegisters_82__13,inputRegisters_82__12,inputRegisters_82__11,
           inputRegisters_82__10,inputRegisters_82__9,inputRegisters_82__8,
           inputRegisters_82__7,inputRegisters_82__6,inputRegisters_82__5,
           inputRegisters_82__4,inputRegisters_82__3,inputRegisters_82__2,
           inputRegisters_82__1,inputRegisters_82__0}), .en (enableRegister_82)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_82__15,
           registerOutputs_82__14,registerOutputs_82__13,registerOutputs_82__12,
           registerOutputs_82__11,registerOutputs_82__10,registerOutputs_82__9,
           registerOutputs_82__8,registerOutputs_82__7,registerOutputs_82__6,
           registerOutputs_82__5,registerOutputs_82__4,registerOutputs_82__3,
           registerOutputs_82__2,registerOutputs_82__1,registerOutputs_82__0})
           ) ;
    Mux2_16 loop1_83_y (.A ({nx35907,nx36049,nx36191,nx36333,nx36475,nx36617,
            nx36759,nx36901,nx37043,nx37185,nx37327,nx37469,nx37611,nx37753,
            nx37895,nx38037}), .B ({nx33663,nx33803,nx33941,nx34079,nx34217,
            nx34355,nx34493,nx34633,nx34775,nx34917,nx35059,nx35201,nx35343,
            nx35485,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35627), .C ({inputRegisters_83__15,inputRegisters_83__14,
            inputRegisters_83__13,inputRegisters_83__12,inputRegisters_83__11,
            inputRegisters_83__10,inputRegisters_83__9,inputRegisters_83__8,
            inputRegisters_83__7,inputRegisters_83__6,inputRegisters_83__5,
            inputRegisters_83__4,inputRegisters_83__3,inputRegisters_83__2,
            inputRegisters_83__1,inputRegisters_83__0})) ;
    Reg_16 loop1_83_x (.D ({inputRegisters_83__15,inputRegisters_83__14,
           inputRegisters_83__13,inputRegisters_83__12,inputRegisters_83__11,
           inputRegisters_83__10,inputRegisters_83__9,inputRegisters_83__8,
           inputRegisters_83__7,inputRegisters_83__6,inputRegisters_83__5,
           inputRegisters_83__4,inputRegisters_83__3,inputRegisters_83__2,
           inputRegisters_83__1,inputRegisters_83__0}), .en (enableRegister_83)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_83__15,
           registerOutputs_83__14,registerOutputs_83__13,registerOutputs_83__12,
           registerOutputs_83__11,registerOutputs_83__10,registerOutputs_83__9,
           registerOutputs_83__8,registerOutputs_83__7,registerOutputs_83__6,
           registerOutputs_83__5,registerOutputs_83__4,registerOutputs_83__3,
           registerOutputs_83__2,registerOutputs_83__1,registerOutputs_83__0})
           ) ;
    Mux2_16 loop1_84_y (.A ({nx35909,nx36051,nx36193,nx36335,nx36477,nx36619,
            nx36761,nx36903,nx37045,nx37187,nx37329,nx37471,nx37613,nx37755,
            nx37897,nx38039}), .B ({nx33665,nx33803,nx33941,nx34079,nx34217,
            nx34355,nx34493,nx34635,nx34777,nx34919,nx35061,nx35203,nx35345,
            nx35487,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35629), .C ({inputRegisters_84__15,inputRegisters_84__14,
            inputRegisters_84__13,inputRegisters_84__12,inputRegisters_84__11,
            inputRegisters_84__10,inputRegisters_84__9,inputRegisters_84__8,
            inputRegisters_84__7,inputRegisters_84__6,inputRegisters_84__5,
            inputRegisters_84__4,inputRegisters_84__3,inputRegisters_84__2,
            inputRegisters_84__1,inputRegisters_84__0})) ;
    Reg_16 loop1_84_x (.D ({inputRegisters_84__15,inputRegisters_84__14,
           inputRegisters_84__13,inputRegisters_84__12,inputRegisters_84__11,
           inputRegisters_84__10,inputRegisters_84__9,inputRegisters_84__8,
           inputRegisters_84__7,inputRegisters_84__6,inputRegisters_84__5,
           inputRegisters_84__4,inputRegisters_84__3,inputRegisters_84__2,
           inputRegisters_84__1,inputRegisters_84__0}), .en (enableRegister_84)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_84__15,
           registerOutputs_84__14,registerOutputs_84__13,registerOutputs_84__12,
           registerOutputs_84__11,registerOutputs_84__10,registerOutputs_84__9,
           registerOutputs_84__8,registerOutputs_84__7,registerOutputs_84__6,
           registerOutputs_84__5,registerOutputs_84__4,registerOutputs_84__3,
           registerOutputs_84__2,registerOutputs_84__1,registerOutputs_84__0})
           ) ;
    Mux2_16 loop1_85_y (.A ({nx35909,nx36051,nx36193,nx36335,nx36477,nx36619,
            nx36761,nx36903,nx37045,nx37187,nx37329,nx37471,nx37613,nx37755,
            nx37897,nx38039}), .B ({nx33665,nx33803,nx33941,nx34079,nx34217,
            nx34355,nx34495,nx34635,nx34777,nx34919,nx35061,nx35203,nx35345,
            nx35487,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35629), .C ({inputRegisters_85__15,inputRegisters_85__14,
            inputRegisters_85__13,inputRegisters_85__12,inputRegisters_85__11,
            inputRegisters_85__10,inputRegisters_85__9,inputRegisters_85__8,
            inputRegisters_85__7,inputRegisters_85__6,inputRegisters_85__5,
            inputRegisters_85__4,inputRegisters_85__3,inputRegisters_85__2,
            inputRegisters_85__1,inputRegisters_85__0})) ;
    Reg_16 loop1_85_x (.D ({inputRegisters_85__15,inputRegisters_85__14,
           inputRegisters_85__13,inputRegisters_85__12,inputRegisters_85__11,
           inputRegisters_85__10,inputRegisters_85__9,inputRegisters_85__8,
           inputRegisters_85__7,inputRegisters_85__6,inputRegisters_85__5,
           inputRegisters_85__4,inputRegisters_85__3,inputRegisters_85__2,
           inputRegisters_85__1,inputRegisters_85__0}), .en (enableRegister_85)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_85__15,
           registerOutputs_85__14,registerOutputs_85__13,registerOutputs_85__12,
           registerOutputs_85__11,registerOutputs_85__10,registerOutputs_85__9,
           registerOutputs_85__8,registerOutputs_85__7,registerOutputs_85__6,
           registerOutputs_85__5,registerOutputs_85__4,registerOutputs_85__3,
           registerOutputs_85__2,registerOutputs_85__1,registerOutputs_85__0})
           ) ;
    Mux2_16 loop1_86_y (.A ({nx35909,nx36051,nx36193,nx36335,nx36477,nx36619,
            nx36761,nx36903,nx37045,nx37187,nx37329,nx37471,nx37613,nx37755,
            nx37897,nx38039}), .B ({nx33665,nx33803,nx33941,nx34079,nx34217,
            nx34357,nx34495,nx34635,nx34777,nx34919,nx35061,nx35203,nx35345,
            nx35487,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35629), .C ({inputRegisters_86__15,inputRegisters_86__14,
            inputRegisters_86__13,inputRegisters_86__12,inputRegisters_86__11,
            inputRegisters_86__10,inputRegisters_86__9,inputRegisters_86__8,
            inputRegisters_86__7,inputRegisters_86__6,inputRegisters_86__5,
            inputRegisters_86__4,inputRegisters_86__3,inputRegisters_86__2,
            inputRegisters_86__1,inputRegisters_86__0})) ;
    Reg_16 loop1_86_x (.D ({inputRegisters_86__15,inputRegisters_86__14,
           inputRegisters_86__13,inputRegisters_86__12,inputRegisters_86__11,
           inputRegisters_86__10,inputRegisters_86__9,inputRegisters_86__8,
           inputRegisters_86__7,inputRegisters_86__6,inputRegisters_86__5,
           inputRegisters_86__4,inputRegisters_86__3,inputRegisters_86__2,
           inputRegisters_86__1,inputRegisters_86__0}), .en (enableRegister_86)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_86__15,
           registerOutputs_86__14,registerOutputs_86__13,registerOutputs_86__12,
           registerOutputs_86__11,registerOutputs_86__10,registerOutputs_86__9,
           registerOutputs_86__8,registerOutputs_86__7,registerOutputs_86__6,
           registerOutputs_86__5,registerOutputs_86__4,registerOutputs_86__3,
           registerOutputs_86__2,registerOutputs_86__1,registerOutputs_86__0})
           ) ;
    Mux2_16 loop1_87_y (.A ({nx35909,nx36051,nx36193,nx36335,nx36477,nx36619,
            nx36761,nx36903,nx37045,nx37187,nx37329,nx37471,nx37613,nx37755,
            nx37897,nx38039}), .B ({nx33665,nx33803,nx33941,nx34079,nx34219,
            nx34357,nx34495,nx34635,nx34777,nx34919,nx35061,nx35203,nx35345,
            nx35487,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35629), .C ({inputRegisters_87__15,inputRegisters_87__14,
            inputRegisters_87__13,inputRegisters_87__12,inputRegisters_87__11,
            inputRegisters_87__10,inputRegisters_87__9,inputRegisters_87__8,
            inputRegisters_87__7,inputRegisters_87__6,inputRegisters_87__5,
            inputRegisters_87__4,inputRegisters_87__3,inputRegisters_87__2,
            inputRegisters_87__1,inputRegisters_87__0})) ;
    Reg_16 loop1_87_x (.D ({inputRegisters_87__15,inputRegisters_87__14,
           inputRegisters_87__13,inputRegisters_87__12,inputRegisters_87__11,
           inputRegisters_87__10,inputRegisters_87__9,inputRegisters_87__8,
           inputRegisters_87__7,inputRegisters_87__6,inputRegisters_87__5,
           inputRegisters_87__4,inputRegisters_87__3,inputRegisters_87__2,
           inputRegisters_87__1,inputRegisters_87__0}), .en (enableRegister_87)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_87__15,
           registerOutputs_87__14,registerOutputs_87__13,registerOutputs_87__12,
           registerOutputs_87__11,registerOutputs_87__10,registerOutputs_87__9,
           registerOutputs_87__8,registerOutputs_87__7,registerOutputs_87__6,
           registerOutputs_87__5,registerOutputs_87__4,registerOutputs_87__3,
           registerOutputs_87__2,registerOutputs_87__1,registerOutputs_87__0})
           ) ;
    Mux2_16 loop1_88_y (.A ({nx35909,nx36051,nx36193,nx36335,nx36477,nx36619,
            nx36761,nx36903,nx37045,nx37187,nx37329,nx37471,nx37613,nx37755,
            nx37897,nx38039}), .B ({nx33665,nx33803,nx33941,nx34081,nx34219,
            nx34357,nx34495,nx34635,nx34777,nx34919,nx35061,nx35203,nx35345,
            nx35487,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35629), .C ({inputRegisters_88__15,inputRegisters_88__14,
            inputRegisters_88__13,inputRegisters_88__12,inputRegisters_88__11,
            inputRegisters_88__10,inputRegisters_88__9,inputRegisters_88__8,
            inputRegisters_88__7,inputRegisters_88__6,inputRegisters_88__5,
            inputRegisters_88__4,inputRegisters_88__3,inputRegisters_88__2,
            inputRegisters_88__1,inputRegisters_88__0})) ;
    Reg_16 loop1_88_x (.D ({inputRegisters_88__15,inputRegisters_88__14,
           inputRegisters_88__13,inputRegisters_88__12,inputRegisters_88__11,
           inputRegisters_88__10,inputRegisters_88__9,inputRegisters_88__8,
           inputRegisters_88__7,inputRegisters_88__6,inputRegisters_88__5,
           inputRegisters_88__4,inputRegisters_88__3,inputRegisters_88__2,
           inputRegisters_88__1,inputRegisters_88__0}), .en (enableRegister_88)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_88__15,
           registerOutputs_88__14,registerOutputs_88__13,registerOutputs_88__12,
           registerOutputs_88__11,registerOutputs_88__10,registerOutputs_88__9,
           registerOutputs_88__8,registerOutputs_88__7,registerOutputs_88__6,
           registerOutputs_88__5,registerOutputs_88__4,registerOutputs_88__3,
           registerOutputs_88__2,registerOutputs_88__1,registerOutputs_88__0})
           ) ;
    Mux2_16 loop1_89_y (.A ({nx35909,nx36051,nx36193,nx36335,nx36477,nx36619,
            nx36761,nx36903,nx37045,nx37187,nx37329,nx37471,nx37613,nx37755,
            nx37897,nx38039}), .B ({nx33665,nx33803,nx33943,nx34081,nx34219,
            nx34357,nx34495,nx34635,nx34777,nx34919,nx35061,nx35203,nx35345,
            nx35487,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35629), .C ({inputRegisters_89__15,inputRegisters_89__14,
            inputRegisters_89__13,inputRegisters_89__12,inputRegisters_89__11,
            inputRegisters_89__10,inputRegisters_89__9,inputRegisters_89__8,
            inputRegisters_89__7,inputRegisters_89__6,inputRegisters_89__5,
            inputRegisters_89__4,inputRegisters_89__3,inputRegisters_89__2,
            inputRegisters_89__1,inputRegisters_89__0})) ;
    Reg_16 loop1_89_x (.D ({inputRegisters_89__15,inputRegisters_89__14,
           inputRegisters_89__13,inputRegisters_89__12,inputRegisters_89__11,
           inputRegisters_89__10,inputRegisters_89__9,inputRegisters_89__8,
           inputRegisters_89__7,inputRegisters_89__6,inputRegisters_89__5,
           inputRegisters_89__4,inputRegisters_89__3,inputRegisters_89__2,
           inputRegisters_89__1,inputRegisters_89__0}), .en (enableRegister_89)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_89__15,
           registerOutputs_89__14,registerOutputs_89__13,registerOutputs_89__12,
           registerOutputs_89__11,registerOutputs_89__10,registerOutputs_89__9,
           registerOutputs_89__8,registerOutputs_89__7,registerOutputs_89__6,
           registerOutputs_89__5,registerOutputs_89__4,registerOutputs_89__3,
           registerOutputs_89__2,registerOutputs_89__1,registerOutputs_89__0})
           ) ;
    Mux2_16 loop1_90_y (.A ({nx35909,nx36051,nx36193,nx36335,nx36477,nx36619,
            nx36761,nx36903,nx37045,nx37187,nx37329,nx37471,nx37613,nx37755,
            nx37897,nx38039}), .B ({nx33665,nx33805,nx33943,nx34081,nx34219,
            nx34357,nx34495,nx34635,nx34777,nx34919,nx35061,nx35203,nx35345,
            nx35487,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35629), .C ({inputRegisters_90__15,inputRegisters_90__14,
            inputRegisters_90__13,inputRegisters_90__12,inputRegisters_90__11,
            inputRegisters_90__10,inputRegisters_90__9,inputRegisters_90__8,
            inputRegisters_90__7,inputRegisters_90__6,inputRegisters_90__5,
            inputRegisters_90__4,inputRegisters_90__3,inputRegisters_90__2,
            inputRegisters_90__1,inputRegisters_90__0})) ;
    Reg_16 loop1_90_x (.D ({inputRegisters_90__15,inputRegisters_90__14,
           inputRegisters_90__13,inputRegisters_90__12,inputRegisters_90__11,
           inputRegisters_90__10,inputRegisters_90__9,inputRegisters_90__8,
           inputRegisters_90__7,inputRegisters_90__6,inputRegisters_90__5,
           inputRegisters_90__4,inputRegisters_90__3,inputRegisters_90__2,
           inputRegisters_90__1,inputRegisters_90__0}), .en (enableRegister_90)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_90__15,
           registerOutputs_90__14,registerOutputs_90__13,registerOutputs_90__12,
           registerOutputs_90__11,registerOutputs_90__10,registerOutputs_90__9,
           registerOutputs_90__8,registerOutputs_90__7,registerOutputs_90__6,
           registerOutputs_90__5,registerOutputs_90__4,registerOutputs_90__3,
           registerOutputs_90__2,registerOutputs_90__1,registerOutputs_90__0})
           ) ;
    Mux2_16 loop1_91_y (.A ({nx35911,nx36053,nx36195,nx36337,nx36479,nx36621,
            nx36763,nx36905,nx37047,nx37189,nx37331,nx37473,nx37615,nx37757,
            nx37899,nx38041}), .B ({nx33667,nx33805,nx33943,nx34081,nx34219,
            nx34357,nx34495,nx34637,nx34779,nx34921,nx35063,nx35205,nx35347,
            nx35489,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35631), .C ({inputRegisters_91__15,inputRegisters_91__14,
            inputRegisters_91__13,inputRegisters_91__12,inputRegisters_91__11,
            inputRegisters_91__10,inputRegisters_91__9,inputRegisters_91__8,
            inputRegisters_91__7,inputRegisters_91__6,inputRegisters_91__5,
            inputRegisters_91__4,inputRegisters_91__3,inputRegisters_91__2,
            inputRegisters_91__1,inputRegisters_91__0})) ;
    Reg_16 loop1_91_x (.D ({inputRegisters_91__15,inputRegisters_91__14,
           inputRegisters_91__13,inputRegisters_91__12,inputRegisters_91__11,
           inputRegisters_91__10,inputRegisters_91__9,inputRegisters_91__8,
           inputRegisters_91__7,inputRegisters_91__6,inputRegisters_91__5,
           inputRegisters_91__4,inputRegisters_91__3,inputRegisters_91__2,
           inputRegisters_91__1,inputRegisters_91__0}), .en (enableRegister_91)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_91__15,
           registerOutputs_91__14,registerOutputs_91__13,registerOutputs_91__12,
           registerOutputs_91__11,registerOutputs_91__10,registerOutputs_91__9,
           registerOutputs_91__8,registerOutputs_91__7,registerOutputs_91__6,
           registerOutputs_91__5,registerOutputs_91__4,registerOutputs_91__3,
           registerOutputs_91__2,registerOutputs_91__1,registerOutputs_91__0})
           ) ;
    Mux2_16 loop1_92_y (.A ({nx35911,nx36053,nx36195,nx36337,nx36479,nx36621,
            nx36763,nx36905,nx37047,nx37189,nx37331,nx37473,nx37615,nx37757,
            nx37899,nx38041}), .B ({nx33667,nx33805,nx33943,nx34081,nx34219,
            nx34357,nx34497,nx34637,nx34779,nx34921,nx35063,nx35205,nx35347,
            nx35489,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35631), .C ({inputRegisters_92__15,inputRegisters_92__14,
            inputRegisters_92__13,inputRegisters_92__12,inputRegisters_92__11,
            inputRegisters_92__10,inputRegisters_92__9,inputRegisters_92__8,
            inputRegisters_92__7,inputRegisters_92__6,inputRegisters_92__5,
            inputRegisters_92__4,inputRegisters_92__3,inputRegisters_92__2,
            inputRegisters_92__1,inputRegisters_92__0})) ;
    Reg_16 loop1_92_x (.D ({inputRegisters_92__15,inputRegisters_92__14,
           inputRegisters_92__13,inputRegisters_92__12,inputRegisters_92__11,
           inputRegisters_92__10,inputRegisters_92__9,inputRegisters_92__8,
           inputRegisters_92__7,inputRegisters_92__6,inputRegisters_92__5,
           inputRegisters_92__4,inputRegisters_92__3,inputRegisters_92__2,
           inputRegisters_92__1,inputRegisters_92__0}), .en (enableRegister_92)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_92__15,
           registerOutputs_92__14,registerOutputs_92__13,registerOutputs_92__12,
           registerOutputs_92__11,registerOutputs_92__10,registerOutputs_92__9,
           registerOutputs_92__8,registerOutputs_92__7,registerOutputs_92__6,
           registerOutputs_92__5,registerOutputs_92__4,registerOutputs_92__3,
           registerOutputs_92__2,registerOutputs_92__1,registerOutputs_92__0})
           ) ;
    Mux2_16 loop1_93_y (.A ({nx35911,nx36053,nx36195,nx36337,nx36479,nx36621,
            nx36763,nx36905,nx37047,nx37189,nx37331,nx37473,nx37615,nx37757,
            nx37899,nx38041}), .B ({nx33667,nx33805,nx33943,nx34081,nx34219,
            nx34359,nx34497,nx34637,nx34779,nx34921,nx35063,nx35205,nx35347,
            nx35489,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35631), .C ({inputRegisters_93__15,inputRegisters_93__14,
            inputRegisters_93__13,inputRegisters_93__12,inputRegisters_93__11,
            inputRegisters_93__10,inputRegisters_93__9,inputRegisters_93__8,
            inputRegisters_93__7,inputRegisters_93__6,inputRegisters_93__5,
            inputRegisters_93__4,inputRegisters_93__3,inputRegisters_93__2,
            inputRegisters_93__1,inputRegisters_93__0})) ;
    Reg_16 loop1_93_x (.D ({inputRegisters_93__15,inputRegisters_93__14,
           inputRegisters_93__13,inputRegisters_93__12,inputRegisters_93__11,
           inputRegisters_93__10,inputRegisters_93__9,inputRegisters_93__8,
           inputRegisters_93__7,inputRegisters_93__6,inputRegisters_93__5,
           inputRegisters_93__4,inputRegisters_93__3,inputRegisters_93__2,
           inputRegisters_93__1,inputRegisters_93__0}), .en (enableRegister_93)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_93__15,
           registerOutputs_93__14,registerOutputs_93__13,registerOutputs_93__12,
           registerOutputs_93__11,registerOutputs_93__10,registerOutputs_93__9,
           registerOutputs_93__8,registerOutputs_93__7,registerOutputs_93__6,
           registerOutputs_93__5,registerOutputs_93__4,registerOutputs_93__3,
           registerOutputs_93__2,registerOutputs_93__1,registerOutputs_93__0})
           ) ;
    Mux2_16 loop1_94_y (.A ({nx35911,nx36053,nx36195,nx36337,nx36479,nx36621,
            nx36763,nx36905,nx37047,nx37189,nx37331,nx37473,nx37615,nx37757,
            nx37899,nx38041}), .B ({nx33667,nx33805,nx33943,nx34081,nx34221,
            nx34359,nx34497,nx34637,nx34779,nx34921,nx35063,nx35205,nx35347,
            nx35489,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35631), .C ({inputRegisters_94__15,inputRegisters_94__14,
            inputRegisters_94__13,inputRegisters_94__12,inputRegisters_94__11,
            inputRegisters_94__10,inputRegisters_94__9,inputRegisters_94__8,
            inputRegisters_94__7,inputRegisters_94__6,inputRegisters_94__5,
            inputRegisters_94__4,inputRegisters_94__3,inputRegisters_94__2,
            inputRegisters_94__1,inputRegisters_94__0})) ;
    Reg_16 loop1_94_x (.D ({inputRegisters_94__15,inputRegisters_94__14,
           inputRegisters_94__13,inputRegisters_94__12,inputRegisters_94__11,
           inputRegisters_94__10,inputRegisters_94__9,inputRegisters_94__8,
           inputRegisters_94__7,inputRegisters_94__6,inputRegisters_94__5,
           inputRegisters_94__4,inputRegisters_94__3,inputRegisters_94__2,
           inputRegisters_94__1,inputRegisters_94__0}), .en (enableRegister_94)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_94__15,
           registerOutputs_94__14,registerOutputs_94__13,registerOutputs_94__12,
           registerOutputs_94__11,registerOutputs_94__10,registerOutputs_94__9,
           registerOutputs_94__8,registerOutputs_94__7,registerOutputs_94__6,
           registerOutputs_94__5,registerOutputs_94__4,registerOutputs_94__3,
           registerOutputs_94__2,registerOutputs_94__1,registerOutputs_94__0})
           ) ;
    Mux2_16 loop1_95_y (.A ({nx35911,nx36053,nx36195,nx36337,nx36479,nx36621,
            nx36763,nx36905,nx37047,nx37189,nx37331,nx37473,nx37615,nx37757,
            nx37899,nx38041}), .B ({nx33667,nx33805,nx33943,nx34083,nx34221,
            nx34359,nx34497,nx34637,nx34779,nx34921,nx35063,nx35205,nx35347,
            nx35489,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35631), .C ({inputRegisters_95__15,inputRegisters_95__14,
            inputRegisters_95__13,inputRegisters_95__12,inputRegisters_95__11,
            inputRegisters_95__10,inputRegisters_95__9,inputRegisters_95__8,
            inputRegisters_95__7,inputRegisters_95__6,inputRegisters_95__5,
            inputRegisters_95__4,inputRegisters_95__3,inputRegisters_95__2,
            inputRegisters_95__1,inputRegisters_95__0})) ;
    Reg_16 loop1_95_x (.D ({inputRegisters_95__15,inputRegisters_95__14,
           inputRegisters_95__13,inputRegisters_95__12,inputRegisters_95__11,
           inputRegisters_95__10,inputRegisters_95__9,inputRegisters_95__8,
           inputRegisters_95__7,inputRegisters_95__6,inputRegisters_95__5,
           inputRegisters_95__4,inputRegisters_95__3,inputRegisters_95__2,
           inputRegisters_95__1,inputRegisters_95__0}), .en (enableRegister_95)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_95__15,
           registerOutputs_95__14,registerOutputs_95__13,registerOutputs_95__12,
           registerOutputs_95__11,registerOutputs_95__10,registerOutputs_95__9,
           registerOutputs_95__8,registerOutputs_95__7,registerOutputs_95__6,
           registerOutputs_95__5,registerOutputs_95__4,registerOutputs_95__3,
           registerOutputs_95__2,registerOutputs_95__1,registerOutputs_95__0})
           ) ;
    Mux2_16 loop1_96_y (.A ({nx35911,nx36053,nx36195,nx36337,nx36479,nx36621,
            nx36763,nx36905,nx37047,nx37189,nx37331,nx37473,nx37615,nx37757,
            nx37899,nx38041}), .B ({nx33667,nx33805,nx33945,nx34083,nx34221,
            nx34359,nx34497,nx34637,nx34779,nx34921,nx35063,nx35205,nx35347,
            nx35489,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35631), .C ({inputRegisters_96__15,inputRegisters_96__14,
            inputRegisters_96__13,inputRegisters_96__12,inputRegisters_96__11,
            inputRegisters_96__10,inputRegisters_96__9,inputRegisters_96__8,
            inputRegisters_96__7,inputRegisters_96__6,inputRegisters_96__5,
            inputRegisters_96__4,inputRegisters_96__3,inputRegisters_96__2,
            inputRegisters_96__1,inputRegisters_96__0})) ;
    Reg_16 loop1_96_x (.D ({inputRegisters_96__15,inputRegisters_96__14,
           inputRegisters_96__13,inputRegisters_96__12,inputRegisters_96__11,
           inputRegisters_96__10,inputRegisters_96__9,inputRegisters_96__8,
           inputRegisters_96__7,inputRegisters_96__6,inputRegisters_96__5,
           inputRegisters_96__4,inputRegisters_96__3,inputRegisters_96__2,
           inputRegisters_96__1,inputRegisters_96__0}), .en (enableRegister_96)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_96__15,
           registerOutputs_96__14,registerOutputs_96__13,registerOutputs_96__12,
           registerOutputs_96__11,registerOutputs_96__10,registerOutputs_96__9,
           registerOutputs_96__8,registerOutputs_96__7,registerOutputs_96__6,
           registerOutputs_96__5,registerOutputs_96__4,registerOutputs_96__3,
           registerOutputs_96__2,registerOutputs_96__1,registerOutputs_96__0})
           ) ;
    Mux2_16 loop1_97_y (.A ({nx35911,nx36053,nx36195,nx36337,nx36479,nx36621,
            nx36763,nx36905,nx37047,nx37189,nx37331,nx37473,nx37615,nx37757,
            nx37899,nx38041}), .B ({nx33667,nx33807,nx33945,nx34083,nx34221,
            nx34359,nx34497,nx34637,nx34779,nx34921,nx35063,nx35205,nx35347,
            nx35489,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35631), .C ({inputRegisters_97__15,inputRegisters_97__14,
            inputRegisters_97__13,inputRegisters_97__12,inputRegisters_97__11,
            inputRegisters_97__10,inputRegisters_97__9,inputRegisters_97__8,
            inputRegisters_97__7,inputRegisters_97__6,inputRegisters_97__5,
            inputRegisters_97__4,inputRegisters_97__3,inputRegisters_97__2,
            inputRegisters_97__1,inputRegisters_97__0})) ;
    Reg_16 loop1_97_x (.D ({inputRegisters_97__15,inputRegisters_97__14,
           inputRegisters_97__13,inputRegisters_97__12,inputRegisters_97__11,
           inputRegisters_97__10,inputRegisters_97__9,inputRegisters_97__8,
           inputRegisters_97__7,inputRegisters_97__6,inputRegisters_97__5,
           inputRegisters_97__4,inputRegisters_97__3,inputRegisters_97__2,
           inputRegisters_97__1,inputRegisters_97__0}), .en (enableRegister_97)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_97__15,
           registerOutputs_97__14,registerOutputs_97__13,registerOutputs_97__12,
           registerOutputs_97__11,registerOutputs_97__10,registerOutputs_97__9,
           registerOutputs_97__8,registerOutputs_97__7,registerOutputs_97__6,
           registerOutputs_97__5,registerOutputs_97__4,registerOutputs_97__3,
           registerOutputs_97__2,registerOutputs_97__1,registerOutputs_97__0})
           ) ;
    Mux2_16 loop1_98_y (.A ({nx35913,nx36055,nx36197,nx36339,nx36481,nx36623,
            nx36765,nx36907,nx37049,nx37191,nx37333,nx37475,nx37617,nx37759,
            nx37901,nx38043}), .B ({nx33669,nx33807,nx33945,nx34083,nx34221,
            nx34359,nx34497,nx34639,nx34781,nx34923,nx35065,nx35207,nx35349,
            nx35491,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35633), .C ({inputRegisters_98__15,inputRegisters_98__14,
            inputRegisters_98__13,inputRegisters_98__12,inputRegisters_98__11,
            inputRegisters_98__10,inputRegisters_98__9,inputRegisters_98__8,
            inputRegisters_98__7,inputRegisters_98__6,inputRegisters_98__5,
            inputRegisters_98__4,inputRegisters_98__3,inputRegisters_98__2,
            inputRegisters_98__1,inputRegisters_98__0})) ;
    Reg_16 loop1_98_x (.D ({inputRegisters_98__15,inputRegisters_98__14,
           inputRegisters_98__13,inputRegisters_98__12,inputRegisters_98__11,
           inputRegisters_98__10,inputRegisters_98__9,inputRegisters_98__8,
           inputRegisters_98__7,inputRegisters_98__6,inputRegisters_98__5,
           inputRegisters_98__4,inputRegisters_98__3,inputRegisters_98__2,
           inputRegisters_98__1,inputRegisters_98__0}), .en (enableRegister_98)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_98__15,
           registerOutputs_98__14,registerOutputs_98__13,registerOutputs_98__12,
           registerOutputs_98__11,registerOutputs_98__10,registerOutputs_98__9,
           registerOutputs_98__8,registerOutputs_98__7,registerOutputs_98__6,
           registerOutputs_98__5,registerOutputs_98__4,registerOutputs_98__3,
           registerOutputs_98__2,registerOutputs_98__1,registerOutputs_98__0})
           ) ;
    Mux2_16 loop1_99_y (.A ({nx35913,nx36055,nx36197,nx36339,nx36481,nx36623,
            nx36765,nx36907,nx37049,nx37191,nx37333,nx37475,nx37617,nx37759,
            nx37901,nx38043}), .B ({nx33669,nx33807,nx33945,nx34083,nx34221,
            nx34359,nx34499,nx34639,nx34781,nx34923,nx35065,nx35207,nx35349,
            nx35491,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35633), .C ({inputRegisters_99__15,inputRegisters_99__14,
            inputRegisters_99__13,inputRegisters_99__12,inputRegisters_99__11,
            inputRegisters_99__10,inputRegisters_99__9,inputRegisters_99__8,
            inputRegisters_99__7,inputRegisters_99__6,inputRegisters_99__5,
            inputRegisters_99__4,inputRegisters_99__3,inputRegisters_99__2,
            inputRegisters_99__1,inputRegisters_99__0})) ;
    Reg_16 loop1_99_x (.D ({inputRegisters_99__15,inputRegisters_99__14,
           inputRegisters_99__13,inputRegisters_99__12,inputRegisters_99__11,
           inputRegisters_99__10,inputRegisters_99__9,inputRegisters_99__8,
           inputRegisters_99__7,inputRegisters_99__6,inputRegisters_99__5,
           inputRegisters_99__4,inputRegisters_99__3,inputRegisters_99__2,
           inputRegisters_99__1,inputRegisters_99__0}), .en (enableRegister_99)
           , .clk (clk), .rst (resetRegisters), .Q ({registerOutputs_99__15,
           registerOutputs_99__14,registerOutputs_99__13,registerOutputs_99__12,
           registerOutputs_99__11,registerOutputs_99__10,registerOutputs_99__9,
           registerOutputs_99__8,registerOutputs_99__7,registerOutputs_99__6,
           registerOutputs_99__5,registerOutputs_99__4,registerOutputs_99__3,
           registerOutputs_99__2,registerOutputs_99__1,registerOutputs_99__0})
           ) ;
    Mux2_16 loop1_100_y (.A ({nx35913,nx36055,nx36197,nx36339,nx36481,nx36623,
            nx36765,nx36907,nx37049,nx37191,nx37333,nx37475,nx37617,nx37759,
            nx37901,nx38043}), .B ({nx33669,nx33807,nx33945,nx34083,nx34221,
            nx34361,nx34499,nx34639,nx34781,nx34923,nx35065,nx35207,nx35349,
            nx35491,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35633), .C ({inputRegisters_100__15,inputRegisters_100__14,
            inputRegisters_100__13,inputRegisters_100__12,inputRegisters_100__11
            ,inputRegisters_100__10,inputRegisters_100__9,inputRegisters_100__8,
            inputRegisters_100__7,inputRegisters_100__6,inputRegisters_100__5,
            inputRegisters_100__4,inputRegisters_100__3,inputRegisters_100__2,
            inputRegisters_100__1,inputRegisters_100__0})) ;
    Reg_16 loop1_100_x (.D ({inputRegisters_100__15,inputRegisters_100__14,
           inputRegisters_100__13,inputRegisters_100__12,inputRegisters_100__11,
           inputRegisters_100__10,inputRegisters_100__9,inputRegisters_100__8,
           inputRegisters_100__7,inputRegisters_100__6,inputRegisters_100__5,
           inputRegisters_100__4,inputRegisters_100__3,inputRegisters_100__2,
           inputRegisters_100__1,inputRegisters_100__0}), .en (
           enableRegister_100), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_100__15,registerOutputs_100__14,
           registerOutputs_100__13,registerOutputs_100__12,
           registerOutputs_100__11,registerOutputs_100__10,
           registerOutputs_100__9,registerOutputs_100__8,registerOutputs_100__7,
           registerOutputs_100__6,registerOutputs_100__5,registerOutputs_100__4,
           registerOutputs_100__3,registerOutputs_100__2,registerOutputs_100__1,
           registerOutputs_100__0})) ;
    Mux2_16 loop1_101_y (.A ({nx35913,nx36055,nx36197,nx36339,nx36481,nx36623,
            nx36765,nx36907,nx37049,nx37191,nx37333,nx37475,nx37617,nx37759,
            nx37901,nx38043}), .B ({nx33669,nx33807,nx33945,nx34083,nx34223,
            nx34361,nx34499,nx34639,nx34781,nx34923,nx35065,nx35207,nx35349,
            nx35491,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35633), .C ({inputRegisters_101__15,inputRegisters_101__14,
            inputRegisters_101__13,inputRegisters_101__12,inputRegisters_101__11
            ,inputRegisters_101__10,inputRegisters_101__9,inputRegisters_101__8,
            inputRegisters_101__7,inputRegisters_101__6,inputRegisters_101__5,
            inputRegisters_101__4,inputRegisters_101__3,inputRegisters_101__2,
            inputRegisters_101__1,inputRegisters_101__0})) ;
    Reg_16 loop1_101_x (.D ({inputRegisters_101__15,inputRegisters_101__14,
           inputRegisters_101__13,inputRegisters_101__12,inputRegisters_101__11,
           inputRegisters_101__10,inputRegisters_101__9,inputRegisters_101__8,
           inputRegisters_101__7,inputRegisters_101__6,inputRegisters_101__5,
           inputRegisters_101__4,inputRegisters_101__3,inputRegisters_101__2,
           inputRegisters_101__1,inputRegisters_101__0}), .en (
           enableRegister_101), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_101__15,registerOutputs_101__14,
           registerOutputs_101__13,registerOutputs_101__12,
           registerOutputs_101__11,registerOutputs_101__10,
           registerOutputs_101__9,registerOutputs_101__8,registerOutputs_101__7,
           registerOutputs_101__6,registerOutputs_101__5,registerOutputs_101__4,
           registerOutputs_101__3,registerOutputs_101__2,registerOutputs_101__1,
           registerOutputs_101__0})) ;
    Mux2_16 loop1_102_y (.A ({nx35913,nx36055,nx36197,nx36339,nx36481,nx36623,
            nx36765,nx36907,nx37049,nx37191,nx37333,nx37475,nx37617,nx37759,
            nx37901,nx38043}), .B ({nx33669,nx33807,nx33945,nx34085,nx34223,
            nx34361,nx34499,nx34639,nx34781,nx34923,nx35065,nx35207,nx35349,
            nx35491,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35633), .C ({inputRegisters_102__15,inputRegisters_102__14,
            inputRegisters_102__13,inputRegisters_102__12,inputRegisters_102__11
            ,inputRegisters_102__10,inputRegisters_102__9,inputRegisters_102__8,
            inputRegisters_102__7,inputRegisters_102__6,inputRegisters_102__5,
            inputRegisters_102__4,inputRegisters_102__3,inputRegisters_102__2,
            inputRegisters_102__1,inputRegisters_102__0})) ;
    Reg_16 loop1_102_x (.D ({inputRegisters_102__15,inputRegisters_102__14,
           inputRegisters_102__13,inputRegisters_102__12,inputRegisters_102__11,
           inputRegisters_102__10,inputRegisters_102__9,inputRegisters_102__8,
           inputRegisters_102__7,inputRegisters_102__6,inputRegisters_102__5,
           inputRegisters_102__4,inputRegisters_102__3,inputRegisters_102__2,
           inputRegisters_102__1,inputRegisters_102__0}), .en (
           enableRegister_102), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_102__15,registerOutputs_102__14,
           registerOutputs_102__13,registerOutputs_102__12,
           registerOutputs_102__11,registerOutputs_102__10,
           registerOutputs_102__9,registerOutputs_102__8,registerOutputs_102__7,
           registerOutputs_102__6,registerOutputs_102__5,registerOutputs_102__4,
           registerOutputs_102__3,registerOutputs_102__2,registerOutputs_102__1,
           registerOutputs_102__0})) ;
    Mux2_16 loop1_103_y (.A ({nx35913,nx36055,nx36197,nx36339,nx36481,nx36623,
            nx36765,nx36907,nx37049,nx37191,nx37333,nx37475,nx37617,nx37759,
            nx37901,nx38043}), .B ({nx33669,nx33807,nx33947,nx34085,nx34223,
            nx34361,nx34499,nx34639,nx34781,nx34923,nx35065,nx35207,nx35349,
            nx35491,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35633), .C ({inputRegisters_103__15,inputRegisters_103__14,
            inputRegisters_103__13,inputRegisters_103__12,inputRegisters_103__11
            ,inputRegisters_103__10,inputRegisters_103__9,inputRegisters_103__8,
            inputRegisters_103__7,inputRegisters_103__6,inputRegisters_103__5,
            inputRegisters_103__4,inputRegisters_103__3,inputRegisters_103__2,
            inputRegisters_103__1,inputRegisters_103__0})) ;
    Reg_16 loop1_103_x (.D ({inputRegisters_103__15,inputRegisters_103__14,
           inputRegisters_103__13,inputRegisters_103__12,inputRegisters_103__11,
           inputRegisters_103__10,inputRegisters_103__9,inputRegisters_103__8,
           inputRegisters_103__7,inputRegisters_103__6,inputRegisters_103__5,
           inputRegisters_103__4,inputRegisters_103__3,inputRegisters_103__2,
           inputRegisters_103__1,inputRegisters_103__0}), .en (
           enableRegister_103), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_103__15,registerOutputs_103__14,
           registerOutputs_103__13,registerOutputs_103__12,
           registerOutputs_103__11,registerOutputs_103__10,
           registerOutputs_103__9,registerOutputs_103__8,registerOutputs_103__7,
           registerOutputs_103__6,registerOutputs_103__5,registerOutputs_103__4,
           registerOutputs_103__3,registerOutputs_103__2,registerOutputs_103__1,
           registerOutputs_103__0})) ;
    Mux2_16 loop1_104_y (.A ({nx35913,nx36055,nx36197,nx36339,nx36481,nx36623,
            nx36765,nx36907,nx37049,nx37191,nx37333,nx37475,nx37617,nx37759,
            nx37901,nx38043}), .B ({nx33669,nx33809,nx33947,nx34085,nx34223,
            nx34361,nx34499,nx34639,nx34781,nx34923,nx35065,nx35207,nx35349,
            nx35491,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35633), .C ({inputRegisters_104__15,inputRegisters_104__14,
            inputRegisters_104__13,inputRegisters_104__12,inputRegisters_104__11
            ,inputRegisters_104__10,inputRegisters_104__9,inputRegisters_104__8,
            inputRegisters_104__7,inputRegisters_104__6,inputRegisters_104__5,
            inputRegisters_104__4,inputRegisters_104__3,inputRegisters_104__2,
            inputRegisters_104__1,inputRegisters_104__0})) ;
    Reg_16 loop1_104_x (.D ({inputRegisters_104__15,inputRegisters_104__14,
           inputRegisters_104__13,inputRegisters_104__12,inputRegisters_104__11,
           inputRegisters_104__10,inputRegisters_104__9,inputRegisters_104__8,
           inputRegisters_104__7,inputRegisters_104__6,inputRegisters_104__5,
           inputRegisters_104__4,inputRegisters_104__3,inputRegisters_104__2,
           inputRegisters_104__1,inputRegisters_104__0}), .en (
           enableRegister_104), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_104__15,registerOutputs_104__14,
           registerOutputs_104__13,registerOutputs_104__12,
           registerOutputs_104__11,registerOutputs_104__10,
           registerOutputs_104__9,registerOutputs_104__8,registerOutputs_104__7,
           registerOutputs_104__6,registerOutputs_104__5,registerOutputs_104__4,
           registerOutputs_104__3,registerOutputs_104__2,registerOutputs_104__1,
           registerOutputs_104__0})) ;
    Mux2_16 loop1_105_y (.A ({nx35915,nx36057,nx36199,nx36341,nx36483,nx36625,
            nx36767,nx36909,nx37051,nx37193,nx37335,nx37477,nx37619,nx37761,
            nx37903,nx38045}), .B ({nx33671,nx33809,nx33947,nx34085,nx34223,
            nx34361,nx34499,nx34641,nx34783,nx34925,nx35067,nx35209,nx35351,
            nx35493,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35635), .C ({inputRegisters_105__15,inputRegisters_105__14,
            inputRegisters_105__13,inputRegisters_105__12,inputRegisters_105__11
            ,inputRegisters_105__10,inputRegisters_105__9,inputRegisters_105__8,
            inputRegisters_105__7,inputRegisters_105__6,inputRegisters_105__5,
            inputRegisters_105__4,inputRegisters_105__3,inputRegisters_105__2,
            inputRegisters_105__1,inputRegisters_105__0})) ;
    Reg_16 loop1_105_x (.D ({inputRegisters_105__15,inputRegisters_105__14,
           inputRegisters_105__13,inputRegisters_105__12,inputRegisters_105__11,
           inputRegisters_105__10,inputRegisters_105__9,inputRegisters_105__8,
           inputRegisters_105__7,inputRegisters_105__6,inputRegisters_105__5,
           inputRegisters_105__4,inputRegisters_105__3,inputRegisters_105__2,
           inputRegisters_105__1,inputRegisters_105__0}), .en (
           enableRegister_105), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_105__15,registerOutputs_105__14,
           registerOutputs_105__13,registerOutputs_105__12,
           registerOutputs_105__11,registerOutputs_105__10,
           registerOutputs_105__9,registerOutputs_105__8,registerOutputs_105__7,
           registerOutputs_105__6,registerOutputs_105__5,registerOutputs_105__4,
           registerOutputs_105__3,registerOutputs_105__2,registerOutputs_105__1,
           registerOutputs_105__0})) ;
    Mux2_16 loop1_106_y (.A ({nx35915,nx36057,nx36199,nx36341,nx36483,nx36625,
            nx36767,nx36909,nx37051,nx37193,nx37335,nx37477,nx37619,nx37761,
            nx37903,nx38045}), .B ({nx33671,nx33809,nx33947,nx34085,nx34223,
            nx34361,nx34501,nx34641,nx34783,nx34925,nx35067,nx35209,nx35351,
            nx35493,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35635), .C ({inputRegisters_106__15,inputRegisters_106__14,
            inputRegisters_106__13,inputRegisters_106__12,inputRegisters_106__11
            ,inputRegisters_106__10,inputRegisters_106__9,inputRegisters_106__8,
            inputRegisters_106__7,inputRegisters_106__6,inputRegisters_106__5,
            inputRegisters_106__4,inputRegisters_106__3,inputRegisters_106__2,
            inputRegisters_106__1,inputRegisters_106__0})) ;
    Reg_16 loop1_106_x (.D ({inputRegisters_106__15,inputRegisters_106__14,
           inputRegisters_106__13,inputRegisters_106__12,inputRegisters_106__11,
           inputRegisters_106__10,inputRegisters_106__9,inputRegisters_106__8,
           inputRegisters_106__7,inputRegisters_106__6,inputRegisters_106__5,
           inputRegisters_106__4,inputRegisters_106__3,inputRegisters_106__2,
           inputRegisters_106__1,inputRegisters_106__0}), .en (
           enableRegister_106), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_106__15,registerOutputs_106__14,
           registerOutputs_106__13,registerOutputs_106__12,
           registerOutputs_106__11,registerOutputs_106__10,
           registerOutputs_106__9,registerOutputs_106__8,registerOutputs_106__7,
           registerOutputs_106__6,registerOutputs_106__5,registerOutputs_106__4,
           registerOutputs_106__3,registerOutputs_106__2,registerOutputs_106__1,
           registerOutputs_106__0})) ;
    Mux2_16 loop1_107_y (.A ({nx35915,nx36057,nx36199,nx36341,nx36483,nx36625,
            nx36767,nx36909,nx37051,nx37193,nx37335,nx37477,nx37619,nx37761,
            nx37903,nx38045}), .B ({nx33671,nx33809,nx33947,nx34085,nx34223,
            nx34363,nx34501,nx34641,nx34783,nx34925,nx35067,nx35209,nx35351,
            nx35493,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35635), .C ({inputRegisters_107__15,inputRegisters_107__14,
            inputRegisters_107__13,inputRegisters_107__12,inputRegisters_107__11
            ,inputRegisters_107__10,inputRegisters_107__9,inputRegisters_107__8,
            inputRegisters_107__7,inputRegisters_107__6,inputRegisters_107__5,
            inputRegisters_107__4,inputRegisters_107__3,inputRegisters_107__2,
            inputRegisters_107__1,inputRegisters_107__0})) ;
    Reg_16 loop1_107_x (.D ({inputRegisters_107__15,inputRegisters_107__14,
           inputRegisters_107__13,inputRegisters_107__12,inputRegisters_107__11,
           inputRegisters_107__10,inputRegisters_107__9,inputRegisters_107__8,
           inputRegisters_107__7,inputRegisters_107__6,inputRegisters_107__5,
           inputRegisters_107__4,inputRegisters_107__3,inputRegisters_107__2,
           inputRegisters_107__1,inputRegisters_107__0}), .en (
           enableRegister_107), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_107__15,registerOutputs_107__14,
           registerOutputs_107__13,registerOutputs_107__12,
           registerOutputs_107__11,registerOutputs_107__10,
           registerOutputs_107__9,registerOutputs_107__8,registerOutputs_107__7,
           registerOutputs_107__6,registerOutputs_107__5,registerOutputs_107__4,
           registerOutputs_107__3,registerOutputs_107__2,registerOutputs_107__1,
           registerOutputs_107__0})) ;
    Mux2_16 loop1_108_y (.A ({nx35915,nx36057,nx36199,nx36341,nx36483,nx36625,
            nx36767,nx36909,nx37051,nx37193,nx37335,nx37477,nx37619,nx37761,
            nx37903,nx38045}), .B ({nx33671,nx33809,nx33947,nx34085,nx34225,
            nx34363,nx34501,nx34641,nx34783,nx34925,nx35067,nx35209,nx35351,
            nx35493,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35635), .C ({inputRegisters_108__15,inputRegisters_108__14,
            inputRegisters_108__13,inputRegisters_108__12,inputRegisters_108__11
            ,inputRegisters_108__10,inputRegisters_108__9,inputRegisters_108__8,
            inputRegisters_108__7,inputRegisters_108__6,inputRegisters_108__5,
            inputRegisters_108__4,inputRegisters_108__3,inputRegisters_108__2,
            inputRegisters_108__1,inputRegisters_108__0})) ;
    Reg_16 loop1_108_x (.D ({inputRegisters_108__15,inputRegisters_108__14,
           inputRegisters_108__13,inputRegisters_108__12,inputRegisters_108__11,
           inputRegisters_108__10,inputRegisters_108__9,inputRegisters_108__8,
           inputRegisters_108__7,inputRegisters_108__6,inputRegisters_108__5,
           inputRegisters_108__4,inputRegisters_108__3,inputRegisters_108__2,
           inputRegisters_108__1,inputRegisters_108__0}), .en (
           enableRegister_108), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_108__15,registerOutputs_108__14,
           registerOutputs_108__13,registerOutputs_108__12,
           registerOutputs_108__11,registerOutputs_108__10,
           registerOutputs_108__9,registerOutputs_108__8,registerOutputs_108__7,
           registerOutputs_108__6,registerOutputs_108__5,registerOutputs_108__4,
           registerOutputs_108__3,registerOutputs_108__2,registerOutputs_108__1,
           registerOutputs_108__0})) ;
    Mux2_16 loop1_109_y (.A ({nx35915,nx36057,nx36199,nx36341,nx36483,nx36625,
            nx36767,nx36909,nx37051,nx37193,nx37335,nx37477,nx37619,nx37761,
            nx37903,nx38045}), .B ({nx33671,nx33809,nx33947,nx34087,nx34225,
            nx34363,nx34501,nx34641,nx34783,nx34925,nx35067,nx35209,nx35351,
            nx35493,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35635), .C ({inputRegisters_109__15,inputRegisters_109__14,
            inputRegisters_109__13,inputRegisters_109__12,inputRegisters_109__11
            ,inputRegisters_109__10,inputRegisters_109__9,inputRegisters_109__8,
            inputRegisters_109__7,inputRegisters_109__6,inputRegisters_109__5,
            inputRegisters_109__4,inputRegisters_109__3,inputRegisters_109__2,
            inputRegisters_109__1,inputRegisters_109__0})) ;
    Reg_16 loop1_109_x (.D ({inputRegisters_109__15,inputRegisters_109__14,
           inputRegisters_109__13,inputRegisters_109__12,inputRegisters_109__11,
           inputRegisters_109__10,inputRegisters_109__9,inputRegisters_109__8,
           inputRegisters_109__7,inputRegisters_109__6,inputRegisters_109__5,
           inputRegisters_109__4,inputRegisters_109__3,inputRegisters_109__2,
           inputRegisters_109__1,inputRegisters_109__0}), .en (
           enableRegister_109), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_109__15,registerOutputs_109__14,
           registerOutputs_109__13,registerOutputs_109__12,
           registerOutputs_109__11,registerOutputs_109__10,
           registerOutputs_109__9,registerOutputs_109__8,registerOutputs_109__7,
           registerOutputs_109__6,registerOutputs_109__5,registerOutputs_109__4,
           registerOutputs_109__3,registerOutputs_109__2,registerOutputs_109__1,
           registerOutputs_109__0})) ;
    Mux2_16 loop1_110_y (.A ({nx35915,nx36057,nx36199,nx36341,nx36483,nx36625,
            nx36767,nx36909,nx37051,nx37193,nx37335,nx37477,nx37619,nx37761,
            nx37903,nx38045}), .B ({nx33671,nx33809,nx33949,nx34087,nx34225,
            nx34363,nx34501,nx34641,nx34783,nx34925,nx35067,nx35209,nx35351,
            nx35493,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35635), .C ({inputRegisters_110__15,inputRegisters_110__14,
            inputRegisters_110__13,inputRegisters_110__12,inputRegisters_110__11
            ,inputRegisters_110__10,inputRegisters_110__9,inputRegisters_110__8,
            inputRegisters_110__7,inputRegisters_110__6,inputRegisters_110__5,
            inputRegisters_110__4,inputRegisters_110__3,inputRegisters_110__2,
            inputRegisters_110__1,inputRegisters_110__0})) ;
    Reg_16 loop1_110_x (.D ({inputRegisters_110__15,inputRegisters_110__14,
           inputRegisters_110__13,inputRegisters_110__12,inputRegisters_110__11,
           inputRegisters_110__10,inputRegisters_110__9,inputRegisters_110__8,
           inputRegisters_110__7,inputRegisters_110__6,inputRegisters_110__5,
           inputRegisters_110__4,inputRegisters_110__3,inputRegisters_110__2,
           inputRegisters_110__1,inputRegisters_110__0}), .en (
           enableRegister_110), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_110__15,registerOutputs_110__14,
           registerOutputs_110__13,registerOutputs_110__12,
           registerOutputs_110__11,registerOutputs_110__10,
           registerOutputs_110__9,registerOutputs_110__8,registerOutputs_110__7,
           registerOutputs_110__6,registerOutputs_110__5,registerOutputs_110__4,
           registerOutputs_110__3,registerOutputs_110__2,registerOutputs_110__1,
           registerOutputs_110__0})) ;
    Mux2_16 loop1_111_y (.A ({nx35915,nx36057,nx36199,nx36341,nx36483,nx36625,
            nx36767,nx36909,nx37051,nx37193,nx37335,nx37477,nx37619,nx37761,
            nx37903,nx38045}), .B ({nx33671,nx33811,nx33949,nx34087,nx34225,
            nx34363,nx34501,nx34641,nx34783,nx34925,nx35067,nx35209,nx35351,
            nx35493,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35635), .C ({inputRegisters_111__15,inputRegisters_111__14,
            inputRegisters_111__13,inputRegisters_111__12,inputRegisters_111__11
            ,inputRegisters_111__10,inputRegisters_111__9,inputRegisters_111__8,
            inputRegisters_111__7,inputRegisters_111__6,inputRegisters_111__5,
            inputRegisters_111__4,inputRegisters_111__3,inputRegisters_111__2,
            inputRegisters_111__1,inputRegisters_111__0})) ;
    Reg_16 loop1_111_x (.D ({inputRegisters_111__15,inputRegisters_111__14,
           inputRegisters_111__13,inputRegisters_111__12,inputRegisters_111__11,
           inputRegisters_111__10,inputRegisters_111__9,inputRegisters_111__8,
           inputRegisters_111__7,inputRegisters_111__6,inputRegisters_111__5,
           inputRegisters_111__4,inputRegisters_111__3,inputRegisters_111__2,
           inputRegisters_111__1,inputRegisters_111__0}), .en (
           enableRegister_111), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_111__15,registerOutputs_111__14,
           registerOutputs_111__13,registerOutputs_111__12,
           registerOutputs_111__11,registerOutputs_111__10,
           registerOutputs_111__9,registerOutputs_111__8,registerOutputs_111__7,
           registerOutputs_111__6,registerOutputs_111__5,registerOutputs_111__4,
           registerOutputs_111__3,registerOutputs_111__2,registerOutputs_111__1,
           registerOutputs_111__0})) ;
    Mux2_16 loop1_112_y (.A ({nx35917,nx36059,nx36201,nx36343,nx36485,nx36627,
            nx36769,nx36911,nx37053,nx37195,nx37337,nx37479,nx37621,nx37763,
            nx37905,nx38047}), .B ({nx33673,nx33811,nx33949,nx34087,nx34225,
            nx34363,nx34501,nx34643,nx34785,nx34927,nx35069,nx35211,nx35353,
            nx35495,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35637), .C ({inputRegisters_112__15,inputRegisters_112__14,
            inputRegisters_112__13,inputRegisters_112__12,inputRegisters_112__11
            ,inputRegisters_112__10,inputRegisters_112__9,inputRegisters_112__8,
            inputRegisters_112__7,inputRegisters_112__6,inputRegisters_112__5,
            inputRegisters_112__4,inputRegisters_112__3,inputRegisters_112__2,
            inputRegisters_112__1,inputRegisters_112__0})) ;
    Reg_16 loop1_112_x (.D ({inputRegisters_112__15,inputRegisters_112__14,
           inputRegisters_112__13,inputRegisters_112__12,inputRegisters_112__11,
           inputRegisters_112__10,inputRegisters_112__9,inputRegisters_112__8,
           inputRegisters_112__7,inputRegisters_112__6,inputRegisters_112__5,
           inputRegisters_112__4,inputRegisters_112__3,inputRegisters_112__2,
           inputRegisters_112__1,inputRegisters_112__0}), .en (
           enableRegister_112), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_112__15,registerOutputs_112__14,
           registerOutputs_112__13,registerOutputs_112__12,
           registerOutputs_112__11,registerOutputs_112__10,
           registerOutputs_112__9,registerOutputs_112__8,registerOutputs_112__7,
           registerOutputs_112__6,registerOutputs_112__5,registerOutputs_112__4,
           registerOutputs_112__3,registerOutputs_112__2,registerOutputs_112__1,
           registerOutputs_112__0})) ;
    Mux2_16 loop1_113_y (.A ({nx35917,nx36059,nx36201,nx36343,nx36485,nx36627,
            nx36769,nx36911,nx37053,nx37195,nx37337,nx37479,nx37621,nx37763,
            nx37905,nx38047}), .B ({nx33673,nx33811,nx33949,nx34087,nx34225,
            nx34363,nx34503,nx34643,nx34785,nx34927,nx35069,nx35211,nx35353,
            nx35495,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35637), .C ({inputRegisters_113__15,inputRegisters_113__14,
            inputRegisters_113__13,inputRegisters_113__12,inputRegisters_113__11
            ,inputRegisters_113__10,inputRegisters_113__9,inputRegisters_113__8,
            inputRegisters_113__7,inputRegisters_113__6,inputRegisters_113__5,
            inputRegisters_113__4,inputRegisters_113__3,inputRegisters_113__2,
            inputRegisters_113__1,inputRegisters_113__0})) ;
    Reg_16 loop1_113_x (.D ({inputRegisters_113__15,inputRegisters_113__14,
           inputRegisters_113__13,inputRegisters_113__12,inputRegisters_113__11,
           inputRegisters_113__10,inputRegisters_113__9,inputRegisters_113__8,
           inputRegisters_113__7,inputRegisters_113__6,inputRegisters_113__5,
           inputRegisters_113__4,inputRegisters_113__3,inputRegisters_113__2,
           inputRegisters_113__1,inputRegisters_113__0}), .en (
           enableRegister_113), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_113__15,registerOutputs_113__14,
           registerOutputs_113__13,registerOutputs_113__12,
           registerOutputs_113__11,registerOutputs_113__10,
           registerOutputs_113__9,registerOutputs_113__8,registerOutputs_113__7,
           registerOutputs_113__6,registerOutputs_113__5,registerOutputs_113__4,
           registerOutputs_113__3,registerOutputs_113__2,registerOutputs_113__1,
           registerOutputs_113__0})) ;
    Mux2_16 loop1_114_y (.A ({nx35917,nx36059,nx36201,nx36343,nx36485,nx36627,
            nx36769,nx36911,nx37053,nx37195,nx37337,nx37479,nx37621,nx37763,
            nx37905,nx38047}), .B ({nx33673,nx33811,nx33949,nx34087,nx34225,
            nx34365,nx34503,nx34643,nx34785,nx34927,nx35069,nx35211,nx35353,
            nx35495,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35637), .C ({inputRegisters_114__15,inputRegisters_114__14,
            inputRegisters_114__13,inputRegisters_114__12,inputRegisters_114__11
            ,inputRegisters_114__10,inputRegisters_114__9,inputRegisters_114__8,
            inputRegisters_114__7,inputRegisters_114__6,inputRegisters_114__5,
            inputRegisters_114__4,inputRegisters_114__3,inputRegisters_114__2,
            inputRegisters_114__1,inputRegisters_114__0})) ;
    Reg_16 loop1_114_x (.D ({inputRegisters_114__15,inputRegisters_114__14,
           inputRegisters_114__13,inputRegisters_114__12,inputRegisters_114__11,
           inputRegisters_114__10,inputRegisters_114__9,inputRegisters_114__8,
           inputRegisters_114__7,inputRegisters_114__6,inputRegisters_114__5,
           inputRegisters_114__4,inputRegisters_114__3,inputRegisters_114__2,
           inputRegisters_114__1,inputRegisters_114__0}), .en (
           enableRegister_114), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_114__15,registerOutputs_114__14,
           registerOutputs_114__13,registerOutputs_114__12,
           registerOutputs_114__11,registerOutputs_114__10,
           registerOutputs_114__9,registerOutputs_114__8,registerOutputs_114__7,
           registerOutputs_114__6,registerOutputs_114__5,registerOutputs_114__4,
           registerOutputs_114__3,registerOutputs_114__2,registerOutputs_114__1,
           registerOutputs_114__0})) ;
    Mux2_16 loop1_115_y (.A ({nx35917,nx36059,nx36201,nx36343,nx36485,nx36627,
            nx36769,nx36911,nx37053,nx37195,nx37337,nx37479,nx37621,nx37763,
            nx37905,nx38047}), .B ({nx33673,nx33811,nx33949,nx34087,nx34227,
            nx34365,nx34503,nx34643,nx34785,nx34927,nx35069,nx35211,nx35353,
            nx35495,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35637), .C ({inputRegisters_115__15,inputRegisters_115__14,
            inputRegisters_115__13,inputRegisters_115__12,inputRegisters_115__11
            ,inputRegisters_115__10,inputRegisters_115__9,inputRegisters_115__8,
            inputRegisters_115__7,inputRegisters_115__6,inputRegisters_115__5,
            inputRegisters_115__4,inputRegisters_115__3,inputRegisters_115__2,
            inputRegisters_115__1,inputRegisters_115__0})) ;
    Reg_16 loop1_115_x (.D ({inputRegisters_115__15,inputRegisters_115__14,
           inputRegisters_115__13,inputRegisters_115__12,inputRegisters_115__11,
           inputRegisters_115__10,inputRegisters_115__9,inputRegisters_115__8,
           inputRegisters_115__7,inputRegisters_115__6,inputRegisters_115__5,
           inputRegisters_115__4,inputRegisters_115__3,inputRegisters_115__2,
           inputRegisters_115__1,inputRegisters_115__0}), .en (
           enableRegister_115), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_115__15,registerOutputs_115__14,
           registerOutputs_115__13,registerOutputs_115__12,
           registerOutputs_115__11,registerOutputs_115__10,
           registerOutputs_115__9,registerOutputs_115__8,registerOutputs_115__7,
           registerOutputs_115__6,registerOutputs_115__5,registerOutputs_115__4,
           registerOutputs_115__3,registerOutputs_115__2,registerOutputs_115__1,
           registerOutputs_115__0})) ;
    Mux2_16 loop1_116_y (.A ({nx35917,nx36059,nx36201,nx36343,nx36485,nx36627,
            nx36769,nx36911,nx37053,nx37195,nx37337,nx37479,nx37621,nx37763,
            nx37905,nx38047}), .B ({nx33673,nx33811,nx33949,nx34089,nx34227,
            nx34365,nx34503,nx34643,nx34785,nx34927,nx35069,nx35211,nx35353,
            nx35495,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35637), .C ({inputRegisters_116__15,inputRegisters_116__14,
            inputRegisters_116__13,inputRegisters_116__12,inputRegisters_116__11
            ,inputRegisters_116__10,inputRegisters_116__9,inputRegisters_116__8,
            inputRegisters_116__7,inputRegisters_116__6,inputRegisters_116__5,
            inputRegisters_116__4,inputRegisters_116__3,inputRegisters_116__2,
            inputRegisters_116__1,inputRegisters_116__0})) ;
    Reg_16 loop1_116_x (.D ({inputRegisters_116__15,inputRegisters_116__14,
           inputRegisters_116__13,inputRegisters_116__12,inputRegisters_116__11,
           inputRegisters_116__10,inputRegisters_116__9,inputRegisters_116__8,
           inputRegisters_116__7,inputRegisters_116__6,inputRegisters_116__5,
           inputRegisters_116__4,inputRegisters_116__3,inputRegisters_116__2,
           inputRegisters_116__1,inputRegisters_116__0}), .en (
           enableRegister_116), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_116__15,registerOutputs_116__14,
           registerOutputs_116__13,registerOutputs_116__12,
           registerOutputs_116__11,registerOutputs_116__10,
           registerOutputs_116__9,registerOutputs_116__8,registerOutputs_116__7,
           registerOutputs_116__6,registerOutputs_116__5,registerOutputs_116__4,
           registerOutputs_116__3,registerOutputs_116__2,registerOutputs_116__1,
           registerOutputs_116__0})) ;
    Mux2_16 loop1_117_y (.A ({nx35917,nx36059,nx36201,nx36343,nx36485,nx36627,
            nx36769,nx36911,nx37053,nx37195,nx37337,nx37479,nx37621,nx37763,
            nx37905,nx38047}), .B ({nx33673,nx33811,nx33951,nx34089,nx34227,
            nx34365,nx34503,nx34643,nx34785,nx34927,nx35069,nx35211,nx35353,
            nx35495,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35637), .C ({inputRegisters_117__15,inputRegisters_117__14,
            inputRegisters_117__13,inputRegisters_117__12,inputRegisters_117__11
            ,inputRegisters_117__10,inputRegisters_117__9,inputRegisters_117__8,
            inputRegisters_117__7,inputRegisters_117__6,inputRegisters_117__5,
            inputRegisters_117__4,inputRegisters_117__3,inputRegisters_117__2,
            inputRegisters_117__1,inputRegisters_117__0})) ;
    Reg_16 loop1_117_x (.D ({inputRegisters_117__15,inputRegisters_117__14,
           inputRegisters_117__13,inputRegisters_117__12,inputRegisters_117__11,
           inputRegisters_117__10,inputRegisters_117__9,inputRegisters_117__8,
           inputRegisters_117__7,inputRegisters_117__6,inputRegisters_117__5,
           inputRegisters_117__4,inputRegisters_117__3,inputRegisters_117__2,
           inputRegisters_117__1,inputRegisters_117__0}), .en (
           enableRegister_117), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_117__15,registerOutputs_117__14,
           registerOutputs_117__13,registerOutputs_117__12,
           registerOutputs_117__11,registerOutputs_117__10,
           registerOutputs_117__9,registerOutputs_117__8,registerOutputs_117__7,
           registerOutputs_117__6,registerOutputs_117__5,registerOutputs_117__4,
           registerOutputs_117__3,registerOutputs_117__2,registerOutputs_117__1,
           registerOutputs_117__0})) ;
    Mux2_16 loop1_118_y (.A ({nx35917,nx36059,nx36201,nx36343,nx36485,nx36627,
            nx36769,nx36911,nx37053,nx37195,nx37337,nx37479,nx37621,nx37763,
            nx37905,nx38047}), .B ({nx33673,nx33813,nx33951,nx34089,nx34227,
            nx34365,nx34503,nx34643,nx34785,nx34927,nx35069,nx35211,nx35353,
            nx35495,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35637), .C ({inputRegisters_118__15,inputRegisters_118__14,
            inputRegisters_118__13,inputRegisters_118__12,inputRegisters_118__11
            ,inputRegisters_118__10,inputRegisters_118__9,inputRegisters_118__8,
            inputRegisters_118__7,inputRegisters_118__6,inputRegisters_118__5,
            inputRegisters_118__4,inputRegisters_118__3,inputRegisters_118__2,
            inputRegisters_118__1,inputRegisters_118__0})) ;
    Reg_16 loop1_118_x (.D ({inputRegisters_118__15,inputRegisters_118__14,
           inputRegisters_118__13,inputRegisters_118__12,inputRegisters_118__11,
           inputRegisters_118__10,inputRegisters_118__9,inputRegisters_118__8,
           inputRegisters_118__7,inputRegisters_118__6,inputRegisters_118__5,
           inputRegisters_118__4,inputRegisters_118__3,inputRegisters_118__2,
           inputRegisters_118__1,inputRegisters_118__0}), .en (
           enableRegister_118), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_118__15,registerOutputs_118__14,
           registerOutputs_118__13,registerOutputs_118__12,
           registerOutputs_118__11,registerOutputs_118__10,
           registerOutputs_118__9,registerOutputs_118__8,registerOutputs_118__7,
           registerOutputs_118__6,registerOutputs_118__5,registerOutputs_118__4,
           registerOutputs_118__3,registerOutputs_118__2,registerOutputs_118__1,
           registerOutputs_118__0})) ;
    Mux2_16 loop1_119_y (.A ({nx35919,nx36061,nx36203,nx36345,nx36487,nx36629,
            nx36771,nx36913,nx37055,nx37197,nx37339,nx37481,nx37623,nx37765,
            nx37907,nx38049}), .B ({nx33675,nx33813,nx33951,nx34089,nx34227,
            nx34365,nx34503,nx34645,nx34787,nx34929,nx35071,nx35213,nx35355,
            nx35497,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35639), .C ({inputRegisters_119__15,inputRegisters_119__14,
            inputRegisters_119__13,inputRegisters_119__12,inputRegisters_119__11
            ,inputRegisters_119__10,inputRegisters_119__9,inputRegisters_119__8,
            inputRegisters_119__7,inputRegisters_119__6,inputRegisters_119__5,
            inputRegisters_119__4,inputRegisters_119__3,inputRegisters_119__2,
            inputRegisters_119__1,inputRegisters_119__0})) ;
    Reg_16 loop1_119_x (.D ({inputRegisters_119__15,inputRegisters_119__14,
           inputRegisters_119__13,inputRegisters_119__12,inputRegisters_119__11,
           inputRegisters_119__10,inputRegisters_119__9,inputRegisters_119__8,
           inputRegisters_119__7,inputRegisters_119__6,inputRegisters_119__5,
           inputRegisters_119__4,inputRegisters_119__3,inputRegisters_119__2,
           inputRegisters_119__1,inputRegisters_119__0}), .en (
           enableRegister_119), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_119__15,registerOutputs_119__14,
           registerOutputs_119__13,registerOutputs_119__12,
           registerOutputs_119__11,registerOutputs_119__10,
           registerOutputs_119__9,registerOutputs_119__8,registerOutputs_119__7,
           registerOutputs_119__6,registerOutputs_119__5,registerOutputs_119__4,
           registerOutputs_119__3,registerOutputs_119__2,registerOutputs_119__1,
           registerOutputs_119__0})) ;
    Mux2_16 loop1_120_y (.A ({nx35919,nx36061,nx36203,nx36345,nx36487,nx36629,
            nx36771,nx36913,nx37055,nx37197,nx37339,nx37481,nx37623,nx37765,
            nx37907,nx38049}), .B ({nx33675,nx33813,nx33951,nx34089,nx34227,
            nx34365,nx34505,nx34645,nx34787,nx34929,nx35071,nx35213,nx35355,
            nx35497,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35639), .C ({inputRegisters_120__15,inputRegisters_120__14,
            inputRegisters_120__13,inputRegisters_120__12,inputRegisters_120__11
            ,inputRegisters_120__10,inputRegisters_120__9,inputRegisters_120__8,
            inputRegisters_120__7,inputRegisters_120__6,inputRegisters_120__5,
            inputRegisters_120__4,inputRegisters_120__3,inputRegisters_120__2,
            inputRegisters_120__1,inputRegisters_120__0})) ;
    Reg_16 loop1_120_x (.D ({inputRegisters_120__15,inputRegisters_120__14,
           inputRegisters_120__13,inputRegisters_120__12,inputRegisters_120__11,
           inputRegisters_120__10,inputRegisters_120__9,inputRegisters_120__8,
           inputRegisters_120__7,inputRegisters_120__6,inputRegisters_120__5,
           inputRegisters_120__4,inputRegisters_120__3,inputRegisters_120__2,
           inputRegisters_120__1,inputRegisters_120__0}), .en (
           enableRegister_120), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_120__15,registerOutputs_120__14,
           registerOutputs_120__13,registerOutputs_120__12,
           registerOutputs_120__11,registerOutputs_120__10,
           registerOutputs_120__9,registerOutputs_120__8,registerOutputs_120__7,
           registerOutputs_120__6,registerOutputs_120__5,registerOutputs_120__4,
           registerOutputs_120__3,registerOutputs_120__2,registerOutputs_120__1,
           registerOutputs_120__0})) ;
    Mux2_16 loop1_121_y (.A ({nx35919,nx36061,nx36203,nx36345,nx36487,nx36629,
            nx36771,nx36913,nx37055,nx37197,nx37339,nx37481,nx37623,nx37765,
            nx37907,nx38049}), .B ({nx33675,nx33813,nx33951,nx34089,nx34227,
            nx34367,nx34505,nx34645,nx34787,nx34929,nx35071,nx35213,nx35355,
            nx35497,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35639), .C ({inputRegisters_121__15,inputRegisters_121__14,
            inputRegisters_121__13,inputRegisters_121__12,inputRegisters_121__11
            ,inputRegisters_121__10,inputRegisters_121__9,inputRegisters_121__8,
            inputRegisters_121__7,inputRegisters_121__6,inputRegisters_121__5,
            inputRegisters_121__4,inputRegisters_121__3,inputRegisters_121__2,
            inputRegisters_121__1,inputRegisters_121__0})) ;
    Reg_16 loop1_121_x (.D ({inputRegisters_121__15,inputRegisters_121__14,
           inputRegisters_121__13,inputRegisters_121__12,inputRegisters_121__11,
           inputRegisters_121__10,inputRegisters_121__9,inputRegisters_121__8,
           inputRegisters_121__7,inputRegisters_121__6,inputRegisters_121__5,
           inputRegisters_121__4,inputRegisters_121__3,inputRegisters_121__2,
           inputRegisters_121__1,inputRegisters_121__0}), .en (
           enableRegister_121), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_121__15,registerOutputs_121__14,
           registerOutputs_121__13,registerOutputs_121__12,
           registerOutputs_121__11,registerOutputs_121__10,
           registerOutputs_121__9,registerOutputs_121__8,registerOutputs_121__7,
           registerOutputs_121__6,registerOutputs_121__5,registerOutputs_121__4,
           registerOutputs_121__3,registerOutputs_121__2,registerOutputs_121__1,
           registerOutputs_121__0})) ;
    Mux2_16 loop1_122_y (.A ({nx35919,nx36061,nx36203,nx36345,nx36487,nx36629,
            nx36771,nx36913,nx37055,nx37197,nx37339,nx37481,nx37623,nx37765,
            nx37907,nx38049}), .B ({nx33675,nx33813,nx33951,nx34089,nx34229,
            nx34367,nx34505,nx34645,nx34787,nx34929,nx35071,nx35213,nx35355,
            nx35497,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35639), .C ({inputRegisters_122__15,inputRegisters_122__14,
            inputRegisters_122__13,inputRegisters_122__12,inputRegisters_122__11
            ,inputRegisters_122__10,inputRegisters_122__9,inputRegisters_122__8,
            inputRegisters_122__7,inputRegisters_122__6,inputRegisters_122__5,
            inputRegisters_122__4,inputRegisters_122__3,inputRegisters_122__2,
            inputRegisters_122__1,inputRegisters_122__0})) ;
    Reg_16 loop1_122_x (.D ({inputRegisters_122__15,inputRegisters_122__14,
           inputRegisters_122__13,inputRegisters_122__12,inputRegisters_122__11,
           inputRegisters_122__10,inputRegisters_122__9,inputRegisters_122__8,
           inputRegisters_122__7,inputRegisters_122__6,inputRegisters_122__5,
           inputRegisters_122__4,inputRegisters_122__3,inputRegisters_122__2,
           inputRegisters_122__1,inputRegisters_122__0}), .en (
           enableRegister_122), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_122__15,registerOutputs_122__14,
           registerOutputs_122__13,registerOutputs_122__12,
           registerOutputs_122__11,registerOutputs_122__10,
           registerOutputs_122__9,registerOutputs_122__8,registerOutputs_122__7,
           registerOutputs_122__6,registerOutputs_122__5,registerOutputs_122__4,
           registerOutputs_122__3,registerOutputs_122__2,registerOutputs_122__1,
           registerOutputs_122__0})) ;
    Mux2_16 loop1_123_y (.A ({nx35919,nx36061,nx36203,nx36345,nx36487,nx36629,
            nx36771,nx36913,nx37055,nx37197,nx37339,nx37481,nx37623,nx37765,
            nx37907,nx38049}), .B ({nx33675,nx33813,nx33951,nx34091,nx34229,
            nx34367,nx34505,nx34645,nx34787,nx34929,nx35071,nx35213,nx35355,
            nx35497,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35639), .C ({inputRegisters_123__15,inputRegisters_123__14,
            inputRegisters_123__13,inputRegisters_123__12,inputRegisters_123__11
            ,inputRegisters_123__10,inputRegisters_123__9,inputRegisters_123__8,
            inputRegisters_123__7,inputRegisters_123__6,inputRegisters_123__5,
            inputRegisters_123__4,inputRegisters_123__3,inputRegisters_123__2,
            inputRegisters_123__1,inputRegisters_123__0})) ;
    Reg_16 loop1_123_x (.D ({inputRegisters_123__15,inputRegisters_123__14,
           inputRegisters_123__13,inputRegisters_123__12,inputRegisters_123__11,
           inputRegisters_123__10,inputRegisters_123__9,inputRegisters_123__8,
           inputRegisters_123__7,inputRegisters_123__6,inputRegisters_123__5,
           inputRegisters_123__4,inputRegisters_123__3,inputRegisters_123__2,
           inputRegisters_123__1,inputRegisters_123__0}), .en (
           enableRegister_123), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_123__15,registerOutputs_123__14,
           registerOutputs_123__13,registerOutputs_123__12,
           registerOutputs_123__11,registerOutputs_123__10,
           registerOutputs_123__9,registerOutputs_123__8,registerOutputs_123__7,
           registerOutputs_123__6,registerOutputs_123__5,registerOutputs_123__4,
           registerOutputs_123__3,registerOutputs_123__2,registerOutputs_123__1,
           registerOutputs_123__0})) ;
    Mux2_16 loop1_124_y (.A ({nx35919,nx36061,nx36203,nx36345,nx36487,nx36629,
            nx36771,nx36913,nx37055,nx37197,nx37339,nx37481,nx37623,nx37765,
            nx37907,nx38049}), .B ({nx33675,nx33813,nx33953,nx34091,nx34229,
            nx34367,nx34505,nx34645,nx34787,nx34929,nx35071,nx35213,nx35355,
            nx35497,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35639), .C ({inputRegisters_124__15,inputRegisters_124__14,
            inputRegisters_124__13,inputRegisters_124__12,inputRegisters_124__11
            ,inputRegisters_124__10,inputRegisters_124__9,inputRegisters_124__8,
            inputRegisters_124__7,inputRegisters_124__6,inputRegisters_124__5,
            inputRegisters_124__4,inputRegisters_124__3,inputRegisters_124__2,
            inputRegisters_124__1,inputRegisters_124__0})) ;
    Reg_16 loop1_124_x (.D ({inputRegisters_124__15,inputRegisters_124__14,
           inputRegisters_124__13,inputRegisters_124__12,inputRegisters_124__11,
           inputRegisters_124__10,inputRegisters_124__9,inputRegisters_124__8,
           inputRegisters_124__7,inputRegisters_124__6,inputRegisters_124__5,
           inputRegisters_124__4,inputRegisters_124__3,inputRegisters_124__2,
           inputRegisters_124__1,inputRegisters_124__0}), .en (
           enableRegister_124), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_124__15,registerOutputs_124__14,
           registerOutputs_124__13,registerOutputs_124__12,
           registerOutputs_124__11,registerOutputs_124__10,
           registerOutputs_124__9,registerOutputs_124__8,registerOutputs_124__7,
           registerOutputs_124__6,registerOutputs_124__5,registerOutputs_124__4,
           registerOutputs_124__3,registerOutputs_124__2,registerOutputs_124__1,
           registerOutputs_124__0})) ;
    Mux2_16 loop1_125_y (.A ({nx35919,nx36061,nx36203,nx36345,nx36487,nx36629,
            nx36771,nx36913,nx37055,nx37197,nx37339,nx37481,nx37623,nx37765,
            nx37907,nx38049}), .B ({nx33675,nx33815,nx33953,nx34091,nx34229,
            nx34367,nx34505,nx34645,nx34787,nx34929,nx35071,nx35213,nx35355,
            nx35497,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35639), .C ({inputRegisters_125__15,inputRegisters_125__14,
            inputRegisters_125__13,inputRegisters_125__12,inputRegisters_125__11
            ,inputRegisters_125__10,inputRegisters_125__9,inputRegisters_125__8,
            inputRegisters_125__7,inputRegisters_125__6,inputRegisters_125__5,
            inputRegisters_125__4,inputRegisters_125__3,inputRegisters_125__2,
            inputRegisters_125__1,inputRegisters_125__0})) ;
    Reg_16 loop1_125_x (.D ({inputRegisters_125__15,inputRegisters_125__14,
           inputRegisters_125__13,inputRegisters_125__12,inputRegisters_125__11,
           inputRegisters_125__10,inputRegisters_125__9,inputRegisters_125__8,
           inputRegisters_125__7,inputRegisters_125__6,inputRegisters_125__5,
           inputRegisters_125__4,inputRegisters_125__3,inputRegisters_125__2,
           inputRegisters_125__1,inputRegisters_125__0}), .en (
           enableRegister_125), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_125__15,registerOutputs_125__14,
           registerOutputs_125__13,registerOutputs_125__12,
           registerOutputs_125__11,registerOutputs_125__10,
           registerOutputs_125__9,registerOutputs_125__8,registerOutputs_125__7,
           registerOutputs_125__6,registerOutputs_125__5,registerOutputs_125__4,
           registerOutputs_125__3,registerOutputs_125__2,registerOutputs_125__1,
           registerOutputs_125__0})) ;
    Mux2_16 loop1_126_y (.A ({nx35921,nx36063,nx36205,nx36347,nx36489,nx36631,
            nx36773,nx36915,nx37057,nx37199,nx37341,nx37483,nx37625,nx37767,
            nx37909,nx38051}), .B ({nx33677,nx33815,nx33953,nx34091,nx34229,
            nx34367,nx34505,nx34647,nx34789,nx34931,nx35073,nx35215,nx35357,
            nx35499,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35641), .C ({inputRegisters_126__15,inputRegisters_126__14,
            inputRegisters_126__13,inputRegisters_126__12,inputRegisters_126__11
            ,inputRegisters_126__10,inputRegisters_126__9,inputRegisters_126__8,
            inputRegisters_126__7,inputRegisters_126__6,inputRegisters_126__5,
            inputRegisters_126__4,inputRegisters_126__3,inputRegisters_126__2,
            inputRegisters_126__1,inputRegisters_126__0})) ;
    Reg_16 loop1_126_x (.D ({inputRegisters_126__15,inputRegisters_126__14,
           inputRegisters_126__13,inputRegisters_126__12,inputRegisters_126__11,
           inputRegisters_126__10,inputRegisters_126__9,inputRegisters_126__8,
           inputRegisters_126__7,inputRegisters_126__6,inputRegisters_126__5,
           inputRegisters_126__4,inputRegisters_126__3,inputRegisters_126__2,
           inputRegisters_126__1,inputRegisters_126__0}), .en (
           enableRegister_126), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_126__15,registerOutputs_126__14,
           registerOutputs_126__13,registerOutputs_126__12,
           registerOutputs_126__11,registerOutputs_126__10,
           registerOutputs_126__9,registerOutputs_126__8,registerOutputs_126__7,
           registerOutputs_126__6,registerOutputs_126__5,registerOutputs_126__4,
           registerOutputs_126__3,registerOutputs_126__2,registerOutputs_126__1,
           registerOutputs_126__0})) ;
    Mux2_16 loop1_127_y (.A ({nx35921,nx36063,nx36205,nx36347,nx36489,nx36631,
            nx36773,nx36915,nx37057,nx37199,nx37341,nx37483,nx37625,nx37767,
            nx37909,nx38051}), .B ({nx33677,nx33815,nx33953,nx34091,nx34229,
            nx34367,nx34507,nx34647,nx34789,nx34931,nx35073,nx35215,nx35357,
            nx35499,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35641), .C ({inputRegisters_127__15,inputRegisters_127__14,
            inputRegisters_127__13,inputRegisters_127__12,inputRegisters_127__11
            ,inputRegisters_127__10,inputRegisters_127__9,inputRegisters_127__8,
            inputRegisters_127__7,inputRegisters_127__6,inputRegisters_127__5,
            inputRegisters_127__4,inputRegisters_127__3,inputRegisters_127__2,
            inputRegisters_127__1,inputRegisters_127__0})) ;
    Reg_16 loop1_127_x (.D ({inputRegisters_127__15,inputRegisters_127__14,
           inputRegisters_127__13,inputRegisters_127__12,inputRegisters_127__11,
           inputRegisters_127__10,inputRegisters_127__9,inputRegisters_127__8,
           inputRegisters_127__7,inputRegisters_127__6,inputRegisters_127__5,
           inputRegisters_127__4,inputRegisters_127__3,inputRegisters_127__2,
           inputRegisters_127__1,inputRegisters_127__0}), .en (
           enableRegister_127), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_127__15,registerOutputs_127__14,
           registerOutputs_127__13,registerOutputs_127__12,
           registerOutputs_127__11,registerOutputs_127__10,
           registerOutputs_127__9,registerOutputs_127__8,registerOutputs_127__7,
           registerOutputs_127__6,registerOutputs_127__5,registerOutputs_127__4,
           registerOutputs_127__3,registerOutputs_127__2,registerOutputs_127__1,
           registerOutputs_127__0})) ;
    Mux2_16 loop1_128_y (.A ({nx35921,nx36063,nx36205,nx36347,nx36489,nx36631,
            nx36773,nx36915,nx37057,nx37199,nx37341,nx37483,nx37625,nx37767,
            nx37909,nx38051}), .B ({nx33677,nx33815,nx33953,nx34091,nx34229,
            nx34369,nx34507,nx34647,nx34789,nx34931,nx35073,nx35215,nx35357,
            nx35499,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35641), .C ({inputRegisters_128__15,inputRegisters_128__14,
            inputRegisters_128__13,inputRegisters_128__12,inputRegisters_128__11
            ,inputRegisters_128__10,inputRegisters_128__9,inputRegisters_128__8,
            inputRegisters_128__7,inputRegisters_128__6,inputRegisters_128__5,
            inputRegisters_128__4,inputRegisters_128__3,inputRegisters_128__2,
            inputRegisters_128__1,inputRegisters_128__0})) ;
    Reg_16 loop1_128_x (.D ({inputRegisters_128__15,inputRegisters_128__14,
           inputRegisters_128__13,inputRegisters_128__12,inputRegisters_128__11,
           inputRegisters_128__10,inputRegisters_128__9,inputRegisters_128__8,
           inputRegisters_128__7,inputRegisters_128__6,inputRegisters_128__5,
           inputRegisters_128__4,inputRegisters_128__3,inputRegisters_128__2,
           inputRegisters_128__1,inputRegisters_128__0}), .en (
           enableRegister_128), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_128__15,registerOutputs_128__14,
           registerOutputs_128__13,registerOutputs_128__12,
           registerOutputs_128__11,registerOutputs_128__10,
           registerOutputs_128__9,registerOutputs_128__8,registerOutputs_128__7,
           registerOutputs_128__6,registerOutputs_128__5,registerOutputs_128__4,
           registerOutputs_128__3,registerOutputs_128__2,registerOutputs_128__1,
           registerOutputs_128__0})) ;
    Mux2_16 loop1_129_y (.A ({nx35921,nx36063,nx36205,nx36347,nx36489,nx36631,
            nx36773,nx36915,nx37057,nx37199,nx37341,nx37483,nx37625,nx37767,
            nx37909,nx38051}), .B ({nx33677,nx33815,nx33953,nx34091,nx34231,
            nx34369,nx34507,nx34647,nx34789,nx34931,nx35073,nx35215,nx35357,
            nx35499,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35641), .C ({inputRegisters_129__15,inputRegisters_129__14,
            inputRegisters_129__13,inputRegisters_129__12,inputRegisters_129__11
            ,inputRegisters_129__10,inputRegisters_129__9,inputRegisters_129__8,
            inputRegisters_129__7,inputRegisters_129__6,inputRegisters_129__5,
            inputRegisters_129__4,inputRegisters_129__3,inputRegisters_129__2,
            inputRegisters_129__1,inputRegisters_129__0})) ;
    Reg_16 loop1_129_x (.D ({inputRegisters_129__15,inputRegisters_129__14,
           inputRegisters_129__13,inputRegisters_129__12,inputRegisters_129__11,
           inputRegisters_129__10,inputRegisters_129__9,inputRegisters_129__8,
           inputRegisters_129__7,inputRegisters_129__6,inputRegisters_129__5,
           inputRegisters_129__4,inputRegisters_129__3,inputRegisters_129__2,
           inputRegisters_129__1,inputRegisters_129__0}), .en (
           enableRegister_129), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_129__15,registerOutputs_129__14,
           registerOutputs_129__13,registerOutputs_129__12,
           registerOutputs_129__11,registerOutputs_129__10,
           registerOutputs_129__9,registerOutputs_129__8,registerOutputs_129__7,
           registerOutputs_129__6,registerOutputs_129__5,registerOutputs_129__4,
           registerOutputs_129__3,registerOutputs_129__2,registerOutputs_129__1,
           registerOutputs_129__0})) ;
    Mux2_16 loop1_130_y (.A ({nx35921,nx36063,nx36205,nx36347,nx36489,nx36631,
            nx36773,nx36915,nx37057,nx37199,nx37341,nx37483,nx37625,nx37767,
            nx37909,nx38051}), .B ({nx33677,nx33815,nx33953,nx34093,nx34231,
            nx34369,nx34507,nx34647,nx34789,nx34931,nx35073,nx35215,nx35357,
            nx35499,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35641), .C ({inputRegisters_130__15,inputRegisters_130__14,
            inputRegisters_130__13,inputRegisters_130__12,inputRegisters_130__11
            ,inputRegisters_130__10,inputRegisters_130__9,inputRegisters_130__8,
            inputRegisters_130__7,inputRegisters_130__6,inputRegisters_130__5,
            inputRegisters_130__4,inputRegisters_130__3,inputRegisters_130__2,
            inputRegisters_130__1,inputRegisters_130__0})) ;
    Reg_16 loop1_130_x (.D ({inputRegisters_130__15,inputRegisters_130__14,
           inputRegisters_130__13,inputRegisters_130__12,inputRegisters_130__11,
           inputRegisters_130__10,inputRegisters_130__9,inputRegisters_130__8,
           inputRegisters_130__7,inputRegisters_130__6,inputRegisters_130__5,
           inputRegisters_130__4,inputRegisters_130__3,inputRegisters_130__2,
           inputRegisters_130__1,inputRegisters_130__0}), .en (
           enableRegister_130), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_130__15,registerOutputs_130__14,
           registerOutputs_130__13,registerOutputs_130__12,
           registerOutputs_130__11,registerOutputs_130__10,
           registerOutputs_130__9,registerOutputs_130__8,registerOutputs_130__7,
           registerOutputs_130__6,registerOutputs_130__5,registerOutputs_130__4,
           registerOutputs_130__3,registerOutputs_130__2,registerOutputs_130__1,
           registerOutputs_130__0})) ;
    Mux2_16 loop1_131_y (.A ({nx35921,nx36063,nx36205,nx36347,nx36489,nx36631,
            nx36773,nx36915,nx37057,nx37199,nx37341,nx37483,nx37625,nx37767,
            nx37909,nx38051}), .B ({nx33677,nx33815,nx33955,nx34093,nx34231,
            nx34369,nx34507,nx34647,nx34789,nx34931,nx35073,nx35215,nx35357,
            nx35499,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35641), .C ({inputRegisters_131__15,inputRegisters_131__14,
            inputRegisters_131__13,inputRegisters_131__12,inputRegisters_131__11
            ,inputRegisters_131__10,inputRegisters_131__9,inputRegisters_131__8,
            inputRegisters_131__7,inputRegisters_131__6,inputRegisters_131__5,
            inputRegisters_131__4,inputRegisters_131__3,inputRegisters_131__2,
            inputRegisters_131__1,inputRegisters_131__0})) ;
    Reg_16 loop1_131_x (.D ({inputRegisters_131__15,inputRegisters_131__14,
           inputRegisters_131__13,inputRegisters_131__12,inputRegisters_131__11,
           inputRegisters_131__10,inputRegisters_131__9,inputRegisters_131__8,
           inputRegisters_131__7,inputRegisters_131__6,inputRegisters_131__5,
           inputRegisters_131__4,inputRegisters_131__3,inputRegisters_131__2,
           inputRegisters_131__1,inputRegisters_131__0}), .en (
           enableRegister_131), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_131__15,registerOutputs_131__14,
           registerOutputs_131__13,registerOutputs_131__12,
           registerOutputs_131__11,registerOutputs_131__10,
           registerOutputs_131__9,registerOutputs_131__8,registerOutputs_131__7,
           registerOutputs_131__6,registerOutputs_131__5,registerOutputs_131__4,
           registerOutputs_131__3,registerOutputs_131__2,registerOutputs_131__1,
           registerOutputs_131__0})) ;
    Mux2_16 loop1_132_y (.A ({nx35921,nx36063,nx36205,nx36347,nx36489,nx36631,
            nx36773,nx36915,nx37057,nx37199,nx37341,nx37483,nx37625,nx37767,
            nx37909,nx38051}), .B ({nx33677,nx33817,nx33955,nx34093,nx34231,
            nx34369,nx34507,nx34647,nx34789,nx34931,nx35073,nx35215,nx35357,
            nx35499,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35641), .C ({inputRegisters_132__15,inputRegisters_132__14,
            inputRegisters_132__13,inputRegisters_132__12,inputRegisters_132__11
            ,inputRegisters_132__10,inputRegisters_132__9,inputRegisters_132__8,
            inputRegisters_132__7,inputRegisters_132__6,inputRegisters_132__5,
            inputRegisters_132__4,inputRegisters_132__3,inputRegisters_132__2,
            inputRegisters_132__1,inputRegisters_132__0})) ;
    Reg_16 loop1_132_x (.D ({inputRegisters_132__15,inputRegisters_132__14,
           inputRegisters_132__13,inputRegisters_132__12,inputRegisters_132__11,
           inputRegisters_132__10,inputRegisters_132__9,inputRegisters_132__8,
           inputRegisters_132__7,inputRegisters_132__6,inputRegisters_132__5,
           inputRegisters_132__4,inputRegisters_132__3,inputRegisters_132__2,
           inputRegisters_132__1,inputRegisters_132__0}), .en (
           enableRegister_132), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_132__15,registerOutputs_132__14,
           registerOutputs_132__13,registerOutputs_132__12,
           registerOutputs_132__11,registerOutputs_132__10,
           registerOutputs_132__9,registerOutputs_132__8,registerOutputs_132__7,
           registerOutputs_132__6,registerOutputs_132__5,registerOutputs_132__4,
           registerOutputs_132__3,registerOutputs_132__2,registerOutputs_132__1,
           registerOutputs_132__0})) ;
    Mux2_16 loop1_133_y (.A ({nx35923,nx36065,nx36207,nx36349,nx36491,nx36633,
            nx36775,nx36917,nx37059,nx37201,nx37343,nx37485,nx37627,nx37769,
            nx37911,nx38053}), .B ({nx33679,nx33817,nx33955,nx34093,nx34231,
            nx34369,nx34507,nx34649,nx34791,nx34933,nx35075,nx35217,nx35359,
            nx35501,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35643), .C ({inputRegisters_133__15,inputRegisters_133__14,
            inputRegisters_133__13,inputRegisters_133__12,inputRegisters_133__11
            ,inputRegisters_133__10,inputRegisters_133__9,inputRegisters_133__8,
            inputRegisters_133__7,inputRegisters_133__6,inputRegisters_133__5,
            inputRegisters_133__4,inputRegisters_133__3,inputRegisters_133__2,
            inputRegisters_133__1,inputRegisters_133__0})) ;
    Reg_16 loop1_133_x (.D ({inputRegisters_133__15,inputRegisters_133__14,
           inputRegisters_133__13,inputRegisters_133__12,inputRegisters_133__11,
           inputRegisters_133__10,inputRegisters_133__9,inputRegisters_133__8,
           inputRegisters_133__7,inputRegisters_133__6,inputRegisters_133__5,
           inputRegisters_133__4,inputRegisters_133__3,inputRegisters_133__2,
           inputRegisters_133__1,inputRegisters_133__0}), .en (
           enableRegister_133), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_133__15,registerOutputs_133__14,
           registerOutputs_133__13,registerOutputs_133__12,
           registerOutputs_133__11,registerOutputs_133__10,
           registerOutputs_133__9,registerOutputs_133__8,registerOutputs_133__7,
           registerOutputs_133__6,registerOutputs_133__5,registerOutputs_133__4,
           registerOutputs_133__3,registerOutputs_133__2,registerOutputs_133__1,
           registerOutputs_133__0})) ;
    Mux2_16 loop1_134_y (.A ({nx35923,nx36065,nx36207,nx36349,nx36491,nx36633,
            nx36775,nx36917,nx37059,nx37201,nx37343,nx37485,nx37627,nx37769,
            nx37911,nx38053}), .B ({nx33679,nx33817,nx33955,nx34093,nx34231,
            nx34369,nx34509,nx34649,nx34791,nx34933,nx35075,nx35217,nx35359,
            nx35501,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35643), .C ({inputRegisters_134__15,inputRegisters_134__14,
            inputRegisters_134__13,inputRegisters_134__12,inputRegisters_134__11
            ,inputRegisters_134__10,inputRegisters_134__9,inputRegisters_134__8,
            inputRegisters_134__7,inputRegisters_134__6,inputRegisters_134__5,
            inputRegisters_134__4,inputRegisters_134__3,inputRegisters_134__2,
            inputRegisters_134__1,inputRegisters_134__0})) ;
    Reg_16 loop1_134_x (.D ({inputRegisters_134__15,inputRegisters_134__14,
           inputRegisters_134__13,inputRegisters_134__12,inputRegisters_134__11,
           inputRegisters_134__10,inputRegisters_134__9,inputRegisters_134__8,
           inputRegisters_134__7,inputRegisters_134__6,inputRegisters_134__5,
           inputRegisters_134__4,inputRegisters_134__3,inputRegisters_134__2,
           inputRegisters_134__1,inputRegisters_134__0}), .en (
           enableRegister_134), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_134__15,registerOutputs_134__14,
           registerOutputs_134__13,registerOutputs_134__12,
           registerOutputs_134__11,registerOutputs_134__10,
           registerOutputs_134__9,registerOutputs_134__8,registerOutputs_134__7,
           registerOutputs_134__6,registerOutputs_134__5,registerOutputs_134__4,
           registerOutputs_134__3,registerOutputs_134__2,registerOutputs_134__1,
           registerOutputs_134__0})) ;
    Mux2_16 loop1_135_y (.A ({nx35923,nx36065,nx36207,nx36349,nx36491,nx36633,
            nx36775,nx36917,nx37059,nx37201,nx37343,nx37485,nx37627,nx37769,
            nx37911,nx38053}), .B ({nx33679,nx33817,nx33955,nx34093,nx34231,
            nx34371,nx34509,nx34649,nx34791,nx34933,nx35075,nx35217,nx35359,
            nx35501,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35643), .C ({inputRegisters_135__15,inputRegisters_135__14,
            inputRegisters_135__13,inputRegisters_135__12,inputRegisters_135__11
            ,inputRegisters_135__10,inputRegisters_135__9,inputRegisters_135__8,
            inputRegisters_135__7,inputRegisters_135__6,inputRegisters_135__5,
            inputRegisters_135__4,inputRegisters_135__3,inputRegisters_135__2,
            inputRegisters_135__1,inputRegisters_135__0})) ;
    Reg_16 loop1_135_x (.D ({inputRegisters_135__15,inputRegisters_135__14,
           inputRegisters_135__13,inputRegisters_135__12,inputRegisters_135__11,
           inputRegisters_135__10,inputRegisters_135__9,inputRegisters_135__8,
           inputRegisters_135__7,inputRegisters_135__6,inputRegisters_135__5,
           inputRegisters_135__4,inputRegisters_135__3,inputRegisters_135__2,
           inputRegisters_135__1,inputRegisters_135__0}), .en (
           enableRegister_135), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_135__15,registerOutputs_135__14,
           registerOutputs_135__13,registerOutputs_135__12,
           registerOutputs_135__11,registerOutputs_135__10,
           registerOutputs_135__9,registerOutputs_135__8,registerOutputs_135__7,
           registerOutputs_135__6,registerOutputs_135__5,registerOutputs_135__4,
           registerOutputs_135__3,registerOutputs_135__2,registerOutputs_135__1,
           registerOutputs_135__0})) ;
    Mux2_16 loop1_136_y (.A ({nx35923,nx36065,nx36207,nx36349,nx36491,nx36633,
            nx36775,nx36917,nx37059,nx37201,nx37343,nx37485,nx37627,nx37769,
            nx37911,nx38053}), .B ({nx33679,nx33817,nx33955,nx34093,nx34233,
            nx34371,nx34509,nx34649,nx34791,nx34933,nx35075,nx35217,nx35359,
            nx35501,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35643), .C ({inputRegisters_136__15,inputRegisters_136__14,
            inputRegisters_136__13,inputRegisters_136__12,inputRegisters_136__11
            ,inputRegisters_136__10,inputRegisters_136__9,inputRegisters_136__8,
            inputRegisters_136__7,inputRegisters_136__6,inputRegisters_136__5,
            inputRegisters_136__4,inputRegisters_136__3,inputRegisters_136__2,
            inputRegisters_136__1,inputRegisters_136__0})) ;
    Reg_16 loop1_136_x (.D ({inputRegisters_136__15,inputRegisters_136__14,
           inputRegisters_136__13,inputRegisters_136__12,inputRegisters_136__11,
           inputRegisters_136__10,inputRegisters_136__9,inputRegisters_136__8,
           inputRegisters_136__7,inputRegisters_136__6,inputRegisters_136__5,
           inputRegisters_136__4,inputRegisters_136__3,inputRegisters_136__2,
           inputRegisters_136__1,inputRegisters_136__0}), .en (
           enableRegister_136), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_136__15,registerOutputs_136__14,
           registerOutputs_136__13,registerOutputs_136__12,
           registerOutputs_136__11,registerOutputs_136__10,
           registerOutputs_136__9,registerOutputs_136__8,registerOutputs_136__7,
           registerOutputs_136__6,registerOutputs_136__5,registerOutputs_136__4,
           registerOutputs_136__3,registerOutputs_136__2,registerOutputs_136__1,
           registerOutputs_136__0})) ;
    Mux2_16 loop1_137_y (.A ({nx35923,nx36065,nx36207,nx36349,nx36491,nx36633,
            nx36775,nx36917,nx37059,nx37201,nx37343,nx37485,nx37627,nx37769,
            nx37911,nx38053}), .B ({nx33679,nx33817,nx33955,nx34095,nx34233,
            nx34371,nx34509,nx34649,nx34791,nx34933,nx35075,nx35217,nx35359,
            nx35501,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35643), .C ({inputRegisters_137__15,inputRegisters_137__14,
            inputRegisters_137__13,inputRegisters_137__12,inputRegisters_137__11
            ,inputRegisters_137__10,inputRegisters_137__9,inputRegisters_137__8,
            inputRegisters_137__7,inputRegisters_137__6,inputRegisters_137__5,
            inputRegisters_137__4,inputRegisters_137__3,inputRegisters_137__2,
            inputRegisters_137__1,inputRegisters_137__0})) ;
    Reg_16 loop1_137_x (.D ({inputRegisters_137__15,inputRegisters_137__14,
           inputRegisters_137__13,inputRegisters_137__12,inputRegisters_137__11,
           inputRegisters_137__10,inputRegisters_137__9,inputRegisters_137__8,
           inputRegisters_137__7,inputRegisters_137__6,inputRegisters_137__5,
           inputRegisters_137__4,inputRegisters_137__3,inputRegisters_137__2,
           inputRegisters_137__1,inputRegisters_137__0}), .en (
           enableRegister_137), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_137__15,registerOutputs_137__14,
           registerOutputs_137__13,registerOutputs_137__12,
           registerOutputs_137__11,registerOutputs_137__10,
           registerOutputs_137__9,registerOutputs_137__8,registerOutputs_137__7,
           registerOutputs_137__6,registerOutputs_137__5,registerOutputs_137__4,
           registerOutputs_137__3,registerOutputs_137__2,registerOutputs_137__1,
           registerOutputs_137__0})) ;
    Mux2_16 loop1_138_y (.A ({nx35923,nx36065,nx36207,nx36349,nx36491,nx36633,
            nx36775,nx36917,nx37059,nx37201,nx37343,nx37485,nx37627,nx37769,
            nx37911,nx38053}), .B ({nx33679,nx33817,nx33957,nx34095,nx34233,
            nx34371,nx34509,nx34649,nx34791,nx34933,nx35075,nx35217,nx35359,
            nx35501,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35643), .C ({inputRegisters_138__15,inputRegisters_138__14,
            inputRegisters_138__13,inputRegisters_138__12,inputRegisters_138__11
            ,inputRegisters_138__10,inputRegisters_138__9,inputRegisters_138__8,
            inputRegisters_138__7,inputRegisters_138__6,inputRegisters_138__5,
            inputRegisters_138__4,inputRegisters_138__3,inputRegisters_138__2,
            inputRegisters_138__1,inputRegisters_138__0})) ;
    Reg_16 loop1_138_x (.D ({inputRegisters_138__15,inputRegisters_138__14,
           inputRegisters_138__13,inputRegisters_138__12,inputRegisters_138__11,
           inputRegisters_138__10,inputRegisters_138__9,inputRegisters_138__8,
           inputRegisters_138__7,inputRegisters_138__6,inputRegisters_138__5,
           inputRegisters_138__4,inputRegisters_138__3,inputRegisters_138__2,
           inputRegisters_138__1,inputRegisters_138__0}), .en (
           enableRegister_138), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_138__15,registerOutputs_138__14,
           registerOutputs_138__13,registerOutputs_138__12,
           registerOutputs_138__11,registerOutputs_138__10,
           registerOutputs_138__9,registerOutputs_138__8,registerOutputs_138__7,
           registerOutputs_138__6,registerOutputs_138__5,registerOutputs_138__4,
           registerOutputs_138__3,registerOutputs_138__2,registerOutputs_138__1,
           registerOutputs_138__0})) ;
    Mux2_16 loop1_139_y (.A ({nx35923,nx36065,nx36207,nx36349,nx36491,nx36633,
            nx36775,nx36917,nx37059,nx37201,nx37343,nx37485,nx37627,nx37769,
            nx37911,nx38053}), .B ({nx33679,nx33819,nx33957,nx34095,nx34233,
            nx34371,nx34509,nx34649,nx34791,nx34933,nx35075,nx35217,nx35359,
            nx35501,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35643), .C ({inputRegisters_139__15,inputRegisters_139__14,
            inputRegisters_139__13,inputRegisters_139__12,inputRegisters_139__11
            ,inputRegisters_139__10,inputRegisters_139__9,inputRegisters_139__8,
            inputRegisters_139__7,inputRegisters_139__6,inputRegisters_139__5,
            inputRegisters_139__4,inputRegisters_139__3,inputRegisters_139__2,
            inputRegisters_139__1,inputRegisters_139__0})) ;
    Reg_16 loop1_139_x (.D ({inputRegisters_139__15,inputRegisters_139__14,
           inputRegisters_139__13,inputRegisters_139__12,inputRegisters_139__11,
           inputRegisters_139__10,inputRegisters_139__9,inputRegisters_139__8,
           inputRegisters_139__7,inputRegisters_139__6,inputRegisters_139__5,
           inputRegisters_139__4,inputRegisters_139__3,inputRegisters_139__2,
           inputRegisters_139__1,inputRegisters_139__0}), .en (
           enableRegister_139), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_139__15,registerOutputs_139__14,
           registerOutputs_139__13,registerOutputs_139__12,
           registerOutputs_139__11,registerOutputs_139__10,
           registerOutputs_139__9,registerOutputs_139__8,registerOutputs_139__7,
           registerOutputs_139__6,registerOutputs_139__5,registerOutputs_139__4,
           registerOutputs_139__3,registerOutputs_139__2,registerOutputs_139__1,
           registerOutputs_139__0})) ;
    Mux2_16 loop1_140_y (.A ({nx35925,nx36067,nx36209,nx36351,nx36493,nx36635,
            nx36777,nx36919,nx37061,nx37203,nx37345,nx37487,nx37629,nx37771,
            nx37913,nx38055}), .B ({nx33681,nx33819,nx33957,nx34095,nx34233,
            nx34371,nx34509,nx34651,nx34793,nx34935,nx35077,nx35219,nx35361,
            nx35503,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35645), .C ({inputRegisters_140__15,inputRegisters_140__14,
            inputRegisters_140__13,inputRegisters_140__12,inputRegisters_140__11
            ,inputRegisters_140__10,inputRegisters_140__9,inputRegisters_140__8,
            inputRegisters_140__7,inputRegisters_140__6,inputRegisters_140__5,
            inputRegisters_140__4,inputRegisters_140__3,inputRegisters_140__2,
            inputRegisters_140__1,inputRegisters_140__0})) ;
    Reg_16 loop1_140_x (.D ({inputRegisters_140__15,inputRegisters_140__14,
           inputRegisters_140__13,inputRegisters_140__12,inputRegisters_140__11,
           inputRegisters_140__10,inputRegisters_140__9,inputRegisters_140__8,
           inputRegisters_140__7,inputRegisters_140__6,inputRegisters_140__5,
           inputRegisters_140__4,inputRegisters_140__3,inputRegisters_140__2,
           inputRegisters_140__1,inputRegisters_140__0}), .en (
           enableRegister_140), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_140__15,registerOutputs_140__14,
           registerOutputs_140__13,registerOutputs_140__12,
           registerOutputs_140__11,registerOutputs_140__10,
           registerOutputs_140__9,registerOutputs_140__8,registerOutputs_140__7,
           registerOutputs_140__6,registerOutputs_140__5,registerOutputs_140__4,
           registerOutputs_140__3,registerOutputs_140__2,registerOutputs_140__1,
           registerOutputs_140__0})) ;
    Mux2_16 loop1_141_y (.A ({nx35925,nx36067,nx36209,nx36351,nx36493,nx36635,
            nx36777,nx36919,nx37061,nx37203,nx37345,nx37487,nx37629,nx37771,
            nx37913,nx38055}), .B ({nx33681,nx33819,nx33957,nx34095,nx34233,
            nx34371,nx34511,nx34651,nx34793,nx34935,nx35077,nx35219,nx35361,
            nx35503,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35645), .C ({inputRegisters_141__15,inputRegisters_141__14,
            inputRegisters_141__13,inputRegisters_141__12,inputRegisters_141__11
            ,inputRegisters_141__10,inputRegisters_141__9,inputRegisters_141__8,
            inputRegisters_141__7,inputRegisters_141__6,inputRegisters_141__5,
            inputRegisters_141__4,inputRegisters_141__3,inputRegisters_141__2,
            inputRegisters_141__1,inputRegisters_141__0})) ;
    Reg_16 loop1_141_x (.D ({inputRegisters_141__15,inputRegisters_141__14,
           inputRegisters_141__13,inputRegisters_141__12,inputRegisters_141__11,
           inputRegisters_141__10,inputRegisters_141__9,inputRegisters_141__8,
           inputRegisters_141__7,inputRegisters_141__6,inputRegisters_141__5,
           inputRegisters_141__4,inputRegisters_141__3,inputRegisters_141__2,
           inputRegisters_141__1,inputRegisters_141__0}), .en (
           enableRegister_141), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_141__15,registerOutputs_141__14,
           registerOutputs_141__13,registerOutputs_141__12,
           registerOutputs_141__11,registerOutputs_141__10,
           registerOutputs_141__9,registerOutputs_141__8,registerOutputs_141__7,
           registerOutputs_141__6,registerOutputs_141__5,registerOutputs_141__4,
           registerOutputs_141__3,registerOutputs_141__2,registerOutputs_141__1,
           registerOutputs_141__0})) ;
    Mux2_16 loop1_142_y (.A ({nx35925,nx36067,nx36209,nx36351,nx36493,nx36635,
            nx36777,nx36919,nx37061,nx37203,nx37345,nx37487,nx37629,nx37771,
            nx37913,nx38055}), .B ({nx33681,nx33819,nx33957,nx34095,nx34233,
            nx34373,nx34511,nx34651,nx34793,nx34935,nx35077,nx35219,nx35361,
            nx35503,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35645), .C ({inputRegisters_142__15,inputRegisters_142__14,
            inputRegisters_142__13,inputRegisters_142__12,inputRegisters_142__11
            ,inputRegisters_142__10,inputRegisters_142__9,inputRegisters_142__8,
            inputRegisters_142__7,inputRegisters_142__6,inputRegisters_142__5,
            inputRegisters_142__4,inputRegisters_142__3,inputRegisters_142__2,
            inputRegisters_142__1,inputRegisters_142__0})) ;
    Reg_16 loop1_142_x (.D ({inputRegisters_142__15,inputRegisters_142__14,
           inputRegisters_142__13,inputRegisters_142__12,inputRegisters_142__11,
           inputRegisters_142__10,inputRegisters_142__9,inputRegisters_142__8,
           inputRegisters_142__7,inputRegisters_142__6,inputRegisters_142__5,
           inputRegisters_142__4,inputRegisters_142__3,inputRegisters_142__2,
           inputRegisters_142__1,inputRegisters_142__0}), .en (
           enableRegister_142), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_142__15,registerOutputs_142__14,
           registerOutputs_142__13,registerOutputs_142__12,
           registerOutputs_142__11,registerOutputs_142__10,
           registerOutputs_142__9,registerOutputs_142__8,registerOutputs_142__7,
           registerOutputs_142__6,registerOutputs_142__5,registerOutputs_142__4,
           registerOutputs_142__3,registerOutputs_142__2,registerOutputs_142__1,
           registerOutputs_142__0})) ;
    Mux2_16 loop1_143_y (.A ({nx35925,nx36067,nx36209,nx36351,nx36493,nx36635,
            nx36777,nx36919,nx37061,nx37203,nx37345,nx37487,nx37629,nx37771,
            nx37913,nx38055}), .B ({nx33681,nx33819,nx33957,nx34095,nx34235,
            nx34373,nx34511,nx34651,nx34793,nx34935,nx35077,nx35219,nx35361,
            nx35503,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35645), .C ({inputRegisters_143__15,inputRegisters_143__14,
            inputRegisters_143__13,inputRegisters_143__12,inputRegisters_143__11
            ,inputRegisters_143__10,inputRegisters_143__9,inputRegisters_143__8,
            inputRegisters_143__7,inputRegisters_143__6,inputRegisters_143__5,
            inputRegisters_143__4,inputRegisters_143__3,inputRegisters_143__2,
            inputRegisters_143__1,inputRegisters_143__0})) ;
    Reg_16 loop1_143_x (.D ({inputRegisters_143__15,inputRegisters_143__14,
           inputRegisters_143__13,inputRegisters_143__12,inputRegisters_143__11,
           inputRegisters_143__10,inputRegisters_143__9,inputRegisters_143__8,
           inputRegisters_143__7,inputRegisters_143__6,inputRegisters_143__5,
           inputRegisters_143__4,inputRegisters_143__3,inputRegisters_143__2,
           inputRegisters_143__1,inputRegisters_143__0}), .en (
           enableRegister_143), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_143__15,registerOutputs_143__14,
           registerOutputs_143__13,registerOutputs_143__12,
           registerOutputs_143__11,registerOutputs_143__10,
           registerOutputs_143__9,registerOutputs_143__8,registerOutputs_143__7,
           registerOutputs_143__6,registerOutputs_143__5,registerOutputs_143__4,
           registerOutputs_143__3,registerOutputs_143__2,registerOutputs_143__1,
           registerOutputs_143__0})) ;
    Mux2_16 loop1_144_y (.A ({nx35925,nx36067,nx36209,nx36351,nx36493,nx36635,
            nx36777,nx36919,nx37061,nx37203,nx37345,nx37487,nx37629,nx37771,
            nx37913,nx38055}), .B ({nx33681,nx33819,nx33957,nx34097,nx34235,
            nx34373,nx34511,nx34651,nx34793,nx34935,nx35077,nx35219,nx35361,
            nx35503,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35645), .C ({inputRegisters_144__15,inputRegisters_144__14,
            inputRegisters_144__13,inputRegisters_144__12,inputRegisters_144__11
            ,inputRegisters_144__10,inputRegisters_144__9,inputRegisters_144__8,
            inputRegisters_144__7,inputRegisters_144__6,inputRegisters_144__5,
            inputRegisters_144__4,inputRegisters_144__3,inputRegisters_144__2,
            inputRegisters_144__1,inputRegisters_144__0})) ;
    Reg_16 loop1_144_x (.D ({inputRegisters_144__15,inputRegisters_144__14,
           inputRegisters_144__13,inputRegisters_144__12,inputRegisters_144__11,
           inputRegisters_144__10,inputRegisters_144__9,inputRegisters_144__8,
           inputRegisters_144__7,inputRegisters_144__6,inputRegisters_144__5,
           inputRegisters_144__4,inputRegisters_144__3,inputRegisters_144__2,
           inputRegisters_144__1,inputRegisters_144__0}), .en (
           enableRegister_144), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_144__15,registerOutputs_144__14,
           registerOutputs_144__13,registerOutputs_144__12,
           registerOutputs_144__11,registerOutputs_144__10,
           registerOutputs_144__9,registerOutputs_144__8,registerOutputs_144__7,
           registerOutputs_144__6,registerOutputs_144__5,registerOutputs_144__4,
           registerOutputs_144__3,registerOutputs_144__2,registerOutputs_144__1,
           registerOutputs_144__0})) ;
    Mux2_16 loop1_145_y (.A ({nx35925,nx36067,nx36209,nx36351,nx36493,nx36635,
            nx36777,nx36919,nx37061,nx37203,nx37345,nx37487,nx37629,nx37771,
            nx37913,nx38055}), .B ({nx33681,nx33819,nx33959,nx34097,nx34235,
            nx34373,nx34511,nx34651,nx34793,nx34935,nx35077,nx35219,nx35361,
            nx35503,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35645), .C ({inputRegisters_145__15,inputRegisters_145__14,
            inputRegisters_145__13,inputRegisters_145__12,inputRegisters_145__11
            ,inputRegisters_145__10,inputRegisters_145__9,inputRegisters_145__8,
            inputRegisters_145__7,inputRegisters_145__6,inputRegisters_145__5,
            inputRegisters_145__4,inputRegisters_145__3,inputRegisters_145__2,
            inputRegisters_145__1,inputRegisters_145__0})) ;
    Reg_16 loop1_145_x (.D ({inputRegisters_145__15,inputRegisters_145__14,
           inputRegisters_145__13,inputRegisters_145__12,inputRegisters_145__11,
           inputRegisters_145__10,inputRegisters_145__9,inputRegisters_145__8,
           inputRegisters_145__7,inputRegisters_145__6,inputRegisters_145__5,
           inputRegisters_145__4,inputRegisters_145__3,inputRegisters_145__2,
           inputRegisters_145__1,inputRegisters_145__0}), .en (
           enableRegister_145), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_145__15,registerOutputs_145__14,
           registerOutputs_145__13,registerOutputs_145__12,
           registerOutputs_145__11,registerOutputs_145__10,
           registerOutputs_145__9,registerOutputs_145__8,registerOutputs_145__7,
           registerOutputs_145__6,registerOutputs_145__5,registerOutputs_145__4,
           registerOutputs_145__3,registerOutputs_145__2,registerOutputs_145__1,
           registerOutputs_145__0})) ;
    Mux2_16 loop1_146_y (.A ({nx35925,nx36067,nx36209,nx36351,nx36493,nx36635,
            nx36777,nx36919,nx37061,nx37203,nx37345,nx37487,nx37629,nx37771,
            nx37913,nx38055}), .B ({nx33681,nx33821,nx33959,nx34097,nx34235,
            nx34373,nx34511,nx34651,nx34793,nx34935,nx35077,nx35219,nx35361,
            nx35503,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35645), .C ({inputRegisters_146__15,inputRegisters_146__14,
            inputRegisters_146__13,inputRegisters_146__12,inputRegisters_146__11
            ,inputRegisters_146__10,inputRegisters_146__9,inputRegisters_146__8,
            inputRegisters_146__7,inputRegisters_146__6,inputRegisters_146__5,
            inputRegisters_146__4,inputRegisters_146__3,inputRegisters_146__2,
            inputRegisters_146__1,inputRegisters_146__0})) ;
    Reg_16 loop1_146_x (.D ({inputRegisters_146__15,inputRegisters_146__14,
           inputRegisters_146__13,inputRegisters_146__12,inputRegisters_146__11,
           inputRegisters_146__10,inputRegisters_146__9,inputRegisters_146__8,
           inputRegisters_146__7,inputRegisters_146__6,inputRegisters_146__5,
           inputRegisters_146__4,inputRegisters_146__3,inputRegisters_146__2,
           inputRegisters_146__1,inputRegisters_146__0}), .en (
           enableRegister_146), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_146__15,registerOutputs_146__14,
           registerOutputs_146__13,registerOutputs_146__12,
           registerOutputs_146__11,registerOutputs_146__10,
           registerOutputs_146__9,registerOutputs_146__8,registerOutputs_146__7,
           registerOutputs_146__6,registerOutputs_146__5,registerOutputs_146__4,
           registerOutputs_146__3,registerOutputs_146__2,registerOutputs_146__1,
           registerOutputs_146__0})) ;
    Mux2_16 loop1_147_y (.A ({nx35927,nx36069,nx36211,nx36353,nx36495,nx36637,
            nx36779,nx36921,nx37063,nx37205,nx37347,nx37489,nx37631,nx37773,
            nx37915,nx38057}), .B ({nx33683,nx33821,nx33959,nx34097,nx34235,
            nx34373,nx34511,nx34653,nx34795,nx34937,nx35079,nx35221,nx35363,
            nx35505,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35647), .C ({inputRegisters_147__15,inputRegisters_147__14,
            inputRegisters_147__13,inputRegisters_147__12,inputRegisters_147__11
            ,inputRegisters_147__10,inputRegisters_147__9,inputRegisters_147__8,
            inputRegisters_147__7,inputRegisters_147__6,inputRegisters_147__5,
            inputRegisters_147__4,inputRegisters_147__3,inputRegisters_147__2,
            inputRegisters_147__1,inputRegisters_147__0})) ;
    Reg_16 loop1_147_x (.D ({inputRegisters_147__15,inputRegisters_147__14,
           inputRegisters_147__13,inputRegisters_147__12,inputRegisters_147__11,
           inputRegisters_147__10,inputRegisters_147__9,inputRegisters_147__8,
           inputRegisters_147__7,inputRegisters_147__6,inputRegisters_147__5,
           inputRegisters_147__4,inputRegisters_147__3,inputRegisters_147__2,
           inputRegisters_147__1,inputRegisters_147__0}), .en (
           enableRegister_147), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_147__15,registerOutputs_147__14,
           registerOutputs_147__13,registerOutputs_147__12,
           registerOutputs_147__11,registerOutputs_147__10,
           registerOutputs_147__9,registerOutputs_147__8,registerOutputs_147__7,
           registerOutputs_147__6,registerOutputs_147__5,registerOutputs_147__4,
           registerOutputs_147__3,registerOutputs_147__2,registerOutputs_147__1,
           registerOutputs_147__0})) ;
    Mux2_16 loop1_148_y (.A ({nx35927,nx36069,nx36211,nx36353,nx36495,nx36637,
            nx36779,nx36921,nx37063,nx37205,nx37347,nx37489,nx37631,nx37773,
            nx37915,nx38057}), .B ({nx33683,nx33821,nx33959,nx34097,nx34235,
            nx34373,nx34513,nx34653,nx34795,nx34937,nx35079,nx35221,nx35363,
            nx35505,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35647), .C ({inputRegisters_148__15,inputRegisters_148__14,
            inputRegisters_148__13,inputRegisters_148__12,inputRegisters_148__11
            ,inputRegisters_148__10,inputRegisters_148__9,inputRegisters_148__8,
            inputRegisters_148__7,inputRegisters_148__6,inputRegisters_148__5,
            inputRegisters_148__4,inputRegisters_148__3,inputRegisters_148__2,
            inputRegisters_148__1,inputRegisters_148__0})) ;
    Reg_16 loop1_148_x (.D ({inputRegisters_148__15,inputRegisters_148__14,
           inputRegisters_148__13,inputRegisters_148__12,inputRegisters_148__11,
           inputRegisters_148__10,inputRegisters_148__9,inputRegisters_148__8,
           inputRegisters_148__7,inputRegisters_148__6,inputRegisters_148__5,
           inputRegisters_148__4,inputRegisters_148__3,inputRegisters_148__2,
           inputRegisters_148__1,inputRegisters_148__0}), .en (
           enableRegister_148), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_148__15,registerOutputs_148__14,
           registerOutputs_148__13,registerOutputs_148__12,
           registerOutputs_148__11,registerOutputs_148__10,
           registerOutputs_148__9,registerOutputs_148__8,registerOutputs_148__7,
           registerOutputs_148__6,registerOutputs_148__5,registerOutputs_148__4,
           registerOutputs_148__3,registerOutputs_148__2,registerOutputs_148__1,
           registerOutputs_148__0})) ;
    Mux2_16 loop1_149_y (.A ({nx35927,nx36069,nx36211,nx36353,nx36495,nx36637,
            nx36779,nx36921,nx37063,nx37205,nx37347,nx37489,nx37631,nx37773,
            nx37915,nx38057}), .B ({nx33683,nx33821,nx33959,nx34097,nx34235,
            nx34375,nx34513,nx34653,nx34795,nx34937,nx35079,nx35221,nx35363,
            nx35505,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35647), .C ({inputRegisters_149__15,inputRegisters_149__14,
            inputRegisters_149__13,inputRegisters_149__12,inputRegisters_149__11
            ,inputRegisters_149__10,inputRegisters_149__9,inputRegisters_149__8,
            inputRegisters_149__7,inputRegisters_149__6,inputRegisters_149__5,
            inputRegisters_149__4,inputRegisters_149__3,inputRegisters_149__2,
            inputRegisters_149__1,inputRegisters_149__0})) ;
    Reg_16 loop1_149_x (.D ({inputRegisters_149__15,inputRegisters_149__14,
           inputRegisters_149__13,inputRegisters_149__12,inputRegisters_149__11,
           inputRegisters_149__10,inputRegisters_149__9,inputRegisters_149__8,
           inputRegisters_149__7,inputRegisters_149__6,inputRegisters_149__5,
           inputRegisters_149__4,inputRegisters_149__3,inputRegisters_149__2,
           inputRegisters_149__1,inputRegisters_149__0}), .en (
           enableRegister_149), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_149__15,registerOutputs_149__14,
           registerOutputs_149__13,registerOutputs_149__12,
           registerOutputs_149__11,registerOutputs_149__10,
           registerOutputs_149__9,registerOutputs_149__8,registerOutputs_149__7,
           registerOutputs_149__6,registerOutputs_149__5,registerOutputs_149__4,
           registerOutputs_149__3,registerOutputs_149__2,registerOutputs_149__1,
           registerOutputs_149__0})) ;
    Mux2_16 loop1_150_y (.A ({nx35927,nx36069,nx36211,nx36353,nx36495,nx36637,
            nx36779,nx36921,nx37063,nx37205,nx37347,nx37489,nx37631,nx37773,
            nx37915,nx38057}), .B ({nx33683,nx33821,nx33959,nx34097,nx34237,
            nx34375,nx34513,nx34653,nx34795,nx34937,nx35079,nx35221,nx35363,
            nx35505,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35647), .C ({inputRegisters_150__15,inputRegisters_150__14,
            inputRegisters_150__13,inputRegisters_150__12,inputRegisters_150__11
            ,inputRegisters_150__10,inputRegisters_150__9,inputRegisters_150__8,
            inputRegisters_150__7,inputRegisters_150__6,inputRegisters_150__5,
            inputRegisters_150__4,inputRegisters_150__3,inputRegisters_150__2,
            inputRegisters_150__1,inputRegisters_150__0})) ;
    Reg_16 loop1_150_x (.D ({inputRegisters_150__15,inputRegisters_150__14,
           inputRegisters_150__13,inputRegisters_150__12,inputRegisters_150__11,
           inputRegisters_150__10,inputRegisters_150__9,inputRegisters_150__8,
           inputRegisters_150__7,inputRegisters_150__6,inputRegisters_150__5,
           inputRegisters_150__4,inputRegisters_150__3,inputRegisters_150__2,
           inputRegisters_150__1,inputRegisters_150__0}), .en (
           enableRegister_150), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_150__15,registerOutputs_150__14,
           registerOutputs_150__13,registerOutputs_150__12,
           registerOutputs_150__11,registerOutputs_150__10,
           registerOutputs_150__9,registerOutputs_150__8,registerOutputs_150__7,
           registerOutputs_150__6,registerOutputs_150__5,registerOutputs_150__4,
           registerOutputs_150__3,registerOutputs_150__2,registerOutputs_150__1,
           registerOutputs_150__0})) ;
    Mux2_16 loop1_151_y (.A ({nx35927,nx36069,nx36211,nx36353,nx36495,nx36637,
            nx36779,nx36921,nx37063,nx37205,nx37347,nx37489,nx37631,nx37773,
            nx37915,nx38057}), .B ({nx33683,nx33821,nx33959,nx34099,nx34237,
            nx34375,nx34513,nx34653,nx34795,nx34937,nx35079,nx35221,nx35363,
            nx35505,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35647), .C ({inputRegisters_151__15,inputRegisters_151__14,
            inputRegisters_151__13,inputRegisters_151__12,inputRegisters_151__11
            ,inputRegisters_151__10,inputRegisters_151__9,inputRegisters_151__8,
            inputRegisters_151__7,inputRegisters_151__6,inputRegisters_151__5,
            inputRegisters_151__4,inputRegisters_151__3,inputRegisters_151__2,
            inputRegisters_151__1,inputRegisters_151__0})) ;
    Reg_16 loop1_151_x (.D ({inputRegisters_151__15,inputRegisters_151__14,
           inputRegisters_151__13,inputRegisters_151__12,inputRegisters_151__11,
           inputRegisters_151__10,inputRegisters_151__9,inputRegisters_151__8,
           inputRegisters_151__7,inputRegisters_151__6,inputRegisters_151__5,
           inputRegisters_151__4,inputRegisters_151__3,inputRegisters_151__2,
           inputRegisters_151__1,inputRegisters_151__0}), .en (
           enableRegister_151), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_151__15,registerOutputs_151__14,
           registerOutputs_151__13,registerOutputs_151__12,
           registerOutputs_151__11,registerOutputs_151__10,
           registerOutputs_151__9,registerOutputs_151__8,registerOutputs_151__7,
           registerOutputs_151__6,registerOutputs_151__5,registerOutputs_151__4,
           registerOutputs_151__3,registerOutputs_151__2,registerOutputs_151__1,
           registerOutputs_151__0})) ;
    Mux2_16 loop1_152_y (.A ({nx35927,nx36069,nx36211,nx36353,nx36495,nx36637,
            nx36779,nx36921,nx37063,nx37205,nx37347,nx37489,nx37631,nx37773,
            nx37915,nx38057}), .B ({nx33683,nx33821,nx33961,nx34099,nx34237,
            nx34375,nx34513,nx34653,nx34795,nx34937,nx35079,nx35221,nx35363,
            nx35505,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35647), .C ({inputRegisters_152__15,inputRegisters_152__14,
            inputRegisters_152__13,inputRegisters_152__12,inputRegisters_152__11
            ,inputRegisters_152__10,inputRegisters_152__9,inputRegisters_152__8,
            inputRegisters_152__7,inputRegisters_152__6,inputRegisters_152__5,
            inputRegisters_152__4,inputRegisters_152__3,inputRegisters_152__2,
            inputRegisters_152__1,inputRegisters_152__0})) ;
    Reg_16 loop1_152_x (.D ({inputRegisters_152__15,inputRegisters_152__14,
           inputRegisters_152__13,inputRegisters_152__12,inputRegisters_152__11,
           inputRegisters_152__10,inputRegisters_152__9,inputRegisters_152__8,
           inputRegisters_152__7,inputRegisters_152__6,inputRegisters_152__5,
           inputRegisters_152__4,inputRegisters_152__3,inputRegisters_152__2,
           inputRegisters_152__1,inputRegisters_152__0}), .en (
           enableRegister_152), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_152__15,registerOutputs_152__14,
           registerOutputs_152__13,registerOutputs_152__12,
           registerOutputs_152__11,registerOutputs_152__10,
           registerOutputs_152__9,registerOutputs_152__8,registerOutputs_152__7,
           registerOutputs_152__6,registerOutputs_152__5,registerOutputs_152__4,
           registerOutputs_152__3,registerOutputs_152__2,registerOutputs_152__1,
           registerOutputs_152__0})) ;
    Mux2_16 loop1_153_y (.A ({nx35927,nx36069,nx36211,nx36353,nx36495,nx36637,
            nx36779,nx36921,nx37063,nx37205,nx37347,nx37489,nx37631,nx37773,
            nx37915,nx38057}), .B ({nx33683,nx33823,nx33961,nx34099,nx34237,
            nx34375,nx34513,nx34653,nx34795,nx34937,nx35079,nx35221,nx35363,
            nx35505,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35647), .C ({inputRegisters_153__15,inputRegisters_153__14,
            inputRegisters_153__13,inputRegisters_153__12,inputRegisters_153__11
            ,inputRegisters_153__10,inputRegisters_153__9,inputRegisters_153__8,
            inputRegisters_153__7,inputRegisters_153__6,inputRegisters_153__5,
            inputRegisters_153__4,inputRegisters_153__3,inputRegisters_153__2,
            inputRegisters_153__1,inputRegisters_153__0})) ;
    Reg_16 loop1_153_x (.D ({inputRegisters_153__15,inputRegisters_153__14,
           inputRegisters_153__13,inputRegisters_153__12,inputRegisters_153__11,
           inputRegisters_153__10,inputRegisters_153__9,inputRegisters_153__8,
           inputRegisters_153__7,inputRegisters_153__6,inputRegisters_153__5,
           inputRegisters_153__4,inputRegisters_153__3,inputRegisters_153__2,
           inputRegisters_153__1,inputRegisters_153__0}), .en (
           enableRegister_153), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_153__15,registerOutputs_153__14,
           registerOutputs_153__13,registerOutputs_153__12,
           registerOutputs_153__11,registerOutputs_153__10,
           registerOutputs_153__9,registerOutputs_153__8,registerOutputs_153__7,
           registerOutputs_153__6,registerOutputs_153__5,registerOutputs_153__4,
           registerOutputs_153__3,registerOutputs_153__2,registerOutputs_153__1,
           registerOutputs_153__0})) ;
    Mux2_16 loop1_154_y (.A ({nx35929,nx36071,nx36213,nx36355,nx36497,nx36639,
            nx36781,nx36923,nx37065,nx37207,nx37349,nx37491,nx37633,nx37775,
            nx37917,nx38059}), .B ({nx33685,nx33823,nx33961,nx34099,nx34237,
            nx34375,nx34513,nx34655,nx34797,nx34939,nx35081,nx35223,nx35365,
            nx35507,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35649), .C ({inputRegisters_154__15,inputRegisters_154__14,
            inputRegisters_154__13,inputRegisters_154__12,inputRegisters_154__11
            ,inputRegisters_154__10,inputRegisters_154__9,inputRegisters_154__8,
            inputRegisters_154__7,inputRegisters_154__6,inputRegisters_154__5,
            inputRegisters_154__4,inputRegisters_154__3,inputRegisters_154__2,
            inputRegisters_154__1,inputRegisters_154__0})) ;
    Reg_16 loop1_154_x (.D ({inputRegisters_154__15,inputRegisters_154__14,
           inputRegisters_154__13,inputRegisters_154__12,inputRegisters_154__11,
           inputRegisters_154__10,inputRegisters_154__9,inputRegisters_154__8,
           inputRegisters_154__7,inputRegisters_154__6,inputRegisters_154__5,
           inputRegisters_154__4,inputRegisters_154__3,inputRegisters_154__2,
           inputRegisters_154__1,inputRegisters_154__0}), .en (
           enableRegister_154), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_154__15,registerOutputs_154__14,
           registerOutputs_154__13,registerOutputs_154__12,
           registerOutputs_154__11,registerOutputs_154__10,
           registerOutputs_154__9,registerOutputs_154__8,registerOutputs_154__7,
           registerOutputs_154__6,registerOutputs_154__5,registerOutputs_154__4,
           registerOutputs_154__3,registerOutputs_154__2,registerOutputs_154__1,
           registerOutputs_154__0})) ;
    Mux2_16 loop1_155_y (.A ({nx35929,nx36071,nx36213,nx36355,nx36497,nx36639,
            nx36781,nx36923,nx37065,nx37207,nx37349,nx37491,nx37633,nx37775,
            nx37917,nx38059}), .B ({nx33685,nx33823,nx33961,nx34099,nx34237,
            nx34375,nx34515,nx34655,nx34797,nx34939,nx35081,nx35223,nx35365,
            nx35507,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35649), .C ({inputRegisters_155__15,inputRegisters_155__14,
            inputRegisters_155__13,inputRegisters_155__12,inputRegisters_155__11
            ,inputRegisters_155__10,inputRegisters_155__9,inputRegisters_155__8,
            inputRegisters_155__7,inputRegisters_155__6,inputRegisters_155__5,
            inputRegisters_155__4,inputRegisters_155__3,inputRegisters_155__2,
            inputRegisters_155__1,inputRegisters_155__0})) ;
    Reg_16 loop1_155_x (.D ({inputRegisters_155__15,inputRegisters_155__14,
           inputRegisters_155__13,inputRegisters_155__12,inputRegisters_155__11,
           inputRegisters_155__10,inputRegisters_155__9,inputRegisters_155__8,
           inputRegisters_155__7,inputRegisters_155__6,inputRegisters_155__5,
           inputRegisters_155__4,inputRegisters_155__3,inputRegisters_155__2,
           inputRegisters_155__1,inputRegisters_155__0}), .en (
           enableRegister_155), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_155__15,registerOutputs_155__14,
           registerOutputs_155__13,registerOutputs_155__12,
           registerOutputs_155__11,registerOutputs_155__10,
           registerOutputs_155__9,registerOutputs_155__8,registerOutputs_155__7,
           registerOutputs_155__6,registerOutputs_155__5,registerOutputs_155__4,
           registerOutputs_155__3,registerOutputs_155__2,registerOutputs_155__1,
           registerOutputs_155__0})) ;
    Mux2_16 loop1_156_y (.A ({nx35929,nx36071,nx36213,nx36355,nx36497,nx36639,
            nx36781,nx36923,nx37065,nx37207,nx37349,nx37491,nx37633,nx37775,
            nx37917,nx38059}), .B ({nx33685,nx33823,nx33961,nx34099,nx34237,
            nx34377,nx34515,nx34655,nx34797,nx34939,nx35081,nx35223,nx35365,
            nx35507,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35649), .C ({inputRegisters_156__15,inputRegisters_156__14,
            inputRegisters_156__13,inputRegisters_156__12,inputRegisters_156__11
            ,inputRegisters_156__10,inputRegisters_156__9,inputRegisters_156__8,
            inputRegisters_156__7,inputRegisters_156__6,inputRegisters_156__5,
            inputRegisters_156__4,inputRegisters_156__3,inputRegisters_156__2,
            inputRegisters_156__1,inputRegisters_156__0})) ;
    Reg_16 loop1_156_x (.D ({inputRegisters_156__15,inputRegisters_156__14,
           inputRegisters_156__13,inputRegisters_156__12,inputRegisters_156__11,
           inputRegisters_156__10,inputRegisters_156__9,inputRegisters_156__8,
           inputRegisters_156__7,inputRegisters_156__6,inputRegisters_156__5,
           inputRegisters_156__4,inputRegisters_156__3,inputRegisters_156__2,
           inputRegisters_156__1,inputRegisters_156__0}), .en (
           enableRegister_156), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_156__15,registerOutputs_156__14,
           registerOutputs_156__13,registerOutputs_156__12,
           registerOutputs_156__11,registerOutputs_156__10,
           registerOutputs_156__9,registerOutputs_156__8,registerOutputs_156__7,
           registerOutputs_156__6,registerOutputs_156__5,registerOutputs_156__4,
           registerOutputs_156__3,registerOutputs_156__2,registerOutputs_156__1,
           registerOutputs_156__0})) ;
    Mux2_16 loop1_157_y (.A ({nx35929,nx36071,nx36213,nx36355,nx36497,nx36639,
            nx36781,nx36923,nx37065,nx37207,nx37349,nx37491,nx37633,nx37775,
            nx37917,nx38059}), .B ({nx33685,nx33823,nx33961,nx34099,nx34239,
            nx34377,nx34515,nx34655,nx34797,nx34939,nx35081,nx35223,nx35365,
            nx35507,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35649), .C ({inputRegisters_157__15,inputRegisters_157__14,
            inputRegisters_157__13,inputRegisters_157__12,inputRegisters_157__11
            ,inputRegisters_157__10,inputRegisters_157__9,inputRegisters_157__8,
            inputRegisters_157__7,inputRegisters_157__6,inputRegisters_157__5,
            inputRegisters_157__4,inputRegisters_157__3,inputRegisters_157__2,
            inputRegisters_157__1,inputRegisters_157__0})) ;
    Reg_16 loop1_157_x (.D ({inputRegisters_157__15,inputRegisters_157__14,
           inputRegisters_157__13,inputRegisters_157__12,inputRegisters_157__11,
           inputRegisters_157__10,inputRegisters_157__9,inputRegisters_157__8,
           inputRegisters_157__7,inputRegisters_157__6,inputRegisters_157__5,
           inputRegisters_157__4,inputRegisters_157__3,inputRegisters_157__2,
           inputRegisters_157__1,inputRegisters_157__0}), .en (
           enableRegister_157), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_157__15,registerOutputs_157__14,
           registerOutputs_157__13,registerOutputs_157__12,
           registerOutputs_157__11,registerOutputs_157__10,
           registerOutputs_157__9,registerOutputs_157__8,registerOutputs_157__7,
           registerOutputs_157__6,registerOutputs_157__5,registerOutputs_157__4,
           registerOutputs_157__3,registerOutputs_157__2,registerOutputs_157__1,
           registerOutputs_157__0})) ;
    Mux2_16 loop1_158_y (.A ({nx35929,nx36071,nx36213,nx36355,nx36497,nx36639,
            nx36781,nx36923,nx37065,nx37207,nx37349,nx37491,nx37633,nx37775,
            nx37917,nx38059}), .B ({nx33685,nx33823,nx33961,nx34101,nx34239,
            nx34377,nx34515,nx34655,nx34797,nx34939,nx35081,nx35223,nx35365,
            nx35507,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35649), .C ({inputRegisters_158__15,inputRegisters_158__14,
            inputRegisters_158__13,inputRegisters_158__12,inputRegisters_158__11
            ,inputRegisters_158__10,inputRegisters_158__9,inputRegisters_158__8,
            inputRegisters_158__7,inputRegisters_158__6,inputRegisters_158__5,
            inputRegisters_158__4,inputRegisters_158__3,inputRegisters_158__2,
            inputRegisters_158__1,inputRegisters_158__0})) ;
    Reg_16 loop1_158_x (.D ({inputRegisters_158__15,inputRegisters_158__14,
           inputRegisters_158__13,inputRegisters_158__12,inputRegisters_158__11,
           inputRegisters_158__10,inputRegisters_158__9,inputRegisters_158__8,
           inputRegisters_158__7,inputRegisters_158__6,inputRegisters_158__5,
           inputRegisters_158__4,inputRegisters_158__3,inputRegisters_158__2,
           inputRegisters_158__1,inputRegisters_158__0}), .en (
           enableRegister_158), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_158__15,registerOutputs_158__14,
           registerOutputs_158__13,registerOutputs_158__12,
           registerOutputs_158__11,registerOutputs_158__10,
           registerOutputs_158__9,registerOutputs_158__8,registerOutputs_158__7,
           registerOutputs_158__6,registerOutputs_158__5,registerOutputs_158__4,
           registerOutputs_158__3,registerOutputs_158__2,registerOutputs_158__1,
           registerOutputs_158__0})) ;
    Mux2_16 loop1_159_y (.A ({nx35929,nx36071,nx36213,nx36355,nx36497,nx36639,
            nx36781,nx36923,nx37065,nx37207,nx37349,nx37491,nx37633,nx37775,
            nx37917,nx38059}), .B ({nx33685,nx33823,nx33963,nx34101,nx34239,
            nx34377,nx34515,nx34655,nx34797,nx34939,nx35081,nx35223,nx35365,
            nx35507,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35649), .C ({inputRegisters_159__15,inputRegisters_159__14,
            inputRegisters_159__13,inputRegisters_159__12,inputRegisters_159__11
            ,inputRegisters_159__10,inputRegisters_159__9,inputRegisters_159__8,
            inputRegisters_159__7,inputRegisters_159__6,inputRegisters_159__5,
            inputRegisters_159__4,inputRegisters_159__3,inputRegisters_159__2,
            inputRegisters_159__1,inputRegisters_159__0})) ;
    Reg_16 loop1_159_x (.D ({inputRegisters_159__15,inputRegisters_159__14,
           inputRegisters_159__13,inputRegisters_159__12,inputRegisters_159__11,
           inputRegisters_159__10,inputRegisters_159__9,inputRegisters_159__8,
           inputRegisters_159__7,inputRegisters_159__6,inputRegisters_159__5,
           inputRegisters_159__4,inputRegisters_159__3,inputRegisters_159__2,
           inputRegisters_159__1,inputRegisters_159__0}), .en (
           enableRegister_159), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_159__15,registerOutputs_159__14,
           registerOutputs_159__13,registerOutputs_159__12,
           registerOutputs_159__11,registerOutputs_159__10,
           registerOutputs_159__9,registerOutputs_159__8,registerOutputs_159__7,
           registerOutputs_159__6,registerOutputs_159__5,registerOutputs_159__4,
           registerOutputs_159__3,registerOutputs_159__2,registerOutputs_159__1,
           registerOutputs_159__0})) ;
    Mux2_16 loop1_160_y (.A ({nx35929,nx36071,nx36213,nx36355,nx36497,nx36639,
            nx36781,nx36923,nx37065,nx37207,nx37349,nx37491,nx37633,nx37775,
            nx37917,nx38059}), .B ({nx33685,nx33825,nx33963,nx34101,nx34239,
            nx34377,nx34515,nx34655,nx34797,nx34939,nx35081,nx35223,nx35365,
            nx35507,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35649), .C ({inputRegisters_160__15,inputRegisters_160__14,
            inputRegisters_160__13,inputRegisters_160__12,inputRegisters_160__11
            ,inputRegisters_160__10,inputRegisters_160__9,inputRegisters_160__8,
            inputRegisters_160__7,inputRegisters_160__6,inputRegisters_160__5,
            inputRegisters_160__4,inputRegisters_160__3,inputRegisters_160__2,
            inputRegisters_160__1,inputRegisters_160__0})) ;
    Reg_16 loop1_160_x (.D ({inputRegisters_160__15,inputRegisters_160__14,
           inputRegisters_160__13,inputRegisters_160__12,inputRegisters_160__11,
           inputRegisters_160__10,inputRegisters_160__9,inputRegisters_160__8,
           inputRegisters_160__7,inputRegisters_160__6,inputRegisters_160__5,
           inputRegisters_160__4,inputRegisters_160__3,inputRegisters_160__2,
           inputRegisters_160__1,inputRegisters_160__0}), .en (
           enableRegister_160), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_160__15,registerOutputs_160__14,
           registerOutputs_160__13,registerOutputs_160__12,
           registerOutputs_160__11,registerOutputs_160__10,
           registerOutputs_160__9,registerOutputs_160__8,registerOutputs_160__7,
           registerOutputs_160__6,registerOutputs_160__5,registerOutputs_160__4,
           registerOutputs_160__3,registerOutputs_160__2,registerOutputs_160__1,
           registerOutputs_160__0})) ;
    Mux2_16 loop1_161_y (.A ({nx35931,nx36073,nx36215,nx36357,nx36499,nx36641,
            nx36783,nx36925,nx37067,nx37209,nx37351,nx37493,nx37635,nx37777,
            nx37919,nx38061}), .B ({nx33687,nx33825,nx33963,nx34101,nx34239,
            nx34377,nx34515,nx34657,nx34799,nx34941,nx35083,nx35225,nx35367,
            nx35509,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35651), .C ({inputRegisters_161__15,inputRegisters_161__14,
            inputRegisters_161__13,inputRegisters_161__12,inputRegisters_161__11
            ,inputRegisters_161__10,inputRegisters_161__9,inputRegisters_161__8,
            inputRegisters_161__7,inputRegisters_161__6,inputRegisters_161__5,
            inputRegisters_161__4,inputRegisters_161__3,inputRegisters_161__2,
            inputRegisters_161__1,inputRegisters_161__0})) ;
    Reg_16 loop1_161_x (.D ({inputRegisters_161__15,inputRegisters_161__14,
           inputRegisters_161__13,inputRegisters_161__12,inputRegisters_161__11,
           inputRegisters_161__10,inputRegisters_161__9,inputRegisters_161__8,
           inputRegisters_161__7,inputRegisters_161__6,inputRegisters_161__5,
           inputRegisters_161__4,inputRegisters_161__3,inputRegisters_161__2,
           inputRegisters_161__1,inputRegisters_161__0}), .en (
           enableRegister_161), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_161__15,registerOutputs_161__14,
           registerOutputs_161__13,registerOutputs_161__12,
           registerOutputs_161__11,registerOutputs_161__10,
           registerOutputs_161__9,registerOutputs_161__8,registerOutputs_161__7,
           registerOutputs_161__6,registerOutputs_161__5,registerOutputs_161__4,
           registerOutputs_161__3,registerOutputs_161__2,registerOutputs_161__1,
           registerOutputs_161__0})) ;
    Mux2_16 loop1_162_y (.A ({nx35931,nx36073,nx36215,nx36357,nx36499,nx36641,
            nx36783,nx36925,nx37067,nx37209,nx37351,nx37493,nx37635,nx37777,
            nx37919,nx38061}), .B ({nx33687,nx33825,nx33963,nx34101,nx34239,
            nx34377,nx34517,nx34657,nx34799,nx34941,nx35083,nx35225,nx35367,
            nx35509,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35651), .C ({inputRegisters_162__15,inputRegisters_162__14,
            inputRegisters_162__13,inputRegisters_162__12,inputRegisters_162__11
            ,inputRegisters_162__10,inputRegisters_162__9,inputRegisters_162__8,
            inputRegisters_162__7,inputRegisters_162__6,inputRegisters_162__5,
            inputRegisters_162__4,inputRegisters_162__3,inputRegisters_162__2,
            inputRegisters_162__1,inputRegisters_162__0})) ;
    Reg_16 loop1_162_x (.D ({inputRegisters_162__15,inputRegisters_162__14,
           inputRegisters_162__13,inputRegisters_162__12,inputRegisters_162__11,
           inputRegisters_162__10,inputRegisters_162__9,inputRegisters_162__8,
           inputRegisters_162__7,inputRegisters_162__6,inputRegisters_162__5,
           inputRegisters_162__4,inputRegisters_162__3,inputRegisters_162__2,
           inputRegisters_162__1,inputRegisters_162__0}), .en (
           enableRegister_162), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_162__15,registerOutputs_162__14,
           registerOutputs_162__13,registerOutputs_162__12,
           registerOutputs_162__11,registerOutputs_162__10,
           registerOutputs_162__9,registerOutputs_162__8,registerOutputs_162__7,
           registerOutputs_162__6,registerOutputs_162__5,registerOutputs_162__4,
           registerOutputs_162__3,registerOutputs_162__2,registerOutputs_162__1,
           registerOutputs_162__0})) ;
    Mux2_16 loop1_163_y (.A ({nx35931,nx36073,nx36215,nx36357,nx36499,nx36641,
            nx36783,nx36925,nx37067,nx37209,nx37351,nx37493,nx37635,nx37777,
            nx37919,nx38061}), .B ({nx33687,nx33825,nx33963,nx34101,nx34239,
            nx34379,nx34517,nx34657,nx34799,nx34941,nx35083,nx35225,nx35367,
            nx35509,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35651), .C ({inputRegisters_163__15,inputRegisters_163__14,
            inputRegisters_163__13,inputRegisters_163__12,inputRegisters_163__11
            ,inputRegisters_163__10,inputRegisters_163__9,inputRegisters_163__8,
            inputRegisters_163__7,inputRegisters_163__6,inputRegisters_163__5,
            inputRegisters_163__4,inputRegisters_163__3,inputRegisters_163__2,
            inputRegisters_163__1,inputRegisters_163__0})) ;
    Reg_16 loop1_163_x (.D ({inputRegisters_163__15,inputRegisters_163__14,
           inputRegisters_163__13,inputRegisters_163__12,inputRegisters_163__11,
           inputRegisters_163__10,inputRegisters_163__9,inputRegisters_163__8,
           inputRegisters_163__7,inputRegisters_163__6,inputRegisters_163__5,
           inputRegisters_163__4,inputRegisters_163__3,inputRegisters_163__2,
           inputRegisters_163__1,inputRegisters_163__0}), .en (
           enableRegister_163), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_163__15,registerOutputs_163__14,
           registerOutputs_163__13,registerOutputs_163__12,
           registerOutputs_163__11,registerOutputs_163__10,
           registerOutputs_163__9,registerOutputs_163__8,registerOutputs_163__7,
           registerOutputs_163__6,registerOutputs_163__5,registerOutputs_163__4,
           registerOutputs_163__3,registerOutputs_163__2,registerOutputs_163__1,
           registerOutputs_163__0})) ;
    Mux2_16 loop1_164_y (.A ({nx35931,nx36073,nx36215,nx36357,nx36499,nx36641,
            nx36783,nx36925,nx37067,nx37209,nx37351,nx37493,nx37635,nx37777,
            nx37919,nx38061}), .B ({nx33687,nx33825,nx33963,nx34101,nx34241,
            nx34379,nx34517,nx34657,nx34799,nx34941,nx35083,nx35225,nx35367,
            nx35509,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35651), .C ({inputRegisters_164__15,inputRegisters_164__14,
            inputRegisters_164__13,inputRegisters_164__12,inputRegisters_164__11
            ,inputRegisters_164__10,inputRegisters_164__9,inputRegisters_164__8,
            inputRegisters_164__7,inputRegisters_164__6,inputRegisters_164__5,
            inputRegisters_164__4,inputRegisters_164__3,inputRegisters_164__2,
            inputRegisters_164__1,inputRegisters_164__0})) ;
    Reg_16 loop1_164_x (.D ({inputRegisters_164__15,inputRegisters_164__14,
           inputRegisters_164__13,inputRegisters_164__12,inputRegisters_164__11,
           inputRegisters_164__10,inputRegisters_164__9,inputRegisters_164__8,
           inputRegisters_164__7,inputRegisters_164__6,inputRegisters_164__5,
           inputRegisters_164__4,inputRegisters_164__3,inputRegisters_164__2,
           inputRegisters_164__1,inputRegisters_164__0}), .en (
           enableRegister_164), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_164__15,registerOutputs_164__14,
           registerOutputs_164__13,registerOutputs_164__12,
           registerOutputs_164__11,registerOutputs_164__10,
           registerOutputs_164__9,registerOutputs_164__8,registerOutputs_164__7,
           registerOutputs_164__6,registerOutputs_164__5,registerOutputs_164__4,
           registerOutputs_164__3,registerOutputs_164__2,registerOutputs_164__1,
           registerOutputs_164__0})) ;
    Mux2_16 loop1_165_y (.A ({nx35931,nx36073,nx36215,nx36357,nx36499,nx36641,
            nx36783,nx36925,nx37067,nx37209,nx37351,nx37493,nx37635,nx37777,
            nx37919,nx38061}), .B ({nx33687,nx33825,nx33963,nx34103,nx34241,
            nx34379,nx34517,nx34657,nx34799,nx34941,nx35083,nx35225,nx35367,
            nx35509,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35651), .C ({inputRegisters_165__15,inputRegisters_165__14,
            inputRegisters_165__13,inputRegisters_165__12,inputRegisters_165__11
            ,inputRegisters_165__10,inputRegisters_165__9,inputRegisters_165__8,
            inputRegisters_165__7,inputRegisters_165__6,inputRegisters_165__5,
            inputRegisters_165__4,inputRegisters_165__3,inputRegisters_165__2,
            inputRegisters_165__1,inputRegisters_165__0})) ;
    Reg_16 loop1_165_x (.D ({inputRegisters_165__15,inputRegisters_165__14,
           inputRegisters_165__13,inputRegisters_165__12,inputRegisters_165__11,
           inputRegisters_165__10,inputRegisters_165__9,inputRegisters_165__8,
           inputRegisters_165__7,inputRegisters_165__6,inputRegisters_165__5,
           inputRegisters_165__4,inputRegisters_165__3,inputRegisters_165__2,
           inputRegisters_165__1,inputRegisters_165__0}), .en (
           enableRegister_165), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_165__15,registerOutputs_165__14,
           registerOutputs_165__13,registerOutputs_165__12,
           registerOutputs_165__11,registerOutputs_165__10,
           registerOutputs_165__9,registerOutputs_165__8,registerOutputs_165__7,
           registerOutputs_165__6,registerOutputs_165__5,registerOutputs_165__4,
           registerOutputs_165__3,registerOutputs_165__2,registerOutputs_165__1,
           registerOutputs_165__0})) ;
    Mux2_16 loop1_166_y (.A ({nx35931,nx36073,nx36215,nx36357,nx36499,nx36641,
            nx36783,nx36925,nx37067,nx37209,nx37351,nx37493,nx37635,nx37777,
            nx37919,nx38061}), .B ({nx33687,nx33825,nx33965,nx34103,nx34241,
            nx34379,nx34517,nx34657,nx34799,nx34941,nx35083,nx35225,nx35367,
            nx35509,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35651), .C ({inputRegisters_166__15,inputRegisters_166__14,
            inputRegisters_166__13,inputRegisters_166__12,inputRegisters_166__11
            ,inputRegisters_166__10,inputRegisters_166__9,inputRegisters_166__8,
            inputRegisters_166__7,inputRegisters_166__6,inputRegisters_166__5,
            inputRegisters_166__4,inputRegisters_166__3,inputRegisters_166__2,
            inputRegisters_166__1,inputRegisters_166__0})) ;
    Reg_16 loop1_166_x (.D ({inputRegisters_166__15,inputRegisters_166__14,
           inputRegisters_166__13,inputRegisters_166__12,inputRegisters_166__11,
           inputRegisters_166__10,inputRegisters_166__9,inputRegisters_166__8,
           inputRegisters_166__7,inputRegisters_166__6,inputRegisters_166__5,
           inputRegisters_166__4,inputRegisters_166__3,inputRegisters_166__2,
           inputRegisters_166__1,inputRegisters_166__0}), .en (
           enableRegister_166), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_166__15,registerOutputs_166__14,
           registerOutputs_166__13,registerOutputs_166__12,
           registerOutputs_166__11,registerOutputs_166__10,
           registerOutputs_166__9,registerOutputs_166__8,registerOutputs_166__7,
           registerOutputs_166__6,registerOutputs_166__5,registerOutputs_166__4,
           registerOutputs_166__3,registerOutputs_166__2,registerOutputs_166__1,
           registerOutputs_166__0})) ;
    Mux2_16 loop1_167_y (.A ({nx35931,nx36073,nx36215,nx36357,nx36499,nx36641,
            nx36783,nx36925,nx37067,nx37209,nx37351,nx37493,nx37635,nx37777,
            nx37919,nx38061}), .B ({nx33687,nx33827,nx33965,nx34103,nx34241,
            nx34379,nx34517,nx34657,nx34799,nx34941,nx35083,nx35225,nx35367,
            nx35509,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35651), .C ({inputRegisters_167__15,inputRegisters_167__14,
            inputRegisters_167__13,inputRegisters_167__12,inputRegisters_167__11
            ,inputRegisters_167__10,inputRegisters_167__9,inputRegisters_167__8,
            inputRegisters_167__7,inputRegisters_167__6,inputRegisters_167__5,
            inputRegisters_167__4,inputRegisters_167__3,inputRegisters_167__2,
            inputRegisters_167__1,inputRegisters_167__0})) ;
    Reg_16 loop1_167_x (.D ({inputRegisters_167__15,inputRegisters_167__14,
           inputRegisters_167__13,inputRegisters_167__12,inputRegisters_167__11,
           inputRegisters_167__10,inputRegisters_167__9,inputRegisters_167__8,
           inputRegisters_167__7,inputRegisters_167__6,inputRegisters_167__5,
           inputRegisters_167__4,inputRegisters_167__3,inputRegisters_167__2,
           inputRegisters_167__1,inputRegisters_167__0}), .en (
           enableRegister_167), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_167__15,registerOutputs_167__14,
           registerOutputs_167__13,registerOutputs_167__12,
           registerOutputs_167__11,registerOutputs_167__10,
           registerOutputs_167__9,registerOutputs_167__8,registerOutputs_167__7,
           registerOutputs_167__6,registerOutputs_167__5,registerOutputs_167__4,
           registerOutputs_167__3,registerOutputs_167__2,registerOutputs_167__1,
           registerOutputs_167__0})) ;
    Mux2_16 loop1_168_y (.A ({nx35933,nx36075,nx36217,nx36359,nx36501,nx36643,
            nx36785,nx36927,nx37069,nx37211,nx37353,nx37495,nx37637,nx37779,
            nx37921,nx38063}), .B ({nx33689,nx33827,nx33965,nx34103,nx34241,
            nx34379,nx34517,nx34659,nx34801,nx34943,nx35085,nx35227,nx35369,
            nx35511,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35653), .C ({inputRegisters_168__15,inputRegisters_168__14,
            inputRegisters_168__13,inputRegisters_168__12,inputRegisters_168__11
            ,inputRegisters_168__10,inputRegisters_168__9,inputRegisters_168__8,
            inputRegisters_168__7,inputRegisters_168__6,inputRegisters_168__5,
            inputRegisters_168__4,inputRegisters_168__3,inputRegisters_168__2,
            inputRegisters_168__1,inputRegisters_168__0})) ;
    Reg_16 loop1_168_x (.D ({inputRegisters_168__15,inputRegisters_168__14,
           inputRegisters_168__13,inputRegisters_168__12,inputRegisters_168__11,
           inputRegisters_168__10,inputRegisters_168__9,inputRegisters_168__8,
           inputRegisters_168__7,inputRegisters_168__6,inputRegisters_168__5,
           inputRegisters_168__4,inputRegisters_168__3,inputRegisters_168__2,
           inputRegisters_168__1,inputRegisters_168__0}), .en (
           enableRegister_168), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_168__15,registerOutputs_168__14,
           registerOutputs_168__13,registerOutputs_168__12,
           registerOutputs_168__11,registerOutputs_168__10,
           registerOutputs_168__9,registerOutputs_168__8,registerOutputs_168__7,
           registerOutputs_168__6,registerOutputs_168__5,registerOutputs_168__4,
           registerOutputs_168__3,registerOutputs_168__2,registerOutputs_168__1,
           registerOutputs_168__0})) ;
    Mux2_16 loop1_169_y (.A ({nx35933,nx36075,nx36217,nx36359,nx36501,nx36643,
            nx36785,nx36927,nx37069,nx37211,nx37353,nx37495,nx37637,nx37779,
            nx37921,nx38063}), .B ({nx33689,nx33827,nx33965,nx34103,nx34241,
            nx34379,nx34519,nx34659,nx34801,nx34943,nx35085,nx35227,nx35369,
            nx35511,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35653), .C ({inputRegisters_169__15,inputRegisters_169__14,
            inputRegisters_169__13,inputRegisters_169__12,inputRegisters_169__11
            ,inputRegisters_169__10,inputRegisters_169__9,inputRegisters_169__8,
            inputRegisters_169__7,inputRegisters_169__6,inputRegisters_169__5,
            inputRegisters_169__4,inputRegisters_169__3,inputRegisters_169__2,
            inputRegisters_169__1,inputRegisters_169__0})) ;
    Reg_16 loop1_169_x (.D ({inputRegisters_169__15,inputRegisters_169__14,
           inputRegisters_169__13,inputRegisters_169__12,inputRegisters_169__11,
           inputRegisters_169__10,inputRegisters_169__9,inputRegisters_169__8,
           inputRegisters_169__7,inputRegisters_169__6,inputRegisters_169__5,
           inputRegisters_169__4,inputRegisters_169__3,inputRegisters_169__2,
           inputRegisters_169__1,inputRegisters_169__0}), .en (
           enableRegister_169), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_169__15,registerOutputs_169__14,
           registerOutputs_169__13,registerOutputs_169__12,
           registerOutputs_169__11,registerOutputs_169__10,
           registerOutputs_169__9,registerOutputs_169__8,registerOutputs_169__7,
           registerOutputs_169__6,registerOutputs_169__5,registerOutputs_169__4,
           registerOutputs_169__3,registerOutputs_169__2,registerOutputs_169__1,
           registerOutputs_169__0})) ;
    Mux2_16 loop1_170_y (.A ({nx35933,nx36075,nx36217,nx36359,nx36501,nx36643,
            nx36785,nx36927,nx37069,nx37211,nx37353,nx37495,nx37637,nx37779,
            nx37921,nx38063}), .B ({nx33689,nx33827,nx33965,nx34103,nx34241,
            nx34381,nx34519,nx34659,nx34801,nx34943,nx35085,nx35227,nx35369,
            nx35511,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35653), .C ({inputRegisters_170__15,inputRegisters_170__14,
            inputRegisters_170__13,inputRegisters_170__12,inputRegisters_170__11
            ,inputRegisters_170__10,inputRegisters_170__9,inputRegisters_170__8,
            inputRegisters_170__7,inputRegisters_170__6,inputRegisters_170__5,
            inputRegisters_170__4,inputRegisters_170__3,inputRegisters_170__2,
            inputRegisters_170__1,inputRegisters_170__0})) ;
    Reg_16 loop1_170_x (.D ({inputRegisters_170__15,inputRegisters_170__14,
           inputRegisters_170__13,inputRegisters_170__12,inputRegisters_170__11,
           inputRegisters_170__10,inputRegisters_170__9,inputRegisters_170__8,
           inputRegisters_170__7,inputRegisters_170__6,inputRegisters_170__5,
           inputRegisters_170__4,inputRegisters_170__3,inputRegisters_170__2,
           inputRegisters_170__1,inputRegisters_170__0}), .en (
           enableRegister_170), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_170__15,registerOutputs_170__14,
           registerOutputs_170__13,registerOutputs_170__12,
           registerOutputs_170__11,registerOutputs_170__10,
           registerOutputs_170__9,registerOutputs_170__8,registerOutputs_170__7,
           registerOutputs_170__6,registerOutputs_170__5,registerOutputs_170__4,
           registerOutputs_170__3,registerOutputs_170__2,registerOutputs_170__1,
           registerOutputs_170__0})) ;
    Mux2_16 loop1_171_y (.A ({nx35933,nx36075,nx36217,nx36359,nx36501,nx36643,
            nx36785,nx36927,nx37069,nx37211,nx37353,nx37495,nx37637,nx37779,
            nx37921,nx38063}), .B ({nx33689,nx33827,nx33965,nx34103,nx34243,
            nx34381,nx34519,nx34659,nx34801,nx34943,nx35085,nx35227,nx35369,
            nx35511,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35653), .C ({inputRegisters_171__15,inputRegisters_171__14,
            inputRegisters_171__13,inputRegisters_171__12,inputRegisters_171__11
            ,inputRegisters_171__10,inputRegisters_171__9,inputRegisters_171__8,
            inputRegisters_171__7,inputRegisters_171__6,inputRegisters_171__5,
            inputRegisters_171__4,inputRegisters_171__3,inputRegisters_171__2,
            inputRegisters_171__1,inputRegisters_171__0})) ;
    Reg_16 loop1_171_x (.D ({inputRegisters_171__15,inputRegisters_171__14,
           inputRegisters_171__13,inputRegisters_171__12,inputRegisters_171__11,
           inputRegisters_171__10,inputRegisters_171__9,inputRegisters_171__8,
           inputRegisters_171__7,inputRegisters_171__6,inputRegisters_171__5,
           inputRegisters_171__4,inputRegisters_171__3,inputRegisters_171__2,
           inputRegisters_171__1,inputRegisters_171__0}), .en (
           enableRegister_171), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_171__15,registerOutputs_171__14,
           registerOutputs_171__13,registerOutputs_171__12,
           registerOutputs_171__11,registerOutputs_171__10,
           registerOutputs_171__9,registerOutputs_171__8,registerOutputs_171__7,
           registerOutputs_171__6,registerOutputs_171__5,registerOutputs_171__4,
           registerOutputs_171__3,registerOutputs_171__2,registerOutputs_171__1,
           registerOutputs_171__0})) ;
    Mux2_16 loop1_172_y (.A ({nx35933,nx36075,nx36217,nx36359,nx36501,nx36643,
            nx36785,nx36927,nx37069,nx37211,nx37353,nx37495,nx37637,nx37779,
            nx37921,nx38063}), .B ({nx33689,nx33827,nx33965,nx34105,nx34243,
            nx34381,nx34519,nx34659,nx34801,nx34943,nx35085,nx35227,nx35369,
            nx35511,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35653), .C ({inputRegisters_172__15,inputRegisters_172__14,
            inputRegisters_172__13,inputRegisters_172__12,inputRegisters_172__11
            ,inputRegisters_172__10,inputRegisters_172__9,inputRegisters_172__8,
            inputRegisters_172__7,inputRegisters_172__6,inputRegisters_172__5,
            inputRegisters_172__4,inputRegisters_172__3,inputRegisters_172__2,
            inputRegisters_172__1,inputRegisters_172__0})) ;
    Reg_16 loop1_172_x (.D ({inputRegisters_172__15,inputRegisters_172__14,
           inputRegisters_172__13,inputRegisters_172__12,inputRegisters_172__11,
           inputRegisters_172__10,inputRegisters_172__9,inputRegisters_172__8,
           inputRegisters_172__7,inputRegisters_172__6,inputRegisters_172__5,
           inputRegisters_172__4,inputRegisters_172__3,inputRegisters_172__2,
           inputRegisters_172__1,inputRegisters_172__0}), .en (
           enableRegister_172), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_172__15,registerOutputs_172__14,
           registerOutputs_172__13,registerOutputs_172__12,
           registerOutputs_172__11,registerOutputs_172__10,
           registerOutputs_172__9,registerOutputs_172__8,registerOutputs_172__7,
           registerOutputs_172__6,registerOutputs_172__5,registerOutputs_172__4,
           registerOutputs_172__3,registerOutputs_172__2,registerOutputs_172__1,
           registerOutputs_172__0})) ;
    Mux2_16 loop1_173_y (.A ({nx35933,nx36075,nx36217,nx36359,nx36501,nx36643,
            nx36785,nx36927,nx37069,nx37211,nx37353,nx37495,nx37637,nx37779,
            nx37921,nx38063}), .B ({nx33689,nx33827,nx33967,nx34105,nx34243,
            nx34381,nx34519,nx34659,nx34801,nx34943,nx35085,nx35227,nx35369,
            nx35511,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35653), .C ({inputRegisters_173__15,inputRegisters_173__14,
            inputRegisters_173__13,inputRegisters_173__12,inputRegisters_173__11
            ,inputRegisters_173__10,inputRegisters_173__9,inputRegisters_173__8,
            inputRegisters_173__7,inputRegisters_173__6,inputRegisters_173__5,
            inputRegisters_173__4,inputRegisters_173__3,inputRegisters_173__2,
            inputRegisters_173__1,inputRegisters_173__0})) ;
    Reg_16 loop1_173_x (.D ({inputRegisters_173__15,inputRegisters_173__14,
           inputRegisters_173__13,inputRegisters_173__12,inputRegisters_173__11,
           inputRegisters_173__10,inputRegisters_173__9,inputRegisters_173__8,
           inputRegisters_173__7,inputRegisters_173__6,inputRegisters_173__5,
           inputRegisters_173__4,inputRegisters_173__3,inputRegisters_173__2,
           inputRegisters_173__1,inputRegisters_173__0}), .en (
           enableRegister_173), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_173__15,registerOutputs_173__14,
           registerOutputs_173__13,registerOutputs_173__12,
           registerOutputs_173__11,registerOutputs_173__10,
           registerOutputs_173__9,registerOutputs_173__8,registerOutputs_173__7,
           registerOutputs_173__6,registerOutputs_173__5,registerOutputs_173__4,
           registerOutputs_173__3,registerOutputs_173__2,registerOutputs_173__1,
           registerOutputs_173__0})) ;
    Mux2_16 loop1_174_y (.A ({nx35933,nx36075,nx36217,nx36359,nx36501,nx36643,
            nx36785,nx36927,nx37069,nx37211,nx37353,nx37495,nx37637,nx37779,
            nx37921,nx38063}), .B ({nx33689,nx33829,nx33967,nx34105,nx34243,
            nx34381,nx34519,nx34659,nx34801,nx34943,nx35085,nx35227,nx35369,
            nx35511,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35653), .C ({inputRegisters_174__15,inputRegisters_174__14,
            inputRegisters_174__13,inputRegisters_174__12,inputRegisters_174__11
            ,inputRegisters_174__10,inputRegisters_174__9,inputRegisters_174__8,
            inputRegisters_174__7,inputRegisters_174__6,inputRegisters_174__5,
            inputRegisters_174__4,inputRegisters_174__3,inputRegisters_174__2,
            inputRegisters_174__1,inputRegisters_174__0})) ;
    Reg_16 loop1_174_x (.D ({inputRegisters_174__15,inputRegisters_174__14,
           inputRegisters_174__13,inputRegisters_174__12,inputRegisters_174__11,
           inputRegisters_174__10,inputRegisters_174__9,inputRegisters_174__8,
           inputRegisters_174__7,inputRegisters_174__6,inputRegisters_174__5,
           inputRegisters_174__4,inputRegisters_174__3,inputRegisters_174__2,
           inputRegisters_174__1,inputRegisters_174__0}), .en (
           enableRegister_174), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_174__15,registerOutputs_174__14,
           registerOutputs_174__13,registerOutputs_174__12,
           registerOutputs_174__11,registerOutputs_174__10,
           registerOutputs_174__9,registerOutputs_174__8,registerOutputs_174__7,
           registerOutputs_174__6,registerOutputs_174__5,registerOutputs_174__4,
           registerOutputs_174__3,registerOutputs_174__2,registerOutputs_174__1,
           registerOutputs_174__0})) ;
    Mux2_16 loop1_175_y (.A ({nx35935,nx36077,nx36219,nx36361,nx36503,nx36645,
            nx36787,nx36929,nx37071,nx37213,nx37355,nx37497,nx37639,nx37781,
            nx37923,nx38065}), .B ({nx33691,nx33829,nx33967,nx34105,nx34243,
            nx34381,nx34519,nx34661,nx34803,nx34945,nx35087,nx35229,nx35371,
            nx35513,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35655), .C ({inputRegisters_175__15,inputRegisters_175__14,
            inputRegisters_175__13,inputRegisters_175__12,inputRegisters_175__11
            ,inputRegisters_175__10,inputRegisters_175__9,inputRegisters_175__8,
            inputRegisters_175__7,inputRegisters_175__6,inputRegisters_175__5,
            inputRegisters_175__4,inputRegisters_175__3,inputRegisters_175__2,
            inputRegisters_175__1,inputRegisters_175__0})) ;
    Reg_16 loop1_175_x (.D ({inputRegisters_175__15,inputRegisters_175__14,
           inputRegisters_175__13,inputRegisters_175__12,inputRegisters_175__11,
           inputRegisters_175__10,inputRegisters_175__9,inputRegisters_175__8,
           inputRegisters_175__7,inputRegisters_175__6,inputRegisters_175__5,
           inputRegisters_175__4,inputRegisters_175__3,inputRegisters_175__2,
           inputRegisters_175__1,inputRegisters_175__0}), .en (
           enableRegister_175), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_175__15,registerOutputs_175__14,
           registerOutputs_175__13,registerOutputs_175__12,
           registerOutputs_175__11,registerOutputs_175__10,
           registerOutputs_175__9,registerOutputs_175__8,registerOutputs_175__7,
           registerOutputs_175__6,registerOutputs_175__5,registerOutputs_175__4,
           registerOutputs_175__3,registerOutputs_175__2,registerOutputs_175__1,
           registerOutputs_175__0})) ;
    Mux2_16 loop1_176_y (.A ({nx35935,nx36077,nx36219,nx36361,nx36503,nx36645,
            nx36787,nx36929,nx37071,nx37213,nx37355,nx37497,nx37639,nx37781,
            nx37923,nx38065}), .B ({nx33691,nx33829,nx33967,nx34105,nx34243,
            nx34381,nx34521,nx34661,nx34803,nx34945,nx35087,nx35229,nx35371,
            nx35513,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35655), .C ({inputRegisters_176__15,inputRegisters_176__14,
            inputRegisters_176__13,inputRegisters_176__12,inputRegisters_176__11
            ,inputRegisters_176__10,inputRegisters_176__9,inputRegisters_176__8,
            inputRegisters_176__7,inputRegisters_176__6,inputRegisters_176__5,
            inputRegisters_176__4,inputRegisters_176__3,inputRegisters_176__2,
            inputRegisters_176__1,inputRegisters_176__0})) ;
    Reg_16 loop1_176_x (.D ({inputRegisters_176__15,inputRegisters_176__14,
           inputRegisters_176__13,inputRegisters_176__12,inputRegisters_176__11,
           inputRegisters_176__10,inputRegisters_176__9,inputRegisters_176__8,
           inputRegisters_176__7,inputRegisters_176__6,inputRegisters_176__5,
           inputRegisters_176__4,inputRegisters_176__3,inputRegisters_176__2,
           inputRegisters_176__1,inputRegisters_176__0}), .en (
           enableRegister_176), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_176__15,registerOutputs_176__14,
           registerOutputs_176__13,registerOutputs_176__12,
           registerOutputs_176__11,registerOutputs_176__10,
           registerOutputs_176__9,registerOutputs_176__8,registerOutputs_176__7,
           registerOutputs_176__6,registerOutputs_176__5,registerOutputs_176__4,
           registerOutputs_176__3,registerOutputs_176__2,registerOutputs_176__1,
           registerOutputs_176__0})) ;
    Mux2_16 loop1_177_y (.A ({nx35935,nx36077,nx36219,nx36361,nx36503,nx36645,
            nx36787,nx36929,nx37071,nx37213,nx37355,nx37497,nx37639,nx37781,
            nx37923,nx38065}), .B ({nx33691,nx33829,nx33967,nx34105,nx34243,
            nx34383,nx34521,nx34661,nx34803,nx34945,nx35087,nx35229,nx35371,
            nx35513,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35655), .C ({inputRegisters_177__15,inputRegisters_177__14,
            inputRegisters_177__13,inputRegisters_177__12,inputRegisters_177__11
            ,inputRegisters_177__10,inputRegisters_177__9,inputRegisters_177__8,
            inputRegisters_177__7,inputRegisters_177__6,inputRegisters_177__5,
            inputRegisters_177__4,inputRegisters_177__3,inputRegisters_177__2,
            inputRegisters_177__1,inputRegisters_177__0})) ;
    Reg_16 loop1_177_x (.D ({inputRegisters_177__15,inputRegisters_177__14,
           inputRegisters_177__13,inputRegisters_177__12,inputRegisters_177__11,
           inputRegisters_177__10,inputRegisters_177__9,inputRegisters_177__8,
           inputRegisters_177__7,inputRegisters_177__6,inputRegisters_177__5,
           inputRegisters_177__4,inputRegisters_177__3,inputRegisters_177__2,
           inputRegisters_177__1,inputRegisters_177__0}), .en (
           enableRegister_177), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_177__15,registerOutputs_177__14,
           registerOutputs_177__13,registerOutputs_177__12,
           registerOutputs_177__11,registerOutputs_177__10,
           registerOutputs_177__9,registerOutputs_177__8,registerOutputs_177__7,
           registerOutputs_177__6,registerOutputs_177__5,registerOutputs_177__4,
           registerOutputs_177__3,registerOutputs_177__2,registerOutputs_177__1,
           registerOutputs_177__0})) ;
    Mux2_16 loop1_178_y (.A ({nx35935,nx36077,nx36219,nx36361,nx36503,nx36645,
            nx36787,nx36929,nx37071,nx37213,nx37355,nx37497,nx37639,nx37781,
            nx37923,nx38065}), .B ({nx33691,nx33829,nx33967,nx34105,nx34245,
            nx34383,nx34521,nx34661,nx34803,nx34945,nx35087,nx35229,nx35371,
            nx35513,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35655), .C ({inputRegisters_178__15,inputRegisters_178__14,
            inputRegisters_178__13,inputRegisters_178__12,inputRegisters_178__11
            ,inputRegisters_178__10,inputRegisters_178__9,inputRegisters_178__8,
            inputRegisters_178__7,inputRegisters_178__6,inputRegisters_178__5,
            inputRegisters_178__4,inputRegisters_178__3,inputRegisters_178__2,
            inputRegisters_178__1,inputRegisters_178__0})) ;
    Reg_16 loop1_178_x (.D ({inputRegisters_178__15,inputRegisters_178__14,
           inputRegisters_178__13,inputRegisters_178__12,inputRegisters_178__11,
           inputRegisters_178__10,inputRegisters_178__9,inputRegisters_178__8,
           inputRegisters_178__7,inputRegisters_178__6,inputRegisters_178__5,
           inputRegisters_178__4,inputRegisters_178__3,inputRegisters_178__2,
           inputRegisters_178__1,inputRegisters_178__0}), .en (
           enableRegister_178), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_178__15,registerOutputs_178__14,
           registerOutputs_178__13,registerOutputs_178__12,
           registerOutputs_178__11,registerOutputs_178__10,
           registerOutputs_178__9,registerOutputs_178__8,registerOutputs_178__7,
           registerOutputs_178__6,registerOutputs_178__5,registerOutputs_178__4,
           registerOutputs_178__3,registerOutputs_178__2,registerOutputs_178__1,
           registerOutputs_178__0})) ;
    Mux2_16 loop1_179_y (.A ({nx35935,nx36077,nx36219,nx36361,nx36503,nx36645,
            nx36787,nx36929,nx37071,nx37213,nx37355,nx37497,nx37639,nx37781,
            nx37923,nx38065}), .B ({nx33691,nx33829,nx33967,nx34107,nx34245,
            nx34383,nx34521,nx34661,nx34803,nx34945,nx35087,nx35229,nx35371,
            nx35513,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35655), .C ({inputRegisters_179__15,inputRegisters_179__14,
            inputRegisters_179__13,inputRegisters_179__12,inputRegisters_179__11
            ,inputRegisters_179__10,inputRegisters_179__9,inputRegisters_179__8,
            inputRegisters_179__7,inputRegisters_179__6,inputRegisters_179__5,
            inputRegisters_179__4,inputRegisters_179__3,inputRegisters_179__2,
            inputRegisters_179__1,inputRegisters_179__0})) ;
    Reg_16 loop1_179_x (.D ({inputRegisters_179__15,inputRegisters_179__14,
           inputRegisters_179__13,inputRegisters_179__12,inputRegisters_179__11,
           inputRegisters_179__10,inputRegisters_179__9,inputRegisters_179__8,
           inputRegisters_179__7,inputRegisters_179__6,inputRegisters_179__5,
           inputRegisters_179__4,inputRegisters_179__3,inputRegisters_179__2,
           inputRegisters_179__1,inputRegisters_179__0}), .en (
           enableRegister_179), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_179__15,registerOutputs_179__14,
           registerOutputs_179__13,registerOutputs_179__12,
           registerOutputs_179__11,registerOutputs_179__10,
           registerOutputs_179__9,registerOutputs_179__8,registerOutputs_179__7,
           registerOutputs_179__6,registerOutputs_179__5,registerOutputs_179__4,
           registerOutputs_179__3,registerOutputs_179__2,registerOutputs_179__1,
           registerOutputs_179__0})) ;
    Mux2_16 loop1_180_y (.A ({nx35935,nx36077,nx36219,nx36361,nx36503,nx36645,
            nx36787,nx36929,nx37071,nx37213,nx37355,nx37497,nx37639,nx37781,
            nx37923,nx38065}), .B ({nx33691,nx33829,nx33969,nx34107,nx34245,
            nx34383,nx34521,nx34661,nx34803,nx34945,nx35087,nx35229,nx35371,
            nx35513,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35655), .C ({inputRegisters_180__15,inputRegisters_180__14,
            inputRegisters_180__13,inputRegisters_180__12,inputRegisters_180__11
            ,inputRegisters_180__10,inputRegisters_180__9,inputRegisters_180__8,
            inputRegisters_180__7,inputRegisters_180__6,inputRegisters_180__5,
            inputRegisters_180__4,inputRegisters_180__3,inputRegisters_180__2,
            inputRegisters_180__1,inputRegisters_180__0})) ;
    Reg_16 loop1_180_x (.D ({inputRegisters_180__15,inputRegisters_180__14,
           inputRegisters_180__13,inputRegisters_180__12,inputRegisters_180__11,
           inputRegisters_180__10,inputRegisters_180__9,inputRegisters_180__8,
           inputRegisters_180__7,inputRegisters_180__6,inputRegisters_180__5,
           inputRegisters_180__4,inputRegisters_180__3,inputRegisters_180__2,
           inputRegisters_180__1,inputRegisters_180__0}), .en (
           enableRegister_180), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_180__15,registerOutputs_180__14,
           registerOutputs_180__13,registerOutputs_180__12,
           registerOutputs_180__11,registerOutputs_180__10,
           registerOutputs_180__9,registerOutputs_180__8,registerOutputs_180__7,
           registerOutputs_180__6,registerOutputs_180__5,registerOutputs_180__4,
           registerOutputs_180__3,registerOutputs_180__2,registerOutputs_180__1,
           registerOutputs_180__0})) ;
    Mux2_16 loop1_181_y (.A ({nx35935,nx36077,nx36219,nx36361,nx36503,nx36645,
            nx36787,nx36929,nx37071,nx37213,nx37355,nx37497,nx37639,nx37781,
            nx37923,nx38065}), .B ({nx33691,nx33831,nx33969,nx34107,nx34245,
            nx34383,nx34521,nx34661,nx34803,nx34945,nx35087,nx35229,nx35371,
            nx35513,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35655), .C ({inputRegisters_181__15,inputRegisters_181__14,
            inputRegisters_181__13,inputRegisters_181__12,inputRegisters_181__11
            ,inputRegisters_181__10,inputRegisters_181__9,inputRegisters_181__8,
            inputRegisters_181__7,inputRegisters_181__6,inputRegisters_181__5,
            inputRegisters_181__4,inputRegisters_181__3,inputRegisters_181__2,
            inputRegisters_181__1,inputRegisters_181__0})) ;
    Reg_16 loop1_181_x (.D ({inputRegisters_181__15,inputRegisters_181__14,
           inputRegisters_181__13,inputRegisters_181__12,inputRegisters_181__11,
           inputRegisters_181__10,inputRegisters_181__9,inputRegisters_181__8,
           inputRegisters_181__7,inputRegisters_181__6,inputRegisters_181__5,
           inputRegisters_181__4,inputRegisters_181__3,inputRegisters_181__2,
           inputRegisters_181__1,inputRegisters_181__0}), .en (
           enableRegister_181), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_181__15,registerOutputs_181__14,
           registerOutputs_181__13,registerOutputs_181__12,
           registerOutputs_181__11,registerOutputs_181__10,
           registerOutputs_181__9,registerOutputs_181__8,registerOutputs_181__7,
           registerOutputs_181__6,registerOutputs_181__5,registerOutputs_181__4,
           registerOutputs_181__3,registerOutputs_181__2,registerOutputs_181__1,
           registerOutputs_181__0})) ;
    Mux2_16 loop1_182_y (.A ({nx35937,nx36079,nx36221,nx36363,nx36505,nx36647,
            nx36789,nx36931,nx37073,nx37215,nx37357,nx37499,nx37641,nx37783,
            nx37925,nx38067}), .B ({nx33693,nx33831,nx33969,nx34107,nx34245,
            nx34383,nx34521,nx34663,nx34805,nx34947,nx35089,nx35231,nx35373,
            nx35515,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35657), .C ({inputRegisters_182__15,inputRegisters_182__14,
            inputRegisters_182__13,inputRegisters_182__12,inputRegisters_182__11
            ,inputRegisters_182__10,inputRegisters_182__9,inputRegisters_182__8,
            inputRegisters_182__7,inputRegisters_182__6,inputRegisters_182__5,
            inputRegisters_182__4,inputRegisters_182__3,inputRegisters_182__2,
            inputRegisters_182__1,inputRegisters_182__0})) ;
    Reg_16 loop1_182_x (.D ({inputRegisters_182__15,inputRegisters_182__14,
           inputRegisters_182__13,inputRegisters_182__12,inputRegisters_182__11,
           inputRegisters_182__10,inputRegisters_182__9,inputRegisters_182__8,
           inputRegisters_182__7,inputRegisters_182__6,inputRegisters_182__5,
           inputRegisters_182__4,inputRegisters_182__3,inputRegisters_182__2,
           inputRegisters_182__1,inputRegisters_182__0}), .en (
           enableRegister_182), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_182__15,registerOutputs_182__14,
           registerOutputs_182__13,registerOutputs_182__12,
           registerOutputs_182__11,registerOutputs_182__10,
           registerOutputs_182__9,registerOutputs_182__8,registerOutputs_182__7,
           registerOutputs_182__6,registerOutputs_182__5,registerOutputs_182__4,
           registerOutputs_182__3,registerOutputs_182__2,registerOutputs_182__1,
           registerOutputs_182__0})) ;
    Mux2_16 loop1_183_y (.A ({nx35937,nx36079,nx36221,nx36363,nx36505,nx36647,
            nx36789,nx36931,nx37073,nx37215,nx37357,nx37499,nx37641,nx37783,
            nx37925,nx38067}), .B ({nx33693,nx33831,nx33969,nx34107,nx34245,
            nx34383,nx34523,nx34663,nx34805,nx34947,nx35089,nx35231,nx35373,
            nx35515,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35657), .C ({inputRegisters_183__15,inputRegisters_183__14,
            inputRegisters_183__13,inputRegisters_183__12,inputRegisters_183__11
            ,inputRegisters_183__10,inputRegisters_183__9,inputRegisters_183__8,
            inputRegisters_183__7,inputRegisters_183__6,inputRegisters_183__5,
            inputRegisters_183__4,inputRegisters_183__3,inputRegisters_183__2,
            inputRegisters_183__1,inputRegisters_183__0})) ;
    Reg_16 loop1_183_x (.D ({inputRegisters_183__15,inputRegisters_183__14,
           inputRegisters_183__13,inputRegisters_183__12,inputRegisters_183__11,
           inputRegisters_183__10,inputRegisters_183__9,inputRegisters_183__8,
           inputRegisters_183__7,inputRegisters_183__6,inputRegisters_183__5,
           inputRegisters_183__4,inputRegisters_183__3,inputRegisters_183__2,
           inputRegisters_183__1,inputRegisters_183__0}), .en (
           enableRegister_183), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_183__15,registerOutputs_183__14,
           registerOutputs_183__13,registerOutputs_183__12,
           registerOutputs_183__11,registerOutputs_183__10,
           registerOutputs_183__9,registerOutputs_183__8,registerOutputs_183__7,
           registerOutputs_183__6,registerOutputs_183__5,registerOutputs_183__4,
           registerOutputs_183__3,registerOutputs_183__2,registerOutputs_183__1,
           registerOutputs_183__0})) ;
    Mux2_16 loop1_184_y (.A ({nx35937,nx36079,nx36221,nx36363,nx36505,nx36647,
            nx36789,nx36931,nx37073,nx37215,nx37357,nx37499,nx37641,nx37783,
            nx37925,nx38067}), .B ({nx33693,nx33831,nx33969,nx34107,nx34245,
            nx34385,nx34523,nx34663,nx34805,nx34947,nx35089,nx35231,nx35373,
            nx35515,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35657), .C ({inputRegisters_184__15,inputRegisters_184__14,
            inputRegisters_184__13,inputRegisters_184__12,inputRegisters_184__11
            ,inputRegisters_184__10,inputRegisters_184__9,inputRegisters_184__8,
            inputRegisters_184__7,inputRegisters_184__6,inputRegisters_184__5,
            inputRegisters_184__4,inputRegisters_184__3,inputRegisters_184__2,
            inputRegisters_184__1,inputRegisters_184__0})) ;
    Reg_16 loop1_184_x (.D ({inputRegisters_184__15,inputRegisters_184__14,
           inputRegisters_184__13,inputRegisters_184__12,inputRegisters_184__11,
           inputRegisters_184__10,inputRegisters_184__9,inputRegisters_184__8,
           inputRegisters_184__7,inputRegisters_184__6,inputRegisters_184__5,
           inputRegisters_184__4,inputRegisters_184__3,inputRegisters_184__2,
           inputRegisters_184__1,inputRegisters_184__0}), .en (
           enableRegister_184), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_184__15,registerOutputs_184__14,
           registerOutputs_184__13,registerOutputs_184__12,
           registerOutputs_184__11,registerOutputs_184__10,
           registerOutputs_184__9,registerOutputs_184__8,registerOutputs_184__7,
           registerOutputs_184__6,registerOutputs_184__5,registerOutputs_184__4,
           registerOutputs_184__3,registerOutputs_184__2,registerOutputs_184__1,
           registerOutputs_184__0})) ;
    Mux2_16 loop1_185_y (.A ({nx35937,nx36079,nx36221,nx36363,nx36505,nx36647,
            nx36789,nx36931,nx37073,nx37215,nx37357,nx37499,nx37641,nx37783,
            nx37925,nx38067}), .B ({nx33693,nx33831,nx33969,nx34107,nx34247,
            nx34385,nx34523,nx34663,nx34805,nx34947,nx35089,nx35231,nx35373,
            nx35515,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35657), .C ({inputRegisters_185__15,inputRegisters_185__14,
            inputRegisters_185__13,inputRegisters_185__12,inputRegisters_185__11
            ,inputRegisters_185__10,inputRegisters_185__9,inputRegisters_185__8,
            inputRegisters_185__7,inputRegisters_185__6,inputRegisters_185__5,
            inputRegisters_185__4,inputRegisters_185__3,inputRegisters_185__2,
            inputRegisters_185__1,inputRegisters_185__0})) ;
    Reg_16 loop1_185_x (.D ({inputRegisters_185__15,inputRegisters_185__14,
           inputRegisters_185__13,inputRegisters_185__12,inputRegisters_185__11,
           inputRegisters_185__10,inputRegisters_185__9,inputRegisters_185__8,
           inputRegisters_185__7,inputRegisters_185__6,inputRegisters_185__5,
           inputRegisters_185__4,inputRegisters_185__3,inputRegisters_185__2,
           inputRegisters_185__1,inputRegisters_185__0}), .en (
           enableRegister_185), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_185__15,registerOutputs_185__14,
           registerOutputs_185__13,registerOutputs_185__12,
           registerOutputs_185__11,registerOutputs_185__10,
           registerOutputs_185__9,registerOutputs_185__8,registerOutputs_185__7,
           registerOutputs_185__6,registerOutputs_185__5,registerOutputs_185__4,
           registerOutputs_185__3,registerOutputs_185__2,registerOutputs_185__1,
           registerOutputs_185__0})) ;
    Mux2_16 loop1_186_y (.A ({nx35937,nx36079,nx36221,nx36363,nx36505,nx36647,
            nx36789,nx36931,nx37073,nx37215,nx37357,nx37499,nx37641,nx37783,
            nx37925,nx38067}), .B ({nx33693,nx33831,nx33969,nx34109,nx34247,
            nx34385,nx34523,nx34663,nx34805,nx34947,nx35089,nx35231,nx35373,
            nx35515,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35657), .C ({inputRegisters_186__15,inputRegisters_186__14,
            inputRegisters_186__13,inputRegisters_186__12,inputRegisters_186__11
            ,inputRegisters_186__10,inputRegisters_186__9,inputRegisters_186__8,
            inputRegisters_186__7,inputRegisters_186__6,inputRegisters_186__5,
            inputRegisters_186__4,inputRegisters_186__3,inputRegisters_186__2,
            inputRegisters_186__1,inputRegisters_186__0})) ;
    Reg_16 loop1_186_x (.D ({inputRegisters_186__15,inputRegisters_186__14,
           inputRegisters_186__13,inputRegisters_186__12,inputRegisters_186__11,
           inputRegisters_186__10,inputRegisters_186__9,inputRegisters_186__8,
           inputRegisters_186__7,inputRegisters_186__6,inputRegisters_186__5,
           inputRegisters_186__4,inputRegisters_186__3,inputRegisters_186__2,
           inputRegisters_186__1,inputRegisters_186__0}), .en (
           enableRegister_186), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_186__15,registerOutputs_186__14,
           registerOutputs_186__13,registerOutputs_186__12,
           registerOutputs_186__11,registerOutputs_186__10,
           registerOutputs_186__9,registerOutputs_186__8,registerOutputs_186__7,
           registerOutputs_186__6,registerOutputs_186__5,registerOutputs_186__4,
           registerOutputs_186__3,registerOutputs_186__2,registerOutputs_186__1,
           registerOutputs_186__0})) ;
    Mux2_16 loop1_187_y (.A ({nx35937,nx36079,nx36221,nx36363,nx36505,nx36647,
            nx36789,nx36931,nx37073,nx37215,nx37357,nx37499,nx37641,nx37783,
            nx37925,nx38067}), .B ({nx33693,nx33831,nx33971,nx34109,nx34247,
            nx34385,nx34523,nx34663,nx34805,nx34947,nx35089,nx35231,nx35373,
            nx35515,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35657), .C ({inputRegisters_187__15,inputRegisters_187__14,
            inputRegisters_187__13,inputRegisters_187__12,inputRegisters_187__11
            ,inputRegisters_187__10,inputRegisters_187__9,inputRegisters_187__8,
            inputRegisters_187__7,inputRegisters_187__6,inputRegisters_187__5,
            inputRegisters_187__4,inputRegisters_187__3,inputRegisters_187__2,
            inputRegisters_187__1,inputRegisters_187__0})) ;
    Reg_16 loop1_187_x (.D ({inputRegisters_187__15,inputRegisters_187__14,
           inputRegisters_187__13,inputRegisters_187__12,inputRegisters_187__11,
           inputRegisters_187__10,inputRegisters_187__9,inputRegisters_187__8,
           inputRegisters_187__7,inputRegisters_187__6,inputRegisters_187__5,
           inputRegisters_187__4,inputRegisters_187__3,inputRegisters_187__2,
           inputRegisters_187__1,inputRegisters_187__0}), .en (
           enableRegister_187), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_187__15,registerOutputs_187__14,
           registerOutputs_187__13,registerOutputs_187__12,
           registerOutputs_187__11,registerOutputs_187__10,
           registerOutputs_187__9,registerOutputs_187__8,registerOutputs_187__7,
           registerOutputs_187__6,registerOutputs_187__5,registerOutputs_187__4,
           registerOutputs_187__3,registerOutputs_187__2,registerOutputs_187__1,
           registerOutputs_187__0})) ;
    Mux2_16 loop1_188_y (.A ({nx35937,nx36079,nx36221,nx36363,nx36505,nx36647,
            nx36789,nx36931,nx37073,nx37215,nx37357,nx37499,nx37641,nx37783,
            nx37925,nx38067}), .B ({nx33693,nx33833,nx33971,nx34109,nx34247,
            nx34385,nx34523,nx34663,nx34805,nx34947,nx35089,nx35231,nx35373,
            nx35515,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35657), .C ({inputRegisters_188__15,inputRegisters_188__14,
            inputRegisters_188__13,inputRegisters_188__12,inputRegisters_188__11
            ,inputRegisters_188__10,inputRegisters_188__9,inputRegisters_188__8,
            inputRegisters_188__7,inputRegisters_188__6,inputRegisters_188__5,
            inputRegisters_188__4,inputRegisters_188__3,inputRegisters_188__2,
            inputRegisters_188__1,inputRegisters_188__0})) ;
    Reg_16 loop1_188_x (.D ({inputRegisters_188__15,inputRegisters_188__14,
           inputRegisters_188__13,inputRegisters_188__12,inputRegisters_188__11,
           inputRegisters_188__10,inputRegisters_188__9,inputRegisters_188__8,
           inputRegisters_188__7,inputRegisters_188__6,inputRegisters_188__5,
           inputRegisters_188__4,inputRegisters_188__3,inputRegisters_188__2,
           inputRegisters_188__1,inputRegisters_188__0}), .en (
           enableRegister_188), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_188__15,registerOutputs_188__14,
           registerOutputs_188__13,registerOutputs_188__12,
           registerOutputs_188__11,registerOutputs_188__10,
           registerOutputs_188__9,registerOutputs_188__8,registerOutputs_188__7,
           registerOutputs_188__6,registerOutputs_188__5,registerOutputs_188__4,
           registerOutputs_188__3,registerOutputs_188__2,registerOutputs_188__1,
           registerOutputs_188__0})) ;
    Mux2_16 loop1_189_y (.A ({nx35939,nx36081,nx36223,nx36365,nx36507,nx36649,
            nx36791,nx36933,nx37075,nx37217,nx37359,nx37501,nx37643,nx37785,
            nx37927,nx38069}), .B ({nx33695,nx33833,nx33971,nx34109,nx34247,
            nx34385,nx34523,nx34665,nx34807,nx34949,nx35091,nx35233,nx35375,
            nx35517,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35659), .C ({inputRegisters_189__15,inputRegisters_189__14,
            inputRegisters_189__13,inputRegisters_189__12,inputRegisters_189__11
            ,inputRegisters_189__10,inputRegisters_189__9,inputRegisters_189__8,
            inputRegisters_189__7,inputRegisters_189__6,inputRegisters_189__5,
            inputRegisters_189__4,inputRegisters_189__3,inputRegisters_189__2,
            inputRegisters_189__1,inputRegisters_189__0})) ;
    Reg_16 loop1_189_x (.D ({inputRegisters_189__15,inputRegisters_189__14,
           inputRegisters_189__13,inputRegisters_189__12,inputRegisters_189__11,
           inputRegisters_189__10,inputRegisters_189__9,inputRegisters_189__8,
           inputRegisters_189__7,inputRegisters_189__6,inputRegisters_189__5,
           inputRegisters_189__4,inputRegisters_189__3,inputRegisters_189__2,
           inputRegisters_189__1,inputRegisters_189__0}), .en (
           enableRegister_189), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_189__15,registerOutputs_189__14,
           registerOutputs_189__13,registerOutputs_189__12,
           registerOutputs_189__11,registerOutputs_189__10,
           registerOutputs_189__9,registerOutputs_189__8,registerOutputs_189__7,
           registerOutputs_189__6,registerOutputs_189__5,registerOutputs_189__4,
           registerOutputs_189__3,registerOutputs_189__2,registerOutputs_189__1,
           registerOutputs_189__0})) ;
    Mux2_16 loop1_190_y (.A ({nx35939,nx36081,nx36223,nx36365,nx36507,nx36649,
            nx36791,nx36933,nx37075,nx37217,nx37359,nx37501,nx37643,nx37785,
            nx37927,nx38069}), .B ({nx33695,nx33833,nx33971,nx34109,nx34247,
            nx34385,nx34525,nx34665,nx34807,nx34949,nx35091,nx35233,nx35375,
            nx35517,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35659), .C ({inputRegisters_190__15,inputRegisters_190__14,
            inputRegisters_190__13,inputRegisters_190__12,inputRegisters_190__11
            ,inputRegisters_190__10,inputRegisters_190__9,inputRegisters_190__8,
            inputRegisters_190__7,inputRegisters_190__6,inputRegisters_190__5,
            inputRegisters_190__4,inputRegisters_190__3,inputRegisters_190__2,
            inputRegisters_190__1,inputRegisters_190__0})) ;
    Reg_16 loop1_190_x (.D ({inputRegisters_190__15,inputRegisters_190__14,
           inputRegisters_190__13,inputRegisters_190__12,inputRegisters_190__11,
           inputRegisters_190__10,inputRegisters_190__9,inputRegisters_190__8,
           inputRegisters_190__7,inputRegisters_190__6,inputRegisters_190__5,
           inputRegisters_190__4,inputRegisters_190__3,inputRegisters_190__2,
           inputRegisters_190__1,inputRegisters_190__0}), .en (
           enableRegister_190), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_190__15,registerOutputs_190__14,
           registerOutputs_190__13,registerOutputs_190__12,
           registerOutputs_190__11,registerOutputs_190__10,
           registerOutputs_190__9,registerOutputs_190__8,registerOutputs_190__7,
           registerOutputs_190__6,registerOutputs_190__5,registerOutputs_190__4,
           registerOutputs_190__3,registerOutputs_190__2,registerOutputs_190__1,
           registerOutputs_190__0})) ;
    Mux2_16 loop1_191_y (.A ({nx35939,nx36081,nx36223,nx36365,nx36507,nx36649,
            nx36791,nx36933,nx37075,nx37217,nx37359,nx37501,nx37643,nx37785,
            nx37927,nx38069}), .B ({nx33695,nx33833,nx33971,nx34109,nx34247,
            nx34387,nx34525,nx34665,nx34807,nx34949,nx35091,nx35233,nx35375,
            nx35517,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35659), .C ({inputRegisters_191__15,inputRegisters_191__14,
            inputRegisters_191__13,inputRegisters_191__12,inputRegisters_191__11
            ,inputRegisters_191__10,inputRegisters_191__9,inputRegisters_191__8,
            inputRegisters_191__7,inputRegisters_191__6,inputRegisters_191__5,
            inputRegisters_191__4,inputRegisters_191__3,inputRegisters_191__2,
            inputRegisters_191__1,inputRegisters_191__0})) ;
    Reg_16 loop1_191_x (.D ({inputRegisters_191__15,inputRegisters_191__14,
           inputRegisters_191__13,inputRegisters_191__12,inputRegisters_191__11,
           inputRegisters_191__10,inputRegisters_191__9,inputRegisters_191__8,
           inputRegisters_191__7,inputRegisters_191__6,inputRegisters_191__5,
           inputRegisters_191__4,inputRegisters_191__3,inputRegisters_191__2,
           inputRegisters_191__1,inputRegisters_191__0}), .en (
           enableRegister_191), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_191__15,registerOutputs_191__14,
           registerOutputs_191__13,registerOutputs_191__12,
           registerOutputs_191__11,registerOutputs_191__10,
           registerOutputs_191__9,registerOutputs_191__8,registerOutputs_191__7,
           registerOutputs_191__6,registerOutputs_191__5,registerOutputs_191__4,
           registerOutputs_191__3,registerOutputs_191__2,registerOutputs_191__1,
           registerOutputs_191__0})) ;
    Mux2_16 loop1_192_y (.A ({nx35939,nx36081,nx36223,nx36365,nx36507,nx36649,
            nx36791,nx36933,nx37075,nx37217,nx37359,nx37501,nx37643,nx37785,
            nx37927,nx38069}), .B ({nx33695,nx33833,nx33971,nx34109,nx34249,
            nx34387,nx34525,nx34665,nx34807,nx34949,nx35091,nx35233,nx35375,
            nx35517,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35659), .C ({inputRegisters_192__15,inputRegisters_192__14,
            inputRegisters_192__13,inputRegisters_192__12,inputRegisters_192__11
            ,inputRegisters_192__10,inputRegisters_192__9,inputRegisters_192__8,
            inputRegisters_192__7,inputRegisters_192__6,inputRegisters_192__5,
            inputRegisters_192__4,inputRegisters_192__3,inputRegisters_192__2,
            inputRegisters_192__1,inputRegisters_192__0})) ;
    Reg_16 loop1_192_x (.D ({inputRegisters_192__15,inputRegisters_192__14,
           inputRegisters_192__13,inputRegisters_192__12,inputRegisters_192__11,
           inputRegisters_192__10,inputRegisters_192__9,inputRegisters_192__8,
           inputRegisters_192__7,inputRegisters_192__6,inputRegisters_192__5,
           inputRegisters_192__4,inputRegisters_192__3,inputRegisters_192__2,
           inputRegisters_192__1,inputRegisters_192__0}), .en (
           enableRegister_192), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_192__15,registerOutputs_192__14,
           registerOutputs_192__13,registerOutputs_192__12,
           registerOutputs_192__11,registerOutputs_192__10,
           registerOutputs_192__9,registerOutputs_192__8,registerOutputs_192__7,
           registerOutputs_192__6,registerOutputs_192__5,registerOutputs_192__4,
           registerOutputs_192__3,registerOutputs_192__2,registerOutputs_192__1,
           registerOutputs_192__0})) ;
    Mux2_16 loop1_193_y (.A ({nx35939,nx36081,nx36223,nx36365,nx36507,nx36649,
            nx36791,nx36933,nx37075,nx37217,nx37359,nx37501,nx37643,nx37785,
            nx37927,nx38069}), .B ({nx33695,nx33833,nx33971,nx34111,nx34249,
            nx34387,nx34525,nx34665,nx34807,nx34949,nx35091,nx35233,nx35375,
            nx35517,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35659), .C ({inputRegisters_193__15,inputRegisters_193__14,
            inputRegisters_193__13,inputRegisters_193__12,inputRegisters_193__11
            ,inputRegisters_193__10,inputRegisters_193__9,inputRegisters_193__8,
            inputRegisters_193__7,inputRegisters_193__6,inputRegisters_193__5,
            inputRegisters_193__4,inputRegisters_193__3,inputRegisters_193__2,
            inputRegisters_193__1,inputRegisters_193__0})) ;
    Reg_16 loop1_193_x (.D ({inputRegisters_193__15,inputRegisters_193__14,
           inputRegisters_193__13,inputRegisters_193__12,inputRegisters_193__11,
           inputRegisters_193__10,inputRegisters_193__9,inputRegisters_193__8,
           inputRegisters_193__7,inputRegisters_193__6,inputRegisters_193__5,
           inputRegisters_193__4,inputRegisters_193__3,inputRegisters_193__2,
           inputRegisters_193__1,inputRegisters_193__0}), .en (
           enableRegister_193), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_193__15,registerOutputs_193__14,
           registerOutputs_193__13,registerOutputs_193__12,
           registerOutputs_193__11,registerOutputs_193__10,
           registerOutputs_193__9,registerOutputs_193__8,registerOutputs_193__7,
           registerOutputs_193__6,registerOutputs_193__5,registerOutputs_193__4,
           registerOutputs_193__3,registerOutputs_193__2,registerOutputs_193__1,
           registerOutputs_193__0})) ;
    Mux2_16 loop1_194_y (.A ({nx35939,nx36081,nx36223,nx36365,nx36507,nx36649,
            nx36791,nx36933,nx37075,nx37217,nx37359,nx37501,nx37643,nx37785,
            nx37927,nx38069}), .B ({nx33695,nx33833,nx33973,nx34111,nx34249,
            nx34387,nx34525,nx34665,nx34807,nx34949,nx35091,nx35233,nx35375,
            nx35517,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35659), .C ({inputRegisters_194__15,inputRegisters_194__14,
            inputRegisters_194__13,inputRegisters_194__12,inputRegisters_194__11
            ,inputRegisters_194__10,inputRegisters_194__9,inputRegisters_194__8,
            inputRegisters_194__7,inputRegisters_194__6,inputRegisters_194__5,
            inputRegisters_194__4,inputRegisters_194__3,inputRegisters_194__2,
            inputRegisters_194__1,inputRegisters_194__0})) ;
    Reg_16 loop1_194_x (.D ({inputRegisters_194__15,inputRegisters_194__14,
           inputRegisters_194__13,inputRegisters_194__12,inputRegisters_194__11,
           inputRegisters_194__10,inputRegisters_194__9,inputRegisters_194__8,
           inputRegisters_194__7,inputRegisters_194__6,inputRegisters_194__5,
           inputRegisters_194__4,inputRegisters_194__3,inputRegisters_194__2,
           inputRegisters_194__1,inputRegisters_194__0}), .en (
           enableRegister_194), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_194__15,registerOutputs_194__14,
           registerOutputs_194__13,registerOutputs_194__12,
           registerOutputs_194__11,registerOutputs_194__10,
           registerOutputs_194__9,registerOutputs_194__8,registerOutputs_194__7,
           registerOutputs_194__6,registerOutputs_194__5,registerOutputs_194__4,
           registerOutputs_194__3,registerOutputs_194__2,registerOutputs_194__1,
           registerOutputs_194__0})) ;
    Mux2_16 loop1_195_y (.A ({nx35939,nx36081,nx36223,nx36365,nx36507,nx36649,
            nx36791,nx36933,nx37075,nx37217,nx37359,nx37501,nx37643,nx37785,
            nx37927,nx38069}), .B ({nx33695,nx33835,nx33973,nx34111,nx34249,
            nx34387,nx34525,nx34665,nx34807,nx34949,nx35091,nx35233,nx35375,
            nx35517,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35659), .C ({inputRegisters_195__15,inputRegisters_195__14,
            inputRegisters_195__13,inputRegisters_195__12,inputRegisters_195__11
            ,inputRegisters_195__10,inputRegisters_195__9,inputRegisters_195__8,
            inputRegisters_195__7,inputRegisters_195__6,inputRegisters_195__5,
            inputRegisters_195__4,inputRegisters_195__3,inputRegisters_195__2,
            inputRegisters_195__1,inputRegisters_195__0})) ;
    Reg_16 loop1_195_x (.D ({inputRegisters_195__15,inputRegisters_195__14,
           inputRegisters_195__13,inputRegisters_195__12,inputRegisters_195__11,
           inputRegisters_195__10,inputRegisters_195__9,inputRegisters_195__8,
           inputRegisters_195__7,inputRegisters_195__6,inputRegisters_195__5,
           inputRegisters_195__4,inputRegisters_195__3,inputRegisters_195__2,
           inputRegisters_195__1,inputRegisters_195__0}), .en (
           enableRegister_195), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_195__15,registerOutputs_195__14,
           registerOutputs_195__13,registerOutputs_195__12,
           registerOutputs_195__11,registerOutputs_195__10,
           registerOutputs_195__9,registerOutputs_195__8,registerOutputs_195__7,
           registerOutputs_195__6,registerOutputs_195__5,registerOutputs_195__4,
           registerOutputs_195__3,registerOutputs_195__2,registerOutputs_195__1,
           registerOutputs_195__0})) ;
    Mux2_16 loop1_196_y (.A ({nx35941,nx36083,nx36225,nx36367,nx36509,nx36651,
            nx36793,nx36935,nx37077,nx37219,nx37361,nx37503,nx37645,nx37787,
            nx37929,nx38071}), .B ({nx33697,nx33835,nx33973,nx34111,nx34249,
            nx34387,nx34525,nx34667,nx34809,nx34951,nx35093,nx35235,nx35377,
            nx35519,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35661), .C ({inputRegisters_196__15,inputRegisters_196__14,
            inputRegisters_196__13,inputRegisters_196__12,inputRegisters_196__11
            ,inputRegisters_196__10,inputRegisters_196__9,inputRegisters_196__8,
            inputRegisters_196__7,inputRegisters_196__6,inputRegisters_196__5,
            inputRegisters_196__4,inputRegisters_196__3,inputRegisters_196__2,
            inputRegisters_196__1,inputRegisters_196__0})) ;
    Reg_16 loop1_196_x (.D ({inputRegisters_196__15,inputRegisters_196__14,
           inputRegisters_196__13,inputRegisters_196__12,inputRegisters_196__11,
           inputRegisters_196__10,inputRegisters_196__9,inputRegisters_196__8,
           inputRegisters_196__7,inputRegisters_196__6,inputRegisters_196__5,
           inputRegisters_196__4,inputRegisters_196__3,inputRegisters_196__2,
           inputRegisters_196__1,inputRegisters_196__0}), .en (
           enableRegister_196), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_196__15,registerOutputs_196__14,
           registerOutputs_196__13,registerOutputs_196__12,
           registerOutputs_196__11,registerOutputs_196__10,
           registerOutputs_196__9,registerOutputs_196__8,registerOutputs_196__7,
           registerOutputs_196__6,registerOutputs_196__5,registerOutputs_196__4,
           registerOutputs_196__3,registerOutputs_196__2,registerOutputs_196__1,
           registerOutputs_196__0})) ;
    Mux2_16 loop1_197_y (.A ({nx35941,nx36083,nx36225,nx36367,nx36509,nx36651,
            nx36793,nx36935,nx37077,nx37219,nx37361,nx37503,nx37645,nx37787,
            nx37929,nx38071}), .B ({nx33697,nx33835,nx33973,nx34111,nx34249,
            nx34387,nx34527,nx34667,nx34809,nx34951,nx35093,nx35235,nx35377,
            nx35519,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35661), .C ({inputRegisters_197__15,inputRegisters_197__14,
            inputRegisters_197__13,inputRegisters_197__12,inputRegisters_197__11
            ,inputRegisters_197__10,inputRegisters_197__9,inputRegisters_197__8,
            inputRegisters_197__7,inputRegisters_197__6,inputRegisters_197__5,
            inputRegisters_197__4,inputRegisters_197__3,inputRegisters_197__2,
            inputRegisters_197__1,inputRegisters_197__0})) ;
    Reg_16 loop1_197_x (.D ({inputRegisters_197__15,inputRegisters_197__14,
           inputRegisters_197__13,inputRegisters_197__12,inputRegisters_197__11,
           inputRegisters_197__10,inputRegisters_197__9,inputRegisters_197__8,
           inputRegisters_197__7,inputRegisters_197__6,inputRegisters_197__5,
           inputRegisters_197__4,inputRegisters_197__3,inputRegisters_197__2,
           inputRegisters_197__1,inputRegisters_197__0}), .en (
           enableRegister_197), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_197__15,registerOutputs_197__14,
           registerOutputs_197__13,registerOutputs_197__12,
           registerOutputs_197__11,registerOutputs_197__10,
           registerOutputs_197__9,registerOutputs_197__8,registerOutputs_197__7,
           registerOutputs_197__6,registerOutputs_197__5,registerOutputs_197__4,
           registerOutputs_197__3,registerOutputs_197__2,registerOutputs_197__1,
           registerOutputs_197__0})) ;
    Mux2_16 loop1_198_y (.A ({nx35941,nx36083,nx36225,nx36367,nx36509,nx36651,
            nx36793,nx36935,nx37077,nx37219,nx37361,nx37503,nx37645,nx37787,
            nx37929,nx38071}), .B ({nx33697,nx33835,nx33973,nx34111,nx34249,
            nx34389,nx34527,nx34667,nx34809,nx34951,nx35093,nx35235,nx35377,
            nx35519,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35661), .C ({inputRegisters_198__15,inputRegisters_198__14,
            inputRegisters_198__13,inputRegisters_198__12,inputRegisters_198__11
            ,inputRegisters_198__10,inputRegisters_198__9,inputRegisters_198__8,
            inputRegisters_198__7,inputRegisters_198__6,inputRegisters_198__5,
            inputRegisters_198__4,inputRegisters_198__3,inputRegisters_198__2,
            inputRegisters_198__1,inputRegisters_198__0})) ;
    Reg_16 loop1_198_x (.D ({inputRegisters_198__15,inputRegisters_198__14,
           inputRegisters_198__13,inputRegisters_198__12,inputRegisters_198__11,
           inputRegisters_198__10,inputRegisters_198__9,inputRegisters_198__8,
           inputRegisters_198__7,inputRegisters_198__6,inputRegisters_198__5,
           inputRegisters_198__4,inputRegisters_198__3,inputRegisters_198__2,
           inputRegisters_198__1,inputRegisters_198__0}), .en (
           enableRegister_198), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_198__15,registerOutputs_198__14,
           registerOutputs_198__13,registerOutputs_198__12,
           registerOutputs_198__11,registerOutputs_198__10,
           registerOutputs_198__9,registerOutputs_198__8,registerOutputs_198__7,
           registerOutputs_198__6,registerOutputs_198__5,registerOutputs_198__4,
           registerOutputs_198__3,registerOutputs_198__2,registerOutputs_198__1,
           registerOutputs_198__0})) ;
    Mux2_16 loop1_199_y (.A ({nx35941,nx36083,nx36225,nx36367,nx36509,nx36651,
            nx36793,nx36935,nx37077,nx37219,nx37361,nx37503,nx37645,nx37787,
            nx37929,nx38071}), .B ({nx33697,nx33835,nx33973,nx34111,nx34251,
            nx34389,nx34527,nx34667,nx34809,nx34951,nx35093,nx35235,nx35377,
            nx35519,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35661), .C ({inputRegisters_199__15,inputRegisters_199__14,
            inputRegisters_199__13,inputRegisters_199__12,inputRegisters_199__11
            ,inputRegisters_199__10,inputRegisters_199__9,inputRegisters_199__8,
            inputRegisters_199__7,inputRegisters_199__6,inputRegisters_199__5,
            inputRegisters_199__4,inputRegisters_199__3,inputRegisters_199__2,
            inputRegisters_199__1,inputRegisters_199__0})) ;
    Reg_16 loop1_199_x (.D ({inputRegisters_199__15,inputRegisters_199__14,
           inputRegisters_199__13,inputRegisters_199__12,inputRegisters_199__11,
           inputRegisters_199__10,inputRegisters_199__9,inputRegisters_199__8,
           inputRegisters_199__7,inputRegisters_199__6,inputRegisters_199__5,
           inputRegisters_199__4,inputRegisters_199__3,inputRegisters_199__2,
           inputRegisters_199__1,inputRegisters_199__0}), .en (
           enableRegister_199), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_199__15,registerOutputs_199__14,
           registerOutputs_199__13,registerOutputs_199__12,
           registerOutputs_199__11,registerOutputs_199__10,
           registerOutputs_199__9,registerOutputs_199__8,registerOutputs_199__7,
           registerOutputs_199__6,registerOutputs_199__5,registerOutputs_199__4,
           registerOutputs_199__3,registerOutputs_199__2,registerOutputs_199__1,
           registerOutputs_199__0})) ;
    Mux2_16 loop1_200_y (.A ({nx35941,nx36083,nx36225,nx36367,nx36509,nx36651,
            nx36793,nx36935,nx37077,nx37219,nx37361,nx37503,nx37645,nx37787,
            nx37929,nx38071}), .B ({nx33697,nx33835,nx33973,nx34113,nx34251,
            nx34389,nx34527,nx34667,nx34809,nx34951,nx35093,nx35235,nx35377,
            nx35519,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35661), .C ({inputRegisters_200__15,inputRegisters_200__14,
            inputRegisters_200__13,inputRegisters_200__12,inputRegisters_200__11
            ,inputRegisters_200__10,inputRegisters_200__9,inputRegisters_200__8,
            inputRegisters_200__7,inputRegisters_200__6,inputRegisters_200__5,
            inputRegisters_200__4,inputRegisters_200__3,inputRegisters_200__2,
            inputRegisters_200__1,inputRegisters_200__0})) ;
    Reg_16 loop1_200_x (.D ({inputRegisters_200__15,inputRegisters_200__14,
           inputRegisters_200__13,inputRegisters_200__12,inputRegisters_200__11,
           inputRegisters_200__10,inputRegisters_200__9,inputRegisters_200__8,
           inputRegisters_200__7,inputRegisters_200__6,inputRegisters_200__5,
           inputRegisters_200__4,inputRegisters_200__3,inputRegisters_200__2,
           inputRegisters_200__1,inputRegisters_200__0}), .en (
           enableRegister_200), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_200__15,registerOutputs_200__14,
           registerOutputs_200__13,registerOutputs_200__12,
           registerOutputs_200__11,registerOutputs_200__10,
           registerOutputs_200__9,registerOutputs_200__8,registerOutputs_200__7,
           registerOutputs_200__6,registerOutputs_200__5,registerOutputs_200__4,
           registerOutputs_200__3,registerOutputs_200__2,registerOutputs_200__1,
           registerOutputs_200__0})) ;
    Mux2_16 loop1_201_y (.A ({nx35941,nx36083,nx36225,nx36367,nx36509,nx36651,
            nx36793,nx36935,nx37077,nx37219,nx37361,nx37503,nx37645,nx37787,
            nx37929,nx38071}), .B ({nx33697,nx33835,nx33975,nx34113,nx34251,
            nx34389,nx34527,nx34667,nx34809,nx34951,nx35093,nx35235,nx35377,
            nx35519,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35661), .C ({inputRegisters_201__15,inputRegisters_201__14,
            inputRegisters_201__13,inputRegisters_201__12,inputRegisters_201__11
            ,inputRegisters_201__10,inputRegisters_201__9,inputRegisters_201__8,
            inputRegisters_201__7,inputRegisters_201__6,inputRegisters_201__5,
            inputRegisters_201__4,inputRegisters_201__3,inputRegisters_201__2,
            inputRegisters_201__1,inputRegisters_201__0})) ;
    Reg_16 loop1_201_x (.D ({inputRegisters_201__15,inputRegisters_201__14,
           inputRegisters_201__13,inputRegisters_201__12,inputRegisters_201__11,
           inputRegisters_201__10,inputRegisters_201__9,inputRegisters_201__8,
           inputRegisters_201__7,inputRegisters_201__6,inputRegisters_201__5,
           inputRegisters_201__4,inputRegisters_201__3,inputRegisters_201__2,
           inputRegisters_201__1,inputRegisters_201__0}), .en (
           enableRegister_201), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_201__15,registerOutputs_201__14,
           registerOutputs_201__13,registerOutputs_201__12,
           registerOutputs_201__11,registerOutputs_201__10,
           registerOutputs_201__9,registerOutputs_201__8,registerOutputs_201__7,
           registerOutputs_201__6,registerOutputs_201__5,registerOutputs_201__4,
           registerOutputs_201__3,registerOutputs_201__2,registerOutputs_201__1,
           registerOutputs_201__0})) ;
    Mux2_16 loop1_202_y (.A ({nx35941,nx36083,nx36225,nx36367,nx36509,nx36651,
            nx36793,nx36935,nx37077,nx37219,nx37361,nx37503,nx37645,nx37787,
            nx37929,nx38071}), .B ({nx33697,nx33837,nx33975,nx34113,nx34251,
            nx34389,nx34527,nx34667,nx34809,nx34951,nx35093,nx35235,nx35377,
            nx35519,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35661), .C ({inputRegisters_202__15,inputRegisters_202__14,
            inputRegisters_202__13,inputRegisters_202__12,inputRegisters_202__11
            ,inputRegisters_202__10,inputRegisters_202__9,inputRegisters_202__8,
            inputRegisters_202__7,inputRegisters_202__6,inputRegisters_202__5,
            inputRegisters_202__4,inputRegisters_202__3,inputRegisters_202__2,
            inputRegisters_202__1,inputRegisters_202__0})) ;
    Reg_16 loop1_202_x (.D ({inputRegisters_202__15,inputRegisters_202__14,
           inputRegisters_202__13,inputRegisters_202__12,inputRegisters_202__11,
           inputRegisters_202__10,inputRegisters_202__9,inputRegisters_202__8,
           inputRegisters_202__7,inputRegisters_202__6,inputRegisters_202__5,
           inputRegisters_202__4,inputRegisters_202__3,inputRegisters_202__2,
           inputRegisters_202__1,inputRegisters_202__0}), .en (
           enableRegister_202), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_202__15,registerOutputs_202__14,
           registerOutputs_202__13,registerOutputs_202__12,
           registerOutputs_202__11,registerOutputs_202__10,
           registerOutputs_202__9,registerOutputs_202__8,registerOutputs_202__7,
           registerOutputs_202__6,registerOutputs_202__5,registerOutputs_202__4,
           registerOutputs_202__3,registerOutputs_202__2,registerOutputs_202__1,
           registerOutputs_202__0})) ;
    Mux2_16 loop1_203_y (.A ({nx35943,nx36085,nx36227,nx36369,nx36511,nx36653,
            nx36795,nx36937,nx37079,nx37221,nx37363,nx37505,nx37647,nx37789,
            nx37931,nx38073}), .B ({nx33699,nx33837,nx33975,nx34113,nx34251,
            nx34389,nx34527,nx34669,nx34811,nx34953,nx35095,nx35237,nx35379,
            nx35521,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35663), .C ({inputRegisters_203__15,inputRegisters_203__14,
            inputRegisters_203__13,inputRegisters_203__12,inputRegisters_203__11
            ,inputRegisters_203__10,inputRegisters_203__9,inputRegisters_203__8,
            inputRegisters_203__7,inputRegisters_203__6,inputRegisters_203__5,
            inputRegisters_203__4,inputRegisters_203__3,inputRegisters_203__2,
            inputRegisters_203__1,inputRegisters_203__0})) ;
    Reg_16 loop1_203_x (.D ({inputRegisters_203__15,inputRegisters_203__14,
           inputRegisters_203__13,inputRegisters_203__12,inputRegisters_203__11,
           inputRegisters_203__10,inputRegisters_203__9,inputRegisters_203__8,
           inputRegisters_203__7,inputRegisters_203__6,inputRegisters_203__5,
           inputRegisters_203__4,inputRegisters_203__3,inputRegisters_203__2,
           inputRegisters_203__1,inputRegisters_203__0}), .en (
           enableRegister_203), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_203__15,registerOutputs_203__14,
           registerOutputs_203__13,registerOutputs_203__12,
           registerOutputs_203__11,registerOutputs_203__10,
           registerOutputs_203__9,registerOutputs_203__8,registerOutputs_203__7,
           registerOutputs_203__6,registerOutputs_203__5,registerOutputs_203__4,
           registerOutputs_203__3,registerOutputs_203__2,registerOutputs_203__1,
           registerOutputs_203__0})) ;
    Mux2_16 loop1_204_y (.A ({nx35943,nx36085,nx36227,nx36369,nx36511,nx36653,
            nx36795,nx36937,nx37079,nx37221,nx37363,nx37505,nx37647,nx37789,
            nx37931,nx38073}), .B ({nx33699,nx33837,nx33975,nx34113,nx34251,
            nx34389,nx34529,nx34669,nx34811,nx34953,nx35095,nx35237,nx35379,
            nx35521,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35663), .C ({inputRegisters_204__15,inputRegisters_204__14,
            inputRegisters_204__13,inputRegisters_204__12,inputRegisters_204__11
            ,inputRegisters_204__10,inputRegisters_204__9,inputRegisters_204__8,
            inputRegisters_204__7,inputRegisters_204__6,inputRegisters_204__5,
            inputRegisters_204__4,inputRegisters_204__3,inputRegisters_204__2,
            inputRegisters_204__1,inputRegisters_204__0})) ;
    Reg_16 loop1_204_x (.D ({inputRegisters_204__15,inputRegisters_204__14,
           inputRegisters_204__13,inputRegisters_204__12,inputRegisters_204__11,
           inputRegisters_204__10,inputRegisters_204__9,inputRegisters_204__8,
           inputRegisters_204__7,inputRegisters_204__6,inputRegisters_204__5,
           inputRegisters_204__4,inputRegisters_204__3,inputRegisters_204__2,
           inputRegisters_204__1,inputRegisters_204__0}), .en (
           enableRegister_204), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_204__15,registerOutputs_204__14,
           registerOutputs_204__13,registerOutputs_204__12,
           registerOutputs_204__11,registerOutputs_204__10,
           registerOutputs_204__9,registerOutputs_204__8,registerOutputs_204__7,
           registerOutputs_204__6,registerOutputs_204__5,registerOutputs_204__4,
           registerOutputs_204__3,registerOutputs_204__2,registerOutputs_204__1,
           registerOutputs_204__0})) ;
    Mux2_16 loop1_205_y (.A ({nx35943,nx36085,nx36227,nx36369,nx36511,nx36653,
            nx36795,nx36937,nx37079,nx37221,nx37363,nx37505,nx37647,nx37789,
            nx37931,nx38073}), .B ({nx33699,nx33837,nx33975,nx34113,nx34251,
            nx34391,nx34529,nx34669,nx34811,nx34953,nx35095,nx35237,nx35379,
            nx35521,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35663), .C ({inputRegisters_205__15,inputRegisters_205__14,
            inputRegisters_205__13,inputRegisters_205__12,inputRegisters_205__11
            ,inputRegisters_205__10,inputRegisters_205__9,inputRegisters_205__8,
            inputRegisters_205__7,inputRegisters_205__6,inputRegisters_205__5,
            inputRegisters_205__4,inputRegisters_205__3,inputRegisters_205__2,
            inputRegisters_205__1,inputRegisters_205__0})) ;
    Reg_16 loop1_205_x (.D ({inputRegisters_205__15,inputRegisters_205__14,
           inputRegisters_205__13,inputRegisters_205__12,inputRegisters_205__11,
           inputRegisters_205__10,inputRegisters_205__9,inputRegisters_205__8,
           inputRegisters_205__7,inputRegisters_205__6,inputRegisters_205__5,
           inputRegisters_205__4,inputRegisters_205__3,inputRegisters_205__2,
           inputRegisters_205__1,inputRegisters_205__0}), .en (
           enableRegister_205), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_205__15,registerOutputs_205__14,
           registerOutputs_205__13,registerOutputs_205__12,
           registerOutputs_205__11,registerOutputs_205__10,
           registerOutputs_205__9,registerOutputs_205__8,registerOutputs_205__7,
           registerOutputs_205__6,registerOutputs_205__5,registerOutputs_205__4,
           registerOutputs_205__3,registerOutputs_205__2,registerOutputs_205__1,
           registerOutputs_205__0})) ;
    Mux2_16 loop1_206_y (.A ({nx35943,nx36085,nx36227,nx36369,nx36511,nx36653,
            nx36795,nx36937,nx37079,nx37221,nx37363,nx37505,nx37647,nx37789,
            nx37931,nx38073}), .B ({nx33699,nx33837,nx33975,nx34113,nx34253,
            nx34391,nx34529,nx34669,nx34811,nx34953,nx35095,nx35237,nx35379,
            nx35521,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35663), .C ({inputRegisters_206__15,inputRegisters_206__14,
            inputRegisters_206__13,inputRegisters_206__12,inputRegisters_206__11
            ,inputRegisters_206__10,inputRegisters_206__9,inputRegisters_206__8,
            inputRegisters_206__7,inputRegisters_206__6,inputRegisters_206__5,
            inputRegisters_206__4,inputRegisters_206__3,inputRegisters_206__2,
            inputRegisters_206__1,inputRegisters_206__0})) ;
    Reg_16 loop1_206_x (.D ({inputRegisters_206__15,inputRegisters_206__14,
           inputRegisters_206__13,inputRegisters_206__12,inputRegisters_206__11,
           inputRegisters_206__10,inputRegisters_206__9,inputRegisters_206__8,
           inputRegisters_206__7,inputRegisters_206__6,inputRegisters_206__5,
           inputRegisters_206__4,inputRegisters_206__3,inputRegisters_206__2,
           inputRegisters_206__1,inputRegisters_206__0}), .en (
           enableRegister_206), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_206__15,registerOutputs_206__14,
           registerOutputs_206__13,registerOutputs_206__12,
           registerOutputs_206__11,registerOutputs_206__10,
           registerOutputs_206__9,registerOutputs_206__8,registerOutputs_206__7,
           registerOutputs_206__6,registerOutputs_206__5,registerOutputs_206__4,
           registerOutputs_206__3,registerOutputs_206__2,registerOutputs_206__1,
           registerOutputs_206__0})) ;
    Mux2_16 loop1_207_y (.A ({nx35943,nx36085,nx36227,nx36369,nx36511,nx36653,
            nx36795,nx36937,nx37079,nx37221,nx37363,nx37505,nx37647,nx37789,
            nx37931,nx38073}), .B ({nx33699,nx33837,nx33975,nx34115,nx34253,
            nx34391,nx34529,nx34669,nx34811,nx34953,nx35095,nx35237,nx35379,
            nx35521,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35663), .C ({inputRegisters_207__15,inputRegisters_207__14,
            inputRegisters_207__13,inputRegisters_207__12,inputRegisters_207__11
            ,inputRegisters_207__10,inputRegisters_207__9,inputRegisters_207__8,
            inputRegisters_207__7,inputRegisters_207__6,inputRegisters_207__5,
            inputRegisters_207__4,inputRegisters_207__3,inputRegisters_207__2,
            inputRegisters_207__1,inputRegisters_207__0})) ;
    Reg_16 loop1_207_x (.D ({inputRegisters_207__15,inputRegisters_207__14,
           inputRegisters_207__13,inputRegisters_207__12,inputRegisters_207__11,
           inputRegisters_207__10,inputRegisters_207__9,inputRegisters_207__8,
           inputRegisters_207__7,inputRegisters_207__6,inputRegisters_207__5,
           inputRegisters_207__4,inputRegisters_207__3,inputRegisters_207__2,
           inputRegisters_207__1,inputRegisters_207__0}), .en (
           enableRegister_207), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_207__15,registerOutputs_207__14,
           registerOutputs_207__13,registerOutputs_207__12,
           registerOutputs_207__11,registerOutputs_207__10,
           registerOutputs_207__9,registerOutputs_207__8,registerOutputs_207__7,
           registerOutputs_207__6,registerOutputs_207__5,registerOutputs_207__4,
           registerOutputs_207__3,registerOutputs_207__2,registerOutputs_207__1,
           registerOutputs_207__0})) ;
    Mux2_16 loop1_208_y (.A ({nx35943,nx36085,nx36227,nx36369,nx36511,nx36653,
            nx36795,nx36937,nx37079,nx37221,nx37363,nx37505,nx37647,nx37789,
            nx37931,nx38073}), .B ({nx33699,nx33837,nx33977,nx34115,nx34253,
            nx34391,nx34529,nx34669,nx34811,nx34953,nx35095,nx35237,nx35379,
            nx35521,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35663), .C ({inputRegisters_208__15,inputRegisters_208__14,
            inputRegisters_208__13,inputRegisters_208__12,inputRegisters_208__11
            ,inputRegisters_208__10,inputRegisters_208__9,inputRegisters_208__8,
            inputRegisters_208__7,inputRegisters_208__6,inputRegisters_208__5,
            inputRegisters_208__4,inputRegisters_208__3,inputRegisters_208__2,
            inputRegisters_208__1,inputRegisters_208__0})) ;
    Reg_16 loop1_208_x (.D ({inputRegisters_208__15,inputRegisters_208__14,
           inputRegisters_208__13,inputRegisters_208__12,inputRegisters_208__11,
           inputRegisters_208__10,inputRegisters_208__9,inputRegisters_208__8,
           inputRegisters_208__7,inputRegisters_208__6,inputRegisters_208__5,
           inputRegisters_208__4,inputRegisters_208__3,inputRegisters_208__2,
           inputRegisters_208__1,inputRegisters_208__0}), .en (
           enableRegister_208), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_208__15,registerOutputs_208__14,
           registerOutputs_208__13,registerOutputs_208__12,
           registerOutputs_208__11,registerOutputs_208__10,
           registerOutputs_208__9,registerOutputs_208__8,registerOutputs_208__7,
           registerOutputs_208__6,registerOutputs_208__5,registerOutputs_208__4,
           registerOutputs_208__3,registerOutputs_208__2,registerOutputs_208__1,
           registerOutputs_208__0})) ;
    Mux2_16 loop1_209_y (.A ({nx35943,nx36085,nx36227,nx36369,nx36511,nx36653,
            nx36795,nx36937,nx37079,nx37221,nx37363,nx37505,nx37647,nx37789,
            nx37931,nx38073}), .B ({nx33699,nx33839,nx33977,nx34115,nx34253,
            nx34391,nx34529,nx34669,nx34811,nx34953,nx35095,nx35237,nx35379,
            nx35521,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35663), .C ({inputRegisters_209__15,inputRegisters_209__14,
            inputRegisters_209__13,inputRegisters_209__12,inputRegisters_209__11
            ,inputRegisters_209__10,inputRegisters_209__9,inputRegisters_209__8,
            inputRegisters_209__7,inputRegisters_209__6,inputRegisters_209__5,
            inputRegisters_209__4,inputRegisters_209__3,inputRegisters_209__2,
            inputRegisters_209__1,inputRegisters_209__0})) ;
    Reg_16 loop1_209_x (.D ({inputRegisters_209__15,inputRegisters_209__14,
           inputRegisters_209__13,inputRegisters_209__12,inputRegisters_209__11,
           inputRegisters_209__10,inputRegisters_209__9,inputRegisters_209__8,
           inputRegisters_209__7,inputRegisters_209__6,inputRegisters_209__5,
           inputRegisters_209__4,inputRegisters_209__3,inputRegisters_209__2,
           inputRegisters_209__1,inputRegisters_209__0}), .en (
           enableRegister_209), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_209__15,registerOutputs_209__14,
           registerOutputs_209__13,registerOutputs_209__12,
           registerOutputs_209__11,registerOutputs_209__10,
           registerOutputs_209__9,registerOutputs_209__8,registerOutputs_209__7,
           registerOutputs_209__6,registerOutputs_209__5,registerOutputs_209__4,
           registerOutputs_209__3,registerOutputs_209__2,registerOutputs_209__1,
           registerOutputs_209__0})) ;
    Mux2_16 loop1_210_y (.A ({nx35945,nx36087,nx36229,nx36371,nx36513,nx36655,
            nx36797,nx36939,nx37081,nx37223,nx37365,nx37507,nx37649,nx37791,
            nx37933,nx38075}), .B ({nx33701,nx33839,nx33977,nx34115,nx34253,
            nx34391,nx34529,nx34671,nx34813,nx34955,nx35097,nx35239,nx35381,
            nx35523,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35665), .C ({inputRegisters_210__15,inputRegisters_210__14,
            inputRegisters_210__13,inputRegisters_210__12,inputRegisters_210__11
            ,inputRegisters_210__10,inputRegisters_210__9,inputRegisters_210__8,
            inputRegisters_210__7,inputRegisters_210__6,inputRegisters_210__5,
            inputRegisters_210__4,inputRegisters_210__3,inputRegisters_210__2,
            inputRegisters_210__1,inputRegisters_210__0})) ;
    Reg_16 loop1_210_x (.D ({inputRegisters_210__15,inputRegisters_210__14,
           inputRegisters_210__13,inputRegisters_210__12,inputRegisters_210__11,
           inputRegisters_210__10,inputRegisters_210__9,inputRegisters_210__8,
           inputRegisters_210__7,inputRegisters_210__6,inputRegisters_210__5,
           inputRegisters_210__4,inputRegisters_210__3,inputRegisters_210__2,
           inputRegisters_210__1,inputRegisters_210__0}), .en (
           enableRegister_210), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_210__15,registerOutputs_210__14,
           registerOutputs_210__13,registerOutputs_210__12,
           registerOutputs_210__11,registerOutputs_210__10,
           registerOutputs_210__9,registerOutputs_210__8,registerOutputs_210__7,
           registerOutputs_210__6,registerOutputs_210__5,registerOutputs_210__4,
           registerOutputs_210__3,registerOutputs_210__2,registerOutputs_210__1,
           registerOutputs_210__0})) ;
    Mux2_16 loop1_211_y (.A ({nx35945,nx36087,nx36229,nx36371,nx36513,nx36655,
            nx36797,nx36939,nx37081,nx37223,nx37365,nx37507,nx37649,nx37791,
            nx37933,nx38075}), .B ({nx33701,nx33839,nx33977,nx34115,nx34253,
            nx34391,nx34531,nx34671,nx34813,nx34955,nx35097,nx35239,nx35381,
            nx35523,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35665), .C ({inputRegisters_211__15,inputRegisters_211__14,
            inputRegisters_211__13,inputRegisters_211__12,inputRegisters_211__11
            ,inputRegisters_211__10,inputRegisters_211__9,inputRegisters_211__8,
            inputRegisters_211__7,inputRegisters_211__6,inputRegisters_211__5,
            inputRegisters_211__4,inputRegisters_211__3,inputRegisters_211__2,
            inputRegisters_211__1,inputRegisters_211__0})) ;
    Reg_16 loop1_211_x (.D ({inputRegisters_211__15,inputRegisters_211__14,
           inputRegisters_211__13,inputRegisters_211__12,inputRegisters_211__11,
           inputRegisters_211__10,inputRegisters_211__9,inputRegisters_211__8,
           inputRegisters_211__7,inputRegisters_211__6,inputRegisters_211__5,
           inputRegisters_211__4,inputRegisters_211__3,inputRegisters_211__2,
           inputRegisters_211__1,inputRegisters_211__0}), .en (
           enableRegister_211), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_211__15,registerOutputs_211__14,
           registerOutputs_211__13,registerOutputs_211__12,
           registerOutputs_211__11,registerOutputs_211__10,
           registerOutputs_211__9,registerOutputs_211__8,registerOutputs_211__7,
           registerOutputs_211__6,registerOutputs_211__5,registerOutputs_211__4,
           registerOutputs_211__3,registerOutputs_211__2,registerOutputs_211__1,
           registerOutputs_211__0})) ;
    Mux2_16 loop1_212_y (.A ({nx35945,nx36087,nx36229,nx36371,nx36513,nx36655,
            nx36797,nx36939,nx37081,nx37223,nx37365,nx37507,nx37649,nx37791,
            nx37933,nx38075}), .B ({nx33701,nx33839,nx33977,nx34115,nx34253,
            nx34393,nx34531,nx34671,nx34813,nx34955,nx35097,nx35239,nx35381,
            nx35523,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35665), .C ({inputRegisters_212__15,inputRegisters_212__14,
            inputRegisters_212__13,inputRegisters_212__12,inputRegisters_212__11
            ,inputRegisters_212__10,inputRegisters_212__9,inputRegisters_212__8,
            inputRegisters_212__7,inputRegisters_212__6,inputRegisters_212__5,
            inputRegisters_212__4,inputRegisters_212__3,inputRegisters_212__2,
            inputRegisters_212__1,inputRegisters_212__0})) ;
    Reg_16 loop1_212_x (.D ({inputRegisters_212__15,inputRegisters_212__14,
           inputRegisters_212__13,inputRegisters_212__12,inputRegisters_212__11,
           inputRegisters_212__10,inputRegisters_212__9,inputRegisters_212__8,
           inputRegisters_212__7,inputRegisters_212__6,inputRegisters_212__5,
           inputRegisters_212__4,inputRegisters_212__3,inputRegisters_212__2,
           inputRegisters_212__1,inputRegisters_212__0}), .en (
           enableRegister_212), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_212__15,registerOutputs_212__14,
           registerOutputs_212__13,registerOutputs_212__12,
           registerOutputs_212__11,registerOutputs_212__10,
           registerOutputs_212__9,registerOutputs_212__8,registerOutputs_212__7,
           registerOutputs_212__6,registerOutputs_212__5,registerOutputs_212__4,
           registerOutputs_212__3,registerOutputs_212__2,registerOutputs_212__1,
           registerOutputs_212__0})) ;
    Mux2_16 loop1_213_y (.A ({nx35945,nx36087,nx36229,nx36371,nx36513,nx36655,
            nx36797,nx36939,nx37081,nx37223,nx37365,nx37507,nx37649,nx37791,
            nx37933,nx38075}), .B ({nx33701,nx33839,nx33977,nx34115,nx34255,
            nx34393,nx34531,nx34671,nx34813,nx34955,nx35097,nx35239,nx35381,
            nx35523,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35665), .C ({inputRegisters_213__15,inputRegisters_213__14,
            inputRegisters_213__13,inputRegisters_213__12,inputRegisters_213__11
            ,inputRegisters_213__10,inputRegisters_213__9,inputRegisters_213__8,
            inputRegisters_213__7,inputRegisters_213__6,inputRegisters_213__5,
            inputRegisters_213__4,inputRegisters_213__3,inputRegisters_213__2,
            inputRegisters_213__1,inputRegisters_213__0})) ;
    Reg_16 loop1_213_x (.D ({inputRegisters_213__15,inputRegisters_213__14,
           inputRegisters_213__13,inputRegisters_213__12,inputRegisters_213__11,
           inputRegisters_213__10,inputRegisters_213__9,inputRegisters_213__8,
           inputRegisters_213__7,inputRegisters_213__6,inputRegisters_213__5,
           inputRegisters_213__4,inputRegisters_213__3,inputRegisters_213__2,
           inputRegisters_213__1,inputRegisters_213__0}), .en (
           enableRegister_213), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_213__15,registerOutputs_213__14,
           registerOutputs_213__13,registerOutputs_213__12,
           registerOutputs_213__11,registerOutputs_213__10,
           registerOutputs_213__9,registerOutputs_213__8,registerOutputs_213__7,
           registerOutputs_213__6,registerOutputs_213__5,registerOutputs_213__4,
           registerOutputs_213__3,registerOutputs_213__2,registerOutputs_213__1,
           registerOutputs_213__0})) ;
    Mux2_16 loop1_214_y (.A ({nx35945,nx36087,nx36229,nx36371,nx36513,nx36655,
            nx36797,nx36939,nx37081,nx37223,nx37365,nx37507,nx37649,nx37791,
            nx37933,nx38075}), .B ({nx33701,nx33839,nx33977,nx34117,nx34255,
            nx34393,nx34531,nx34671,nx34813,nx34955,nx35097,nx35239,nx35381,
            nx35523,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35665), .C ({inputRegisters_214__15,inputRegisters_214__14,
            inputRegisters_214__13,inputRegisters_214__12,inputRegisters_214__11
            ,inputRegisters_214__10,inputRegisters_214__9,inputRegisters_214__8,
            inputRegisters_214__7,inputRegisters_214__6,inputRegisters_214__5,
            inputRegisters_214__4,inputRegisters_214__3,inputRegisters_214__2,
            inputRegisters_214__1,inputRegisters_214__0})) ;
    Reg_16 loop1_214_x (.D ({inputRegisters_214__15,inputRegisters_214__14,
           inputRegisters_214__13,inputRegisters_214__12,inputRegisters_214__11,
           inputRegisters_214__10,inputRegisters_214__9,inputRegisters_214__8,
           inputRegisters_214__7,inputRegisters_214__6,inputRegisters_214__5,
           inputRegisters_214__4,inputRegisters_214__3,inputRegisters_214__2,
           inputRegisters_214__1,inputRegisters_214__0}), .en (
           enableRegister_214), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_214__15,registerOutputs_214__14,
           registerOutputs_214__13,registerOutputs_214__12,
           registerOutputs_214__11,registerOutputs_214__10,
           registerOutputs_214__9,registerOutputs_214__8,registerOutputs_214__7,
           registerOutputs_214__6,registerOutputs_214__5,registerOutputs_214__4,
           registerOutputs_214__3,registerOutputs_214__2,registerOutputs_214__1,
           registerOutputs_214__0})) ;
    Mux2_16 loop1_215_y (.A ({nx35945,nx36087,nx36229,nx36371,nx36513,nx36655,
            nx36797,nx36939,nx37081,nx37223,nx37365,nx37507,nx37649,nx37791,
            nx37933,nx38075}), .B ({nx33701,nx33839,nx33979,nx34117,nx34255,
            nx34393,nx34531,nx34671,nx34813,nx34955,nx35097,nx35239,nx35381,
            nx35523,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35665), .C ({inputRegisters_215__15,inputRegisters_215__14,
            inputRegisters_215__13,inputRegisters_215__12,inputRegisters_215__11
            ,inputRegisters_215__10,inputRegisters_215__9,inputRegisters_215__8,
            inputRegisters_215__7,inputRegisters_215__6,inputRegisters_215__5,
            inputRegisters_215__4,inputRegisters_215__3,inputRegisters_215__2,
            inputRegisters_215__1,inputRegisters_215__0})) ;
    Reg_16 loop1_215_x (.D ({inputRegisters_215__15,inputRegisters_215__14,
           inputRegisters_215__13,inputRegisters_215__12,inputRegisters_215__11,
           inputRegisters_215__10,inputRegisters_215__9,inputRegisters_215__8,
           inputRegisters_215__7,inputRegisters_215__6,inputRegisters_215__5,
           inputRegisters_215__4,inputRegisters_215__3,inputRegisters_215__2,
           inputRegisters_215__1,inputRegisters_215__0}), .en (
           enableRegister_215), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_215__15,registerOutputs_215__14,
           registerOutputs_215__13,registerOutputs_215__12,
           registerOutputs_215__11,registerOutputs_215__10,
           registerOutputs_215__9,registerOutputs_215__8,registerOutputs_215__7,
           registerOutputs_215__6,registerOutputs_215__5,registerOutputs_215__4,
           registerOutputs_215__3,registerOutputs_215__2,registerOutputs_215__1,
           registerOutputs_215__0})) ;
    Mux2_16 loop1_216_y (.A ({nx35945,nx36087,nx36229,nx36371,nx36513,nx36655,
            nx36797,nx36939,nx37081,nx37223,nx37365,nx37507,nx37649,nx37791,
            nx37933,nx38075}), .B ({nx33701,nx33841,nx33979,nx34117,nx34255,
            nx34393,nx34531,nx34671,nx34813,nx34955,nx35097,nx35239,nx35381,
            nx35523,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35665), .C ({inputRegisters_216__15,inputRegisters_216__14,
            inputRegisters_216__13,inputRegisters_216__12,inputRegisters_216__11
            ,inputRegisters_216__10,inputRegisters_216__9,inputRegisters_216__8,
            inputRegisters_216__7,inputRegisters_216__6,inputRegisters_216__5,
            inputRegisters_216__4,inputRegisters_216__3,inputRegisters_216__2,
            inputRegisters_216__1,inputRegisters_216__0})) ;
    Reg_16 loop1_216_x (.D ({inputRegisters_216__15,inputRegisters_216__14,
           inputRegisters_216__13,inputRegisters_216__12,inputRegisters_216__11,
           inputRegisters_216__10,inputRegisters_216__9,inputRegisters_216__8,
           inputRegisters_216__7,inputRegisters_216__6,inputRegisters_216__5,
           inputRegisters_216__4,inputRegisters_216__3,inputRegisters_216__2,
           inputRegisters_216__1,inputRegisters_216__0}), .en (
           enableRegister_216), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_216__15,registerOutputs_216__14,
           registerOutputs_216__13,registerOutputs_216__12,
           registerOutputs_216__11,registerOutputs_216__10,
           registerOutputs_216__9,registerOutputs_216__8,registerOutputs_216__7,
           registerOutputs_216__6,registerOutputs_216__5,registerOutputs_216__4,
           registerOutputs_216__3,registerOutputs_216__2,registerOutputs_216__1,
           registerOutputs_216__0})) ;
    Mux2_16 loop1_217_y (.A ({nx35947,nx36089,nx36231,nx36373,nx36515,nx36657,
            nx36799,nx36941,nx37083,nx37225,nx37367,nx37509,nx37651,nx37793,
            nx37935,nx38077}), .B ({nx33703,nx33841,nx33979,nx34117,nx34255,
            nx34393,nx34531,nx34673,nx34815,nx34957,nx35099,nx35241,nx35383,
            nx35525,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35667), .C ({inputRegisters_217__15,inputRegisters_217__14,
            inputRegisters_217__13,inputRegisters_217__12,inputRegisters_217__11
            ,inputRegisters_217__10,inputRegisters_217__9,inputRegisters_217__8,
            inputRegisters_217__7,inputRegisters_217__6,inputRegisters_217__5,
            inputRegisters_217__4,inputRegisters_217__3,inputRegisters_217__2,
            inputRegisters_217__1,inputRegisters_217__0})) ;
    Reg_16 loop1_217_x (.D ({inputRegisters_217__15,inputRegisters_217__14,
           inputRegisters_217__13,inputRegisters_217__12,inputRegisters_217__11,
           inputRegisters_217__10,inputRegisters_217__9,inputRegisters_217__8,
           inputRegisters_217__7,inputRegisters_217__6,inputRegisters_217__5,
           inputRegisters_217__4,inputRegisters_217__3,inputRegisters_217__2,
           inputRegisters_217__1,inputRegisters_217__0}), .en (
           enableRegister_217), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_217__15,registerOutputs_217__14,
           registerOutputs_217__13,registerOutputs_217__12,
           registerOutputs_217__11,registerOutputs_217__10,
           registerOutputs_217__9,registerOutputs_217__8,registerOutputs_217__7,
           registerOutputs_217__6,registerOutputs_217__5,registerOutputs_217__4,
           registerOutputs_217__3,registerOutputs_217__2,registerOutputs_217__1,
           registerOutputs_217__0})) ;
    Mux2_16 loop1_218_y (.A ({nx35947,nx36089,nx36231,nx36373,nx36515,nx36657,
            nx36799,nx36941,nx37083,nx37225,nx37367,nx37509,nx37651,nx37793,
            nx37935,nx38077}), .B ({nx33703,nx33841,nx33979,nx34117,nx34255,
            nx34393,nx34533,nx34673,nx34815,nx34957,nx35099,nx35241,nx35383,
            nx35525,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35667), .C ({inputRegisters_218__15,inputRegisters_218__14,
            inputRegisters_218__13,inputRegisters_218__12,inputRegisters_218__11
            ,inputRegisters_218__10,inputRegisters_218__9,inputRegisters_218__8,
            inputRegisters_218__7,inputRegisters_218__6,inputRegisters_218__5,
            inputRegisters_218__4,inputRegisters_218__3,inputRegisters_218__2,
            inputRegisters_218__1,inputRegisters_218__0})) ;
    Reg_16 loop1_218_x (.D ({inputRegisters_218__15,inputRegisters_218__14,
           inputRegisters_218__13,inputRegisters_218__12,inputRegisters_218__11,
           inputRegisters_218__10,inputRegisters_218__9,inputRegisters_218__8,
           inputRegisters_218__7,inputRegisters_218__6,inputRegisters_218__5,
           inputRegisters_218__4,inputRegisters_218__3,inputRegisters_218__2,
           inputRegisters_218__1,inputRegisters_218__0}), .en (
           enableRegister_218), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_218__15,registerOutputs_218__14,
           registerOutputs_218__13,registerOutputs_218__12,
           registerOutputs_218__11,registerOutputs_218__10,
           registerOutputs_218__9,registerOutputs_218__8,registerOutputs_218__7,
           registerOutputs_218__6,registerOutputs_218__5,registerOutputs_218__4,
           registerOutputs_218__3,registerOutputs_218__2,registerOutputs_218__1,
           registerOutputs_218__0})) ;
    Mux2_16 loop1_219_y (.A ({nx35947,nx36089,nx36231,nx36373,nx36515,nx36657,
            nx36799,nx36941,nx37083,nx37225,nx37367,nx37509,nx37651,nx37793,
            nx37935,nx38077}), .B ({nx33703,nx33841,nx33979,nx34117,nx34255,
            nx34395,nx34533,nx34673,nx34815,nx34957,nx35099,nx35241,nx35383,
            nx35525,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35667), .C ({inputRegisters_219__15,inputRegisters_219__14,
            inputRegisters_219__13,inputRegisters_219__12,inputRegisters_219__11
            ,inputRegisters_219__10,inputRegisters_219__9,inputRegisters_219__8,
            inputRegisters_219__7,inputRegisters_219__6,inputRegisters_219__5,
            inputRegisters_219__4,inputRegisters_219__3,inputRegisters_219__2,
            inputRegisters_219__1,inputRegisters_219__0})) ;
    Reg_16 loop1_219_x (.D ({inputRegisters_219__15,inputRegisters_219__14,
           inputRegisters_219__13,inputRegisters_219__12,inputRegisters_219__11,
           inputRegisters_219__10,inputRegisters_219__9,inputRegisters_219__8,
           inputRegisters_219__7,inputRegisters_219__6,inputRegisters_219__5,
           inputRegisters_219__4,inputRegisters_219__3,inputRegisters_219__2,
           inputRegisters_219__1,inputRegisters_219__0}), .en (
           enableRegister_219), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_219__15,registerOutputs_219__14,
           registerOutputs_219__13,registerOutputs_219__12,
           registerOutputs_219__11,registerOutputs_219__10,
           registerOutputs_219__9,registerOutputs_219__8,registerOutputs_219__7,
           registerOutputs_219__6,registerOutputs_219__5,registerOutputs_219__4,
           registerOutputs_219__3,registerOutputs_219__2,registerOutputs_219__1,
           registerOutputs_219__0})) ;
    Mux2_16 loop1_220_y (.A ({nx35947,nx36089,nx36231,nx36373,nx36515,nx36657,
            nx36799,nx36941,nx37083,nx37225,nx37367,nx37509,nx37651,nx37793,
            nx37935,nx38077}), .B ({nx33703,nx33841,nx33979,nx34117,nx34257,
            nx34395,nx34533,nx34673,nx34815,nx34957,nx35099,nx35241,nx35383,
            nx35525,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35667), .C ({inputRegisters_220__15,inputRegisters_220__14,
            inputRegisters_220__13,inputRegisters_220__12,inputRegisters_220__11
            ,inputRegisters_220__10,inputRegisters_220__9,inputRegisters_220__8,
            inputRegisters_220__7,inputRegisters_220__6,inputRegisters_220__5,
            inputRegisters_220__4,inputRegisters_220__3,inputRegisters_220__2,
            inputRegisters_220__1,inputRegisters_220__0})) ;
    Reg_16 loop1_220_x (.D ({inputRegisters_220__15,inputRegisters_220__14,
           inputRegisters_220__13,inputRegisters_220__12,inputRegisters_220__11,
           inputRegisters_220__10,inputRegisters_220__9,inputRegisters_220__8,
           inputRegisters_220__7,inputRegisters_220__6,inputRegisters_220__5,
           inputRegisters_220__4,inputRegisters_220__3,inputRegisters_220__2,
           inputRegisters_220__1,inputRegisters_220__0}), .en (
           enableRegister_220), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_220__15,registerOutputs_220__14,
           registerOutputs_220__13,registerOutputs_220__12,
           registerOutputs_220__11,registerOutputs_220__10,
           registerOutputs_220__9,registerOutputs_220__8,registerOutputs_220__7,
           registerOutputs_220__6,registerOutputs_220__5,registerOutputs_220__4,
           registerOutputs_220__3,registerOutputs_220__2,registerOutputs_220__1,
           registerOutputs_220__0})) ;
    Mux2_16 loop1_221_y (.A ({nx35947,nx36089,nx36231,nx36373,nx36515,nx36657,
            nx36799,nx36941,nx37083,nx37225,nx37367,nx37509,nx37651,nx37793,
            nx37935,nx38077}), .B ({nx33703,nx33841,nx33979,nx34119,nx34257,
            nx34395,nx34533,nx34673,nx34815,nx34957,nx35099,nx35241,nx35383,
            nx35525,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35667), .C ({inputRegisters_221__15,inputRegisters_221__14,
            inputRegisters_221__13,inputRegisters_221__12,inputRegisters_221__11
            ,inputRegisters_221__10,inputRegisters_221__9,inputRegisters_221__8,
            inputRegisters_221__7,inputRegisters_221__6,inputRegisters_221__5,
            inputRegisters_221__4,inputRegisters_221__3,inputRegisters_221__2,
            inputRegisters_221__1,inputRegisters_221__0})) ;
    Reg_16 loop1_221_x (.D ({inputRegisters_221__15,inputRegisters_221__14,
           inputRegisters_221__13,inputRegisters_221__12,inputRegisters_221__11,
           inputRegisters_221__10,inputRegisters_221__9,inputRegisters_221__8,
           inputRegisters_221__7,inputRegisters_221__6,inputRegisters_221__5,
           inputRegisters_221__4,inputRegisters_221__3,inputRegisters_221__2,
           inputRegisters_221__1,inputRegisters_221__0}), .en (
           enableRegister_221), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_221__15,registerOutputs_221__14,
           registerOutputs_221__13,registerOutputs_221__12,
           registerOutputs_221__11,registerOutputs_221__10,
           registerOutputs_221__9,registerOutputs_221__8,registerOutputs_221__7,
           registerOutputs_221__6,registerOutputs_221__5,registerOutputs_221__4,
           registerOutputs_221__3,registerOutputs_221__2,registerOutputs_221__1,
           registerOutputs_221__0})) ;
    Mux2_16 loop1_222_y (.A ({nx35947,nx36089,nx36231,nx36373,nx36515,nx36657,
            nx36799,nx36941,nx37083,nx37225,nx37367,nx37509,nx37651,nx37793,
            nx37935,nx38077}), .B ({nx33703,nx33841,nx33981,nx34119,nx34257,
            nx34395,nx34533,nx34673,nx34815,nx34957,nx35099,nx35241,nx35383,
            nx35525,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35667), .C ({inputRegisters_222__15,inputRegisters_222__14,
            inputRegisters_222__13,inputRegisters_222__12,inputRegisters_222__11
            ,inputRegisters_222__10,inputRegisters_222__9,inputRegisters_222__8,
            inputRegisters_222__7,inputRegisters_222__6,inputRegisters_222__5,
            inputRegisters_222__4,inputRegisters_222__3,inputRegisters_222__2,
            inputRegisters_222__1,inputRegisters_222__0})) ;
    Reg_16 loop1_222_x (.D ({inputRegisters_222__15,inputRegisters_222__14,
           inputRegisters_222__13,inputRegisters_222__12,inputRegisters_222__11,
           inputRegisters_222__10,inputRegisters_222__9,inputRegisters_222__8,
           inputRegisters_222__7,inputRegisters_222__6,inputRegisters_222__5,
           inputRegisters_222__4,inputRegisters_222__3,inputRegisters_222__2,
           inputRegisters_222__1,inputRegisters_222__0}), .en (
           enableRegister_222), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_222__15,registerOutputs_222__14,
           registerOutputs_222__13,registerOutputs_222__12,
           registerOutputs_222__11,registerOutputs_222__10,
           registerOutputs_222__9,registerOutputs_222__8,registerOutputs_222__7,
           registerOutputs_222__6,registerOutputs_222__5,registerOutputs_222__4,
           registerOutputs_222__3,registerOutputs_222__2,registerOutputs_222__1,
           registerOutputs_222__0})) ;
    Mux2_16 loop1_223_y (.A ({nx35947,nx36089,nx36231,nx36373,nx36515,nx36657,
            nx36799,nx36941,nx37083,nx37225,nx37367,nx37509,nx37651,nx37793,
            nx37935,nx38077}), .B ({nx33703,nx33843,nx33981,nx34119,nx34257,
            nx34395,nx34533,nx34673,nx34815,nx34957,nx35099,nx35241,nx35383,
            nx35525,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35667), .C ({inputRegisters_223__15,inputRegisters_223__14,
            inputRegisters_223__13,inputRegisters_223__12,inputRegisters_223__11
            ,inputRegisters_223__10,inputRegisters_223__9,inputRegisters_223__8,
            inputRegisters_223__7,inputRegisters_223__6,inputRegisters_223__5,
            inputRegisters_223__4,inputRegisters_223__3,inputRegisters_223__2,
            inputRegisters_223__1,inputRegisters_223__0})) ;
    Reg_16 loop1_223_x (.D ({inputRegisters_223__15,inputRegisters_223__14,
           inputRegisters_223__13,inputRegisters_223__12,inputRegisters_223__11,
           inputRegisters_223__10,inputRegisters_223__9,inputRegisters_223__8,
           inputRegisters_223__7,inputRegisters_223__6,inputRegisters_223__5,
           inputRegisters_223__4,inputRegisters_223__3,inputRegisters_223__2,
           inputRegisters_223__1,inputRegisters_223__0}), .en (
           enableRegister_223), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_223__15,registerOutputs_223__14,
           registerOutputs_223__13,registerOutputs_223__12,
           registerOutputs_223__11,registerOutputs_223__10,
           registerOutputs_223__9,registerOutputs_223__8,registerOutputs_223__7,
           registerOutputs_223__6,registerOutputs_223__5,registerOutputs_223__4,
           registerOutputs_223__3,registerOutputs_223__2,registerOutputs_223__1,
           registerOutputs_223__0})) ;
    Mux2_16 loop1_224_y (.A ({nx35949,nx36091,nx36233,nx36375,nx36517,nx36659,
            nx36801,nx36943,nx37085,nx37227,nx37369,nx37511,nx37653,nx37795,
            nx37937,nx38079}), .B ({nx33705,nx33843,nx33981,nx34119,nx34257,
            nx34395,nx34533,nx34675,nx34817,nx34959,nx35101,nx35243,nx35385,
            nx35527,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35669), .C ({inputRegisters_224__15,inputRegisters_224__14,
            inputRegisters_224__13,inputRegisters_224__12,inputRegisters_224__11
            ,inputRegisters_224__10,inputRegisters_224__9,inputRegisters_224__8,
            inputRegisters_224__7,inputRegisters_224__6,inputRegisters_224__5,
            inputRegisters_224__4,inputRegisters_224__3,inputRegisters_224__2,
            inputRegisters_224__1,inputRegisters_224__0})) ;
    Reg_16 loop1_224_x (.D ({inputRegisters_224__15,inputRegisters_224__14,
           inputRegisters_224__13,inputRegisters_224__12,inputRegisters_224__11,
           inputRegisters_224__10,inputRegisters_224__9,inputRegisters_224__8,
           inputRegisters_224__7,inputRegisters_224__6,inputRegisters_224__5,
           inputRegisters_224__4,inputRegisters_224__3,inputRegisters_224__2,
           inputRegisters_224__1,inputRegisters_224__0}), .en (
           enableRegister_224), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_224__15,registerOutputs_224__14,
           registerOutputs_224__13,registerOutputs_224__12,
           registerOutputs_224__11,registerOutputs_224__10,
           registerOutputs_224__9,registerOutputs_224__8,registerOutputs_224__7,
           registerOutputs_224__6,registerOutputs_224__5,registerOutputs_224__4,
           registerOutputs_224__3,registerOutputs_224__2,registerOutputs_224__1,
           registerOutputs_224__0})) ;
    Mux2_16 loop1_225_y (.A ({nx35949,nx36091,nx36233,nx36375,nx36517,nx36659,
            nx36801,nx36943,nx37085,nx37227,nx37369,nx37511,nx37653,nx37795,
            nx37937,nx38079}), .B ({nx33705,nx33843,nx33981,nx34119,nx34257,
            nx34395,nx34535,nx34675,nx34817,nx34959,nx35101,nx35243,nx35385,
            nx35527,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35669), .C ({inputRegisters_225__15,inputRegisters_225__14,
            inputRegisters_225__13,inputRegisters_225__12,inputRegisters_225__11
            ,inputRegisters_225__10,inputRegisters_225__9,inputRegisters_225__8,
            inputRegisters_225__7,inputRegisters_225__6,inputRegisters_225__5,
            inputRegisters_225__4,inputRegisters_225__3,inputRegisters_225__2,
            inputRegisters_225__1,inputRegisters_225__0})) ;
    Reg_16 loop1_225_x (.D ({inputRegisters_225__15,inputRegisters_225__14,
           inputRegisters_225__13,inputRegisters_225__12,inputRegisters_225__11,
           inputRegisters_225__10,inputRegisters_225__9,inputRegisters_225__8,
           inputRegisters_225__7,inputRegisters_225__6,inputRegisters_225__5,
           inputRegisters_225__4,inputRegisters_225__3,inputRegisters_225__2,
           inputRegisters_225__1,inputRegisters_225__0}), .en (
           enableRegister_225), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_225__15,registerOutputs_225__14,
           registerOutputs_225__13,registerOutputs_225__12,
           registerOutputs_225__11,registerOutputs_225__10,
           registerOutputs_225__9,registerOutputs_225__8,registerOutputs_225__7,
           registerOutputs_225__6,registerOutputs_225__5,registerOutputs_225__4,
           registerOutputs_225__3,registerOutputs_225__2,registerOutputs_225__1,
           registerOutputs_225__0})) ;
    Mux2_16 loop1_226_y (.A ({nx35949,nx36091,nx36233,nx36375,nx36517,nx36659,
            nx36801,nx36943,nx37085,nx37227,nx37369,nx37511,nx37653,nx37795,
            nx37937,nx38079}), .B ({nx33705,nx33843,nx33981,nx34119,nx34257,
            nx34397,nx34535,nx34675,nx34817,nx34959,nx35101,nx35243,nx35385,
            nx35527,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35669), .C ({inputRegisters_226__15,inputRegisters_226__14,
            inputRegisters_226__13,inputRegisters_226__12,inputRegisters_226__11
            ,inputRegisters_226__10,inputRegisters_226__9,inputRegisters_226__8,
            inputRegisters_226__7,inputRegisters_226__6,inputRegisters_226__5,
            inputRegisters_226__4,inputRegisters_226__3,inputRegisters_226__2,
            inputRegisters_226__1,inputRegisters_226__0})) ;
    Reg_16 loop1_226_x (.D ({inputRegisters_226__15,inputRegisters_226__14,
           inputRegisters_226__13,inputRegisters_226__12,inputRegisters_226__11,
           inputRegisters_226__10,inputRegisters_226__9,inputRegisters_226__8,
           inputRegisters_226__7,inputRegisters_226__6,inputRegisters_226__5,
           inputRegisters_226__4,inputRegisters_226__3,inputRegisters_226__2,
           inputRegisters_226__1,inputRegisters_226__0}), .en (
           enableRegister_226), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_226__15,registerOutputs_226__14,
           registerOutputs_226__13,registerOutputs_226__12,
           registerOutputs_226__11,registerOutputs_226__10,
           registerOutputs_226__9,registerOutputs_226__8,registerOutputs_226__7,
           registerOutputs_226__6,registerOutputs_226__5,registerOutputs_226__4,
           registerOutputs_226__3,registerOutputs_226__2,registerOutputs_226__1,
           registerOutputs_226__0})) ;
    Mux2_16 loop1_227_y (.A ({nx35949,nx36091,nx36233,nx36375,nx36517,nx36659,
            nx36801,nx36943,nx37085,nx37227,nx37369,nx37511,nx37653,nx37795,
            nx37937,nx38079}), .B ({nx33705,nx33843,nx33981,nx34119,nx34259,
            nx34397,nx34535,nx34675,nx34817,nx34959,nx35101,nx35243,nx35385,
            nx35527,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35669), .C ({inputRegisters_227__15,inputRegisters_227__14,
            inputRegisters_227__13,inputRegisters_227__12,inputRegisters_227__11
            ,inputRegisters_227__10,inputRegisters_227__9,inputRegisters_227__8,
            inputRegisters_227__7,inputRegisters_227__6,inputRegisters_227__5,
            inputRegisters_227__4,inputRegisters_227__3,inputRegisters_227__2,
            inputRegisters_227__1,inputRegisters_227__0})) ;
    Reg_16 loop1_227_x (.D ({inputRegisters_227__15,inputRegisters_227__14,
           inputRegisters_227__13,inputRegisters_227__12,inputRegisters_227__11,
           inputRegisters_227__10,inputRegisters_227__9,inputRegisters_227__8,
           inputRegisters_227__7,inputRegisters_227__6,inputRegisters_227__5,
           inputRegisters_227__4,inputRegisters_227__3,inputRegisters_227__2,
           inputRegisters_227__1,inputRegisters_227__0}), .en (
           enableRegister_227), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_227__15,registerOutputs_227__14,
           registerOutputs_227__13,registerOutputs_227__12,
           registerOutputs_227__11,registerOutputs_227__10,
           registerOutputs_227__9,registerOutputs_227__8,registerOutputs_227__7,
           registerOutputs_227__6,registerOutputs_227__5,registerOutputs_227__4,
           registerOutputs_227__3,registerOutputs_227__2,registerOutputs_227__1,
           registerOutputs_227__0})) ;
    Mux2_16 loop1_228_y (.A ({nx35949,nx36091,nx36233,nx36375,nx36517,nx36659,
            nx36801,nx36943,nx37085,nx37227,nx37369,nx37511,nx37653,nx37795,
            nx37937,nx38079}), .B ({nx33705,nx33843,nx33981,nx34121,nx34259,
            nx34397,nx34535,nx34675,nx34817,nx34959,nx35101,nx35243,nx35385,
            nx35527,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35669), .C ({inputRegisters_228__15,inputRegisters_228__14,
            inputRegisters_228__13,inputRegisters_228__12,inputRegisters_228__11
            ,inputRegisters_228__10,inputRegisters_228__9,inputRegisters_228__8,
            inputRegisters_228__7,inputRegisters_228__6,inputRegisters_228__5,
            inputRegisters_228__4,inputRegisters_228__3,inputRegisters_228__2,
            inputRegisters_228__1,inputRegisters_228__0})) ;
    Reg_16 loop1_228_x (.D ({inputRegisters_228__15,inputRegisters_228__14,
           inputRegisters_228__13,inputRegisters_228__12,inputRegisters_228__11,
           inputRegisters_228__10,inputRegisters_228__9,inputRegisters_228__8,
           inputRegisters_228__7,inputRegisters_228__6,inputRegisters_228__5,
           inputRegisters_228__4,inputRegisters_228__3,inputRegisters_228__2,
           inputRegisters_228__1,inputRegisters_228__0}), .en (
           enableRegister_228), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_228__15,registerOutputs_228__14,
           registerOutputs_228__13,registerOutputs_228__12,
           registerOutputs_228__11,registerOutputs_228__10,
           registerOutputs_228__9,registerOutputs_228__8,registerOutputs_228__7,
           registerOutputs_228__6,registerOutputs_228__5,registerOutputs_228__4,
           registerOutputs_228__3,registerOutputs_228__2,registerOutputs_228__1,
           registerOutputs_228__0})) ;
    Mux2_16 loop1_229_y (.A ({nx35949,nx36091,nx36233,nx36375,nx36517,nx36659,
            nx36801,nx36943,nx37085,nx37227,nx37369,nx37511,nx37653,nx37795,
            nx37937,nx38079}), .B ({nx33705,nx33843,nx33983,nx34121,nx34259,
            nx34397,nx34535,nx34675,nx34817,nx34959,nx35101,nx35243,nx35385,
            nx35527,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35669), .C ({inputRegisters_229__15,inputRegisters_229__14,
            inputRegisters_229__13,inputRegisters_229__12,inputRegisters_229__11
            ,inputRegisters_229__10,inputRegisters_229__9,inputRegisters_229__8,
            inputRegisters_229__7,inputRegisters_229__6,inputRegisters_229__5,
            inputRegisters_229__4,inputRegisters_229__3,inputRegisters_229__2,
            inputRegisters_229__1,inputRegisters_229__0})) ;
    Reg_16 loop1_229_x (.D ({inputRegisters_229__15,inputRegisters_229__14,
           inputRegisters_229__13,inputRegisters_229__12,inputRegisters_229__11,
           inputRegisters_229__10,inputRegisters_229__9,inputRegisters_229__8,
           inputRegisters_229__7,inputRegisters_229__6,inputRegisters_229__5,
           inputRegisters_229__4,inputRegisters_229__3,inputRegisters_229__2,
           inputRegisters_229__1,inputRegisters_229__0}), .en (
           enableRegister_229), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_229__15,registerOutputs_229__14,
           registerOutputs_229__13,registerOutputs_229__12,
           registerOutputs_229__11,registerOutputs_229__10,
           registerOutputs_229__9,registerOutputs_229__8,registerOutputs_229__7,
           registerOutputs_229__6,registerOutputs_229__5,registerOutputs_229__4,
           registerOutputs_229__3,registerOutputs_229__2,registerOutputs_229__1,
           registerOutputs_229__0})) ;
    Mux2_16 loop1_230_y (.A ({nx35949,nx36091,nx36233,nx36375,nx36517,nx36659,
            nx36801,nx36943,nx37085,nx37227,nx37369,nx37511,nx37653,nx37795,
            nx37937,nx38079}), .B ({nx33705,nx33845,nx33983,nx34121,nx34259,
            nx34397,nx34535,nx34675,nx34817,nx34959,nx35101,nx35243,nx35385,
            nx35527,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35669), .C ({inputRegisters_230__15,inputRegisters_230__14,
            inputRegisters_230__13,inputRegisters_230__12,inputRegisters_230__11
            ,inputRegisters_230__10,inputRegisters_230__9,inputRegisters_230__8,
            inputRegisters_230__7,inputRegisters_230__6,inputRegisters_230__5,
            inputRegisters_230__4,inputRegisters_230__3,inputRegisters_230__2,
            inputRegisters_230__1,inputRegisters_230__0})) ;
    Reg_16 loop1_230_x (.D ({inputRegisters_230__15,inputRegisters_230__14,
           inputRegisters_230__13,inputRegisters_230__12,inputRegisters_230__11,
           inputRegisters_230__10,inputRegisters_230__9,inputRegisters_230__8,
           inputRegisters_230__7,inputRegisters_230__6,inputRegisters_230__5,
           inputRegisters_230__4,inputRegisters_230__3,inputRegisters_230__2,
           inputRegisters_230__1,inputRegisters_230__0}), .en (
           enableRegister_230), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_230__15,registerOutputs_230__14,
           registerOutputs_230__13,registerOutputs_230__12,
           registerOutputs_230__11,registerOutputs_230__10,
           registerOutputs_230__9,registerOutputs_230__8,registerOutputs_230__7,
           registerOutputs_230__6,registerOutputs_230__5,registerOutputs_230__4,
           registerOutputs_230__3,registerOutputs_230__2,registerOutputs_230__1,
           registerOutputs_230__0})) ;
    Mux2_16 loop1_231_y (.A ({nx35951,nx36093,nx36235,nx36377,nx36519,nx36661,
            nx36803,nx36945,nx37087,nx37229,nx37371,nx37513,nx37655,nx37797,
            nx37939,nx38081}), .B ({nx33707,nx33845,nx33983,nx34121,nx34259,
            nx34397,nx34535,nx34677,nx34819,nx34961,nx35103,nx35245,nx35387,
            nx35529,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35671), .C ({inputRegisters_231__15,inputRegisters_231__14,
            inputRegisters_231__13,inputRegisters_231__12,inputRegisters_231__11
            ,inputRegisters_231__10,inputRegisters_231__9,inputRegisters_231__8,
            inputRegisters_231__7,inputRegisters_231__6,inputRegisters_231__5,
            inputRegisters_231__4,inputRegisters_231__3,inputRegisters_231__2,
            inputRegisters_231__1,inputRegisters_231__0})) ;
    Reg_16 loop1_231_x (.D ({inputRegisters_231__15,inputRegisters_231__14,
           inputRegisters_231__13,inputRegisters_231__12,inputRegisters_231__11,
           inputRegisters_231__10,inputRegisters_231__9,inputRegisters_231__8,
           inputRegisters_231__7,inputRegisters_231__6,inputRegisters_231__5,
           inputRegisters_231__4,inputRegisters_231__3,inputRegisters_231__2,
           inputRegisters_231__1,inputRegisters_231__0}), .en (
           enableRegister_231), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_231__15,registerOutputs_231__14,
           registerOutputs_231__13,registerOutputs_231__12,
           registerOutputs_231__11,registerOutputs_231__10,
           registerOutputs_231__9,registerOutputs_231__8,registerOutputs_231__7,
           registerOutputs_231__6,registerOutputs_231__5,registerOutputs_231__4,
           registerOutputs_231__3,registerOutputs_231__2,registerOutputs_231__1,
           registerOutputs_231__0})) ;
    Mux2_16 loop1_232_y (.A ({nx35951,nx36093,nx36235,nx36377,nx36519,nx36661,
            nx36803,nx36945,nx37087,nx37229,nx37371,nx37513,nx37655,nx37797,
            nx37939,nx38081}), .B ({nx33707,nx33845,nx33983,nx34121,nx34259,
            nx34397,nx34537,nx34677,nx34819,nx34961,nx35103,nx35245,nx35387,
            nx35529,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35671), .C ({inputRegisters_232__15,inputRegisters_232__14,
            inputRegisters_232__13,inputRegisters_232__12,inputRegisters_232__11
            ,inputRegisters_232__10,inputRegisters_232__9,inputRegisters_232__8,
            inputRegisters_232__7,inputRegisters_232__6,inputRegisters_232__5,
            inputRegisters_232__4,inputRegisters_232__3,inputRegisters_232__2,
            inputRegisters_232__1,inputRegisters_232__0})) ;
    Reg_16 loop1_232_x (.D ({inputRegisters_232__15,inputRegisters_232__14,
           inputRegisters_232__13,inputRegisters_232__12,inputRegisters_232__11,
           inputRegisters_232__10,inputRegisters_232__9,inputRegisters_232__8,
           inputRegisters_232__7,inputRegisters_232__6,inputRegisters_232__5,
           inputRegisters_232__4,inputRegisters_232__3,inputRegisters_232__2,
           inputRegisters_232__1,inputRegisters_232__0}), .en (
           enableRegister_232), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_232__15,registerOutputs_232__14,
           registerOutputs_232__13,registerOutputs_232__12,
           registerOutputs_232__11,registerOutputs_232__10,
           registerOutputs_232__9,registerOutputs_232__8,registerOutputs_232__7,
           registerOutputs_232__6,registerOutputs_232__5,registerOutputs_232__4,
           registerOutputs_232__3,registerOutputs_232__2,registerOutputs_232__1,
           registerOutputs_232__0})) ;
    Mux2_16 loop1_233_y (.A ({nx35951,nx36093,nx36235,nx36377,nx36519,nx36661,
            nx36803,nx36945,nx37087,nx37229,nx37371,nx37513,nx37655,nx37797,
            nx37939,nx38081}), .B ({nx33707,nx33845,nx33983,nx34121,nx34259,
            nx34399,nx34537,nx34677,nx34819,nx34961,nx35103,nx35245,nx35387,
            nx35529,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35671), .C ({inputRegisters_233__15,inputRegisters_233__14,
            inputRegisters_233__13,inputRegisters_233__12,inputRegisters_233__11
            ,inputRegisters_233__10,inputRegisters_233__9,inputRegisters_233__8,
            inputRegisters_233__7,inputRegisters_233__6,inputRegisters_233__5,
            inputRegisters_233__4,inputRegisters_233__3,inputRegisters_233__2,
            inputRegisters_233__1,inputRegisters_233__0})) ;
    Reg_16 loop1_233_x (.D ({inputRegisters_233__15,inputRegisters_233__14,
           inputRegisters_233__13,inputRegisters_233__12,inputRegisters_233__11,
           inputRegisters_233__10,inputRegisters_233__9,inputRegisters_233__8,
           inputRegisters_233__7,inputRegisters_233__6,inputRegisters_233__5,
           inputRegisters_233__4,inputRegisters_233__3,inputRegisters_233__2,
           inputRegisters_233__1,inputRegisters_233__0}), .en (
           enableRegister_233), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_233__15,registerOutputs_233__14,
           registerOutputs_233__13,registerOutputs_233__12,
           registerOutputs_233__11,registerOutputs_233__10,
           registerOutputs_233__9,registerOutputs_233__8,registerOutputs_233__7,
           registerOutputs_233__6,registerOutputs_233__5,registerOutputs_233__4,
           registerOutputs_233__3,registerOutputs_233__2,registerOutputs_233__1,
           registerOutputs_233__0})) ;
    Mux2_16 loop1_234_y (.A ({nx35951,nx36093,nx36235,nx36377,nx36519,nx36661,
            nx36803,nx36945,nx37087,nx37229,nx37371,nx37513,nx37655,nx37797,
            nx37939,nx38081}), .B ({nx33707,nx33845,nx33983,nx34121,nx34261,
            nx34399,nx34537,nx34677,nx34819,nx34961,nx35103,nx35245,nx35387,
            nx35529,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35671), .C ({inputRegisters_234__15,inputRegisters_234__14,
            inputRegisters_234__13,inputRegisters_234__12,inputRegisters_234__11
            ,inputRegisters_234__10,inputRegisters_234__9,inputRegisters_234__8,
            inputRegisters_234__7,inputRegisters_234__6,inputRegisters_234__5,
            inputRegisters_234__4,inputRegisters_234__3,inputRegisters_234__2,
            inputRegisters_234__1,inputRegisters_234__0})) ;
    Reg_16 loop1_234_x (.D ({inputRegisters_234__15,inputRegisters_234__14,
           inputRegisters_234__13,inputRegisters_234__12,inputRegisters_234__11,
           inputRegisters_234__10,inputRegisters_234__9,inputRegisters_234__8,
           inputRegisters_234__7,inputRegisters_234__6,inputRegisters_234__5,
           inputRegisters_234__4,inputRegisters_234__3,inputRegisters_234__2,
           inputRegisters_234__1,inputRegisters_234__0}), .en (
           enableRegister_234), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_234__15,registerOutputs_234__14,
           registerOutputs_234__13,registerOutputs_234__12,
           registerOutputs_234__11,registerOutputs_234__10,
           registerOutputs_234__9,registerOutputs_234__8,registerOutputs_234__7,
           registerOutputs_234__6,registerOutputs_234__5,registerOutputs_234__4,
           registerOutputs_234__3,registerOutputs_234__2,registerOutputs_234__1,
           registerOutputs_234__0})) ;
    Mux2_16 loop1_235_y (.A ({nx35951,nx36093,nx36235,nx36377,nx36519,nx36661,
            nx36803,nx36945,nx37087,nx37229,nx37371,nx37513,nx37655,nx37797,
            nx37939,nx38081}), .B ({nx33707,nx33845,nx33983,nx34123,nx34261,
            nx34399,nx34537,nx34677,nx34819,nx34961,nx35103,nx35245,nx35387,
            nx35529,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35671), .C ({inputRegisters_235__15,inputRegisters_235__14,
            inputRegisters_235__13,inputRegisters_235__12,inputRegisters_235__11
            ,inputRegisters_235__10,inputRegisters_235__9,inputRegisters_235__8,
            inputRegisters_235__7,inputRegisters_235__6,inputRegisters_235__5,
            inputRegisters_235__4,inputRegisters_235__3,inputRegisters_235__2,
            inputRegisters_235__1,inputRegisters_235__0})) ;
    Reg_16 loop1_235_x (.D ({inputRegisters_235__15,inputRegisters_235__14,
           inputRegisters_235__13,inputRegisters_235__12,inputRegisters_235__11,
           inputRegisters_235__10,inputRegisters_235__9,inputRegisters_235__8,
           inputRegisters_235__7,inputRegisters_235__6,inputRegisters_235__5,
           inputRegisters_235__4,inputRegisters_235__3,inputRegisters_235__2,
           inputRegisters_235__1,inputRegisters_235__0}), .en (
           enableRegister_235), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_235__15,registerOutputs_235__14,
           registerOutputs_235__13,registerOutputs_235__12,
           registerOutputs_235__11,registerOutputs_235__10,
           registerOutputs_235__9,registerOutputs_235__8,registerOutputs_235__7,
           registerOutputs_235__6,registerOutputs_235__5,registerOutputs_235__4,
           registerOutputs_235__3,registerOutputs_235__2,registerOutputs_235__1,
           registerOutputs_235__0})) ;
    Mux2_16 loop1_236_y (.A ({nx35951,nx36093,nx36235,nx36377,nx36519,nx36661,
            nx36803,nx36945,nx37087,nx37229,nx37371,nx37513,nx37655,nx37797,
            nx37939,nx38081}), .B ({nx33707,nx33845,nx33985,nx34123,nx34261,
            nx34399,nx34537,nx34677,nx34819,nx34961,nx35103,nx35245,nx35387,
            nx35529,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35671), .C ({inputRegisters_236__15,inputRegisters_236__14,
            inputRegisters_236__13,inputRegisters_236__12,inputRegisters_236__11
            ,inputRegisters_236__10,inputRegisters_236__9,inputRegisters_236__8,
            inputRegisters_236__7,inputRegisters_236__6,inputRegisters_236__5,
            inputRegisters_236__4,inputRegisters_236__3,inputRegisters_236__2,
            inputRegisters_236__1,inputRegisters_236__0})) ;
    Reg_16 loop1_236_x (.D ({inputRegisters_236__15,inputRegisters_236__14,
           inputRegisters_236__13,inputRegisters_236__12,inputRegisters_236__11,
           inputRegisters_236__10,inputRegisters_236__9,inputRegisters_236__8,
           inputRegisters_236__7,inputRegisters_236__6,inputRegisters_236__5,
           inputRegisters_236__4,inputRegisters_236__3,inputRegisters_236__2,
           inputRegisters_236__1,inputRegisters_236__0}), .en (
           enableRegister_236), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_236__15,registerOutputs_236__14,
           registerOutputs_236__13,registerOutputs_236__12,
           registerOutputs_236__11,registerOutputs_236__10,
           registerOutputs_236__9,registerOutputs_236__8,registerOutputs_236__7,
           registerOutputs_236__6,registerOutputs_236__5,registerOutputs_236__4,
           registerOutputs_236__3,registerOutputs_236__2,registerOutputs_236__1,
           registerOutputs_236__0})) ;
    Mux2_16 loop1_237_y (.A ({nx35951,nx36093,nx36235,nx36377,nx36519,nx36661,
            nx36803,nx36945,nx37087,nx37229,nx37371,nx37513,nx37655,nx37797,
            nx37939,nx38081}), .B ({nx33707,nx33847,nx33985,nx34123,nx34261,
            nx34399,nx34537,nx34677,nx34819,nx34961,nx35103,nx35245,nx35387,
            nx35529,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35671), .C ({inputRegisters_237__15,inputRegisters_237__14,
            inputRegisters_237__13,inputRegisters_237__12,inputRegisters_237__11
            ,inputRegisters_237__10,inputRegisters_237__9,inputRegisters_237__8,
            inputRegisters_237__7,inputRegisters_237__6,inputRegisters_237__5,
            inputRegisters_237__4,inputRegisters_237__3,inputRegisters_237__2,
            inputRegisters_237__1,inputRegisters_237__0})) ;
    Reg_16 loop1_237_x (.D ({inputRegisters_237__15,inputRegisters_237__14,
           inputRegisters_237__13,inputRegisters_237__12,inputRegisters_237__11,
           inputRegisters_237__10,inputRegisters_237__9,inputRegisters_237__8,
           inputRegisters_237__7,inputRegisters_237__6,inputRegisters_237__5,
           inputRegisters_237__4,inputRegisters_237__3,inputRegisters_237__2,
           inputRegisters_237__1,inputRegisters_237__0}), .en (
           enableRegister_237), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_237__15,registerOutputs_237__14,
           registerOutputs_237__13,registerOutputs_237__12,
           registerOutputs_237__11,registerOutputs_237__10,
           registerOutputs_237__9,registerOutputs_237__8,registerOutputs_237__7,
           registerOutputs_237__6,registerOutputs_237__5,registerOutputs_237__4,
           registerOutputs_237__3,registerOutputs_237__2,registerOutputs_237__1,
           registerOutputs_237__0})) ;
    Mux2_16 loop1_238_y (.A ({nx35953,nx36095,nx36237,nx36379,nx36521,nx36663,
            nx36805,nx36947,nx37089,nx37231,nx37373,nx37515,nx37657,nx37799,
            nx37941,nx38083}), .B ({nx33709,nx33847,nx33985,nx34123,nx34261,
            nx34399,nx34537,nx34679,nx34821,nx34963,nx35105,nx35247,nx35389,
            nx35531,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35673), .C ({inputRegisters_238__15,inputRegisters_238__14,
            inputRegisters_238__13,inputRegisters_238__12,inputRegisters_238__11
            ,inputRegisters_238__10,inputRegisters_238__9,inputRegisters_238__8,
            inputRegisters_238__7,inputRegisters_238__6,inputRegisters_238__5,
            inputRegisters_238__4,inputRegisters_238__3,inputRegisters_238__2,
            inputRegisters_238__1,inputRegisters_238__0})) ;
    Reg_16 loop1_238_x (.D ({inputRegisters_238__15,inputRegisters_238__14,
           inputRegisters_238__13,inputRegisters_238__12,inputRegisters_238__11,
           inputRegisters_238__10,inputRegisters_238__9,inputRegisters_238__8,
           inputRegisters_238__7,inputRegisters_238__6,inputRegisters_238__5,
           inputRegisters_238__4,inputRegisters_238__3,inputRegisters_238__2,
           inputRegisters_238__1,inputRegisters_238__0}), .en (
           enableRegister_238), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_238__15,registerOutputs_238__14,
           registerOutputs_238__13,registerOutputs_238__12,
           registerOutputs_238__11,registerOutputs_238__10,
           registerOutputs_238__9,registerOutputs_238__8,registerOutputs_238__7,
           registerOutputs_238__6,registerOutputs_238__5,registerOutputs_238__4,
           registerOutputs_238__3,registerOutputs_238__2,registerOutputs_238__1,
           registerOutputs_238__0})) ;
    Mux2_16 loop1_239_y (.A ({nx35953,nx36095,nx36237,nx36379,nx36521,nx36663,
            nx36805,nx36947,nx37089,nx37231,nx37373,nx37515,nx37657,nx37799,
            nx37941,nx38083}), .B ({nx33709,nx33847,nx33985,nx34123,nx34261,
            nx34399,nx34539,nx34679,nx34821,nx34963,nx35105,nx35247,nx35389,
            nx35531,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35673), .C ({inputRegisters_239__15,inputRegisters_239__14,
            inputRegisters_239__13,inputRegisters_239__12,inputRegisters_239__11
            ,inputRegisters_239__10,inputRegisters_239__9,inputRegisters_239__8,
            inputRegisters_239__7,inputRegisters_239__6,inputRegisters_239__5,
            inputRegisters_239__4,inputRegisters_239__3,inputRegisters_239__2,
            inputRegisters_239__1,inputRegisters_239__0})) ;
    Reg_16 loop1_239_x (.D ({inputRegisters_239__15,inputRegisters_239__14,
           inputRegisters_239__13,inputRegisters_239__12,inputRegisters_239__11,
           inputRegisters_239__10,inputRegisters_239__9,inputRegisters_239__8,
           inputRegisters_239__7,inputRegisters_239__6,inputRegisters_239__5,
           inputRegisters_239__4,inputRegisters_239__3,inputRegisters_239__2,
           inputRegisters_239__1,inputRegisters_239__0}), .en (
           enableRegister_239), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_239__15,registerOutputs_239__14,
           registerOutputs_239__13,registerOutputs_239__12,
           registerOutputs_239__11,registerOutputs_239__10,
           registerOutputs_239__9,registerOutputs_239__8,registerOutputs_239__7,
           registerOutputs_239__6,registerOutputs_239__5,registerOutputs_239__4,
           registerOutputs_239__3,registerOutputs_239__2,registerOutputs_239__1,
           registerOutputs_239__0})) ;
    Mux2_16 loop1_240_y (.A ({nx35953,nx36095,nx36237,nx36379,nx36521,nx36663,
            nx36805,nx36947,nx37089,nx37231,nx37373,nx37515,nx37657,nx37799,
            nx37941,nx38083}), .B ({nx33709,nx33847,nx33985,nx34123,nx34261,
            nx34401,nx34539,nx34679,nx34821,nx34963,nx35105,nx35247,nx35389,
            nx35531,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35673), .C ({inputRegisters_240__15,inputRegisters_240__14,
            inputRegisters_240__13,inputRegisters_240__12,inputRegisters_240__11
            ,inputRegisters_240__10,inputRegisters_240__9,inputRegisters_240__8,
            inputRegisters_240__7,inputRegisters_240__6,inputRegisters_240__5,
            inputRegisters_240__4,inputRegisters_240__3,inputRegisters_240__2,
            inputRegisters_240__1,inputRegisters_240__0})) ;
    Reg_16 loop1_240_x (.D ({inputRegisters_240__15,inputRegisters_240__14,
           inputRegisters_240__13,inputRegisters_240__12,inputRegisters_240__11,
           inputRegisters_240__10,inputRegisters_240__9,inputRegisters_240__8,
           inputRegisters_240__7,inputRegisters_240__6,inputRegisters_240__5,
           inputRegisters_240__4,inputRegisters_240__3,inputRegisters_240__2,
           inputRegisters_240__1,inputRegisters_240__0}), .en (
           enableRegister_240), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_240__15,registerOutputs_240__14,
           registerOutputs_240__13,registerOutputs_240__12,
           registerOutputs_240__11,registerOutputs_240__10,
           registerOutputs_240__9,registerOutputs_240__8,registerOutputs_240__7,
           registerOutputs_240__6,registerOutputs_240__5,registerOutputs_240__4,
           registerOutputs_240__3,registerOutputs_240__2,registerOutputs_240__1,
           registerOutputs_240__0})) ;
    Mux2_16 loop1_241_y (.A ({nx35953,nx36095,nx36237,nx36379,nx36521,nx36663,
            nx36805,nx36947,nx37089,nx37231,nx37373,nx37515,nx37657,nx37799,
            nx37941,nx38083}), .B ({nx33709,nx33847,nx33985,nx34123,nx34263,
            nx34401,nx34539,nx34679,nx34821,nx34963,nx35105,nx35247,nx35389,
            nx35531,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35673), .C ({inputRegisters_241__15,inputRegisters_241__14,
            inputRegisters_241__13,inputRegisters_241__12,inputRegisters_241__11
            ,inputRegisters_241__10,inputRegisters_241__9,inputRegisters_241__8,
            inputRegisters_241__7,inputRegisters_241__6,inputRegisters_241__5,
            inputRegisters_241__4,inputRegisters_241__3,inputRegisters_241__2,
            inputRegisters_241__1,inputRegisters_241__0})) ;
    Reg_16 loop1_241_x (.D ({inputRegisters_241__15,inputRegisters_241__14,
           inputRegisters_241__13,inputRegisters_241__12,inputRegisters_241__11,
           inputRegisters_241__10,inputRegisters_241__9,inputRegisters_241__8,
           inputRegisters_241__7,inputRegisters_241__6,inputRegisters_241__5,
           inputRegisters_241__4,inputRegisters_241__3,inputRegisters_241__2,
           inputRegisters_241__1,inputRegisters_241__0}), .en (
           enableRegister_241), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_241__15,registerOutputs_241__14,
           registerOutputs_241__13,registerOutputs_241__12,
           registerOutputs_241__11,registerOutputs_241__10,
           registerOutputs_241__9,registerOutputs_241__8,registerOutputs_241__7,
           registerOutputs_241__6,registerOutputs_241__5,registerOutputs_241__4,
           registerOutputs_241__3,registerOutputs_241__2,registerOutputs_241__1,
           registerOutputs_241__0})) ;
    Mux2_16 loop1_242_y (.A ({nx35953,nx36095,nx36237,nx36379,nx36521,nx36663,
            nx36805,nx36947,nx37089,nx37231,nx37373,nx37515,nx37657,nx37799,
            nx37941,nx38083}), .B ({nx33709,nx33847,nx33985,nx34125,nx34263,
            nx34401,nx34539,nx34679,nx34821,nx34963,nx35105,nx35247,nx35389,
            nx35531,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35673), .C ({inputRegisters_242__15,inputRegisters_242__14,
            inputRegisters_242__13,inputRegisters_242__12,inputRegisters_242__11
            ,inputRegisters_242__10,inputRegisters_242__9,inputRegisters_242__8,
            inputRegisters_242__7,inputRegisters_242__6,inputRegisters_242__5,
            inputRegisters_242__4,inputRegisters_242__3,inputRegisters_242__2,
            inputRegisters_242__1,inputRegisters_242__0})) ;
    Reg_16 loop1_242_x (.D ({inputRegisters_242__15,inputRegisters_242__14,
           inputRegisters_242__13,inputRegisters_242__12,inputRegisters_242__11,
           inputRegisters_242__10,inputRegisters_242__9,inputRegisters_242__8,
           inputRegisters_242__7,inputRegisters_242__6,inputRegisters_242__5,
           inputRegisters_242__4,inputRegisters_242__3,inputRegisters_242__2,
           inputRegisters_242__1,inputRegisters_242__0}), .en (
           enableRegister_242), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_242__15,registerOutputs_242__14,
           registerOutputs_242__13,registerOutputs_242__12,
           registerOutputs_242__11,registerOutputs_242__10,
           registerOutputs_242__9,registerOutputs_242__8,registerOutputs_242__7,
           registerOutputs_242__6,registerOutputs_242__5,registerOutputs_242__4,
           registerOutputs_242__3,registerOutputs_242__2,registerOutputs_242__1,
           registerOutputs_242__0})) ;
    Mux2_16 loop1_243_y (.A ({nx35953,nx36095,nx36237,nx36379,nx36521,nx36663,
            nx36805,nx36947,nx37089,nx37231,nx37373,nx37515,nx37657,nx37799,
            nx37941,nx38083}), .B ({nx33709,nx33847,nx33987,nx34125,nx34263,
            nx34401,nx34539,nx34679,nx34821,nx34963,nx35105,nx35247,nx35389,
            nx35531,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35673), .C ({inputRegisters_243__15,inputRegisters_243__14,
            inputRegisters_243__13,inputRegisters_243__12,inputRegisters_243__11
            ,inputRegisters_243__10,inputRegisters_243__9,inputRegisters_243__8,
            inputRegisters_243__7,inputRegisters_243__6,inputRegisters_243__5,
            inputRegisters_243__4,inputRegisters_243__3,inputRegisters_243__2,
            inputRegisters_243__1,inputRegisters_243__0})) ;
    Reg_16 loop1_243_x (.D ({inputRegisters_243__15,inputRegisters_243__14,
           inputRegisters_243__13,inputRegisters_243__12,inputRegisters_243__11,
           inputRegisters_243__10,inputRegisters_243__9,inputRegisters_243__8,
           inputRegisters_243__7,inputRegisters_243__6,inputRegisters_243__5,
           inputRegisters_243__4,inputRegisters_243__3,inputRegisters_243__2,
           inputRegisters_243__1,inputRegisters_243__0}), .en (
           enableRegister_243), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_243__15,registerOutputs_243__14,
           registerOutputs_243__13,registerOutputs_243__12,
           registerOutputs_243__11,registerOutputs_243__10,
           registerOutputs_243__9,registerOutputs_243__8,registerOutputs_243__7,
           registerOutputs_243__6,registerOutputs_243__5,registerOutputs_243__4,
           registerOutputs_243__3,registerOutputs_243__2,registerOutputs_243__1,
           registerOutputs_243__0})) ;
    Mux2_16 loop1_244_y (.A ({nx35953,nx36095,nx36237,nx36379,nx36521,nx36663,
            nx36805,nx36947,nx37089,nx37231,nx37373,nx37515,nx37657,nx37799,
            nx37941,nx38083}), .B ({nx33709,nx33849,nx33987,nx34125,nx34263,
            nx34401,nx34539,nx34679,nx34821,nx34963,nx35105,nx35247,nx35389,
            nx35531,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35673), .C ({inputRegisters_244__15,inputRegisters_244__14,
            inputRegisters_244__13,inputRegisters_244__12,inputRegisters_244__11
            ,inputRegisters_244__10,inputRegisters_244__9,inputRegisters_244__8,
            inputRegisters_244__7,inputRegisters_244__6,inputRegisters_244__5,
            inputRegisters_244__4,inputRegisters_244__3,inputRegisters_244__2,
            inputRegisters_244__1,inputRegisters_244__0})) ;
    Reg_16 loop1_244_x (.D ({inputRegisters_244__15,inputRegisters_244__14,
           inputRegisters_244__13,inputRegisters_244__12,inputRegisters_244__11,
           inputRegisters_244__10,inputRegisters_244__9,inputRegisters_244__8,
           inputRegisters_244__7,inputRegisters_244__6,inputRegisters_244__5,
           inputRegisters_244__4,inputRegisters_244__3,inputRegisters_244__2,
           inputRegisters_244__1,inputRegisters_244__0}), .en (
           enableRegister_244), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_244__15,registerOutputs_244__14,
           registerOutputs_244__13,registerOutputs_244__12,
           registerOutputs_244__11,registerOutputs_244__10,
           registerOutputs_244__9,registerOutputs_244__8,registerOutputs_244__7,
           registerOutputs_244__6,registerOutputs_244__5,registerOutputs_244__4,
           registerOutputs_244__3,registerOutputs_244__2,registerOutputs_244__1,
           registerOutputs_244__0})) ;
    Mux2_16 loop1_245_y (.A ({nx35955,nx36097,nx36239,nx36381,nx36523,nx36665,
            nx36807,nx36949,nx37091,nx37233,nx37375,nx37517,nx37659,nx37801,
            nx37943,nx38085}), .B ({nx33711,nx33849,nx33987,nx34125,nx34263,
            nx34401,nx34539,nx34681,nx34823,nx34965,nx35107,nx35249,nx35391,
            nx35533,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35675), .C ({inputRegisters_245__15,inputRegisters_245__14,
            inputRegisters_245__13,inputRegisters_245__12,inputRegisters_245__11
            ,inputRegisters_245__10,inputRegisters_245__9,inputRegisters_245__8,
            inputRegisters_245__7,inputRegisters_245__6,inputRegisters_245__5,
            inputRegisters_245__4,inputRegisters_245__3,inputRegisters_245__2,
            inputRegisters_245__1,inputRegisters_245__0})) ;
    Reg_16 loop1_245_x (.D ({inputRegisters_245__15,inputRegisters_245__14,
           inputRegisters_245__13,inputRegisters_245__12,inputRegisters_245__11,
           inputRegisters_245__10,inputRegisters_245__9,inputRegisters_245__8,
           inputRegisters_245__7,inputRegisters_245__6,inputRegisters_245__5,
           inputRegisters_245__4,inputRegisters_245__3,inputRegisters_245__2,
           inputRegisters_245__1,inputRegisters_245__0}), .en (
           enableRegister_245), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_245__15,registerOutputs_245__14,
           registerOutputs_245__13,registerOutputs_245__12,
           registerOutputs_245__11,registerOutputs_245__10,
           registerOutputs_245__9,registerOutputs_245__8,registerOutputs_245__7,
           registerOutputs_245__6,registerOutputs_245__5,registerOutputs_245__4,
           registerOutputs_245__3,registerOutputs_245__2,registerOutputs_245__1,
           registerOutputs_245__0})) ;
    Mux2_16 loop1_246_y (.A ({nx35955,nx36097,nx36239,nx36381,nx36523,nx36665,
            nx36807,nx36949,nx37091,nx37233,nx37375,nx37517,nx37659,nx37801,
            nx37943,nx38085}), .B ({nx33711,nx33849,nx33987,nx34125,nx34263,
            nx34401,nx34541,nx34681,nx34823,nx34965,nx35107,nx35249,nx35391,
            nx35533,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35675), .C ({inputRegisters_246__15,inputRegisters_246__14,
            inputRegisters_246__13,inputRegisters_246__12,inputRegisters_246__11
            ,inputRegisters_246__10,inputRegisters_246__9,inputRegisters_246__8,
            inputRegisters_246__7,inputRegisters_246__6,inputRegisters_246__5,
            inputRegisters_246__4,inputRegisters_246__3,inputRegisters_246__2,
            inputRegisters_246__1,inputRegisters_246__0})) ;
    Reg_16 loop1_246_x (.D ({inputRegisters_246__15,inputRegisters_246__14,
           inputRegisters_246__13,inputRegisters_246__12,inputRegisters_246__11,
           inputRegisters_246__10,inputRegisters_246__9,inputRegisters_246__8,
           inputRegisters_246__7,inputRegisters_246__6,inputRegisters_246__5,
           inputRegisters_246__4,inputRegisters_246__3,inputRegisters_246__2,
           inputRegisters_246__1,inputRegisters_246__0}), .en (
           enableRegister_246), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_246__15,registerOutputs_246__14,
           registerOutputs_246__13,registerOutputs_246__12,
           registerOutputs_246__11,registerOutputs_246__10,
           registerOutputs_246__9,registerOutputs_246__8,registerOutputs_246__7,
           registerOutputs_246__6,registerOutputs_246__5,registerOutputs_246__4,
           registerOutputs_246__3,registerOutputs_246__2,registerOutputs_246__1,
           registerOutputs_246__0})) ;
    Mux2_16 loop1_247_y (.A ({nx35955,nx36097,nx36239,nx36381,nx36523,nx36665,
            nx36807,nx36949,nx37091,nx37233,nx37375,nx37517,nx37659,nx37801,
            nx37943,nx38085}), .B ({nx33711,nx33849,nx33987,nx34125,nx34263,
            nx34403,nx34541,nx34681,nx34823,nx34965,nx35107,nx35249,nx35391,
            nx35533,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35675), .C ({inputRegisters_247__15,inputRegisters_247__14,
            inputRegisters_247__13,inputRegisters_247__12,inputRegisters_247__11
            ,inputRegisters_247__10,inputRegisters_247__9,inputRegisters_247__8,
            inputRegisters_247__7,inputRegisters_247__6,inputRegisters_247__5,
            inputRegisters_247__4,inputRegisters_247__3,inputRegisters_247__2,
            inputRegisters_247__1,inputRegisters_247__0})) ;
    Reg_16 loop1_247_x (.D ({inputRegisters_247__15,inputRegisters_247__14,
           inputRegisters_247__13,inputRegisters_247__12,inputRegisters_247__11,
           inputRegisters_247__10,inputRegisters_247__9,inputRegisters_247__8,
           inputRegisters_247__7,inputRegisters_247__6,inputRegisters_247__5,
           inputRegisters_247__4,inputRegisters_247__3,inputRegisters_247__2,
           inputRegisters_247__1,inputRegisters_247__0}), .en (
           enableRegister_247), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_247__15,registerOutputs_247__14,
           registerOutputs_247__13,registerOutputs_247__12,
           registerOutputs_247__11,registerOutputs_247__10,
           registerOutputs_247__9,registerOutputs_247__8,registerOutputs_247__7,
           registerOutputs_247__6,registerOutputs_247__5,registerOutputs_247__4,
           registerOutputs_247__3,registerOutputs_247__2,registerOutputs_247__1,
           registerOutputs_247__0})) ;
    Mux2_16 loop1_248_y (.A ({nx35955,nx36097,nx36239,nx36381,nx36523,nx36665,
            nx36807,nx36949,nx37091,nx37233,nx37375,nx37517,nx37659,nx37801,
            nx37943,nx38085}), .B ({nx33711,nx33849,nx33987,nx34125,nx34265,
            nx34403,nx34541,nx34681,nx34823,nx34965,nx35107,nx35249,nx35391,
            nx35533,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35675), .C ({inputRegisters_248__15,inputRegisters_248__14,
            inputRegisters_248__13,inputRegisters_248__12,inputRegisters_248__11
            ,inputRegisters_248__10,inputRegisters_248__9,inputRegisters_248__8,
            inputRegisters_248__7,inputRegisters_248__6,inputRegisters_248__5,
            inputRegisters_248__4,inputRegisters_248__3,inputRegisters_248__2,
            inputRegisters_248__1,inputRegisters_248__0})) ;
    Reg_16 loop1_248_x (.D ({inputRegisters_248__15,inputRegisters_248__14,
           inputRegisters_248__13,inputRegisters_248__12,inputRegisters_248__11,
           inputRegisters_248__10,inputRegisters_248__9,inputRegisters_248__8,
           inputRegisters_248__7,inputRegisters_248__6,inputRegisters_248__5,
           inputRegisters_248__4,inputRegisters_248__3,inputRegisters_248__2,
           inputRegisters_248__1,inputRegisters_248__0}), .en (
           enableRegister_248), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_248__15,registerOutputs_248__14,
           registerOutputs_248__13,registerOutputs_248__12,
           registerOutputs_248__11,registerOutputs_248__10,
           registerOutputs_248__9,registerOutputs_248__8,registerOutputs_248__7,
           registerOutputs_248__6,registerOutputs_248__5,registerOutputs_248__4,
           registerOutputs_248__3,registerOutputs_248__2,registerOutputs_248__1,
           registerOutputs_248__0})) ;
    Mux2_16 loop1_249_y (.A ({nx35955,nx36097,nx36239,nx36381,nx36523,nx36665,
            nx36807,nx36949,nx37091,nx37233,nx37375,nx37517,nx37659,nx37801,
            nx37943,nx38085}), .B ({nx33711,nx33849,nx33987,nx34127,nx34265,
            nx34403,nx34541,nx34681,nx34823,nx34965,nx35107,nx35249,nx35391,
            nx35533,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35675), .C ({inputRegisters_249__15,inputRegisters_249__14,
            inputRegisters_249__13,inputRegisters_249__12,inputRegisters_249__11
            ,inputRegisters_249__10,inputRegisters_249__9,inputRegisters_249__8,
            inputRegisters_249__7,inputRegisters_249__6,inputRegisters_249__5,
            inputRegisters_249__4,inputRegisters_249__3,inputRegisters_249__2,
            inputRegisters_249__1,inputRegisters_249__0})) ;
    Reg_16 loop1_249_x (.D ({inputRegisters_249__15,inputRegisters_249__14,
           inputRegisters_249__13,inputRegisters_249__12,inputRegisters_249__11,
           inputRegisters_249__10,inputRegisters_249__9,inputRegisters_249__8,
           inputRegisters_249__7,inputRegisters_249__6,inputRegisters_249__5,
           inputRegisters_249__4,inputRegisters_249__3,inputRegisters_249__2,
           inputRegisters_249__1,inputRegisters_249__0}), .en (
           enableRegister_249), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_249__15,registerOutputs_249__14,
           registerOutputs_249__13,registerOutputs_249__12,
           registerOutputs_249__11,registerOutputs_249__10,
           registerOutputs_249__9,registerOutputs_249__8,registerOutputs_249__7,
           registerOutputs_249__6,registerOutputs_249__5,registerOutputs_249__4,
           registerOutputs_249__3,registerOutputs_249__2,registerOutputs_249__1,
           registerOutputs_249__0})) ;
    Mux2_16 loop1_250_y (.A ({nx35955,nx36097,nx36239,nx36381,nx36523,nx36665,
            nx36807,nx36949,nx37091,nx37233,nx37375,nx37517,nx37659,nx37801,
            nx37943,nx38085}), .B ({nx33711,nx33849,nx33989,nx34127,nx34265,
            nx34403,nx34541,nx34681,nx34823,nx34965,nx35107,nx35249,nx35391,
            nx35533,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35675), .C ({inputRegisters_250__15,inputRegisters_250__14,
            inputRegisters_250__13,inputRegisters_250__12,inputRegisters_250__11
            ,inputRegisters_250__10,inputRegisters_250__9,inputRegisters_250__8,
            inputRegisters_250__7,inputRegisters_250__6,inputRegisters_250__5,
            inputRegisters_250__4,inputRegisters_250__3,inputRegisters_250__2,
            inputRegisters_250__1,inputRegisters_250__0})) ;
    Reg_16 loop1_250_x (.D ({inputRegisters_250__15,inputRegisters_250__14,
           inputRegisters_250__13,inputRegisters_250__12,inputRegisters_250__11,
           inputRegisters_250__10,inputRegisters_250__9,inputRegisters_250__8,
           inputRegisters_250__7,inputRegisters_250__6,inputRegisters_250__5,
           inputRegisters_250__4,inputRegisters_250__3,inputRegisters_250__2,
           inputRegisters_250__1,inputRegisters_250__0}), .en (
           enableRegister_250), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_250__15,registerOutputs_250__14,
           registerOutputs_250__13,registerOutputs_250__12,
           registerOutputs_250__11,registerOutputs_250__10,
           registerOutputs_250__9,registerOutputs_250__8,registerOutputs_250__7,
           registerOutputs_250__6,registerOutputs_250__5,registerOutputs_250__4,
           registerOutputs_250__3,registerOutputs_250__2,registerOutputs_250__1,
           registerOutputs_250__0})) ;
    Mux2_16 loop1_251_y (.A ({nx35955,nx36097,nx36239,nx36381,nx36523,nx36665,
            nx36807,nx36949,nx37091,nx37233,nx37375,nx37517,nx37659,nx37801,
            nx37943,nx38085}), .B ({nx33711,nx33851,nx33989,nx34127,nx34265,
            nx34403,nx34541,nx34681,nx34823,nx34965,nx35107,nx35249,nx35391,
            nx35533,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35675), .C ({inputRegisters_251__15,inputRegisters_251__14,
            inputRegisters_251__13,inputRegisters_251__12,inputRegisters_251__11
            ,inputRegisters_251__10,inputRegisters_251__9,inputRegisters_251__8,
            inputRegisters_251__7,inputRegisters_251__6,inputRegisters_251__5,
            inputRegisters_251__4,inputRegisters_251__3,inputRegisters_251__2,
            inputRegisters_251__1,inputRegisters_251__0})) ;
    Reg_16 loop1_251_x (.D ({inputRegisters_251__15,inputRegisters_251__14,
           inputRegisters_251__13,inputRegisters_251__12,inputRegisters_251__11,
           inputRegisters_251__10,inputRegisters_251__9,inputRegisters_251__8,
           inputRegisters_251__7,inputRegisters_251__6,inputRegisters_251__5,
           inputRegisters_251__4,inputRegisters_251__3,inputRegisters_251__2,
           inputRegisters_251__1,inputRegisters_251__0}), .en (
           enableRegister_251), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_251__15,registerOutputs_251__14,
           registerOutputs_251__13,registerOutputs_251__12,
           registerOutputs_251__11,registerOutputs_251__10,
           registerOutputs_251__9,registerOutputs_251__8,registerOutputs_251__7,
           registerOutputs_251__6,registerOutputs_251__5,registerOutputs_251__4,
           registerOutputs_251__3,registerOutputs_251__2,registerOutputs_251__1,
           registerOutputs_251__0})) ;
    Mux2_16 loop1_252_y (.A ({nx35957,nx36099,nx36241,nx36383,nx36525,nx36667,
            nx36809,nx36951,nx37093,nx37235,nx37377,nx37519,nx37661,nx37803,
            nx37945,nx38087}), .B ({nx33713,nx33851,nx33989,nx34127,nx34265,
            nx34403,nx34541,nx34683,nx34825,nx34967,nx35109,nx35251,nx35393,
            nx35535,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35677), .C ({inputRegisters_252__15,inputRegisters_252__14,
            inputRegisters_252__13,inputRegisters_252__12,inputRegisters_252__11
            ,inputRegisters_252__10,inputRegisters_252__9,inputRegisters_252__8,
            inputRegisters_252__7,inputRegisters_252__6,inputRegisters_252__5,
            inputRegisters_252__4,inputRegisters_252__3,inputRegisters_252__2,
            inputRegisters_252__1,inputRegisters_252__0})) ;
    Reg_16 loop1_252_x (.D ({inputRegisters_252__15,inputRegisters_252__14,
           inputRegisters_252__13,inputRegisters_252__12,inputRegisters_252__11,
           inputRegisters_252__10,inputRegisters_252__9,inputRegisters_252__8,
           inputRegisters_252__7,inputRegisters_252__6,inputRegisters_252__5,
           inputRegisters_252__4,inputRegisters_252__3,inputRegisters_252__2,
           inputRegisters_252__1,inputRegisters_252__0}), .en (
           enableRegister_252), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_252__15,registerOutputs_252__14,
           registerOutputs_252__13,registerOutputs_252__12,
           registerOutputs_252__11,registerOutputs_252__10,
           registerOutputs_252__9,registerOutputs_252__8,registerOutputs_252__7,
           registerOutputs_252__6,registerOutputs_252__5,registerOutputs_252__4,
           registerOutputs_252__3,registerOutputs_252__2,registerOutputs_252__1,
           registerOutputs_252__0})) ;
    Mux2_16 loop1_253_y (.A ({nx35957,nx36099,nx36241,nx36383,nx36525,nx36667,
            nx36809,nx36951,nx37093,nx37235,nx37377,nx37519,nx37661,nx37803,
            nx37945,nx38087}), .B ({nx33713,nx33851,nx33989,nx34127,nx34265,
            nx34403,nx34543,nx34683,nx34825,nx34967,nx35109,nx35251,nx35393,
            nx35535,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35677), .C ({inputRegisters_253__15,inputRegisters_253__14,
            inputRegisters_253__13,inputRegisters_253__12,inputRegisters_253__11
            ,inputRegisters_253__10,inputRegisters_253__9,inputRegisters_253__8,
            inputRegisters_253__7,inputRegisters_253__6,inputRegisters_253__5,
            inputRegisters_253__4,inputRegisters_253__3,inputRegisters_253__2,
            inputRegisters_253__1,inputRegisters_253__0})) ;
    Reg_16 loop1_253_x (.D ({inputRegisters_253__15,inputRegisters_253__14,
           inputRegisters_253__13,inputRegisters_253__12,inputRegisters_253__11,
           inputRegisters_253__10,inputRegisters_253__9,inputRegisters_253__8,
           inputRegisters_253__7,inputRegisters_253__6,inputRegisters_253__5,
           inputRegisters_253__4,inputRegisters_253__3,inputRegisters_253__2,
           inputRegisters_253__1,inputRegisters_253__0}), .en (
           enableRegister_253), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_253__15,registerOutputs_253__14,
           registerOutputs_253__13,registerOutputs_253__12,
           registerOutputs_253__11,registerOutputs_253__10,
           registerOutputs_253__9,registerOutputs_253__8,registerOutputs_253__7,
           registerOutputs_253__6,registerOutputs_253__5,registerOutputs_253__4,
           registerOutputs_253__3,registerOutputs_253__2,registerOutputs_253__1,
           registerOutputs_253__0})) ;
    Mux2_16 loop1_254_y (.A ({nx35957,nx36099,nx36241,nx36383,nx36525,nx36667,
            nx36809,nx36951,nx37093,nx37235,nx37377,nx37519,nx37661,nx37803,
            nx37945,nx38087}), .B ({nx33713,nx33851,nx33989,nx34127,nx34265,
            nx34405,nx34543,nx34683,nx34825,nx34967,nx35109,nx35251,nx35393,
            nx35535,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35677), .C ({inputRegisters_254__15,inputRegisters_254__14,
            inputRegisters_254__13,inputRegisters_254__12,inputRegisters_254__11
            ,inputRegisters_254__10,inputRegisters_254__9,inputRegisters_254__8,
            inputRegisters_254__7,inputRegisters_254__6,inputRegisters_254__5,
            inputRegisters_254__4,inputRegisters_254__3,inputRegisters_254__2,
            inputRegisters_254__1,inputRegisters_254__0})) ;
    Reg_16 loop1_254_x (.D ({inputRegisters_254__15,inputRegisters_254__14,
           inputRegisters_254__13,inputRegisters_254__12,inputRegisters_254__11,
           inputRegisters_254__10,inputRegisters_254__9,inputRegisters_254__8,
           inputRegisters_254__7,inputRegisters_254__6,inputRegisters_254__5,
           inputRegisters_254__4,inputRegisters_254__3,inputRegisters_254__2,
           inputRegisters_254__1,inputRegisters_254__0}), .en (
           enableRegister_254), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_254__15,registerOutputs_254__14,
           registerOutputs_254__13,registerOutputs_254__12,
           registerOutputs_254__11,registerOutputs_254__10,
           registerOutputs_254__9,registerOutputs_254__8,registerOutputs_254__7,
           registerOutputs_254__6,registerOutputs_254__5,registerOutputs_254__4,
           registerOutputs_254__3,registerOutputs_254__2,registerOutputs_254__1,
           registerOutputs_254__0})) ;
    Mux2_16 loop1_255_y (.A ({nx35957,nx36099,nx36241,nx36383,nx36525,nx36667,
            nx36809,nx36951,nx37093,nx37235,nx37377,nx37519,nx37661,nx37803,
            nx37945,nx38087}), .B ({nx33713,nx33851,nx33989,nx34127,nx34267,
            nx34405,nx34543,nx34683,nx34825,nx34967,nx35109,nx35251,nx35393,
            nx35535,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35677), .C ({inputRegisters_255__15,inputRegisters_255__14,
            inputRegisters_255__13,inputRegisters_255__12,inputRegisters_255__11
            ,inputRegisters_255__10,inputRegisters_255__9,inputRegisters_255__8,
            inputRegisters_255__7,inputRegisters_255__6,inputRegisters_255__5,
            inputRegisters_255__4,inputRegisters_255__3,inputRegisters_255__2,
            inputRegisters_255__1,inputRegisters_255__0})) ;
    Reg_16 loop1_255_x (.D ({inputRegisters_255__15,inputRegisters_255__14,
           inputRegisters_255__13,inputRegisters_255__12,inputRegisters_255__11,
           inputRegisters_255__10,inputRegisters_255__9,inputRegisters_255__8,
           inputRegisters_255__7,inputRegisters_255__6,inputRegisters_255__5,
           inputRegisters_255__4,inputRegisters_255__3,inputRegisters_255__2,
           inputRegisters_255__1,inputRegisters_255__0}), .en (
           enableRegister_255), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_255__15,registerOutputs_255__14,
           registerOutputs_255__13,registerOutputs_255__12,
           registerOutputs_255__11,registerOutputs_255__10,
           registerOutputs_255__9,registerOutputs_255__8,registerOutputs_255__7,
           registerOutputs_255__6,registerOutputs_255__5,registerOutputs_255__4,
           registerOutputs_255__3,registerOutputs_255__2,registerOutputs_255__1,
           registerOutputs_255__0})) ;
    Mux2_16 loop1_256_y (.A ({nx35957,nx36099,nx36241,nx36383,nx36525,nx36667,
            nx36809,nx36951,nx37093,nx37235,nx37377,nx37519,nx37661,nx37803,
            nx37945,nx38087}), .B ({nx33713,nx33851,nx33989,nx34129,nx34267,
            nx34405,nx34543,nx34683,nx34825,nx34967,nx35109,nx35251,nx35393,
            nx35535,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35677), .C ({inputRegisters_256__15,inputRegisters_256__14,
            inputRegisters_256__13,inputRegisters_256__12,inputRegisters_256__11
            ,inputRegisters_256__10,inputRegisters_256__9,inputRegisters_256__8,
            inputRegisters_256__7,inputRegisters_256__6,inputRegisters_256__5,
            inputRegisters_256__4,inputRegisters_256__3,inputRegisters_256__2,
            inputRegisters_256__1,inputRegisters_256__0})) ;
    Reg_16 loop1_256_x (.D ({inputRegisters_256__15,inputRegisters_256__14,
           inputRegisters_256__13,inputRegisters_256__12,inputRegisters_256__11,
           inputRegisters_256__10,inputRegisters_256__9,inputRegisters_256__8,
           inputRegisters_256__7,inputRegisters_256__6,inputRegisters_256__5,
           inputRegisters_256__4,inputRegisters_256__3,inputRegisters_256__2,
           inputRegisters_256__1,inputRegisters_256__0}), .en (
           enableRegister_256), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_256__15,registerOutputs_256__14,
           registerOutputs_256__13,registerOutputs_256__12,
           registerOutputs_256__11,registerOutputs_256__10,
           registerOutputs_256__9,registerOutputs_256__8,registerOutputs_256__7,
           registerOutputs_256__6,registerOutputs_256__5,registerOutputs_256__4,
           registerOutputs_256__3,registerOutputs_256__2,registerOutputs_256__1,
           registerOutputs_256__0})) ;
    Mux2_16 loop1_257_y (.A ({nx35957,nx36099,nx36241,nx36383,nx36525,nx36667,
            nx36809,nx36951,nx37093,nx37235,nx37377,nx37519,nx37661,nx37803,
            nx37945,nx38087}), .B ({nx33713,nx33851,nx33991,nx34129,nx34267,
            nx34405,nx34543,nx34683,nx34825,nx34967,nx35109,nx35251,nx35393,
            nx35535,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35677), .C ({inputRegisters_257__15,inputRegisters_257__14,
            inputRegisters_257__13,inputRegisters_257__12,inputRegisters_257__11
            ,inputRegisters_257__10,inputRegisters_257__9,inputRegisters_257__8,
            inputRegisters_257__7,inputRegisters_257__6,inputRegisters_257__5,
            inputRegisters_257__4,inputRegisters_257__3,inputRegisters_257__2,
            inputRegisters_257__1,inputRegisters_257__0})) ;
    Reg_16 loop1_257_x (.D ({inputRegisters_257__15,inputRegisters_257__14,
           inputRegisters_257__13,inputRegisters_257__12,inputRegisters_257__11,
           inputRegisters_257__10,inputRegisters_257__9,inputRegisters_257__8,
           inputRegisters_257__7,inputRegisters_257__6,inputRegisters_257__5,
           inputRegisters_257__4,inputRegisters_257__3,inputRegisters_257__2,
           inputRegisters_257__1,inputRegisters_257__0}), .en (
           enableRegister_257), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_257__15,registerOutputs_257__14,
           registerOutputs_257__13,registerOutputs_257__12,
           registerOutputs_257__11,registerOutputs_257__10,
           registerOutputs_257__9,registerOutputs_257__8,registerOutputs_257__7,
           registerOutputs_257__6,registerOutputs_257__5,registerOutputs_257__4,
           registerOutputs_257__3,registerOutputs_257__2,registerOutputs_257__1,
           registerOutputs_257__0})) ;
    Mux2_16 loop1_258_y (.A ({nx35957,nx36099,nx36241,nx36383,nx36525,nx36667,
            nx36809,nx36951,nx37093,nx37235,nx37377,nx37519,nx37661,nx37803,
            nx37945,nx38087}), .B ({nx33713,nx33853,nx33991,nx34129,nx34267,
            nx34405,nx34543,nx34683,nx34825,nx34967,nx35109,nx35251,nx35393,
            nx35535,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35677), .C ({inputRegisters_258__15,inputRegisters_258__14,
            inputRegisters_258__13,inputRegisters_258__12,inputRegisters_258__11
            ,inputRegisters_258__10,inputRegisters_258__9,inputRegisters_258__8,
            inputRegisters_258__7,inputRegisters_258__6,inputRegisters_258__5,
            inputRegisters_258__4,inputRegisters_258__3,inputRegisters_258__2,
            inputRegisters_258__1,inputRegisters_258__0})) ;
    Reg_16 loop1_258_x (.D ({inputRegisters_258__15,inputRegisters_258__14,
           inputRegisters_258__13,inputRegisters_258__12,inputRegisters_258__11,
           inputRegisters_258__10,inputRegisters_258__9,inputRegisters_258__8,
           inputRegisters_258__7,inputRegisters_258__6,inputRegisters_258__5,
           inputRegisters_258__4,inputRegisters_258__3,inputRegisters_258__2,
           inputRegisters_258__1,inputRegisters_258__0}), .en (
           enableRegister_258), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_258__15,registerOutputs_258__14,
           registerOutputs_258__13,registerOutputs_258__12,
           registerOutputs_258__11,registerOutputs_258__10,
           registerOutputs_258__9,registerOutputs_258__8,registerOutputs_258__7,
           registerOutputs_258__6,registerOutputs_258__5,registerOutputs_258__4,
           registerOutputs_258__3,registerOutputs_258__2,registerOutputs_258__1,
           registerOutputs_258__0})) ;
    Mux2_16 loop1_259_y (.A ({nx35959,nx36101,nx36243,nx36385,nx36527,nx36669,
            nx36811,nx36953,nx37095,nx37237,nx37379,nx37521,nx37663,nx37805,
            nx37947,nx38089}), .B ({nx33715,nx33853,nx33991,nx34129,nx34267,
            nx34405,nx34543,nx34685,nx34827,nx34969,nx35111,nx35253,nx35395,
            nx35537,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35679), .C ({inputRegisters_259__15,inputRegisters_259__14,
            inputRegisters_259__13,inputRegisters_259__12,inputRegisters_259__11
            ,inputRegisters_259__10,inputRegisters_259__9,inputRegisters_259__8,
            inputRegisters_259__7,inputRegisters_259__6,inputRegisters_259__5,
            inputRegisters_259__4,inputRegisters_259__3,inputRegisters_259__2,
            inputRegisters_259__1,inputRegisters_259__0})) ;
    Reg_16 loop1_259_x (.D ({inputRegisters_259__15,inputRegisters_259__14,
           inputRegisters_259__13,inputRegisters_259__12,inputRegisters_259__11,
           inputRegisters_259__10,inputRegisters_259__9,inputRegisters_259__8,
           inputRegisters_259__7,inputRegisters_259__6,inputRegisters_259__5,
           inputRegisters_259__4,inputRegisters_259__3,inputRegisters_259__2,
           inputRegisters_259__1,inputRegisters_259__0}), .en (
           enableRegister_259), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_259__15,registerOutputs_259__14,
           registerOutputs_259__13,registerOutputs_259__12,
           registerOutputs_259__11,registerOutputs_259__10,
           registerOutputs_259__9,registerOutputs_259__8,registerOutputs_259__7,
           registerOutputs_259__6,registerOutputs_259__5,registerOutputs_259__4,
           registerOutputs_259__3,registerOutputs_259__2,registerOutputs_259__1,
           registerOutputs_259__0})) ;
    Mux2_16 loop1_260_y (.A ({nx35959,nx36101,nx36243,nx36385,nx36527,nx36669,
            nx36811,nx36953,nx37095,nx37237,nx37379,nx37521,nx37663,nx37805,
            nx37947,nx38089}), .B ({nx33715,nx33853,nx33991,nx34129,nx34267,
            nx34405,nx34545,nx34685,nx34827,nx34969,nx35111,nx35253,nx35395,
            nx35537,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35679), .C ({inputRegisters_260__15,inputRegisters_260__14,
            inputRegisters_260__13,inputRegisters_260__12,inputRegisters_260__11
            ,inputRegisters_260__10,inputRegisters_260__9,inputRegisters_260__8,
            inputRegisters_260__7,inputRegisters_260__6,inputRegisters_260__5,
            inputRegisters_260__4,inputRegisters_260__3,inputRegisters_260__2,
            inputRegisters_260__1,inputRegisters_260__0})) ;
    Reg_16 loop1_260_x (.D ({inputRegisters_260__15,inputRegisters_260__14,
           inputRegisters_260__13,inputRegisters_260__12,inputRegisters_260__11,
           inputRegisters_260__10,inputRegisters_260__9,inputRegisters_260__8,
           inputRegisters_260__7,inputRegisters_260__6,inputRegisters_260__5,
           inputRegisters_260__4,inputRegisters_260__3,inputRegisters_260__2,
           inputRegisters_260__1,inputRegisters_260__0}), .en (
           enableRegister_260), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_260__15,registerOutputs_260__14,
           registerOutputs_260__13,registerOutputs_260__12,
           registerOutputs_260__11,registerOutputs_260__10,
           registerOutputs_260__9,registerOutputs_260__8,registerOutputs_260__7,
           registerOutputs_260__6,registerOutputs_260__5,registerOutputs_260__4,
           registerOutputs_260__3,registerOutputs_260__2,registerOutputs_260__1,
           registerOutputs_260__0})) ;
    Mux2_16 loop1_261_y (.A ({nx35959,nx36101,nx36243,nx36385,nx36527,nx36669,
            nx36811,nx36953,nx37095,nx37237,nx37379,nx37521,nx37663,nx37805,
            nx37947,nx38089}), .B ({nx33715,nx33853,nx33991,nx34129,nx34267,
            nx34407,nx34545,nx34685,nx34827,nx34969,nx35111,nx35253,nx35395,
            nx35537,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35679), .C ({inputRegisters_261__15,inputRegisters_261__14,
            inputRegisters_261__13,inputRegisters_261__12,inputRegisters_261__11
            ,inputRegisters_261__10,inputRegisters_261__9,inputRegisters_261__8,
            inputRegisters_261__7,inputRegisters_261__6,inputRegisters_261__5,
            inputRegisters_261__4,inputRegisters_261__3,inputRegisters_261__2,
            inputRegisters_261__1,inputRegisters_261__0})) ;
    Reg_16 loop1_261_x (.D ({inputRegisters_261__15,inputRegisters_261__14,
           inputRegisters_261__13,inputRegisters_261__12,inputRegisters_261__11,
           inputRegisters_261__10,inputRegisters_261__9,inputRegisters_261__8,
           inputRegisters_261__7,inputRegisters_261__6,inputRegisters_261__5,
           inputRegisters_261__4,inputRegisters_261__3,inputRegisters_261__2,
           inputRegisters_261__1,inputRegisters_261__0}), .en (
           enableRegister_261), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_261__15,registerOutputs_261__14,
           registerOutputs_261__13,registerOutputs_261__12,
           registerOutputs_261__11,registerOutputs_261__10,
           registerOutputs_261__9,registerOutputs_261__8,registerOutputs_261__7,
           registerOutputs_261__6,registerOutputs_261__5,registerOutputs_261__4,
           registerOutputs_261__3,registerOutputs_261__2,registerOutputs_261__1,
           registerOutputs_261__0})) ;
    Mux2_16 loop1_262_y (.A ({nx35959,nx36101,nx36243,nx36385,nx36527,nx36669,
            nx36811,nx36953,nx37095,nx37237,nx37379,nx37521,nx37663,nx37805,
            nx37947,nx38089}), .B ({nx33715,nx33853,nx33991,nx34129,nx34269,
            nx34407,nx34545,nx34685,nx34827,nx34969,nx35111,nx35253,nx35395,
            nx35537,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35679), .C ({inputRegisters_262__15,inputRegisters_262__14,
            inputRegisters_262__13,inputRegisters_262__12,inputRegisters_262__11
            ,inputRegisters_262__10,inputRegisters_262__9,inputRegisters_262__8,
            inputRegisters_262__7,inputRegisters_262__6,inputRegisters_262__5,
            inputRegisters_262__4,inputRegisters_262__3,inputRegisters_262__2,
            inputRegisters_262__1,inputRegisters_262__0})) ;
    Reg_16 loop1_262_x (.D ({inputRegisters_262__15,inputRegisters_262__14,
           inputRegisters_262__13,inputRegisters_262__12,inputRegisters_262__11,
           inputRegisters_262__10,inputRegisters_262__9,inputRegisters_262__8,
           inputRegisters_262__7,inputRegisters_262__6,inputRegisters_262__5,
           inputRegisters_262__4,inputRegisters_262__3,inputRegisters_262__2,
           inputRegisters_262__1,inputRegisters_262__0}), .en (
           enableRegister_262), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_262__15,registerOutputs_262__14,
           registerOutputs_262__13,registerOutputs_262__12,
           registerOutputs_262__11,registerOutputs_262__10,
           registerOutputs_262__9,registerOutputs_262__8,registerOutputs_262__7,
           registerOutputs_262__6,registerOutputs_262__5,registerOutputs_262__4,
           registerOutputs_262__3,registerOutputs_262__2,registerOutputs_262__1,
           registerOutputs_262__0})) ;
    Mux2_16 loop1_263_y (.A ({nx35959,nx36101,nx36243,nx36385,nx36527,nx36669,
            nx36811,nx36953,nx37095,nx37237,nx37379,nx37521,nx37663,nx37805,
            nx37947,nx38089}), .B ({nx33715,nx33853,nx33991,nx34131,nx34269,
            nx34407,nx34545,nx34685,nx34827,nx34969,nx35111,nx35253,nx35395,
            nx35537,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35679), .C ({inputRegisters_263__15,inputRegisters_263__14,
            inputRegisters_263__13,inputRegisters_263__12,inputRegisters_263__11
            ,inputRegisters_263__10,inputRegisters_263__9,inputRegisters_263__8,
            inputRegisters_263__7,inputRegisters_263__6,inputRegisters_263__5,
            inputRegisters_263__4,inputRegisters_263__3,inputRegisters_263__2,
            inputRegisters_263__1,inputRegisters_263__0})) ;
    Reg_16 loop1_263_x (.D ({inputRegisters_263__15,inputRegisters_263__14,
           inputRegisters_263__13,inputRegisters_263__12,inputRegisters_263__11,
           inputRegisters_263__10,inputRegisters_263__9,inputRegisters_263__8,
           inputRegisters_263__7,inputRegisters_263__6,inputRegisters_263__5,
           inputRegisters_263__4,inputRegisters_263__3,inputRegisters_263__2,
           inputRegisters_263__1,inputRegisters_263__0}), .en (
           enableRegister_263), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_263__15,registerOutputs_263__14,
           registerOutputs_263__13,registerOutputs_263__12,
           registerOutputs_263__11,registerOutputs_263__10,
           registerOutputs_263__9,registerOutputs_263__8,registerOutputs_263__7,
           registerOutputs_263__6,registerOutputs_263__5,registerOutputs_263__4,
           registerOutputs_263__3,registerOutputs_263__2,registerOutputs_263__1,
           registerOutputs_263__0})) ;
    Mux2_16 loop1_264_y (.A ({nx35959,nx36101,nx36243,nx36385,nx36527,nx36669,
            nx36811,nx36953,nx37095,nx37237,nx37379,nx37521,nx37663,nx37805,
            nx37947,nx38089}), .B ({nx33715,nx33853,nx33993,nx34131,nx34269,
            nx34407,nx34545,nx34685,nx34827,nx34969,nx35111,nx35253,nx35395,
            nx35537,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35679), .C ({inputRegisters_264__15,inputRegisters_264__14,
            inputRegisters_264__13,inputRegisters_264__12,inputRegisters_264__11
            ,inputRegisters_264__10,inputRegisters_264__9,inputRegisters_264__8,
            inputRegisters_264__7,inputRegisters_264__6,inputRegisters_264__5,
            inputRegisters_264__4,inputRegisters_264__3,inputRegisters_264__2,
            inputRegisters_264__1,inputRegisters_264__0})) ;
    Reg_16 loop1_264_x (.D ({inputRegisters_264__15,inputRegisters_264__14,
           inputRegisters_264__13,inputRegisters_264__12,inputRegisters_264__11,
           inputRegisters_264__10,inputRegisters_264__9,inputRegisters_264__8,
           inputRegisters_264__7,inputRegisters_264__6,inputRegisters_264__5,
           inputRegisters_264__4,inputRegisters_264__3,inputRegisters_264__2,
           inputRegisters_264__1,inputRegisters_264__0}), .en (
           enableRegister_264), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_264__15,registerOutputs_264__14,
           registerOutputs_264__13,registerOutputs_264__12,
           registerOutputs_264__11,registerOutputs_264__10,
           registerOutputs_264__9,registerOutputs_264__8,registerOutputs_264__7,
           registerOutputs_264__6,registerOutputs_264__5,registerOutputs_264__4,
           registerOutputs_264__3,registerOutputs_264__2,registerOutputs_264__1,
           registerOutputs_264__0})) ;
    Mux2_16 loop1_265_y (.A ({nx35959,nx36101,nx36243,nx36385,nx36527,nx36669,
            nx36811,nx36953,nx37095,nx37237,nx37379,nx37521,nx37663,nx37805,
            nx37947,nx38089}), .B ({nx33715,nx33855,nx33993,nx34131,nx34269,
            nx34407,nx34545,nx34685,nx34827,nx34969,nx35111,nx35253,nx35395,
            nx35537,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35679), .C ({inputRegisters_265__15,inputRegisters_265__14,
            inputRegisters_265__13,inputRegisters_265__12,inputRegisters_265__11
            ,inputRegisters_265__10,inputRegisters_265__9,inputRegisters_265__8,
            inputRegisters_265__7,inputRegisters_265__6,inputRegisters_265__5,
            inputRegisters_265__4,inputRegisters_265__3,inputRegisters_265__2,
            inputRegisters_265__1,inputRegisters_265__0})) ;
    Reg_16 loop1_265_x (.D ({inputRegisters_265__15,inputRegisters_265__14,
           inputRegisters_265__13,inputRegisters_265__12,inputRegisters_265__11,
           inputRegisters_265__10,inputRegisters_265__9,inputRegisters_265__8,
           inputRegisters_265__7,inputRegisters_265__6,inputRegisters_265__5,
           inputRegisters_265__4,inputRegisters_265__3,inputRegisters_265__2,
           inputRegisters_265__1,inputRegisters_265__0}), .en (
           enableRegister_265), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_265__15,registerOutputs_265__14,
           registerOutputs_265__13,registerOutputs_265__12,
           registerOutputs_265__11,registerOutputs_265__10,
           registerOutputs_265__9,registerOutputs_265__8,registerOutputs_265__7,
           registerOutputs_265__6,registerOutputs_265__5,registerOutputs_265__4,
           registerOutputs_265__3,registerOutputs_265__2,registerOutputs_265__1,
           registerOutputs_265__0})) ;
    Mux2_16 loop1_266_y (.A ({nx35961,nx36103,nx36245,nx36387,nx36529,nx36671,
            nx36813,nx36955,nx37097,nx37239,nx37381,nx37523,nx37665,nx37807,
            nx37949,nx38091}), .B ({nx33717,nx33855,nx33993,nx34131,nx34269,
            nx34407,nx34545,nx34687,nx34829,nx34971,nx35113,nx35255,nx35397,
            nx35539,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35681), .C ({inputRegisters_266__15,inputRegisters_266__14,
            inputRegisters_266__13,inputRegisters_266__12,inputRegisters_266__11
            ,inputRegisters_266__10,inputRegisters_266__9,inputRegisters_266__8,
            inputRegisters_266__7,inputRegisters_266__6,inputRegisters_266__5,
            inputRegisters_266__4,inputRegisters_266__3,inputRegisters_266__2,
            inputRegisters_266__1,inputRegisters_266__0})) ;
    Reg_16 loop1_266_x (.D ({inputRegisters_266__15,inputRegisters_266__14,
           inputRegisters_266__13,inputRegisters_266__12,inputRegisters_266__11,
           inputRegisters_266__10,inputRegisters_266__9,inputRegisters_266__8,
           inputRegisters_266__7,inputRegisters_266__6,inputRegisters_266__5,
           inputRegisters_266__4,inputRegisters_266__3,inputRegisters_266__2,
           inputRegisters_266__1,inputRegisters_266__0}), .en (
           enableRegister_266), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_266__15,registerOutputs_266__14,
           registerOutputs_266__13,registerOutputs_266__12,
           registerOutputs_266__11,registerOutputs_266__10,
           registerOutputs_266__9,registerOutputs_266__8,registerOutputs_266__7,
           registerOutputs_266__6,registerOutputs_266__5,registerOutputs_266__4,
           registerOutputs_266__3,registerOutputs_266__2,registerOutputs_266__1,
           registerOutputs_266__0})) ;
    Mux2_16 loop1_267_y (.A ({nx35961,nx36103,nx36245,nx36387,nx36529,nx36671,
            nx36813,nx36955,nx37097,nx37239,nx37381,nx37523,nx37665,nx37807,
            nx37949,nx38091}), .B ({nx33717,nx33855,nx33993,nx34131,nx34269,
            nx34407,nx34547,nx34687,nx34829,nx34971,nx35113,nx35255,nx35397,
            nx35539,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35681), .C ({inputRegisters_267__15,inputRegisters_267__14,
            inputRegisters_267__13,inputRegisters_267__12,inputRegisters_267__11
            ,inputRegisters_267__10,inputRegisters_267__9,inputRegisters_267__8,
            inputRegisters_267__7,inputRegisters_267__6,inputRegisters_267__5,
            inputRegisters_267__4,inputRegisters_267__3,inputRegisters_267__2,
            inputRegisters_267__1,inputRegisters_267__0})) ;
    Reg_16 loop1_267_x (.D ({inputRegisters_267__15,inputRegisters_267__14,
           inputRegisters_267__13,inputRegisters_267__12,inputRegisters_267__11,
           inputRegisters_267__10,inputRegisters_267__9,inputRegisters_267__8,
           inputRegisters_267__7,inputRegisters_267__6,inputRegisters_267__5,
           inputRegisters_267__4,inputRegisters_267__3,inputRegisters_267__2,
           inputRegisters_267__1,inputRegisters_267__0}), .en (
           enableRegister_267), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_267__15,registerOutputs_267__14,
           registerOutputs_267__13,registerOutputs_267__12,
           registerOutputs_267__11,registerOutputs_267__10,
           registerOutputs_267__9,registerOutputs_267__8,registerOutputs_267__7,
           registerOutputs_267__6,registerOutputs_267__5,registerOutputs_267__4,
           registerOutputs_267__3,registerOutputs_267__2,registerOutputs_267__1,
           registerOutputs_267__0})) ;
    Mux2_16 loop1_268_y (.A ({nx35961,nx36103,nx36245,nx36387,nx36529,nx36671,
            nx36813,nx36955,nx37097,nx37239,nx37381,nx37523,nx37665,nx37807,
            nx37949,nx38091}), .B ({nx33717,nx33855,nx33993,nx34131,nx34269,
            nx34409,nx34547,nx34687,nx34829,nx34971,nx35113,nx35255,nx35397,
            nx35539,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35681), .C ({inputRegisters_268__15,inputRegisters_268__14,
            inputRegisters_268__13,inputRegisters_268__12,inputRegisters_268__11
            ,inputRegisters_268__10,inputRegisters_268__9,inputRegisters_268__8,
            inputRegisters_268__7,inputRegisters_268__6,inputRegisters_268__5,
            inputRegisters_268__4,inputRegisters_268__3,inputRegisters_268__2,
            inputRegisters_268__1,inputRegisters_268__0})) ;
    Reg_16 loop1_268_x (.D ({inputRegisters_268__15,inputRegisters_268__14,
           inputRegisters_268__13,inputRegisters_268__12,inputRegisters_268__11,
           inputRegisters_268__10,inputRegisters_268__9,inputRegisters_268__8,
           inputRegisters_268__7,inputRegisters_268__6,inputRegisters_268__5,
           inputRegisters_268__4,inputRegisters_268__3,inputRegisters_268__2,
           inputRegisters_268__1,inputRegisters_268__0}), .en (
           enableRegister_268), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_268__15,registerOutputs_268__14,
           registerOutputs_268__13,registerOutputs_268__12,
           registerOutputs_268__11,registerOutputs_268__10,
           registerOutputs_268__9,registerOutputs_268__8,registerOutputs_268__7,
           registerOutputs_268__6,registerOutputs_268__5,registerOutputs_268__4,
           registerOutputs_268__3,registerOutputs_268__2,registerOutputs_268__1,
           registerOutputs_268__0})) ;
    Mux2_16 loop1_269_y (.A ({nx35961,nx36103,nx36245,nx36387,nx36529,nx36671,
            nx36813,nx36955,nx37097,nx37239,nx37381,nx37523,nx37665,nx37807,
            nx37949,nx38091}), .B ({nx33717,nx33855,nx33993,nx34131,nx34271,
            nx34409,nx34547,nx34687,nx34829,nx34971,nx35113,nx35255,nx35397,
            nx35539,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35681), .C ({inputRegisters_269__15,inputRegisters_269__14,
            inputRegisters_269__13,inputRegisters_269__12,inputRegisters_269__11
            ,inputRegisters_269__10,inputRegisters_269__9,inputRegisters_269__8,
            inputRegisters_269__7,inputRegisters_269__6,inputRegisters_269__5,
            inputRegisters_269__4,inputRegisters_269__3,inputRegisters_269__2,
            inputRegisters_269__1,inputRegisters_269__0})) ;
    Reg_16 loop1_269_x (.D ({inputRegisters_269__15,inputRegisters_269__14,
           inputRegisters_269__13,inputRegisters_269__12,inputRegisters_269__11,
           inputRegisters_269__10,inputRegisters_269__9,inputRegisters_269__8,
           inputRegisters_269__7,inputRegisters_269__6,inputRegisters_269__5,
           inputRegisters_269__4,inputRegisters_269__3,inputRegisters_269__2,
           inputRegisters_269__1,inputRegisters_269__0}), .en (
           enableRegister_269), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_269__15,registerOutputs_269__14,
           registerOutputs_269__13,registerOutputs_269__12,
           registerOutputs_269__11,registerOutputs_269__10,
           registerOutputs_269__9,registerOutputs_269__8,registerOutputs_269__7,
           registerOutputs_269__6,registerOutputs_269__5,registerOutputs_269__4,
           registerOutputs_269__3,registerOutputs_269__2,registerOutputs_269__1,
           registerOutputs_269__0})) ;
    Mux2_16 loop1_270_y (.A ({nx35961,nx36103,nx36245,nx36387,nx36529,nx36671,
            nx36813,nx36955,nx37097,nx37239,nx37381,nx37523,nx37665,nx37807,
            nx37949,nx38091}), .B ({nx33717,nx33855,nx33993,nx34133,nx34271,
            nx34409,nx34547,nx34687,nx34829,nx34971,nx35113,nx35255,nx35397,
            nx35539,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35681), .C ({inputRegisters_270__15,inputRegisters_270__14,
            inputRegisters_270__13,inputRegisters_270__12,inputRegisters_270__11
            ,inputRegisters_270__10,inputRegisters_270__9,inputRegisters_270__8,
            inputRegisters_270__7,inputRegisters_270__6,inputRegisters_270__5,
            inputRegisters_270__4,inputRegisters_270__3,inputRegisters_270__2,
            inputRegisters_270__1,inputRegisters_270__0})) ;
    Reg_16 loop1_270_x (.D ({inputRegisters_270__15,inputRegisters_270__14,
           inputRegisters_270__13,inputRegisters_270__12,inputRegisters_270__11,
           inputRegisters_270__10,inputRegisters_270__9,inputRegisters_270__8,
           inputRegisters_270__7,inputRegisters_270__6,inputRegisters_270__5,
           inputRegisters_270__4,inputRegisters_270__3,inputRegisters_270__2,
           inputRegisters_270__1,inputRegisters_270__0}), .en (
           enableRegister_270), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_270__15,registerOutputs_270__14,
           registerOutputs_270__13,registerOutputs_270__12,
           registerOutputs_270__11,registerOutputs_270__10,
           registerOutputs_270__9,registerOutputs_270__8,registerOutputs_270__7,
           registerOutputs_270__6,registerOutputs_270__5,registerOutputs_270__4,
           registerOutputs_270__3,registerOutputs_270__2,registerOutputs_270__1,
           registerOutputs_270__0})) ;
    Mux2_16 loop1_271_y (.A ({nx35961,nx36103,nx36245,nx36387,nx36529,nx36671,
            nx36813,nx36955,nx37097,nx37239,nx37381,nx37523,nx37665,nx37807,
            nx37949,nx38091}), .B ({nx33717,nx33855,nx33995,nx34133,nx34271,
            nx34409,nx34547,nx34687,nx34829,nx34971,nx35113,nx35255,nx35397,
            nx35539,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35681), .C ({inputRegisters_271__15,inputRegisters_271__14,
            inputRegisters_271__13,inputRegisters_271__12,inputRegisters_271__11
            ,inputRegisters_271__10,inputRegisters_271__9,inputRegisters_271__8,
            inputRegisters_271__7,inputRegisters_271__6,inputRegisters_271__5,
            inputRegisters_271__4,inputRegisters_271__3,inputRegisters_271__2,
            inputRegisters_271__1,inputRegisters_271__0})) ;
    Reg_16 loop1_271_x (.D ({inputRegisters_271__15,inputRegisters_271__14,
           inputRegisters_271__13,inputRegisters_271__12,inputRegisters_271__11,
           inputRegisters_271__10,inputRegisters_271__9,inputRegisters_271__8,
           inputRegisters_271__7,inputRegisters_271__6,inputRegisters_271__5,
           inputRegisters_271__4,inputRegisters_271__3,inputRegisters_271__2,
           inputRegisters_271__1,inputRegisters_271__0}), .en (
           enableRegister_271), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_271__15,registerOutputs_271__14,
           registerOutputs_271__13,registerOutputs_271__12,
           registerOutputs_271__11,registerOutputs_271__10,
           registerOutputs_271__9,registerOutputs_271__8,registerOutputs_271__7,
           registerOutputs_271__6,registerOutputs_271__5,registerOutputs_271__4,
           registerOutputs_271__3,registerOutputs_271__2,registerOutputs_271__1,
           registerOutputs_271__0})) ;
    Mux2_16 loop1_272_y (.A ({nx35961,nx36103,nx36245,nx36387,nx36529,nx36671,
            nx36813,nx36955,nx37097,nx37239,nx37381,nx37523,nx37665,nx37807,
            nx37949,nx38091}), .B ({nx33717,nx33857,nx33995,nx34133,nx34271,
            nx34409,nx34547,nx34687,nx34829,nx34971,nx35113,nx35255,nx35397,
            nx35539,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35681), .C ({inputRegisters_272__15,inputRegisters_272__14,
            inputRegisters_272__13,inputRegisters_272__12,inputRegisters_272__11
            ,inputRegisters_272__10,inputRegisters_272__9,inputRegisters_272__8,
            inputRegisters_272__7,inputRegisters_272__6,inputRegisters_272__5,
            inputRegisters_272__4,inputRegisters_272__3,inputRegisters_272__2,
            inputRegisters_272__1,inputRegisters_272__0})) ;
    Reg_16 loop1_272_x (.D ({inputRegisters_272__15,inputRegisters_272__14,
           inputRegisters_272__13,inputRegisters_272__12,inputRegisters_272__11,
           inputRegisters_272__10,inputRegisters_272__9,inputRegisters_272__8,
           inputRegisters_272__7,inputRegisters_272__6,inputRegisters_272__5,
           inputRegisters_272__4,inputRegisters_272__3,inputRegisters_272__2,
           inputRegisters_272__1,inputRegisters_272__0}), .en (
           enableRegister_272), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_272__15,registerOutputs_272__14,
           registerOutputs_272__13,registerOutputs_272__12,
           registerOutputs_272__11,registerOutputs_272__10,
           registerOutputs_272__9,registerOutputs_272__8,registerOutputs_272__7,
           registerOutputs_272__6,registerOutputs_272__5,registerOutputs_272__4,
           registerOutputs_272__3,registerOutputs_272__2,registerOutputs_272__1,
           registerOutputs_272__0})) ;
    Mux2_16 loop1_273_y (.A ({nx35963,nx36105,nx36247,nx36389,nx36531,nx36673,
            nx36815,nx36957,nx37099,nx37241,nx37383,nx37525,nx37667,nx37809,
            nx37951,nx38093}), .B ({nx33719,nx33857,nx33995,nx34133,nx34271,
            nx34409,nx34547,nx34689,nx34831,nx34973,nx35115,nx35257,nx35399,
            nx35541,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35683), .C ({inputRegisters_273__15,inputRegisters_273__14,
            inputRegisters_273__13,inputRegisters_273__12,inputRegisters_273__11
            ,inputRegisters_273__10,inputRegisters_273__9,inputRegisters_273__8,
            inputRegisters_273__7,inputRegisters_273__6,inputRegisters_273__5,
            inputRegisters_273__4,inputRegisters_273__3,inputRegisters_273__2,
            inputRegisters_273__1,inputRegisters_273__0})) ;
    Reg_16 loop1_273_x (.D ({inputRegisters_273__15,inputRegisters_273__14,
           inputRegisters_273__13,inputRegisters_273__12,inputRegisters_273__11,
           inputRegisters_273__10,inputRegisters_273__9,inputRegisters_273__8,
           inputRegisters_273__7,inputRegisters_273__6,inputRegisters_273__5,
           inputRegisters_273__4,inputRegisters_273__3,inputRegisters_273__2,
           inputRegisters_273__1,inputRegisters_273__0}), .en (
           enableRegister_273), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_273__15,registerOutputs_273__14,
           registerOutputs_273__13,registerOutputs_273__12,
           registerOutputs_273__11,registerOutputs_273__10,
           registerOutputs_273__9,registerOutputs_273__8,registerOutputs_273__7,
           registerOutputs_273__6,registerOutputs_273__5,registerOutputs_273__4,
           registerOutputs_273__3,registerOutputs_273__2,registerOutputs_273__1,
           registerOutputs_273__0})) ;
    Mux2_16 loop1_274_y (.A ({nx35963,nx36105,nx36247,nx36389,nx36531,nx36673,
            nx36815,nx36957,nx37099,nx37241,nx37383,nx37525,nx37667,nx37809,
            nx37951,nx38093}), .B ({nx33719,nx33857,nx33995,nx34133,nx34271,
            nx34409,nx34549,nx34689,nx34831,nx34973,nx35115,nx35257,nx35399,
            nx35541,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35683), .C ({inputRegisters_274__15,inputRegisters_274__14,
            inputRegisters_274__13,inputRegisters_274__12,inputRegisters_274__11
            ,inputRegisters_274__10,inputRegisters_274__9,inputRegisters_274__8,
            inputRegisters_274__7,inputRegisters_274__6,inputRegisters_274__5,
            inputRegisters_274__4,inputRegisters_274__3,inputRegisters_274__2,
            inputRegisters_274__1,inputRegisters_274__0})) ;
    Reg_16 loop1_274_x (.D ({inputRegisters_274__15,inputRegisters_274__14,
           inputRegisters_274__13,inputRegisters_274__12,inputRegisters_274__11,
           inputRegisters_274__10,inputRegisters_274__9,inputRegisters_274__8,
           inputRegisters_274__7,inputRegisters_274__6,inputRegisters_274__5,
           inputRegisters_274__4,inputRegisters_274__3,inputRegisters_274__2,
           inputRegisters_274__1,inputRegisters_274__0}), .en (
           enableRegister_274), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_274__15,registerOutputs_274__14,
           registerOutputs_274__13,registerOutputs_274__12,
           registerOutputs_274__11,registerOutputs_274__10,
           registerOutputs_274__9,registerOutputs_274__8,registerOutputs_274__7,
           registerOutputs_274__6,registerOutputs_274__5,registerOutputs_274__4,
           registerOutputs_274__3,registerOutputs_274__2,registerOutputs_274__1,
           registerOutputs_274__0})) ;
    Mux2_16 loop1_275_y (.A ({nx35963,nx36105,nx36247,nx36389,nx36531,nx36673,
            nx36815,nx36957,nx37099,nx37241,nx37383,nx37525,nx37667,nx37809,
            nx37951,nx38093}), .B ({nx33719,nx33857,nx33995,nx34133,nx34271,
            nx34411,nx34549,nx34689,nx34831,nx34973,nx35115,nx35257,nx35399,
            nx35541,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35683), .C ({inputRegisters_275__15,inputRegisters_275__14,
            inputRegisters_275__13,inputRegisters_275__12,inputRegisters_275__11
            ,inputRegisters_275__10,inputRegisters_275__9,inputRegisters_275__8,
            inputRegisters_275__7,inputRegisters_275__6,inputRegisters_275__5,
            inputRegisters_275__4,inputRegisters_275__3,inputRegisters_275__2,
            inputRegisters_275__1,inputRegisters_275__0})) ;
    Reg_16 loop1_275_x (.D ({inputRegisters_275__15,inputRegisters_275__14,
           inputRegisters_275__13,inputRegisters_275__12,inputRegisters_275__11,
           inputRegisters_275__10,inputRegisters_275__9,inputRegisters_275__8,
           inputRegisters_275__7,inputRegisters_275__6,inputRegisters_275__5,
           inputRegisters_275__4,inputRegisters_275__3,inputRegisters_275__2,
           inputRegisters_275__1,inputRegisters_275__0}), .en (
           enableRegister_275), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_275__15,registerOutputs_275__14,
           registerOutputs_275__13,registerOutputs_275__12,
           registerOutputs_275__11,registerOutputs_275__10,
           registerOutputs_275__9,registerOutputs_275__8,registerOutputs_275__7,
           registerOutputs_275__6,registerOutputs_275__5,registerOutputs_275__4,
           registerOutputs_275__3,registerOutputs_275__2,registerOutputs_275__1,
           registerOutputs_275__0})) ;
    Mux2_16 loop1_276_y (.A ({nx35963,nx36105,nx36247,nx36389,nx36531,nx36673,
            nx36815,nx36957,nx37099,nx37241,nx37383,nx37525,nx37667,nx37809,
            nx37951,nx38093}), .B ({nx33719,nx33857,nx33995,nx34133,nx34273,
            nx34411,nx34549,nx34689,nx34831,nx34973,nx35115,nx35257,nx35399,
            nx35541,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35683), .C ({inputRegisters_276__15,inputRegisters_276__14,
            inputRegisters_276__13,inputRegisters_276__12,inputRegisters_276__11
            ,inputRegisters_276__10,inputRegisters_276__9,inputRegisters_276__8,
            inputRegisters_276__7,inputRegisters_276__6,inputRegisters_276__5,
            inputRegisters_276__4,inputRegisters_276__3,inputRegisters_276__2,
            inputRegisters_276__1,inputRegisters_276__0})) ;
    Reg_16 loop1_276_x (.D ({inputRegisters_276__15,inputRegisters_276__14,
           inputRegisters_276__13,inputRegisters_276__12,inputRegisters_276__11,
           inputRegisters_276__10,inputRegisters_276__9,inputRegisters_276__8,
           inputRegisters_276__7,inputRegisters_276__6,inputRegisters_276__5,
           inputRegisters_276__4,inputRegisters_276__3,inputRegisters_276__2,
           inputRegisters_276__1,inputRegisters_276__0}), .en (
           enableRegister_276), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_276__15,registerOutputs_276__14,
           registerOutputs_276__13,registerOutputs_276__12,
           registerOutputs_276__11,registerOutputs_276__10,
           registerOutputs_276__9,registerOutputs_276__8,registerOutputs_276__7,
           registerOutputs_276__6,registerOutputs_276__5,registerOutputs_276__4,
           registerOutputs_276__3,registerOutputs_276__2,registerOutputs_276__1,
           registerOutputs_276__0})) ;
    Mux2_16 loop1_277_y (.A ({nx35963,nx36105,nx36247,nx36389,nx36531,nx36673,
            nx36815,nx36957,nx37099,nx37241,nx37383,nx37525,nx37667,nx37809,
            nx37951,nx38093}), .B ({nx33719,nx33857,nx33995,nx34135,nx34273,
            nx34411,nx34549,nx34689,nx34831,nx34973,nx35115,nx35257,nx35399,
            nx35541,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35683), .C ({inputRegisters_277__15,inputRegisters_277__14,
            inputRegisters_277__13,inputRegisters_277__12,inputRegisters_277__11
            ,inputRegisters_277__10,inputRegisters_277__9,inputRegisters_277__8,
            inputRegisters_277__7,inputRegisters_277__6,inputRegisters_277__5,
            inputRegisters_277__4,inputRegisters_277__3,inputRegisters_277__2,
            inputRegisters_277__1,inputRegisters_277__0})) ;
    Reg_16 loop1_277_x (.D ({inputRegisters_277__15,inputRegisters_277__14,
           inputRegisters_277__13,inputRegisters_277__12,inputRegisters_277__11,
           inputRegisters_277__10,inputRegisters_277__9,inputRegisters_277__8,
           inputRegisters_277__7,inputRegisters_277__6,inputRegisters_277__5,
           inputRegisters_277__4,inputRegisters_277__3,inputRegisters_277__2,
           inputRegisters_277__1,inputRegisters_277__0}), .en (
           enableRegister_277), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_277__15,registerOutputs_277__14,
           registerOutputs_277__13,registerOutputs_277__12,
           registerOutputs_277__11,registerOutputs_277__10,
           registerOutputs_277__9,registerOutputs_277__8,registerOutputs_277__7,
           registerOutputs_277__6,registerOutputs_277__5,registerOutputs_277__4,
           registerOutputs_277__3,registerOutputs_277__2,registerOutputs_277__1,
           registerOutputs_277__0})) ;
    Mux2_16 loop1_278_y (.A ({nx35963,nx36105,nx36247,nx36389,nx36531,nx36673,
            nx36815,nx36957,nx37099,nx37241,nx37383,nx37525,nx37667,nx37809,
            nx37951,nx38093}), .B ({nx33719,nx33857,nx33997,nx34135,nx34273,
            nx34411,nx34549,nx34689,nx34831,nx34973,nx35115,nx35257,nx35399,
            nx35541,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35683), .C ({inputRegisters_278__15,inputRegisters_278__14,
            inputRegisters_278__13,inputRegisters_278__12,inputRegisters_278__11
            ,inputRegisters_278__10,inputRegisters_278__9,inputRegisters_278__8,
            inputRegisters_278__7,inputRegisters_278__6,inputRegisters_278__5,
            inputRegisters_278__4,inputRegisters_278__3,inputRegisters_278__2,
            inputRegisters_278__1,inputRegisters_278__0})) ;
    Reg_16 loop1_278_x (.D ({inputRegisters_278__15,inputRegisters_278__14,
           inputRegisters_278__13,inputRegisters_278__12,inputRegisters_278__11,
           inputRegisters_278__10,inputRegisters_278__9,inputRegisters_278__8,
           inputRegisters_278__7,inputRegisters_278__6,inputRegisters_278__5,
           inputRegisters_278__4,inputRegisters_278__3,inputRegisters_278__2,
           inputRegisters_278__1,inputRegisters_278__0}), .en (
           enableRegister_278), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_278__15,registerOutputs_278__14,
           registerOutputs_278__13,registerOutputs_278__12,
           registerOutputs_278__11,registerOutputs_278__10,
           registerOutputs_278__9,registerOutputs_278__8,registerOutputs_278__7,
           registerOutputs_278__6,registerOutputs_278__5,registerOutputs_278__4,
           registerOutputs_278__3,registerOutputs_278__2,registerOutputs_278__1,
           registerOutputs_278__0})) ;
    Mux2_16 loop1_279_y (.A ({nx35963,nx36105,nx36247,nx36389,nx36531,nx36673,
            nx36815,nx36957,nx37099,nx37241,nx37383,nx37525,nx37667,nx37809,
            nx37951,nx38093}), .B ({nx33719,nx33859,nx33997,nx34135,nx34273,
            nx34411,nx34549,nx34689,nx34831,nx34973,nx35115,nx35257,nx35399,
            nx35541,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35683), .C ({inputRegisters_279__15,inputRegisters_279__14,
            inputRegisters_279__13,inputRegisters_279__12,inputRegisters_279__11
            ,inputRegisters_279__10,inputRegisters_279__9,inputRegisters_279__8,
            inputRegisters_279__7,inputRegisters_279__6,inputRegisters_279__5,
            inputRegisters_279__4,inputRegisters_279__3,inputRegisters_279__2,
            inputRegisters_279__1,inputRegisters_279__0})) ;
    Reg_16 loop1_279_x (.D ({inputRegisters_279__15,inputRegisters_279__14,
           inputRegisters_279__13,inputRegisters_279__12,inputRegisters_279__11,
           inputRegisters_279__10,inputRegisters_279__9,inputRegisters_279__8,
           inputRegisters_279__7,inputRegisters_279__6,inputRegisters_279__5,
           inputRegisters_279__4,inputRegisters_279__3,inputRegisters_279__2,
           inputRegisters_279__1,inputRegisters_279__0}), .en (
           enableRegister_279), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_279__15,registerOutputs_279__14,
           registerOutputs_279__13,registerOutputs_279__12,
           registerOutputs_279__11,registerOutputs_279__10,
           registerOutputs_279__9,registerOutputs_279__8,registerOutputs_279__7,
           registerOutputs_279__6,registerOutputs_279__5,registerOutputs_279__4,
           registerOutputs_279__3,registerOutputs_279__2,registerOutputs_279__1,
           registerOutputs_279__0})) ;
    Mux2_16 loop1_280_y (.A ({nx35965,nx36107,nx36249,nx36391,nx36533,nx36675,
            nx36817,nx36959,nx37101,nx37243,nx37385,nx37527,nx37669,nx37811,
            nx37953,nx38095}), .B ({nx33721,nx33859,nx33997,nx34135,nx34273,
            nx34411,nx34549,nx34691,nx34833,nx34975,nx35117,nx35259,nx35401,
            nx35543,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35685), .C ({inputRegisters_280__15,inputRegisters_280__14,
            inputRegisters_280__13,inputRegisters_280__12,inputRegisters_280__11
            ,inputRegisters_280__10,inputRegisters_280__9,inputRegisters_280__8,
            inputRegisters_280__7,inputRegisters_280__6,inputRegisters_280__5,
            inputRegisters_280__4,inputRegisters_280__3,inputRegisters_280__2,
            inputRegisters_280__1,inputRegisters_280__0})) ;
    Reg_16 loop1_280_x (.D ({inputRegisters_280__15,inputRegisters_280__14,
           inputRegisters_280__13,inputRegisters_280__12,inputRegisters_280__11,
           inputRegisters_280__10,inputRegisters_280__9,inputRegisters_280__8,
           inputRegisters_280__7,inputRegisters_280__6,inputRegisters_280__5,
           inputRegisters_280__4,inputRegisters_280__3,inputRegisters_280__2,
           inputRegisters_280__1,inputRegisters_280__0}), .en (
           enableRegister_280), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_280__15,registerOutputs_280__14,
           registerOutputs_280__13,registerOutputs_280__12,
           registerOutputs_280__11,registerOutputs_280__10,
           registerOutputs_280__9,registerOutputs_280__8,registerOutputs_280__7,
           registerOutputs_280__6,registerOutputs_280__5,registerOutputs_280__4,
           registerOutputs_280__3,registerOutputs_280__2,registerOutputs_280__1,
           registerOutputs_280__0})) ;
    Mux2_16 loop1_281_y (.A ({nx35965,nx36107,nx36249,nx36391,nx36533,nx36675,
            nx36817,nx36959,nx37101,nx37243,nx37385,nx37527,nx37669,nx37811,
            nx37953,nx38095}), .B ({nx33721,nx33859,nx33997,nx34135,nx34273,
            nx34411,nx34551,nx34691,nx34833,nx34975,nx35117,nx35259,nx35401,
            nx35543,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35685), .C ({inputRegisters_281__15,inputRegisters_281__14,
            inputRegisters_281__13,inputRegisters_281__12,inputRegisters_281__11
            ,inputRegisters_281__10,inputRegisters_281__9,inputRegisters_281__8,
            inputRegisters_281__7,inputRegisters_281__6,inputRegisters_281__5,
            inputRegisters_281__4,inputRegisters_281__3,inputRegisters_281__2,
            inputRegisters_281__1,inputRegisters_281__0})) ;
    Reg_16 loop1_281_x (.D ({inputRegisters_281__15,inputRegisters_281__14,
           inputRegisters_281__13,inputRegisters_281__12,inputRegisters_281__11,
           inputRegisters_281__10,inputRegisters_281__9,inputRegisters_281__8,
           inputRegisters_281__7,inputRegisters_281__6,inputRegisters_281__5,
           inputRegisters_281__4,inputRegisters_281__3,inputRegisters_281__2,
           inputRegisters_281__1,inputRegisters_281__0}), .en (
           enableRegister_281), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_281__15,registerOutputs_281__14,
           registerOutputs_281__13,registerOutputs_281__12,
           registerOutputs_281__11,registerOutputs_281__10,
           registerOutputs_281__9,registerOutputs_281__8,registerOutputs_281__7,
           registerOutputs_281__6,registerOutputs_281__5,registerOutputs_281__4,
           registerOutputs_281__3,registerOutputs_281__2,registerOutputs_281__1,
           registerOutputs_281__0})) ;
    Mux2_16 loop1_282_y (.A ({nx35965,nx36107,nx36249,nx36391,nx36533,nx36675,
            nx36817,nx36959,nx37101,nx37243,nx37385,nx37527,nx37669,nx37811,
            nx37953,nx38095}), .B ({nx33721,nx33859,nx33997,nx34135,nx34273,
            nx34413,nx34551,nx34691,nx34833,nx34975,nx35117,nx35259,nx35401,
            nx35543,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35685), .C ({inputRegisters_282__15,inputRegisters_282__14,
            inputRegisters_282__13,inputRegisters_282__12,inputRegisters_282__11
            ,inputRegisters_282__10,inputRegisters_282__9,inputRegisters_282__8,
            inputRegisters_282__7,inputRegisters_282__6,inputRegisters_282__5,
            inputRegisters_282__4,inputRegisters_282__3,inputRegisters_282__2,
            inputRegisters_282__1,inputRegisters_282__0})) ;
    Reg_16 loop1_282_x (.D ({inputRegisters_282__15,inputRegisters_282__14,
           inputRegisters_282__13,inputRegisters_282__12,inputRegisters_282__11,
           inputRegisters_282__10,inputRegisters_282__9,inputRegisters_282__8,
           inputRegisters_282__7,inputRegisters_282__6,inputRegisters_282__5,
           inputRegisters_282__4,inputRegisters_282__3,inputRegisters_282__2,
           inputRegisters_282__1,inputRegisters_282__0}), .en (
           enableRegister_282), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_282__15,registerOutputs_282__14,
           registerOutputs_282__13,registerOutputs_282__12,
           registerOutputs_282__11,registerOutputs_282__10,
           registerOutputs_282__9,registerOutputs_282__8,registerOutputs_282__7,
           registerOutputs_282__6,registerOutputs_282__5,registerOutputs_282__4,
           registerOutputs_282__3,registerOutputs_282__2,registerOutputs_282__1,
           registerOutputs_282__0})) ;
    Mux2_16 loop1_283_y (.A ({nx35965,nx36107,nx36249,nx36391,nx36533,nx36675,
            nx36817,nx36959,nx37101,nx37243,nx37385,nx37527,nx37669,nx37811,
            nx37953,nx38095}), .B ({nx33721,nx33859,nx33997,nx34135,nx34275,
            nx34413,nx34551,nx34691,nx34833,nx34975,nx35117,nx35259,nx35401,
            nx35543,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35685), .C ({inputRegisters_283__15,inputRegisters_283__14,
            inputRegisters_283__13,inputRegisters_283__12,inputRegisters_283__11
            ,inputRegisters_283__10,inputRegisters_283__9,inputRegisters_283__8,
            inputRegisters_283__7,inputRegisters_283__6,inputRegisters_283__5,
            inputRegisters_283__4,inputRegisters_283__3,inputRegisters_283__2,
            inputRegisters_283__1,inputRegisters_283__0})) ;
    Reg_16 loop1_283_x (.D ({inputRegisters_283__15,inputRegisters_283__14,
           inputRegisters_283__13,inputRegisters_283__12,inputRegisters_283__11,
           inputRegisters_283__10,inputRegisters_283__9,inputRegisters_283__8,
           inputRegisters_283__7,inputRegisters_283__6,inputRegisters_283__5,
           inputRegisters_283__4,inputRegisters_283__3,inputRegisters_283__2,
           inputRegisters_283__1,inputRegisters_283__0}), .en (
           enableRegister_283), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_283__15,registerOutputs_283__14,
           registerOutputs_283__13,registerOutputs_283__12,
           registerOutputs_283__11,registerOutputs_283__10,
           registerOutputs_283__9,registerOutputs_283__8,registerOutputs_283__7,
           registerOutputs_283__6,registerOutputs_283__5,registerOutputs_283__4,
           registerOutputs_283__3,registerOutputs_283__2,registerOutputs_283__1,
           registerOutputs_283__0})) ;
    Mux2_16 loop1_284_y (.A ({nx35965,nx36107,nx36249,nx36391,nx36533,nx36675,
            nx36817,nx36959,nx37101,nx37243,nx37385,nx37527,nx37669,nx37811,
            nx37953,nx38095}), .B ({nx33721,nx33859,nx33997,nx34137,nx34275,
            nx34413,nx34551,nx34691,nx34833,nx34975,nx35117,nx35259,nx35401,
            nx35543,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35685), .C ({inputRegisters_284__15,inputRegisters_284__14,
            inputRegisters_284__13,inputRegisters_284__12,inputRegisters_284__11
            ,inputRegisters_284__10,inputRegisters_284__9,inputRegisters_284__8,
            inputRegisters_284__7,inputRegisters_284__6,inputRegisters_284__5,
            inputRegisters_284__4,inputRegisters_284__3,inputRegisters_284__2,
            inputRegisters_284__1,inputRegisters_284__0})) ;
    Reg_16 loop1_284_x (.D ({inputRegisters_284__15,inputRegisters_284__14,
           inputRegisters_284__13,inputRegisters_284__12,inputRegisters_284__11,
           inputRegisters_284__10,inputRegisters_284__9,inputRegisters_284__8,
           inputRegisters_284__7,inputRegisters_284__6,inputRegisters_284__5,
           inputRegisters_284__4,inputRegisters_284__3,inputRegisters_284__2,
           inputRegisters_284__1,inputRegisters_284__0}), .en (
           enableRegister_284), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_284__15,registerOutputs_284__14,
           registerOutputs_284__13,registerOutputs_284__12,
           registerOutputs_284__11,registerOutputs_284__10,
           registerOutputs_284__9,registerOutputs_284__8,registerOutputs_284__7,
           registerOutputs_284__6,registerOutputs_284__5,registerOutputs_284__4,
           registerOutputs_284__3,registerOutputs_284__2,registerOutputs_284__1,
           registerOutputs_284__0})) ;
    Mux2_16 loop1_285_y (.A ({nx35965,nx36107,nx36249,nx36391,nx36533,nx36675,
            nx36817,nx36959,nx37101,nx37243,nx37385,nx37527,nx37669,nx37811,
            nx37953,nx38095}), .B ({nx33721,nx33859,nx33999,nx34137,nx34275,
            nx34413,nx34551,nx34691,nx34833,nx34975,nx35117,nx35259,nx35401,
            nx35543,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35685), .C ({inputRegisters_285__15,inputRegisters_285__14,
            inputRegisters_285__13,inputRegisters_285__12,inputRegisters_285__11
            ,inputRegisters_285__10,inputRegisters_285__9,inputRegisters_285__8,
            inputRegisters_285__7,inputRegisters_285__6,inputRegisters_285__5,
            inputRegisters_285__4,inputRegisters_285__3,inputRegisters_285__2,
            inputRegisters_285__1,inputRegisters_285__0})) ;
    Reg_16 loop1_285_x (.D ({inputRegisters_285__15,inputRegisters_285__14,
           inputRegisters_285__13,inputRegisters_285__12,inputRegisters_285__11,
           inputRegisters_285__10,inputRegisters_285__9,inputRegisters_285__8,
           inputRegisters_285__7,inputRegisters_285__6,inputRegisters_285__5,
           inputRegisters_285__4,inputRegisters_285__3,inputRegisters_285__2,
           inputRegisters_285__1,inputRegisters_285__0}), .en (
           enableRegister_285), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_285__15,registerOutputs_285__14,
           registerOutputs_285__13,registerOutputs_285__12,
           registerOutputs_285__11,registerOutputs_285__10,
           registerOutputs_285__9,registerOutputs_285__8,registerOutputs_285__7,
           registerOutputs_285__6,registerOutputs_285__5,registerOutputs_285__4,
           registerOutputs_285__3,registerOutputs_285__2,registerOutputs_285__1,
           registerOutputs_285__0})) ;
    Mux2_16 loop1_286_y (.A ({nx35965,nx36107,nx36249,nx36391,nx36533,nx36675,
            nx36817,nx36959,nx37101,nx37243,nx37385,nx37527,nx37669,nx37811,
            nx37953,nx38095}), .B ({nx33721,nx33861,nx33999,nx34137,nx34275,
            nx34413,nx34551,nx34691,nx34833,nx34975,nx35117,nx35259,nx35401,
            nx35543,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35685), .C ({inputRegisters_286__15,inputRegisters_286__14,
            inputRegisters_286__13,inputRegisters_286__12,inputRegisters_286__11
            ,inputRegisters_286__10,inputRegisters_286__9,inputRegisters_286__8,
            inputRegisters_286__7,inputRegisters_286__6,inputRegisters_286__5,
            inputRegisters_286__4,inputRegisters_286__3,inputRegisters_286__2,
            inputRegisters_286__1,inputRegisters_286__0})) ;
    Reg_16 loop1_286_x (.D ({inputRegisters_286__15,inputRegisters_286__14,
           inputRegisters_286__13,inputRegisters_286__12,inputRegisters_286__11,
           inputRegisters_286__10,inputRegisters_286__9,inputRegisters_286__8,
           inputRegisters_286__7,inputRegisters_286__6,inputRegisters_286__5,
           inputRegisters_286__4,inputRegisters_286__3,inputRegisters_286__2,
           inputRegisters_286__1,inputRegisters_286__0}), .en (
           enableRegister_286), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_286__15,registerOutputs_286__14,
           registerOutputs_286__13,registerOutputs_286__12,
           registerOutputs_286__11,registerOutputs_286__10,
           registerOutputs_286__9,registerOutputs_286__8,registerOutputs_286__7,
           registerOutputs_286__6,registerOutputs_286__5,registerOutputs_286__4,
           registerOutputs_286__3,registerOutputs_286__2,registerOutputs_286__1,
           registerOutputs_286__0})) ;
    Mux2_16 loop1_287_y (.A ({nx35967,nx36109,nx36251,nx36393,nx36535,nx36677,
            nx36819,nx36961,nx37103,nx37245,nx37387,nx37529,nx37671,nx37813,
            nx37955,nx38097}), .B ({nx33723,nx33861,nx33999,nx34137,nx34275,
            nx34413,nx34551,nx34693,nx34835,nx34977,nx35119,nx35261,nx35403,
            nx35545,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35687), .C ({inputRegisters_287__15,inputRegisters_287__14,
            inputRegisters_287__13,inputRegisters_287__12,inputRegisters_287__11
            ,inputRegisters_287__10,inputRegisters_287__9,inputRegisters_287__8,
            inputRegisters_287__7,inputRegisters_287__6,inputRegisters_287__5,
            inputRegisters_287__4,inputRegisters_287__3,inputRegisters_287__2,
            inputRegisters_287__1,inputRegisters_287__0})) ;
    Reg_16 loop1_287_x (.D ({inputRegisters_287__15,inputRegisters_287__14,
           inputRegisters_287__13,inputRegisters_287__12,inputRegisters_287__11,
           inputRegisters_287__10,inputRegisters_287__9,inputRegisters_287__8,
           inputRegisters_287__7,inputRegisters_287__6,inputRegisters_287__5,
           inputRegisters_287__4,inputRegisters_287__3,inputRegisters_287__2,
           inputRegisters_287__1,inputRegisters_287__0}), .en (
           enableRegister_287), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_287__15,registerOutputs_287__14,
           registerOutputs_287__13,registerOutputs_287__12,
           registerOutputs_287__11,registerOutputs_287__10,
           registerOutputs_287__9,registerOutputs_287__8,registerOutputs_287__7,
           registerOutputs_287__6,registerOutputs_287__5,registerOutputs_287__4,
           registerOutputs_287__3,registerOutputs_287__2,registerOutputs_287__1,
           registerOutputs_287__0})) ;
    Mux2_16 loop1_288_y (.A ({nx35967,nx36109,nx36251,nx36393,nx36535,nx36677,
            nx36819,nx36961,nx37103,nx37245,nx37387,nx37529,nx37671,nx37813,
            nx37955,nx38097}), .B ({nx33723,nx33861,nx33999,nx34137,nx34275,
            nx34413,nx34553,nx34693,nx34835,nx34977,nx35119,nx35261,nx35403,
            nx35545,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35687), .C ({inputRegisters_288__15,inputRegisters_288__14,
            inputRegisters_288__13,inputRegisters_288__12,inputRegisters_288__11
            ,inputRegisters_288__10,inputRegisters_288__9,inputRegisters_288__8,
            inputRegisters_288__7,inputRegisters_288__6,inputRegisters_288__5,
            inputRegisters_288__4,inputRegisters_288__3,inputRegisters_288__2,
            inputRegisters_288__1,inputRegisters_288__0})) ;
    Reg_16 loop1_288_x (.D ({inputRegisters_288__15,inputRegisters_288__14,
           inputRegisters_288__13,inputRegisters_288__12,inputRegisters_288__11,
           inputRegisters_288__10,inputRegisters_288__9,inputRegisters_288__8,
           inputRegisters_288__7,inputRegisters_288__6,inputRegisters_288__5,
           inputRegisters_288__4,inputRegisters_288__3,inputRegisters_288__2,
           inputRegisters_288__1,inputRegisters_288__0}), .en (
           enableRegister_288), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_288__15,registerOutputs_288__14,
           registerOutputs_288__13,registerOutputs_288__12,
           registerOutputs_288__11,registerOutputs_288__10,
           registerOutputs_288__9,registerOutputs_288__8,registerOutputs_288__7,
           registerOutputs_288__6,registerOutputs_288__5,registerOutputs_288__4,
           registerOutputs_288__3,registerOutputs_288__2,registerOutputs_288__1,
           registerOutputs_288__0})) ;
    Mux2_16 loop1_289_y (.A ({nx35967,nx36109,nx36251,nx36393,nx36535,nx36677,
            nx36819,nx36961,nx37103,nx37245,nx37387,nx37529,nx37671,nx37813,
            nx37955,nx38097}), .B ({nx33723,nx33861,nx33999,nx34137,nx34275,
            nx34415,nx34553,nx34693,nx34835,nx34977,nx35119,nx35261,nx35403,
            nx35545,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35687), .C ({inputRegisters_289__15,inputRegisters_289__14,
            inputRegisters_289__13,inputRegisters_289__12,inputRegisters_289__11
            ,inputRegisters_289__10,inputRegisters_289__9,inputRegisters_289__8,
            inputRegisters_289__7,inputRegisters_289__6,inputRegisters_289__5,
            inputRegisters_289__4,inputRegisters_289__3,inputRegisters_289__2,
            inputRegisters_289__1,inputRegisters_289__0})) ;
    Reg_16 loop1_289_x (.D ({inputRegisters_289__15,inputRegisters_289__14,
           inputRegisters_289__13,inputRegisters_289__12,inputRegisters_289__11,
           inputRegisters_289__10,inputRegisters_289__9,inputRegisters_289__8,
           inputRegisters_289__7,inputRegisters_289__6,inputRegisters_289__5,
           inputRegisters_289__4,inputRegisters_289__3,inputRegisters_289__2,
           inputRegisters_289__1,inputRegisters_289__0}), .en (
           enableRegister_289), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_289__15,registerOutputs_289__14,
           registerOutputs_289__13,registerOutputs_289__12,
           registerOutputs_289__11,registerOutputs_289__10,
           registerOutputs_289__9,registerOutputs_289__8,registerOutputs_289__7,
           registerOutputs_289__6,registerOutputs_289__5,registerOutputs_289__4,
           registerOutputs_289__3,registerOutputs_289__2,registerOutputs_289__1,
           registerOutputs_289__0})) ;
    Mux2_16 loop1_290_y (.A ({nx35967,nx36109,nx36251,nx36393,nx36535,nx36677,
            nx36819,nx36961,nx37103,nx37245,nx37387,nx37529,nx37671,nx37813,
            nx37955,nx38097}), .B ({nx33723,nx33861,nx33999,nx34137,nx34277,
            nx34415,nx34553,nx34693,nx34835,nx34977,nx35119,nx35261,nx35403,
            nx35545,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35687), .C ({inputRegisters_290__15,inputRegisters_290__14,
            inputRegisters_290__13,inputRegisters_290__12,inputRegisters_290__11
            ,inputRegisters_290__10,inputRegisters_290__9,inputRegisters_290__8,
            inputRegisters_290__7,inputRegisters_290__6,inputRegisters_290__5,
            inputRegisters_290__4,inputRegisters_290__3,inputRegisters_290__2,
            inputRegisters_290__1,inputRegisters_290__0})) ;
    Reg_16 loop1_290_x (.D ({inputRegisters_290__15,inputRegisters_290__14,
           inputRegisters_290__13,inputRegisters_290__12,inputRegisters_290__11,
           inputRegisters_290__10,inputRegisters_290__9,inputRegisters_290__8,
           inputRegisters_290__7,inputRegisters_290__6,inputRegisters_290__5,
           inputRegisters_290__4,inputRegisters_290__3,inputRegisters_290__2,
           inputRegisters_290__1,inputRegisters_290__0}), .en (
           enableRegister_290), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_290__15,registerOutputs_290__14,
           registerOutputs_290__13,registerOutputs_290__12,
           registerOutputs_290__11,registerOutputs_290__10,
           registerOutputs_290__9,registerOutputs_290__8,registerOutputs_290__7,
           registerOutputs_290__6,registerOutputs_290__5,registerOutputs_290__4,
           registerOutputs_290__3,registerOutputs_290__2,registerOutputs_290__1,
           registerOutputs_290__0})) ;
    Mux2_16 loop1_291_y (.A ({nx35967,nx36109,nx36251,nx36393,nx36535,nx36677,
            nx36819,nx36961,nx37103,nx37245,nx37387,nx37529,nx37671,nx37813,
            nx37955,nx38097}), .B ({nx33723,nx33861,nx33999,nx34139,nx34277,
            nx34415,nx34553,nx34693,nx34835,nx34977,nx35119,nx35261,nx35403,
            nx35545,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35687), .C ({inputRegisters_291__15,inputRegisters_291__14,
            inputRegisters_291__13,inputRegisters_291__12,inputRegisters_291__11
            ,inputRegisters_291__10,inputRegisters_291__9,inputRegisters_291__8,
            inputRegisters_291__7,inputRegisters_291__6,inputRegisters_291__5,
            inputRegisters_291__4,inputRegisters_291__3,inputRegisters_291__2,
            inputRegisters_291__1,inputRegisters_291__0})) ;
    Reg_16 loop1_291_x (.D ({inputRegisters_291__15,inputRegisters_291__14,
           inputRegisters_291__13,inputRegisters_291__12,inputRegisters_291__11,
           inputRegisters_291__10,inputRegisters_291__9,inputRegisters_291__8,
           inputRegisters_291__7,inputRegisters_291__6,inputRegisters_291__5,
           inputRegisters_291__4,inputRegisters_291__3,inputRegisters_291__2,
           inputRegisters_291__1,inputRegisters_291__0}), .en (
           enableRegister_291), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_291__15,registerOutputs_291__14,
           registerOutputs_291__13,registerOutputs_291__12,
           registerOutputs_291__11,registerOutputs_291__10,
           registerOutputs_291__9,registerOutputs_291__8,registerOutputs_291__7,
           registerOutputs_291__6,registerOutputs_291__5,registerOutputs_291__4,
           registerOutputs_291__3,registerOutputs_291__2,registerOutputs_291__1,
           registerOutputs_291__0})) ;
    Mux2_16 loop1_292_y (.A ({nx35967,nx36109,nx36251,nx36393,nx36535,nx36677,
            nx36819,nx36961,nx37103,nx37245,nx37387,nx37529,nx37671,nx37813,
            nx37955,nx38097}), .B ({nx33723,nx33861,nx34001,nx34139,nx34277,
            nx34415,nx34553,nx34693,nx34835,nx34977,nx35119,nx35261,nx35403,
            nx35545,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35687), .C ({inputRegisters_292__15,inputRegisters_292__14,
            inputRegisters_292__13,inputRegisters_292__12,inputRegisters_292__11
            ,inputRegisters_292__10,inputRegisters_292__9,inputRegisters_292__8,
            inputRegisters_292__7,inputRegisters_292__6,inputRegisters_292__5,
            inputRegisters_292__4,inputRegisters_292__3,inputRegisters_292__2,
            inputRegisters_292__1,inputRegisters_292__0})) ;
    Reg_16 loop1_292_x (.D ({inputRegisters_292__15,inputRegisters_292__14,
           inputRegisters_292__13,inputRegisters_292__12,inputRegisters_292__11,
           inputRegisters_292__10,inputRegisters_292__9,inputRegisters_292__8,
           inputRegisters_292__7,inputRegisters_292__6,inputRegisters_292__5,
           inputRegisters_292__4,inputRegisters_292__3,inputRegisters_292__2,
           inputRegisters_292__1,inputRegisters_292__0}), .en (
           enableRegister_292), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_292__15,registerOutputs_292__14,
           registerOutputs_292__13,registerOutputs_292__12,
           registerOutputs_292__11,registerOutputs_292__10,
           registerOutputs_292__9,registerOutputs_292__8,registerOutputs_292__7,
           registerOutputs_292__6,registerOutputs_292__5,registerOutputs_292__4,
           registerOutputs_292__3,registerOutputs_292__2,registerOutputs_292__1,
           registerOutputs_292__0})) ;
    Mux2_16 loop1_293_y (.A ({nx35967,nx36109,nx36251,nx36393,nx36535,nx36677,
            nx36819,nx36961,nx37103,nx37245,nx37387,nx37529,nx37671,nx37813,
            nx37955,nx38097}), .B ({nx33723,nx33863,nx34001,nx34139,nx34277,
            nx34415,nx34553,nx34693,nx34835,nx34977,nx35119,nx35261,nx35403,
            nx35545,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35687), .C ({inputRegisters_293__15,inputRegisters_293__14,
            inputRegisters_293__13,inputRegisters_293__12,inputRegisters_293__11
            ,inputRegisters_293__10,inputRegisters_293__9,inputRegisters_293__8,
            inputRegisters_293__7,inputRegisters_293__6,inputRegisters_293__5,
            inputRegisters_293__4,inputRegisters_293__3,inputRegisters_293__2,
            inputRegisters_293__1,inputRegisters_293__0})) ;
    Reg_16 loop1_293_x (.D ({inputRegisters_293__15,inputRegisters_293__14,
           inputRegisters_293__13,inputRegisters_293__12,inputRegisters_293__11,
           inputRegisters_293__10,inputRegisters_293__9,inputRegisters_293__8,
           inputRegisters_293__7,inputRegisters_293__6,inputRegisters_293__5,
           inputRegisters_293__4,inputRegisters_293__3,inputRegisters_293__2,
           inputRegisters_293__1,inputRegisters_293__0}), .en (
           enableRegister_293), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_293__15,registerOutputs_293__14,
           registerOutputs_293__13,registerOutputs_293__12,
           registerOutputs_293__11,registerOutputs_293__10,
           registerOutputs_293__9,registerOutputs_293__8,registerOutputs_293__7,
           registerOutputs_293__6,registerOutputs_293__5,registerOutputs_293__4,
           registerOutputs_293__3,registerOutputs_293__2,registerOutputs_293__1,
           registerOutputs_293__0})) ;
    Mux2_16 loop1_294_y (.A ({nx35969,nx36111,nx36253,nx36395,nx36537,nx36679,
            nx36821,nx36963,nx37105,nx37247,nx37389,nx37531,nx37673,nx37815,
            nx37957,nx38099}), .B ({nx33725,nx33863,nx34001,nx34139,nx34277,
            nx34415,nx34553,nx34695,nx34837,nx34979,nx35121,nx35263,nx35405,
            nx35547,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35689), .C ({inputRegisters_294__15,inputRegisters_294__14,
            inputRegisters_294__13,inputRegisters_294__12,inputRegisters_294__11
            ,inputRegisters_294__10,inputRegisters_294__9,inputRegisters_294__8,
            inputRegisters_294__7,inputRegisters_294__6,inputRegisters_294__5,
            inputRegisters_294__4,inputRegisters_294__3,inputRegisters_294__2,
            inputRegisters_294__1,inputRegisters_294__0})) ;
    Reg_16 loop1_294_x (.D ({inputRegisters_294__15,inputRegisters_294__14,
           inputRegisters_294__13,inputRegisters_294__12,inputRegisters_294__11,
           inputRegisters_294__10,inputRegisters_294__9,inputRegisters_294__8,
           inputRegisters_294__7,inputRegisters_294__6,inputRegisters_294__5,
           inputRegisters_294__4,inputRegisters_294__3,inputRegisters_294__2,
           inputRegisters_294__1,inputRegisters_294__0}), .en (
           enableRegister_294), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_294__15,registerOutputs_294__14,
           registerOutputs_294__13,registerOutputs_294__12,
           registerOutputs_294__11,registerOutputs_294__10,
           registerOutputs_294__9,registerOutputs_294__8,registerOutputs_294__7,
           registerOutputs_294__6,registerOutputs_294__5,registerOutputs_294__4,
           registerOutputs_294__3,registerOutputs_294__2,registerOutputs_294__1,
           registerOutputs_294__0})) ;
    Mux2_16 loop1_295_y (.A ({nx35969,nx36111,nx36253,nx36395,nx36537,nx36679,
            nx36821,nx36963,nx37105,nx37247,nx37389,nx37531,nx37673,nx37815,
            nx37957,nx38099}), .B ({nx33725,nx33863,nx34001,nx34139,nx34277,
            nx34415,nx34555,nx34695,nx34837,nx34979,nx35121,nx35263,nx35405,
            nx35547,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35689), .C ({inputRegisters_295__15,inputRegisters_295__14,
            inputRegisters_295__13,inputRegisters_295__12,inputRegisters_295__11
            ,inputRegisters_295__10,inputRegisters_295__9,inputRegisters_295__8,
            inputRegisters_295__7,inputRegisters_295__6,inputRegisters_295__5,
            inputRegisters_295__4,inputRegisters_295__3,inputRegisters_295__2,
            inputRegisters_295__1,inputRegisters_295__0})) ;
    Reg_16 loop1_295_x (.D ({inputRegisters_295__15,inputRegisters_295__14,
           inputRegisters_295__13,inputRegisters_295__12,inputRegisters_295__11,
           inputRegisters_295__10,inputRegisters_295__9,inputRegisters_295__8,
           inputRegisters_295__7,inputRegisters_295__6,inputRegisters_295__5,
           inputRegisters_295__4,inputRegisters_295__3,inputRegisters_295__2,
           inputRegisters_295__1,inputRegisters_295__0}), .en (
           enableRegister_295), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_295__15,registerOutputs_295__14,
           registerOutputs_295__13,registerOutputs_295__12,
           registerOutputs_295__11,registerOutputs_295__10,
           registerOutputs_295__9,registerOutputs_295__8,registerOutputs_295__7,
           registerOutputs_295__6,registerOutputs_295__5,registerOutputs_295__4,
           registerOutputs_295__3,registerOutputs_295__2,registerOutputs_295__1,
           registerOutputs_295__0})) ;
    Mux2_16 loop1_296_y (.A ({nx35969,nx36111,nx36253,nx36395,nx36537,nx36679,
            nx36821,nx36963,nx37105,nx37247,nx37389,nx37531,nx37673,nx37815,
            nx37957,nx38099}), .B ({nx33725,nx33863,nx34001,nx34139,nx34277,
            nx34417,nx34555,nx34695,nx34837,nx34979,nx35121,nx35263,nx35405,
            nx35547,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35689), .C ({inputRegisters_296__15,inputRegisters_296__14,
            inputRegisters_296__13,inputRegisters_296__12,inputRegisters_296__11
            ,inputRegisters_296__10,inputRegisters_296__9,inputRegisters_296__8,
            inputRegisters_296__7,inputRegisters_296__6,inputRegisters_296__5,
            inputRegisters_296__4,inputRegisters_296__3,inputRegisters_296__2,
            inputRegisters_296__1,inputRegisters_296__0})) ;
    Reg_16 loop1_296_x (.D ({inputRegisters_296__15,inputRegisters_296__14,
           inputRegisters_296__13,inputRegisters_296__12,inputRegisters_296__11,
           inputRegisters_296__10,inputRegisters_296__9,inputRegisters_296__8,
           inputRegisters_296__7,inputRegisters_296__6,inputRegisters_296__5,
           inputRegisters_296__4,inputRegisters_296__3,inputRegisters_296__2,
           inputRegisters_296__1,inputRegisters_296__0}), .en (
           enableRegister_296), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_296__15,registerOutputs_296__14,
           registerOutputs_296__13,registerOutputs_296__12,
           registerOutputs_296__11,registerOutputs_296__10,
           registerOutputs_296__9,registerOutputs_296__8,registerOutputs_296__7,
           registerOutputs_296__6,registerOutputs_296__5,registerOutputs_296__4,
           registerOutputs_296__3,registerOutputs_296__2,registerOutputs_296__1,
           registerOutputs_296__0})) ;
    Mux2_16 loop1_297_y (.A ({nx35969,nx36111,nx36253,nx36395,nx36537,nx36679,
            nx36821,nx36963,nx37105,nx37247,nx37389,nx37531,nx37673,nx37815,
            nx37957,nx38099}), .B ({nx33725,nx33863,nx34001,nx34139,nx34279,
            nx34417,nx34555,nx34695,nx34837,nx34979,nx35121,nx35263,nx35405,
            nx35547,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35689), .C ({inputRegisters_297__15,inputRegisters_297__14,
            inputRegisters_297__13,inputRegisters_297__12,inputRegisters_297__11
            ,inputRegisters_297__10,inputRegisters_297__9,inputRegisters_297__8,
            inputRegisters_297__7,inputRegisters_297__6,inputRegisters_297__5,
            inputRegisters_297__4,inputRegisters_297__3,inputRegisters_297__2,
            inputRegisters_297__1,inputRegisters_297__0})) ;
    Reg_16 loop1_297_x (.D ({inputRegisters_297__15,inputRegisters_297__14,
           inputRegisters_297__13,inputRegisters_297__12,inputRegisters_297__11,
           inputRegisters_297__10,inputRegisters_297__9,inputRegisters_297__8,
           inputRegisters_297__7,inputRegisters_297__6,inputRegisters_297__5,
           inputRegisters_297__4,inputRegisters_297__3,inputRegisters_297__2,
           inputRegisters_297__1,inputRegisters_297__0}), .en (
           enableRegister_297), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_297__15,registerOutputs_297__14,
           registerOutputs_297__13,registerOutputs_297__12,
           registerOutputs_297__11,registerOutputs_297__10,
           registerOutputs_297__9,registerOutputs_297__8,registerOutputs_297__7,
           registerOutputs_297__6,registerOutputs_297__5,registerOutputs_297__4,
           registerOutputs_297__3,registerOutputs_297__2,registerOutputs_297__1,
           registerOutputs_297__0})) ;
    Mux2_16 loop1_298_y (.A ({nx35969,nx36111,nx36253,nx36395,nx36537,nx36679,
            nx36821,nx36963,nx37105,nx37247,nx37389,nx37531,nx37673,nx37815,
            nx37957,nx38099}), .B ({nx33725,nx33863,nx34001,nx34141,nx34279,
            nx34417,nx34555,nx34695,nx34837,nx34979,nx35121,nx35263,nx35405,
            nx35547,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35689), .C ({inputRegisters_298__15,inputRegisters_298__14,
            inputRegisters_298__13,inputRegisters_298__12,inputRegisters_298__11
            ,inputRegisters_298__10,inputRegisters_298__9,inputRegisters_298__8,
            inputRegisters_298__7,inputRegisters_298__6,inputRegisters_298__5,
            inputRegisters_298__4,inputRegisters_298__3,inputRegisters_298__2,
            inputRegisters_298__1,inputRegisters_298__0})) ;
    Reg_16 loop1_298_x (.D ({inputRegisters_298__15,inputRegisters_298__14,
           inputRegisters_298__13,inputRegisters_298__12,inputRegisters_298__11,
           inputRegisters_298__10,inputRegisters_298__9,inputRegisters_298__8,
           inputRegisters_298__7,inputRegisters_298__6,inputRegisters_298__5,
           inputRegisters_298__4,inputRegisters_298__3,inputRegisters_298__2,
           inputRegisters_298__1,inputRegisters_298__0}), .en (
           enableRegister_298), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_298__15,registerOutputs_298__14,
           registerOutputs_298__13,registerOutputs_298__12,
           registerOutputs_298__11,registerOutputs_298__10,
           registerOutputs_298__9,registerOutputs_298__8,registerOutputs_298__7,
           registerOutputs_298__6,registerOutputs_298__5,registerOutputs_298__4,
           registerOutputs_298__3,registerOutputs_298__2,registerOutputs_298__1,
           registerOutputs_298__0})) ;
    Mux2_16 loop1_299_y (.A ({nx35969,nx36111,nx36253,nx36395,nx36537,nx36679,
            nx36821,nx36963,nx37105,nx37247,nx37389,nx37531,nx37673,nx37815,
            nx37957,nx38099}), .B ({nx33725,nx33863,nx34003,nx34141,nx34279,
            nx34417,nx34555,nx34695,nx34837,nx34979,nx35121,nx35263,nx35405,
            nx35547,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35689), .C ({inputRegisters_299__15,inputRegisters_299__14,
            inputRegisters_299__13,inputRegisters_299__12,inputRegisters_299__11
            ,inputRegisters_299__10,inputRegisters_299__9,inputRegisters_299__8,
            inputRegisters_299__7,inputRegisters_299__6,inputRegisters_299__5,
            inputRegisters_299__4,inputRegisters_299__3,inputRegisters_299__2,
            inputRegisters_299__1,inputRegisters_299__0})) ;
    Reg_16 loop1_299_x (.D ({inputRegisters_299__15,inputRegisters_299__14,
           inputRegisters_299__13,inputRegisters_299__12,inputRegisters_299__11,
           inputRegisters_299__10,inputRegisters_299__9,inputRegisters_299__8,
           inputRegisters_299__7,inputRegisters_299__6,inputRegisters_299__5,
           inputRegisters_299__4,inputRegisters_299__3,inputRegisters_299__2,
           inputRegisters_299__1,inputRegisters_299__0}), .en (
           enableRegister_299), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_299__15,registerOutputs_299__14,
           registerOutputs_299__13,registerOutputs_299__12,
           registerOutputs_299__11,registerOutputs_299__10,
           registerOutputs_299__9,registerOutputs_299__8,registerOutputs_299__7,
           registerOutputs_299__6,registerOutputs_299__5,registerOutputs_299__4,
           registerOutputs_299__3,registerOutputs_299__2,registerOutputs_299__1,
           registerOutputs_299__0})) ;
    Mux2_16 loop1_300_y (.A ({nx35969,nx36111,nx36253,nx36395,nx36537,nx36679,
            nx36821,nx36963,nx37105,nx37247,nx37389,nx37531,nx37673,nx37815,
            nx37957,nx38099}), .B ({nx33725,nx33865,nx34003,nx34141,nx34279,
            nx34417,nx34555,nx34695,nx34837,nx34979,nx35121,nx35263,nx35405,
            nx35547,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35689), .C ({inputRegisters_300__15,inputRegisters_300__14,
            inputRegisters_300__13,inputRegisters_300__12,inputRegisters_300__11
            ,inputRegisters_300__10,inputRegisters_300__9,inputRegisters_300__8,
            inputRegisters_300__7,inputRegisters_300__6,inputRegisters_300__5,
            inputRegisters_300__4,inputRegisters_300__3,inputRegisters_300__2,
            inputRegisters_300__1,inputRegisters_300__0})) ;
    Reg_16 loop1_300_x (.D ({inputRegisters_300__15,inputRegisters_300__14,
           inputRegisters_300__13,inputRegisters_300__12,inputRegisters_300__11,
           inputRegisters_300__10,inputRegisters_300__9,inputRegisters_300__8,
           inputRegisters_300__7,inputRegisters_300__6,inputRegisters_300__5,
           inputRegisters_300__4,inputRegisters_300__3,inputRegisters_300__2,
           inputRegisters_300__1,inputRegisters_300__0}), .en (
           enableRegister_300), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_300__15,registerOutputs_300__14,
           registerOutputs_300__13,registerOutputs_300__12,
           registerOutputs_300__11,registerOutputs_300__10,
           registerOutputs_300__9,registerOutputs_300__8,registerOutputs_300__7,
           registerOutputs_300__6,registerOutputs_300__5,registerOutputs_300__4,
           registerOutputs_300__3,registerOutputs_300__2,registerOutputs_300__1,
           registerOutputs_300__0})) ;
    Mux2_16 loop1_301_y (.A ({nx35971,nx36113,nx36255,nx36397,nx36539,nx36681,
            nx36823,nx36965,nx37107,nx37249,nx37391,nx37533,nx37675,nx37817,
            nx37959,nx38101}), .B ({nx33727,nx33865,nx34003,nx34141,nx34279,
            nx34417,nx34555,nx34697,nx34839,nx34981,nx35123,nx35265,nx35407,
            nx35549,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35691), .C ({inputRegisters_301__15,inputRegisters_301__14,
            inputRegisters_301__13,inputRegisters_301__12,inputRegisters_301__11
            ,inputRegisters_301__10,inputRegisters_301__9,inputRegisters_301__8,
            inputRegisters_301__7,inputRegisters_301__6,inputRegisters_301__5,
            inputRegisters_301__4,inputRegisters_301__3,inputRegisters_301__2,
            inputRegisters_301__1,inputRegisters_301__0})) ;
    Reg_16 loop1_301_x (.D ({inputRegisters_301__15,inputRegisters_301__14,
           inputRegisters_301__13,inputRegisters_301__12,inputRegisters_301__11,
           inputRegisters_301__10,inputRegisters_301__9,inputRegisters_301__8,
           inputRegisters_301__7,inputRegisters_301__6,inputRegisters_301__5,
           inputRegisters_301__4,inputRegisters_301__3,inputRegisters_301__2,
           inputRegisters_301__1,inputRegisters_301__0}), .en (
           enableRegister_301), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_301__15,registerOutputs_301__14,
           registerOutputs_301__13,registerOutputs_301__12,
           registerOutputs_301__11,registerOutputs_301__10,
           registerOutputs_301__9,registerOutputs_301__8,registerOutputs_301__7,
           registerOutputs_301__6,registerOutputs_301__5,registerOutputs_301__4,
           registerOutputs_301__3,registerOutputs_301__2,registerOutputs_301__1,
           registerOutputs_301__0})) ;
    Mux2_16 loop1_302_y (.A ({nx35971,nx36113,nx36255,nx36397,nx36539,nx36681,
            nx36823,nx36965,nx37107,nx37249,nx37391,nx37533,nx37675,nx37817,
            nx37959,nx38101}), .B ({nx33727,nx33865,nx34003,nx34141,nx34279,
            nx34417,nx34557,nx34697,nx34839,nx34981,nx35123,nx35265,nx35407,
            nx35549,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35691), .C ({inputRegisters_302__15,inputRegisters_302__14,
            inputRegisters_302__13,inputRegisters_302__12,inputRegisters_302__11
            ,inputRegisters_302__10,inputRegisters_302__9,inputRegisters_302__8,
            inputRegisters_302__7,inputRegisters_302__6,inputRegisters_302__5,
            inputRegisters_302__4,inputRegisters_302__3,inputRegisters_302__2,
            inputRegisters_302__1,inputRegisters_302__0})) ;
    Reg_16 loop1_302_x (.D ({inputRegisters_302__15,inputRegisters_302__14,
           inputRegisters_302__13,inputRegisters_302__12,inputRegisters_302__11,
           inputRegisters_302__10,inputRegisters_302__9,inputRegisters_302__8,
           inputRegisters_302__7,inputRegisters_302__6,inputRegisters_302__5,
           inputRegisters_302__4,inputRegisters_302__3,inputRegisters_302__2,
           inputRegisters_302__1,inputRegisters_302__0}), .en (
           enableRegister_302), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_302__15,registerOutputs_302__14,
           registerOutputs_302__13,registerOutputs_302__12,
           registerOutputs_302__11,registerOutputs_302__10,
           registerOutputs_302__9,registerOutputs_302__8,registerOutputs_302__7,
           registerOutputs_302__6,registerOutputs_302__5,registerOutputs_302__4,
           registerOutputs_302__3,registerOutputs_302__2,registerOutputs_302__1,
           registerOutputs_302__0})) ;
    Mux2_16 loop1_303_y (.A ({nx35971,nx36113,nx36255,nx36397,nx36539,nx36681,
            nx36823,nx36965,nx37107,nx37249,nx37391,nx37533,nx37675,nx37817,
            nx37959,nx38101}), .B ({nx33727,nx33865,nx34003,nx34141,nx34279,
            nx34419,nx34557,nx34697,nx34839,nx34981,nx35123,nx35265,nx35407,
            nx35549,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35691), .C ({inputRegisters_303__15,inputRegisters_303__14,
            inputRegisters_303__13,inputRegisters_303__12,inputRegisters_303__11
            ,inputRegisters_303__10,inputRegisters_303__9,inputRegisters_303__8,
            inputRegisters_303__7,inputRegisters_303__6,inputRegisters_303__5,
            inputRegisters_303__4,inputRegisters_303__3,inputRegisters_303__2,
            inputRegisters_303__1,inputRegisters_303__0})) ;
    Reg_16 loop1_303_x (.D ({inputRegisters_303__15,inputRegisters_303__14,
           inputRegisters_303__13,inputRegisters_303__12,inputRegisters_303__11,
           inputRegisters_303__10,inputRegisters_303__9,inputRegisters_303__8,
           inputRegisters_303__7,inputRegisters_303__6,inputRegisters_303__5,
           inputRegisters_303__4,inputRegisters_303__3,inputRegisters_303__2,
           inputRegisters_303__1,inputRegisters_303__0}), .en (
           enableRegister_303), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_303__15,registerOutputs_303__14,
           registerOutputs_303__13,registerOutputs_303__12,
           registerOutputs_303__11,registerOutputs_303__10,
           registerOutputs_303__9,registerOutputs_303__8,registerOutputs_303__7,
           registerOutputs_303__6,registerOutputs_303__5,registerOutputs_303__4,
           registerOutputs_303__3,registerOutputs_303__2,registerOutputs_303__1,
           registerOutputs_303__0})) ;
    Mux2_16 loop1_304_y (.A ({nx35971,nx36113,nx36255,nx36397,nx36539,nx36681,
            nx36823,nx36965,nx37107,nx37249,nx37391,nx37533,nx37675,nx37817,
            nx37959,nx38101}), .B ({nx33727,nx33865,nx34003,nx34141,nx34281,
            nx34419,nx34557,nx34697,nx34839,nx34981,nx35123,nx35265,nx35407,
            nx35549,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35691), .C ({inputRegisters_304__15,inputRegisters_304__14,
            inputRegisters_304__13,inputRegisters_304__12,inputRegisters_304__11
            ,inputRegisters_304__10,inputRegisters_304__9,inputRegisters_304__8,
            inputRegisters_304__7,inputRegisters_304__6,inputRegisters_304__5,
            inputRegisters_304__4,inputRegisters_304__3,inputRegisters_304__2,
            inputRegisters_304__1,inputRegisters_304__0})) ;
    Reg_16 loop1_304_x (.D ({inputRegisters_304__15,inputRegisters_304__14,
           inputRegisters_304__13,inputRegisters_304__12,inputRegisters_304__11,
           inputRegisters_304__10,inputRegisters_304__9,inputRegisters_304__8,
           inputRegisters_304__7,inputRegisters_304__6,inputRegisters_304__5,
           inputRegisters_304__4,inputRegisters_304__3,inputRegisters_304__2,
           inputRegisters_304__1,inputRegisters_304__0}), .en (
           enableRegister_304), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_304__15,registerOutputs_304__14,
           registerOutputs_304__13,registerOutputs_304__12,
           registerOutputs_304__11,registerOutputs_304__10,
           registerOutputs_304__9,registerOutputs_304__8,registerOutputs_304__7,
           registerOutputs_304__6,registerOutputs_304__5,registerOutputs_304__4,
           registerOutputs_304__3,registerOutputs_304__2,registerOutputs_304__1,
           registerOutputs_304__0})) ;
    Mux2_16 loop1_305_y (.A ({nx35971,nx36113,nx36255,nx36397,nx36539,nx36681,
            nx36823,nx36965,nx37107,nx37249,nx37391,nx37533,nx37675,nx37817,
            nx37959,nx38101}), .B ({nx33727,nx33865,nx34003,nx34143,nx34281,
            nx34419,nx34557,nx34697,nx34839,nx34981,nx35123,nx35265,nx35407,
            nx35549,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35691), .C ({inputRegisters_305__15,inputRegisters_305__14,
            inputRegisters_305__13,inputRegisters_305__12,inputRegisters_305__11
            ,inputRegisters_305__10,inputRegisters_305__9,inputRegisters_305__8,
            inputRegisters_305__7,inputRegisters_305__6,inputRegisters_305__5,
            inputRegisters_305__4,inputRegisters_305__3,inputRegisters_305__2,
            inputRegisters_305__1,inputRegisters_305__0})) ;
    Reg_16 loop1_305_x (.D ({inputRegisters_305__15,inputRegisters_305__14,
           inputRegisters_305__13,inputRegisters_305__12,inputRegisters_305__11,
           inputRegisters_305__10,inputRegisters_305__9,inputRegisters_305__8,
           inputRegisters_305__7,inputRegisters_305__6,inputRegisters_305__5,
           inputRegisters_305__4,inputRegisters_305__3,inputRegisters_305__2,
           inputRegisters_305__1,inputRegisters_305__0}), .en (
           enableRegister_305), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_305__15,registerOutputs_305__14,
           registerOutputs_305__13,registerOutputs_305__12,
           registerOutputs_305__11,registerOutputs_305__10,
           registerOutputs_305__9,registerOutputs_305__8,registerOutputs_305__7,
           registerOutputs_305__6,registerOutputs_305__5,registerOutputs_305__4,
           registerOutputs_305__3,registerOutputs_305__2,registerOutputs_305__1,
           registerOutputs_305__0})) ;
    Mux2_16 loop1_306_y (.A ({nx35971,nx36113,nx36255,nx36397,nx36539,nx36681,
            nx36823,nx36965,nx37107,nx37249,nx37391,nx37533,nx37675,nx37817,
            nx37959,nx38101}), .B ({nx33727,nx33865,nx34005,nx34143,nx34281,
            nx34419,nx34557,nx34697,nx34839,nx34981,nx35123,nx35265,nx35407,
            nx35549,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35691), .C ({inputRegisters_306__15,inputRegisters_306__14,
            inputRegisters_306__13,inputRegisters_306__12,inputRegisters_306__11
            ,inputRegisters_306__10,inputRegisters_306__9,inputRegisters_306__8,
            inputRegisters_306__7,inputRegisters_306__6,inputRegisters_306__5,
            inputRegisters_306__4,inputRegisters_306__3,inputRegisters_306__2,
            inputRegisters_306__1,inputRegisters_306__0})) ;
    Reg_16 loop1_306_x (.D ({inputRegisters_306__15,inputRegisters_306__14,
           inputRegisters_306__13,inputRegisters_306__12,inputRegisters_306__11,
           inputRegisters_306__10,inputRegisters_306__9,inputRegisters_306__8,
           inputRegisters_306__7,inputRegisters_306__6,inputRegisters_306__5,
           inputRegisters_306__4,inputRegisters_306__3,inputRegisters_306__2,
           inputRegisters_306__1,inputRegisters_306__0}), .en (
           enableRegister_306), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_306__15,registerOutputs_306__14,
           registerOutputs_306__13,registerOutputs_306__12,
           registerOutputs_306__11,registerOutputs_306__10,
           registerOutputs_306__9,registerOutputs_306__8,registerOutputs_306__7,
           registerOutputs_306__6,registerOutputs_306__5,registerOutputs_306__4,
           registerOutputs_306__3,registerOutputs_306__2,registerOutputs_306__1,
           registerOutputs_306__0})) ;
    Mux2_16 loop1_307_y (.A ({nx35971,nx36113,nx36255,nx36397,nx36539,nx36681,
            nx36823,nx36965,nx37107,nx37249,nx37391,nx37533,nx37675,nx37817,
            nx37959,nx38101}), .B ({nx33727,nx33867,nx34005,nx34143,nx34281,
            nx34419,nx34557,nx34697,nx34839,nx34981,nx35123,nx35265,nx35407,
            nx35549,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35691), .C ({inputRegisters_307__15,inputRegisters_307__14,
            inputRegisters_307__13,inputRegisters_307__12,inputRegisters_307__11
            ,inputRegisters_307__10,inputRegisters_307__9,inputRegisters_307__8,
            inputRegisters_307__7,inputRegisters_307__6,inputRegisters_307__5,
            inputRegisters_307__4,inputRegisters_307__3,inputRegisters_307__2,
            inputRegisters_307__1,inputRegisters_307__0})) ;
    Reg_16 loop1_307_x (.D ({inputRegisters_307__15,inputRegisters_307__14,
           inputRegisters_307__13,inputRegisters_307__12,inputRegisters_307__11,
           inputRegisters_307__10,inputRegisters_307__9,inputRegisters_307__8,
           inputRegisters_307__7,inputRegisters_307__6,inputRegisters_307__5,
           inputRegisters_307__4,inputRegisters_307__3,inputRegisters_307__2,
           inputRegisters_307__1,inputRegisters_307__0}), .en (
           enableRegister_307), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_307__15,registerOutputs_307__14,
           registerOutputs_307__13,registerOutputs_307__12,
           registerOutputs_307__11,registerOutputs_307__10,
           registerOutputs_307__9,registerOutputs_307__8,registerOutputs_307__7,
           registerOutputs_307__6,registerOutputs_307__5,registerOutputs_307__4,
           registerOutputs_307__3,registerOutputs_307__2,registerOutputs_307__1,
           registerOutputs_307__0})) ;
    Mux2_16 loop1_308_y (.A ({nx35973,nx36115,nx36257,nx36399,nx36541,nx36683,
            nx36825,nx36967,nx37109,nx37251,nx37393,nx37535,nx37677,nx37819,
            nx37961,nx38103}), .B ({nx33729,nx33867,nx34005,nx34143,nx34281,
            nx34419,nx34557,nx34699,nx34841,nx34983,nx35125,nx35267,nx35409,
            nx35551,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35693), .C ({inputRegisters_308__15,inputRegisters_308__14,
            inputRegisters_308__13,inputRegisters_308__12,inputRegisters_308__11
            ,inputRegisters_308__10,inputRegisters_308__9,inputRegisters_308__8,
            inputRegisters_308__7,inputRegisters_308__6,inputRegisters_308__5,
            inputRegisters_308__4,inputRegisters_308__3,inputRegisters_308__2,
            inputRegisters_308__1,inputRegisters_308__0})) ;
    Reg_16 loop1_308_x (.D ({inputRegisters_308__15,inputRegisters_308__14,
           inputRegisters_308__13,inputRegisters_308__12,inputRegisters_308__11,
           inputRegisters_308__10,inputRegisters_308__9,inputRegisters_308__8,
           inputRegisters_308__7,inputRegisters_308__6,inputRegisters_308__5,
           inputRegisters_308__4,inputRegisters_308__3,inputRegisters_308__2,
           inputRegisters_308__1,inputRegisters_308__0}), .en (
           enableRegister_308), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_308__15,registerOutputs_308__14,
           registerOutputs_308__13,registerOutputs_308__12,
           registerOutputs_308__11,registerOutputs_308__10,
           registerOutputs_308__9,registerOutputs_308__8,registerOutputs_308__7,
           registerOutputs_308__6,registerOutputs_308__5,registerOutputs_308__4,
           registerOutputs_308__3,registerOutputs_308__2,registerOutputs_308__1,
           registerOutputs_308__0})) ;
    Mux2_16 loop1_309_y (.A ({nx35973,nx36115,nx36257,nx36399,nx36541,nx36683,
            nx36825,nx36967,nx37109,nx37251,nx37393,nx37535,nx37677,nx37819,
            nx37961,nx38103}), .B ({nx33729,nx33867,nx34005,nx34143,nx34281,
            nx34419,nx34559,nx34699,nx34841,nx34983,nx35125,nx35267,nx35409,
            nx35551,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35693), .C ({inputRegisters_309__15,inputRegisters_309__14,
            inputRegisters_309__13,inputRegisters_309__12,inputRegisters_309__11
            ,inputRegisters_309__10,inputRegisters_309__9,inputRegisters_309__8,
            inputRegisters_309__7,inputRegisters_309__6,inputRegisters_309__5,
            inputRegisters_309__4,inputRegisters_309__3,inputRegisters_309__2,
            inputRegisters_309__1,inputRegisters_309__0})) ;
    Reg_16 loop1_309_x (.D ({inputRegisters_309__15,inputRegisters_309__14,
           inputRegisters_309__13,inputRegisters_309__12,inputRegisters_309__11,
           inputRegisters_309__10,inputRegisters_309__9,inputRegisters_309__8,
           inputRegisters_309__7,inputRegisters_309__6,inputRegisters_309__5,
           inputRegisters_309__4,inputRegisters_309__3,inputRegisters_309__2,
           inputRegisters_309__1,inputRegisters_309__0}), .en (
           enableRegister_309), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_309__15,registerOutputs_309__14,
           registerOutputs_309__13,registerOutputs_309__12,
           registerOutputs_309__11,registerOutputs_309__10,
           registerOutputs_309__9,registerOutputs_309__8,registerOutputs_309__7,
           registerOutputs_309__6,registerOutputs_309__5,registerOutputs_309__4,
           registerOutputs_309__3,registerOutputs_309__2,registerOutputs_309__1,
           registerOutputs_309__0})) ;
    Mux2_16 loop1_310_y (.A ({nx35973,nx36115,nx36257,nx36399,nx36541,nx36683,
            nx36825,nx36967,nx37109,nx37251,nx37393,nx37535,nx37677,nx37819,
            nx37961,nx38103}), .B ({nx33729,nx33867,nx34005,nx34143,nx34281,
            nx34421,nx34559,nx34699,nx34841,nx34983,nx35125,nx35267,nx35409,
            nx35551,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35693), .C ({inputRegisters_310__15,inputRegisters_310__14,
            inputRegisters_310__13,inputRegisters_310__12,inputRegisters_310__11
            ,inputRegisters_310__10,inputRegisters_310__9,inputRegisters_310__8,
            inputRegisters_310__7,inputRegisters_310__6,inputRegisters_310__5,
            inputRegisters_310__4,inputRegisters_310__3,inputRegisters_310__2,
            inputRegisters_310__1,inputRegisters_310__0})) ;
    Reg_16 loop1_310_x (.D ({inputRegisters_310__15,inputRegisters_310__14,
           inputRegisters_310__13,inputRegisters_310__12,inputRegisters_310__11,
           inputRegisters_310__10,inputRegisters_310__9,inputRegisters_310__8,
           inputRegisters_310__7,inputRegisters_310__6,inputRegisters_310__5,
           inputRegisters_310__4,inputRegisters_310__3,inputRegisters_310__2,
           inputRegisters_310__1,inputRegisters_310__0}), .en (
           enableRegister_310), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_310__15,registerOutputs_310__14,
           registerOutputs_310__13,registerOutputs_310__12,
           registerOutputs_310__11,registerOutputs_310__10,
           registerOutputs_310__9,registerOutputs_310__8,registerOutputs_310__7,
           registerOutputs_310__6,registerOutputs_310__5,registerOutputs_310__4,
           registerOutputs_310__3,registerOutputs_310__2,registerOutputs_310__1,
           registerOutputs_310__0})) ;
    Mux2_16 loop1_311_y (.A ({nx35973,nx36115,nx36257,nx36399,nx36541,nx36683,
            nx36825,nx36967,nx37109,nx37251,nx37393,nx37535,nx37677,nx37819,
            nx37961,nx38103}), .B ({nx33729,nx33867,nx34005,nx34143,nx34283,
            nx34421,nx34559,nx34699,nx34841,nx34983,nx35125,nx35267,nx35409,
            nx35551,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35693), .C ({inputRegisters_311__15,inputRegisters_311__14,
            inputRegisters_311__13,inputRegisters_311__12,inputRegisters_311__11
            ,inputRegisters_311__10,inputRegisters_311__9,inputRegisters_311__8,
            inputRegisters_311__7,inputRegisters_311__6,inputRegisters_311__5,
            inputRegisters_311__4,inputRegisters_311__3,inputRegisters_311__2,
            inputRegisters_311__1,inputRegisters_311__0})) ;
    Reg_16 loop1_311_x (.D ({inputRegisters_311__15,inputRegisters_311__14,
           inputRegisters_311__13,inputRegisters_311__12,inputRegisters_311__11,
           inputRegisters_311__10,inputRegisters_311__9,inputRegisters_311__8,
           inputRegisters_311__7,inputRegisters_311__6,inputRegisters_311__5,
           inputRegisters_311__4,inputRegisters_311__3,inputRegisters_311__2,
           inputRegisters_311__1,inputRegisters_311__0}), .en (
           enableRegister_311), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_311__15,registerOutputs_311__14,
           registerOutputs_311__13,registerOutputs_311__12,
           registerOutputs_311__11,registerOutputs_311__10,
           registerOutputs_311__9,registerOutputs_311__8,registerOutputs_311__7,
           registerOutputs_311__6,registerOutputs_311__5,registerOutputs_311__4,
           registerOutputs_311__3,registerOutputs_311__2,registerOutputs_311__1,
           registerOutputs_311__0})) ;
    Mux2_16 loop1_312_y (.A ({nx35973,nx36115,nx36257,nx36399,nx36541,nx36683,
            nx36825,nx36967,nx37109,nx37251,nx37393,nx37535,nx37677,nx37819,
            nx37961,nx38103}), .B ({nx33729,nx33867,nx34005,nx34145,nx34283,
            nx34421,nx34559,nx34699,nx34841,nx34983,nx35125,nx35267,nx35409,
            nx35551,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35693), .C ({inputRegisters_312__15,inputRegisters_312__14,
            inputRegisters_312__13,inputRegisters_312__12,inputRegisters_312__11
            ,inputRegisters_312__10,inputRegisters_312__9,inputRegisters_312__8,
            inputRegisters_312__7,inputRegisters_312__6,inputRegisters_312__5,
            inputRegisters_312__4,inputRegisters_312__3,inputRegisters_312__2,
            inputRegisters_312__1,inputRegisters_312__0})) ;
    Reg_16 loop1_312_x (.D ({inputRegisters_312__15,inputRegisters_312__14,
           inputRegisters_312__13,inputRegisters_312__12,inputRegisters_312__11,
           inputRegisters_312__10,inputRegisters_312__9,inputRegisters_312__8,
           inputRegisters_312__7,inputRegisters_312__6,inputRegisters_312__5,
           inputRegisters_312__4,inputRegisters_312__3,inputRegisters_312__2,
           inputRegisters_312__1,inputRegisters_312__0}), .en (
           enableRegister_312), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_312__15,registerOutputs_312__14,
           registerOutputs_312__13,registerOutputs_312__12,
           registerOutputs_312__11,registerOutputs_312__10,
           registerOutputs_312__9,registerOutputs_312__8,registerOutputs_312__7,
           registerOutputs_312__6,registerOutputs_312__5,registerOutputs_312__4,
           registerOutputs_312__3,registerOutputs_312__2,registerOutputs_312__1,
           registerOutputs_312__0})) ;
    Mux2_16 loop1_313_y (.A ({nx35973,nx36115,nx36257,nx36399,nx36541,nx36683,
            nx36825,nx36967,nx37109,nx37251,nx37393,nx37535,nx37677,nx37819,
            nx37961,nx38103}), .B ({nx33729,nx33867,nx34007,nx34145,nx34283,
            nx34421,nx34559,nx34699,nx34841,nx34983,nx35125,nx35267,nx35409,
            nx35551,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35693), .C ({inputRegisters_313__15,inputRegisters_313__14,
            inputRegisters_313__13,inputRegisters_313__12,inputRegisters_313__11
            ,inputRegisters_313__10,inputRegisters_313__9,inputRegisters_313__8,
            inputRegisters_313__7,inputRegisters_313__6,inputRegisters_313__5,
            inputRegisters_313__4,inputRegisters_313__3,inputRegisters_313__2,
            inputRegisters_313__1,inputRegisters_313__0})) ;
    Reg_16 loop1_313_x (.D ({inputRegisters_313__15,inputRegisters_313__14,
           inputRegisters_313__13,inputRegisters_313__12,inputRegisters_313__11,
           inputRegisters_313__10,inputRegisters_313__9,inputRegisters_313__8,
           inputRegisters_313__7,inputRegisters_313__6,inputRegisters_313__5,
           inputRegisters_313__4,inputRegisters_313__3,inputRegisters_313__2,
           inputRegisters_313__1,inputRegisters_313__0}), .en (
           enableRegister_313), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_313__15,registerOutputs_313__14,
           registerOutputs_313__13,registerOutputs_313__12,
           registerOutputs_313__11,registerOutputs_313__10,
           registerOutputs_313__9,registerOutputs_313__8,registerOutputs_313__7,
           registerOutputs_313__6,registerOutputs_313__5,registerOutputs_313__4,
           registerOutputs_313__3,registerOutputs_313__2,registerOutputs_313__1,
           registerOutputs_313__0})) ;
    Mux2_16 loop1_314_y (.A ({nx35973,nx36115,nx36257,nx36399,nx36541,nx36683,
            nx36825,nx36967,nx37109,nx37251,nx37393,nx37535,nx37677,nx37819,
            nx37961,nx38103}), .B ({nx33729,nx33869,nx34007,nx34145,nx34283,
            nx34421,nx34559,nx34699,nx34841,nx34983,nx35125,nx35267,nx35409,
            nx35551,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35693), .C ({inputRegisters_314__15,inputRegisters_314__14,
            inputRegisters_314__13,inputRegisters_314__12,inputRegisters_314__11
            ,inputRegisters_314__10,inputRegisters_314__9,inputRegisters_314__8,
            inputRegisters_314__7,inputRegisters_314__6,inputRegisters_314__5,
            inputRegisters_314__4,inputRegisters_314__3,inputRegisters_314__2,
            inputRegisters_314__1,inputRegisters_314__0})) ;
    Reg_16 loop1_314_x (.D ({inputRegisters_314__15,inputRegisters_314__14,
           inputRegisters_314__13,inputRegisters_314__12,inputRegisters_314__11,
           inputRegisters_314__10,inputRegisters_314__9,inputRegisters_314__8,
           inputRegisters_314__7,inputRegisters_314__6,inputRegisters_314__5,
           inputRegisters_314__4,inputRegisters_314__3,inputRegisters_314__2,
           inputRegisters_314__1,inputRegisters_314__0}), .en (
           enableRegister_314), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_314__15,registerOutputs_314__14,
           registerOutputs_314__13,registerOutputs_314__12,
           registerOutputs_314__11,registerOutputs_314__10,
           registerOutputs_314__9,registerOutputs_314__8,registerOutputs_314__7,
           registerOutputs_314__6,registerOutputs_314__5,registerOutputs_314__4,
           registerOutputs_314__3,registerOutputs_314__2,registerOutputs_314__1,
           registerOutputs_314__0})) ;
    Mux2_16 loop1_315_y (.A ({nx35975,nx36117,nx36259,nx36401,nx36543,nx36685,
            nx36827,nx36969,nx37111,nx37253,nx37395,nx37537,nx37679,nx37821,
            nx37963,nx38105}), .B ({nx33731,nx33869,nx34007,nx34145,nx34283,
            nx34421,nx34559,nx34701,nx34843,nx34985,nx35127,nx35269,nx35411,
            nx35553,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35695), .C ({inputRegisters_315__15,inputRegisters_315__14,
            inputRegisters_315__13,inputRegisters_315__12,inputRegisters_315__11
            ,inputRegisters_315__10,inputRegisters_315__9,inputRegisters_315__8,
            inputRegisters_315__7,inputRegisters_315__6,inputRegisters_315__5,
            inputRegisters_315__4,inputRegisters_315__3,inputRegisters_315__2,
            inputRegisters_315__1,inputRegisters_315__0})) ;
    Reg_16 loop1_315_x (.D ({inputRegisters_315__15,inputRegisters_315__14,
           inputRegisters_315__13,inputRegisters_315__12,inputRegisters_315__11,
           inputRegisters_315__10,inputRegisters_315__9,inputRegisters_315__8,
           inputRegisters_315__7,inputRegisters_315__6,inputRegisters_315__5,
           inputRegisters_315__4,inputRegisters_315__3,inputRegisters_315__2,
           inputRegisters_315__1,inputRegisters_315__0}), .en (
           enableRegister_315), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_315__15,registerOutputs_315__14,
           registerOutputs_315__13,registerOutputs_315__12,
           registerOutputs_315__11,registerOutputs_315__10,
           registerOutputs_315__9,registerOutputs_315__8,registerOutputs_315__7,
           registerOutputs_315__6,registerOutputs_315__5,registerOutputs_315__4,
           registerOutputs_315__3,registerOutputs_315__2,registerOutputs_315__1,
           registerOutputs_315__0})) ;
    Mux2_16 loop1_316_y (.A ({nx35975,nx36117,nx36259,nx36401,nx36543,nx36685,
            nx36827,nx36969,nx37111,nx37253,nx37395,nx37537,nx37679,nx37821,
            nx37963,nx38105}), .B ({nx33731,nx33869,nx34007,nx34145,nx34283,
            nx34421,nx34561,nx34701,nx34843,nx34985,nx35127,nx35269,nx35411,
            nx35553,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35695), .C ({inputRegisters_316__15,inputRegisters_316__14,
            inputRegisters_316__13,inputRegisters_316__12,inputRegisters_316__11
            ,inputRegisters_316__10,inputRegisters_316__9,inputRegisters_316__8,
            inputRegisters_316__7,inputRegisters_316__6,inputRegisters_316__5,
            inputRegisters_316__4,inputRegisters_316__3,inputRegisters_316__2,
            inputRegisters_316__1,inputRegisters_316__0})) ;
    Reg_16 loop1_316_x (.D ({inputRegisters_316__15,inputRegisters_316__14,
           inputRegisters_316__13,inputRegisters_316__12,inputRegisters_316__11,
           inputRegisters_316__10,inputRegisters_316__9,inputRegisters_316__8,
           inputRegisters_316__7,inputRegisters_316__6,inputRegisters_316__5,
           inputRegisters_316__4,inputRegisters_316__3,inputRegisters_316__2,
           inputRegisters_316__1,inputRegisters_316__0}), .en (
           enableRegister_316), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_316__15,registerOutputs_316__14,
           registerOutputs_316__13,registerOutputs_316__12,
           registerOutputs_316__11,registerOutputs_316__10,
           registerOutputs_316__9,registerOutputs_316__8,registerOutputs_316__7,
           registerOutputs_316__6,registerOutputs_316__5,registerOutputs_316__4,
           registerOutputs_316__3,registerOutputs_316__2,registerOutputs_316__1,
           registerOutputs_316__0})) ;
    Mux2_16 loop1_317_y (.A ({nx35975,nx36117,nx36259,nx36401,nx36543,nx36685,
            nx36827,nx36969,nx37111,nx37253,nx37395,nx37537,nx37679,nx37821,
            nx37963,nx38105}), .B ({nx33731,nx33869,nx34007,nx34145,nx34283,
            nx34423,nx34561,nx34701,nx34843,nx34985,nx35127,nx35269,nx35411,
            nx35553,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35695), .C ({inputRegisters_317__15,inputRegisters_317__14,
            inputRegisters_317__13,inputRegisters_317__12,inputRegisters_317__11
            ,inputRegisters_317__10,inputRegisters_317__9,inputRegisters_317__8,
            inputRegisters_317__7,inputRegisters_317__6,inputRegisters_317__5,
            inputRegisters_317__4,inputRegisters_317__3,inputRegisters_317__2,
            inputRegisters_317__1,inputRegisters_317__0})) ;
    Reg_16 loop1_317_x (.D ({inputRegisters_317__15,inputRegisters_317__14,
           inputRegisters_317__13,inputRegisters_317__12,inputRegisters_317__11,
           inputRegisters_317__10,inputRegisters_317__9,inputRegisters_317__8,
           inputRegisters_317__7,inputRegisters_317__6,inputRegisters_317__5,
           inputRegisters_317__4,inputRegisters_317__3,inputRegisters_317__2,
           inputRegisters_317__1,inputRegisters_317__0}), .en (
           enableRegister_317), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_317__15,registerOutputs_317__14,
           registerOutputs_317__13,registerOutputs_317__12,
           registerOutputs_317__11,registerOutputs_317__10,
           registerOutputs_317__9,registerOutputs_317__8,registerOutputs_317__7,
           registerOutputs_317__6,registerOutputs_317__5,registerOutputs_317__4,
           registerOutputs_317__3,registerOutputs_317__2,registerOutputs_317__1,
           registerOutputs_317__0})) ;
    Mux2_16 loop1_318_y (.A ({nx35975,nx36117,nx36259,nx36401,nx36543,nx36685,
            nx36827,nx36969,nx37111,nx37253,nx37395,nx37537,nx37679,nx37821,
            nx37963,nx38105}), .B ({nx33731,nx33869,nx34007,nx34145,nx34285,
            nx34423,nx34561,nx34701,nx34843,nx34985,nx35127,nx35269,nx35411,
            nx35553,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35695), .C ({inputRegisters_318__15,inputRegisters_318__14,
            inputRegisters_318__13,inputRegisters_318__12,inputRegisters_318__11
            ,inputRegisters_318__10,inputRegisters_318__9,inputRegisters_318__8,
            inputRegisters_318__7,inputRegisters_318__6,inputRegisters_318__5,
            inputRegisters_318__4,inputRegisters_318__3,inputRegisters_318__2,
            inputRegisters_318__1,inputRegisters_318__0})) ;
    Reg_16 loop1_318_x (.D ({inputRegisters_318__15,inputRegisters_318__14,
           inputRegisters_318__13,inputRegisters_318__12,inputRegisters_318__11,
           inputRegisters_318__10,inputRegisters_318__9,inputRegisters_318__8,
           inputRegisters_318__7,inputRegisters_318__6,inputRegisters_318__5,
           inputRegisters_318__4,inputRegisters_318__3,inputRegisters_318__2,
           inputRegisters_318__1,inputRegisters_318__0}), .en (
           enableRegister_318), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_318__15,registerOutputs_318__14,
           registerOutputs_318__13,registerOutputs_318__12,
           registerOutputs_318__11,registerOutputs_318__10,
           registerOutputs_318__9,registerOutputs_318__8,registerOutputs_318__7,
           registerOutputs_318__6,registerOutputs_318__5,registerOutputs_318__4,
           registerOutputs_318__3,registerOutputs_318__2,registerOutputs_318__1,
           registerOutputs_318__0})) ;
    Mux2_16 loop1_319_y (.A ({nx35975,nx36117,nx36259,nx36401,nx36543,nx36685,
            nx36827,nx36969,nx37111,nx37253,nx37395,nx37537,nx37679,nx37821,
            nx37963,nx38105}), .B ({nx33731,nx33869,nx34007,nx34147,nx34285,
            nx34423,nx34561,nx34701,nx34843,nx34985,nx35127,nx35269,nx35411,
            nx35553,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35695), .C ({inputRegisters_319__15,inputRegisters_319__14,
            inputRegisters_319__13,inputRegisters_319__12,inputRegisters_319__11
            ,inputRegisters_319__10,inputRegisters_319__9,inputRegisters_319__8,
            inputRegisters_319__7,inputRegisters_319__6,inputRegisters_319__5,
            inputRegisters_319__4,inputRegisters_319__3,inputRegisters_319__2,
            inputRegisters_319__1,inputRegisters_319__0})) ;
    Reg_16 loop1_319_x (.D ({inputRegisters_319__15,inputRegisters_319__14,
           inputRegisters_319__13,inputRegisters_319__12,inputRegisters_319__11,
           inputRegisters_319__10,inputRegisters_319__9,inputRegisters_319__8,
           inputRegisters_319__7,inputRegisters_319__6,inputRegisters_319__5,
           inputRegisters_319__4,inputRegisters_319__3,inputRegisters_319__2,
           inputRegisters_319__1,inputRegisters_319__0}), .en (
           enableRegister_319), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_319__15,registerOutputs_319__14,
           registerOutputs_319__13,registerOutputs_319__12,
           registerOutputs_319__11,registerOutputs_319__10,
           registerOutputs_319__9,registerOutputs_319__8,registerOutputs_319__7,
           registerOutputs_319__6,registerOutputs_319__5,registerOutputs_319__4,
           registerOutputs_319__3,registerOutputs_319__2,registerOutputs_319__1,
           registerOutputs_319__0})) ;
    Mux2_16 loop1_320_y (.A ({nx35975,nx36117,nx36259,nx36401,nx36543,nx36685,
            nx36827,nx36969,nx37111,nx37253,nx37395,nx37537,nx37679,nx37821,
            nx37963,nx38105}), .B ({nx33731,nx33869,nx34009,nx34147,nx34285,
            nx34423,nx34561,nx34701,nx34843,nx34985,nx35127,nx35269,nx35411,
            nx35553,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35695), .C ({inputRegisters_320__15,inputRegisters_320__14,
            inputRegisters_320__13,inputRegisters_320__12,inputRegisters_320__11
            ,inputRegisters_320__10,inputRegisters_320__9,inputRegisters_320__8,
            inputRegisters_320__7,inputRegisters_320__6,inputRegisters_320__5,
            inputRegisters_320__4,inputRegisters_320__3,inputRegisters_320__2,
            inputRegisters_320__1,inputRegisters_320__0})) ;
    Reg_16 loop1_320_x (.D ({inputRegisters_320__15,inputRegisters_320__14,
           inputRegisters_320__13,inputRegisters_320__12,inputRegisters_320__11,
           inputRegisters_320__10,inputRegisters_320__9,inputRegisters_320__8,
           inputRegisters_320__7,inputRegisters_320__6,inputRegisters_320__5,
           inputRegisters_320__4,inputRegisters_320__3,inputRegisters_320__2,
           inputRegisters_320__1,inputRegisters_320__0}), .en (
           enableRegister_320), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_320__15,registerOutputs_320__14,
           registerOutputs_320__13,registerOutputs_320__12,
           registerOutputs_320__11,registerOutputs_320__10,
           registerOutputs_320__9,registerOutputs_320__8,registerOutputs_320__7,
           registerOutputs_320__6,registerOutputs_320__5,registerOutputs_320__4,
           registerOutputs_320__3,registerOutputs_320__2,registerOutputs_320__1,
           registerOutputs_320__0})) ;
    Mux2_16 loop1_321_y (.A ({nx35975,nx36117,nx36259,nx36401,nx36543,nx36685,
            nx36827,nx36969,nx37111,nx37253,nx37395,nx37537,nx37679,nx37821,
            nx37963,nx38105}), .B ({nx33731,nx33871,nx34009,nx34147,nx34285,
            nx34423,nx34561,nx34701,nx34843,nx34985,nx35127,nx35269,nx35411,
            nx35553,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35695), .C ({inputRegisters_321__15,inputRegisters_321__14,
            inputRegisters_321__13,inputRegisters_321__12,inputRegisters_321__11
            ,inputRegisters_321__10,inputRegisters_321__9,inputRegisters_321__8,
            inputRegisters_321__7,inputRegisters_321__6,inputRegisters_321__5,
            inputRegisters_321__4,inputRegisters_321__3,inputRegisters_321__2,
            inputRegisters_321__1,inputRegisters_321__0})) ;
    Reg_16 loop1_321_x (.D ({inputRegisters_321__15,inputRegisters_321__14,
           inputRegisters_321__13,inputRegisters_321__12,inputRegisters_321__11,
           inputRegisters_321__10,inputRegisters_321__9,inputRegisters_321__8,
           inputRegisters_321__7,inputRegisters_321__6,inputRegisters_321__5,
           inputRegisters_321__4,inputRegisters_321__3,inputRegisters_321__2,
           inputRegisters_321__1,inputRegisters_321__0}), .en (
           enableRegister_321), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_321__15,registerOutputs_321__14,
           registerOutputs_321__13,registerOutputs_321__12,
           registerOutputs_321__11,registerOutputs_321__10,
           registerOutputs_321__9,registerOutputs_321__8,registerOutputs_321__7,
           registerOutputs_321__6,registerOutputs_321__5,registerOutputs_321__4,
           registerOutputs_321__3,registerOutputs_321__2,registerOutputs_321__1,
           registerOutputs_321__0})) ;
    Mux2_16 loop1_322_y (.A ({nx35977,nx36119,nx36261,nx36403,nx36545,nx36687,
            nx36829,nx36971,nx37113,nx37255,nx37397,nx37539,nx37681,nx37823,
            nx37965,nx38107}), .B ({nx33733,nx33871,nx34009,nx34147,nx34285,
            nx34423,nx34561,nx34703,nx34845,nx34987,nx35129,nx35271,nx35413,
            nx35555,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35697), .C ({inputRegisters_322__15,inputRegisters_322__14,
            inputRegisters_322__13,inputRegisters_322__12,inputRegisters_322__11
            ,inputRegisters_322__10,inputRegisters_322__9,inputRegisters_322__8,
            inputRegisters_322__7,inputRegisters_322__6,inputRegisters_322__5,
            inputRegisters_322__4,inputRegisters_322__3,inputRegisters_322__2,
            inputRegisters_322__1,inputRegisters_322__0})) ;
    Reg_16 loop1_322_x (.D ({inputRegisters_322__15,inputRegisters_322__14,
           inputRegisters_322__13,inputRegisters_322__12,inputRegisters_322__11,
           inputRegisters_322__10,inputRegisters_322__9,inputRegisters_322__8,
           inputRegisters_322__7,inputRegisters_322__6,inputRegisters_322__5,
           inputRegisters_322__4,inputRegisters_322__3,inputRegisters_322__2,
           inputRegisters_322__1,inputRegisters_322__0}), .en (
           enableRegister_322), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_322__15,registerOutputs_322__14,
           registerOutputs_322__13,registerOutputs_322__12,
           registerOutputs_322__11,registerOutputs_322__10,
           registerOutputs_322__9,registerOutputs_322__8,registerOutputs_322__7,
           registerOutputs_322__6,registerOutputs_322__5,registerOutputs_322__4,
           registerOutputs_322__3,registerOutputs_322__2,registerOutputs_322__1,
           registerOutputs_322__0})) ;
    Mux2_16 loop1_323_y (.A ({nx35977,nx36119,nx36261,nx36403,nx36545,nx36687,
            nx36829,nx36971,nx37113,nx37255,nx37397,nx37539,nx37681,nx37823,
            nx37965,nx38107}), .B ({nx33733,nx33871,nx34009,nx34147,nx34285,
            nx34423,nx34563,nx34703,nx34845,nx34987,nx35129,nx35271,nx35413,
            nx35555,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35697), .C ({inputRegisters_323__15,inputRegisters_323__14,
            inputRegisters_323__13,inputRegisters_323__12,inputRegisters_323__11
            ,inputRegisters_323__10,inputRegisters_323__9,inputRegisters_323__8,
            inputRegisters_323__7,inputRegisters_323__6,inputRegisters_323__5,
            inputRegisters_323__4,inputRegisters_323__3,inputRegisters_323__2,
            inputRegisters_323__1,inputRegisters_323__0})) ;
    Reg_16 loop1_323_x (.D ({inputRegisters_323__15,inputRegisters_323__14,
           inputRegisters_323__13,inputRegisters_323__12,inputRegisters_323__11,
           inputRegisters_323__10,inputRegisters_323__9,inputRegisters_323__8,
           inputRegisters_323__7,inputRegisters_323__6,inputRegisters_323__5,
           inputRegisters_323__4,inputRegisters_323__3,inputRegisters_323__2,
           inputRegisters_323__1,inputRegisters_323__0}), .en (
           enableRegister_323), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_323__15,registerOutputs_323__14,
           registerOutputs_323__13,registerOutputs_323__12,
           registerOutputs_323__11,registerOutputs_323__10,
           registerOutputs_323__9,registerOutputs_323__8,registerOutputs_323__7,
           registerOutputs_323__6,registerOutputs_323__5,registerOutputs_323__4,
           registerOutputs_323__3,registerOutputs_323__2,registerOutputs_323__1,
           registerOutputs_323__0})) ;
    Mux2_16 loop1_324_y (.A ({nx35977,nx36119,nx36261,nx36403,nx36545,nx36687,
            nx36829,nx36971,nx37113,nx37255,nx37397,nx37539,nx37681,nx37823,
            nx37965,nx38107}), .B ({nx33733,nx33871,nx34009,nx34147,nx34285,
            nx34425,nx34563,nx34703,nx34845,nx34987,nx35129,nx35271,nx35413,
            nx35555,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35697), .C ({inputRegisters_324__15,inputRegisters_324__14,
            inputRegisters_324__13,inputRegisters_324__12,inputRegisters_324__11
            ,inputRegisters_324__10,inputRegisters_324__9,inputRegisters_324__8,
            inputRegisters_324__7,inputRegisters_324__6,inputRegisters_324__5,
            inputRegisters_324__4,inputRegisters_324__3,inputRegisters_324__2,
            inputRegisters_324__1,inputRegisters_324__0})) ;
    Reg_16 loop1_324_x (.D ({inputRegisters_324__15,inputRegisters_324__14,
           inputRegisters_324__13,inputRegisters_324__12,inputRegisters_324__11,
           inputRegisters_324__10,inputRegisters_324__9,inputRegisters_324__8,
           inputRegisters_324__7,inputRegisters_324__6,inputRegisters_324__5,
           inputRegisters_324__4,inputRegisters_324__3,inputRegisters_324__2,
           inputRegisters_324__1,inputRegisters_324__0}), .en (
           enableRegister_324), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_324__15,registerOutputs_324__14,
           registerOutputs_324__13,registerOutputs_324__12,
           registerOutputs_324__11,registerOutputs_324__10,
           registerOutputs_324__9,registerOutputs_324__8,registerOutputs_324__7,
           registerOutputs_324__6,registerOutputs_324__5,registerOutputs_324__4,
           registerOutputs_324__3,registerOutputs_324__2,registerOutputs_324__1,
           registerOutputs_324__0})) ;
    Mux2_16 loop1_325_y (.A ({nx35977,nx36119,nx36261,nx36403,nx36545,nx36687,
            nx36829,nx36971,nx37113,nx37255,nx37397,nx37539,nx37681,nx37823,
            nx37965,nx38107}), .B ({nx33733,nx33871,nx34009,nx34147,nx34287,
            nx34425,nx34563,nx34703,nx34845,nx34987,nx35129,nx35271,nx35413,
            nx35555,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35697), .C ({inputRegisters_325__15,inputRegisters_325__14,
            inputRegisters_325__13,inputRegisters_325__12,inputRegisters_325__11
            ,inputRegisters_325__10,inputRegisters_325__9,inputRegisters_325__8,
            inputRegisters_325__7,inputRegisters_325__6,inputRegisters_325__5,
            inputRegisters_325__4,inputRegisters_325__3,inputRegisters_325__2,
            inputRegisters_325__1,inputRegisters_325__0})) ;
    Reg_16 loop1_325_x (.D ({inputRegisters_325__15,inputRegisters_325__14,
           inputRegisters_325__13,inputRegisters_325__12,inputRegisters_325__11,
           inputRegisters_325__10,inputRegisters_325__9,inputRegisters_325__8,
           inputRegisters_325__7,inputRegisters_325__6,inputRegisters_325__5,
           inputRegisters_325__4,inputRegisters_325__3,inputRegisters_325__2,
           inputRegisters_325__1,inputRegisters_325__0}), .en (
           enableRegister_325), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_325__15,registerOutputs_325__14,
           registerOutputs_325__13,registerOutputs_325__12,
           registerOutputs_325__11,registerOutputs_325__10,
           registerOutputs_325__9,registerOutputs_325__8,registerOutputs_325__7,
           registerOutputs_325__6,registerOutputs_325__5,registerOutputs_325__4,
           registerOutputs_325__3,registerOutputs_325__2,registerOutputs_325__1,
           registerOutputs_325__0})) ;
    Mux2_16 loop1_326_y (.A ({nx35977,nx36119,nx36261,nx36403,nx36545,nx36687,
            nx36829,nx36971,nx37113,nx37255,nx37397,nx37539,nx37681,nx37823,
            nx37965,nx38107}), .B ({nx33733,nx33871,nx34009,nx34149,nx34287,
            nx34425,nx34563,nx34703,nx34845,nx34987,nx35129,nx35271,nx35413,
            nx35555,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35697), .C ({inputRegisters_326__15,inputRegisters_326__14,
            inputRegisters_326__13,inputRegisters_326__12,inputRegisters_326__11
            ,inputRegisters_326__10,inputRegisters_326__9,inputRegisters_326__8,
            inputRegisters_326__7,inputRegisters_326__6,inputRegisters_326__5,
            inputRegisters_326__4,inputRegisters_326__3,inputRegisters_326__2,
            inputRegisters_326__1,inputRegisters_326__0})) ;
    Reg_16 loop1_326_x (.D ({inputRegisters_326__15,inputRegisters_326__14,
           inputRegisters_326__13,inputRegisters_326__12,inputRegisters_326__11,
           inputRegisters_326__10,inputRegisters_326__9,inputRegisters_326__8,
           inputRegisters_326__7,inputRegisters_326__6,inputRegisters_326__5,
           inputRegisters_326__4,inputRegisters_326__3,inputRegisters_326__2,
           inputRegisters_326__1,inputRegisters_326__0}), .en (
           enableRegister_326), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_326__15,registerOutputs_326__14,
           registerOutputs_326__13,registerOutputs_326__12,
           registerOutputs_326__11,registerOutputs_326__10,
           registerOutputs_326__9,registerOutputs_326__8,registerOutputs_326__7,
           registerOutputs_326__6,registerOutputs_326__5,registerOutputs_326__4,
           registerOutputs_326__3,registerOutputs_326__2,registerOutputs_326__1,
           registerOutputs_326__0})) ;
    Mux2_16 loop1_327_y (.A ({nx35977,nx36119,nx36261,nx36403,nx36545,nx36687,
            nx36829,nx36971,nx37113,nx37255,nx37397,nx37539,nx37681,nx37823,
            nx37965,nx38107}), .B ({nx33733,nx33871,nx34011,nx34149,nx34287,
            nx34425,nx34563,nx34703,nx34845,nx34987,nx35129,nx35271,nx35413,
            nx35555,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35697), .C ({inputRegisters_327__15,inputRegisters_327__14,
            inputRegisters_327__13,inputRegisters_327__12,inputRegisters_327__11
            ,inputRegisters_327__10,inputRegisters_327__9,inputRegisters_327__8,
            inputRegisters_327__7,inputRegisters_327__6,inputRegisters_327__5,
            inputRegisters_327__4,inputRegisters_327__3,inputRegisters_327__2,
            inputRegisters_327__1,inputRegisters_327__0})) ;
    Reg_16 loop1_327_x (.D ({inputRegisters_327__15,inputRegisters_327__14,
           inputRegisters_327__13,inputRegisters_327__12,inputRegisters_327__11,
           inputRegisters_327__10,inputRegisters_327__9,inputRegisters_327__8,
           inputRegisters_327__7,inputRegisters_327__6,inputRegisters_327__5,
           inputRegisters_327__4,inputRegisters_327__3,inputRegisters_327__2,
           inputRegisters_327__1,inputRegisters_327__0}), .en (
           enableRegister_327), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_327__15,registerOutputs_327__14,
           registerOutputs_327__13,registerOutputs_327__12,
           registerOutputs_327__11,registerOutputs_327__10,
           registerOutputs_327__9,registerOutputs_327__8,registerOutputs_327__7,
           registerOutputs_327__6,registerOutputs_327__5,registerOutputs_327__4,
           registerOutputs_327__3,registerOutputs_327__2,registerOutputs_327__1,
           registerOutputs_327__0})) ;
    Mux2_16 loop1_328_y (.A ({nx35977,nx36119,nx36261,nx36403,nx36545,nx36687,
            nx36829,nx36971,nx37113,nx37255,nx37397,nx37539,nx37681,nx37823,
            nx37965,nx38107}), .B ({nx33733,nx33873,nx34011,nx34149,nx34287,
            nx34425,nx34563,nx34703,nx34845,nx34987,nx35129,nx35271,nx35413,
            nx35555,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35697), .C ({inputRegisters_328__15,inputRegisters_328__14,
            inputRegisters_328__13,inputRegisters_328__12,inputRegisters_328__11
            ,inputRegisters_328__10,inputRegisters_328__9,inputRegisters_328__8,
            inputRegisters_328__7,inputRegisters_328__6,inputRegisters_328__5,
            inputRegisters_328__4,inputRegisters_328__3,inputRegisters_328__2,
            inputRegisters_328__1,inputRegisters_328__0})) ;
    Reg_16 loop1_328_x (.D ({inputRegisters_328__15,inputRegisters_328__14,
           inputRegisters_328__13,inputRegisters_328__12,inputRegisters_328__11,
           inputRegisters_328__10,inputRegisters_328__9,inputRegisters_328__8,
           inputRegisters_328__7,inputRegisters_328__6,inputRegisters_328__5,
           inputRegisters_328__4,inputRegisters_328__3,inputRegisters_328__2,
           inputRegisters_328__1,inputRegisters_328__0}), .en (
           enableRegister_328), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_328__15,registerOutputs_328__14,
           registerOutputs_328__13,registerOutputs_328__12,
           registerOutputs_328__11,registerOutputs_328__10,
           registerOutputs_328__9,registerOutputs_328__8,registerOutputs_328__7,
           registerOutputs_328__6,registerOutputs_328__5,registerOutputs_328__4,
           registerOutputs_328__3,registerOutputs_328__2,registerOutputs_328__1,
           registerOutputs_328__0})) ;
    Mux2_16 loop1_329_y (.A ({nx35979,nx36121,nx36263,nx36405,nx36547,nx36689,
            nx36831,nx36973,nx37115,nx37257,nx37399,nx37541,nx37683,nx37825,
            nx37967,nx38109}), .B ({nx33735,nx33873,nx34011,nx34149,nx34287,
            nx34425,nx34563,nx34705,nx34847,nx34989,nx35131,nx35273,nx35415,
            nx35557,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35699), .C ({inputRegisters_329__15,inputRegisters_329__14,
            inputRegisters_329__13,inputRegisters_329__12,inputRegisters_329__11
            ,inputRegisters_329__10,inputRegisters_329__9,inputRegisters_329__8,
            inputRegisters_329__7,inputRegisters_329__6,inputRegisters_329__5,
            inputRegisters_329__4,inputRegisters_329__3,inputRegisters_329__2,
            inputRegisters_329__1,inputRegisters_329__0})) ;
    Reg_16 loop1_329_x (.D ({inputRegisters_329__15,inputRegisters_329__14,
           inputRegisters_329__13,inputRegisters_329__12,inputRegisters_329__11,
           inputRegisters_329__10,inputRegisters_329__9,inputRegisters_329__8,
           inputRegisters_329__7,inputRegisters_329__6,inputRegisters_329__5,
           inputRegisters_329__4,inputRegisters_329__3,inputRegisters_329__2,
           inputRegisters_329__1,inputRegisters_329__0}), .en (
           enableRegister_329), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_329__15,registerOutputs_329__14,
           registerOutputs_329__13,registerOutputs_329__12,
           registerOutputs_329__11,registerOutputs_329__10,
           registerOutputs_329__9,registerOutputs_329__8,registerOutputs_329__7,
           registerOutputs_329__6,registerOutputs_329__5,registerOutputs_329__4,
           registerOutputs_329__3,registerOutputs_329__2,registerOutputs_329__1,
           registerOutputs_329__0})) ;
    Mux2_16 loop1_330_y (.A ({nx35979,nx36121,nx36263,nx36405,nx36547,nx36689,
            nx36831,nx36973,nx37115,nx37257,nx37399,nx37541,nx37683,nx37825,
            nx37967,nx38109}), .B ({nx33735,nx33873,nx34011,nx34149,nx34287,
            nx34425,nx34565,nx34705,nx34847,nx34989,nx35131,nx35273,nx35415,
            nx35557,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35699), .C ({inputRegisters_330__15,inputRegisters_330__14,
            inputRegisters_330__13,inputRegisters_330__12,inputRegisters_330__11
            ,inputRegisters_330__10,inputRegisters_330__9,inputRegisters_330__8,
            inputRegisters_330__7,inputRegisters_330__6,inputRegisters_330__5,
            inputRegisters_330__4,inputRegisters_330__3,inputRegisters_330__2,
            inputRegisters_330__1,inputRegisters_330__0})) ;
    Reg_16 loop1_330_x (.D ({inputRegisters_330__15,inputRegisters_330__14,
           inputRegisters_330__13,inputRegisters_330__12,inputRegisters_330__11,
           inputRegisters_330__10,inputRegisters_330__9,inputRegisters_330__8,
           inputRegisters_330__7,inputRegisters_330__6,inputRegisters_330__5,
           inputRegisters_330__4,inputRegisters_330__3,inputRegisters_330__2,
           inputRegisters_330__1,inputRegisters_330__0}), .en (
           enableRegister_330), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_330__15,registerOutputs_330__14,
           registerOutputs_330__13,registerOutputs_330__12,
           registerOutputs_330__11,registerOutputs_330__10,
           registerOutputs_330__9,registerOutputs_330__8,registerOutputs_330__7,
           registerOutputs_330__6,registerOutputs_330__5,registerOutputs_330__4,
           registerOutputs_330__3,registerOutputs_330__2,registerOutputs_330__1,
           registerOutputs_330__0})) ;
    Mux2_16 loop1_331_y (.A ({nx35979,nx36121,nx36263,nx36405,nx36547,nx36689,
            nx36831,nx36973,nx37115,nx37257,nx37399,nx37541,nx37683,nx37825,
            nx37967,nx38109}), .B ({nx33735,nx33873,nx34011,nx34149,nx34287,
            nx34427,nx34565,nx34705,nx34847,nx34989,nx35131,nx35273,nx35415,
            nx35557,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35699), .C ({inputRegisters_331__15,inputRegisters_331__14,
            inputRegisters_331__13,inputRegisters_331__12,inputRegisters_331__11
            ,inputRegisters_331__10,inputRegisters_331__9,inputRegisters_331__8,
            inputRegisters_331__7,inputRegisters_331__6,inputRegisters_331__5,
            inputRegisters_331__4,inputRegisters_331__3,inputRegisters_331__2,
            inputRegisters_331__1,inputRegisters_331__0})) ;
    Reg_16 loop1_331_x (.D ({inputRegisters_331__15,inputRegisters_331__14,
           inputRegisters_331__13,inputRegisters_331__12,inputRegisters_331__11,
           inputRegisters_331__10,inputRegisters_331__9,inputRegisters_331__8,
           inputRegisters_331__7,inputRegisters_331__6,inputRegisters_331__5,
           inputRegisters_331__4,inputRegisters_331__3,inputRegisters_331__2,
           inputRegisters_331__1,inputRegisters_331__0}), .en (
           enableRegister_331), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_331__15,registerOutputs_331__14,
           registerOutputs_331__13,registerOutputs_331__12,
           registerOutputs_331__11,registerOutputs_331__10,
           registerOutputs_331__9,registerOutputs_331__8,registerOutputs_331__7,
           registerOutputs_331__6,registerOutputs_331__5,registerOutputs_331__4,
           registerOutputs_331__3,registerOutputs_331__2,registerOutputs_331__1,
           registerOutputs_331__0})) ;
    Mux2_16 loop1_332_y (.A ({nx35979,nx36121,nx36263,nx36405,nx36547,nx36689,
            nx36831,nx36973,nx37115,nx37257,nx37399,nx37541,nx37683,nx37825,
            nx37967,nx38109}), .B ({nx33735,nx33873,nx34011,nx34149,nx34289,
            nx34427,nx34565,nx34705,nx34847,nx34989,nx35131,nx35273,nx35415,
            nx35557,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35699), .C ({inputRegisters_332__15,inputRegisters_332__14,
            inputRegisters_332__13,inputRegisters_332__12,inputRegisters_332__11
            ,inputRegisters_332__10,inputRegisters_332__9,inputRegisters_332__8,
            inputRegisters_332__7,inputRegisters_332__6,inputRegisters_332__5,
            inputRegisters_332__4,inputRegisters_332__3,inputRegisters_332__2,
            inputRegisters_332__1,inputRegisters_332__0})) ;
    Reg_16 loop1_332_x (.D ({inputRegisters_332__15,inputRegisters_332__14,
           inputRegisters_332__13,inputRegisters_332__12,inputRegisters_332__11,
           inputRegisters_332__10,inputRegisters_332__9,inputRegisters_332__8,
           inputRegisters_332__7,inputRegisters_332__6,inputRegisters_332__5,
           inputRegisters_332__4,inputRegisters_332__3,inputRegisters_332__2,
           inputRegisters_332__1,inputRegisters_332__0}), .en (
           enableRegister_332), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_332__15,registerOutputs_332__14,
           registerOutputs_332__13,registerOutputs_332__12,
           registerOutputs_332__11,registerOutputs_332__10,
           registerOutputs_332__9,registerOutputs_332__8,registerOutputs_332__7,
           registerOutputs_332__6,registerOutputs_332__5,registerOutputs_332__4,
           registerOutputs_332__3,registerOutputs_332__2,registerOutputs_332__1,
           registerOutputs_332__0})) ;
    Mux2_16 loop1_333_y (.A ({nx35979,nx36121,nx36263,nx36405,nx36547,nx36689,
            nx36831,nx36973,nx37115,nx37257,nx37399,nx37541,nx37683,nx37825,
            nx37967,nx38109}), .B ({nx33735,nx33873,nx34011,nx34151,nx34289,
            nx34427,nx34565,nx34705,nx34847,nx34989,nx35131,nx35273,nx35415,
            nx35557,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35699), .C ({inputRegisters_333__15,inputRegisters_333__14,
            inputRegisters_333__13,inputRegisters_333__12,inputRegisters_333__11
            ,inputRegisters_333__10,inputRegisters_333__9,inputRegisters_333__8,
            inputRegisters_333__7,inputRegisters_333__6,inputRegisters_333__5,
            inputRegisters_333__4,inputRegisters_333__3,inputRegisters_333__2,
            inputRegisters_333__1,inputRegisters_333__0})) ;
    Reg_16 loop1_333_x (.D ({inputRegisters_333__15,inputRegisters_333__14,
           inputRegisters_333__13,inputRegisters_333__12,inputRegisters_333__11,
           inputRegisters_333__10,inputRegisters_333__9,inputRegisters_333__8,
           inputRegisters_333__7,inputRegisters_333__6,inputRegisters_333__5,
           inputRegisters_333__4,inputRegisters_333__3,inputRegisters_333__2,
           inputRegisters_333__1,inputRegisters_333__0}), .en (
           enableRegister_333), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_333__15,registerOutputs_333__14,
           registerOutputs_333__13,registerOutputs_333__12,
           registerOutputs_333__11,registerOutputs_333__10,
           registerOutputs_333__9,registerOutputs_333__8,registerOutputs_333__7,
           registerOutputs_333__6,registerOutputs_333__5,registerOutputs_333__4,
           registerOutputs_333__3,registerOutputs_333__2,registerOutputs_333__1,
           registerOutputs_333__0})) ;
    Mux2_16 loop1_334_y (.A ({nx35979,nx36121,nx36263,nx36405,nx36547,nx36689,
            nx36831,nx36973,nx37115,nx37257,nx37399,nx37541,nx37683,nx37825,
            nx37967,nx38109}), .B ({nx33735,nx33873,nx34013,nx34151,nx34289,
            nx34427,nx34565,nx34705,nx34847,nx34989,nx35131,nx35273,nx35415,
            nx35557,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35699), .C ({inputRegisters_334__15,inputRegisters_334__14,
            inputRegisters_334__13,inputRegisters_334__12,inputRegisters_334__11
            ,inputRegisters_334__10,inputRegisters_334__9,inputRegisters_334__8,
            inputRegisters_334__7,inputRegisters_334__6,inputRegisters_334__5,
            inputRegisters_334__4,inputRegisters_334__3,inputRegisters_334__2,
            inputRegisters_334__1,inputRegisters_334__0})) ;
    Reg_16 loop1_334_x (.D ({inputRegisters_334__15,inputRegisters_334__14,
           inputRegisters_334__13,inputRegisters_334__12,inputRegisters_334__11,
           inputRegisters_334__10,inputRegisters_334__9,inputRegisters_334__8,
           inputRegisters_334__7,inputRegisters_334__6,inputRegisters_334__5,
           inputRegisters_334__4,inputRegisters_334__3,inputRegisters_334__2,
           inputRegisters_334__1,inputRegisters_334__0}), .en (
           enableRegister_334), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_334__15,registerOutputs_334__14,
           registerOutputs_334__13,registerOutputs_334__12,
           registerOutputs_334__11,registerOutputs_334__10,
           registerOutputs_334__9,registerOutputs_334__8,registerOutputs_334__7,
           registerOutputs_334__6,registerOutputs_334__5,registerOutputs_334__4,
           registerOutputs_334__3,registerOutputs_334__2,registerOutputs_334__1,
           registerOutputs_334__0})) ;
    Mux2_16 loop1_335_y (.A ({nx35979,nx36121,nx36263,nx36405,nx36547,nx36689,
            nx36831,nx36973,nx37115,nx37257,nx37399,nx37541,nx37683,nx37825,
            nx37967,nx38109}), .B ({nx33735,nx33875,nx34013,nx34151,nx34289,
            nx34427,nx34565,nx34705,nx34847,nx34989,nx35131,nx35273,nx35415,
            nx35557,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35699), .C ({inputRegisters_335__15,inputRegisters_335__14,
            inputRegisters_335__13,inputRegisters_335__12,inputRegisters_335__11
            ,inputRegisters_335__10,inputRegisters_335__9,inputRegisters_335__8,
            inputRegisters_335__7,inputRegisters_335__6,inputRegisters_335__5,
            inputRegisters_335__4,inputRegisters_335__3,inputRegisters_335__2,
            inputRegisters_335__1,inputRegisters_335__0})) ;
    Reg_16 loop1_335_x (.D ({inputRegisters_335__15,inputRegisters_335__14,
           inputRegisters_335__13,inputRegisters_335__12,inputRegisters_335__11,
           inputRegisters_335__10,inputRegisters_335__9,inputRegisters_335__8,
           inputRegisters_335__7,inputRegisters_335__6,inputRegisters_335__5,
           inputRegisters_335__4,inputRegisters_335__3,inputRegisters_335__2,
           inputRegisters_335__1,inputRegisters_335__0}), .en (
           enableRegister_335), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_335__15,registerOutputs_335__14,
           registerOutputs_335__13,registerOutputs_335__12,
           registerOutputs_335__11,registerOutputs_335__10,
           registerOutputs_335__9,registerOutputs_335__8,registerOutputs_335__7,
           registerOutputs_335__6,registerOutputs_335__5,registerOutputs_335__4,
           registerOutputs_335__3,registerOutputs_335__2,registerOutputs_335__1,
           registerOutputs_335__0})) ;
    Mux2_16 loop1_336_y (.A ({nx35981,nx36123,nx36265,nx36407,nx36549,nx36691,
            nx36833,nx36975,nx37117,nx37259,nx37401,nx37543,nx37685,nx37827,
            nx37969,nx38111}), .B ({nx33737,nx33875,nx34013,nx34151,nx34289,
            nx34427,nx34565,nx34707,nx34849,nx34991,nx35133,nx35275,nx35417,
            nx35559,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35701), .C ({inputRegisters_336__15,inputRegisters_336__14,
            inputRegisters_336__13,inputRegisters_336__12,inputRegisters_336__11
            ,inputRegisters_336__10,inputRegisters_336__9,inputRegisters_336__8,
            inputRegisters_336__7,inputRegisters_336__6,inputRegisters_336__5,
            inputRegisters_336__4,inputRegisters_336__3,inputRegisters_336__2,
            inputRegisters_336__1,inputRegisters_336__0})) ;
    Reg_16 loop1_336_x (.D ({inputRegisters_336__15,inputRegisters_336__14,
           inputRegisters_336__13,inputRegisters_336__12,inputRegisters_336__11,
           inputRegisters_336__10,inputRegisters_336__9,inputRegisters_336__8,
           inputRegisters_336__7,inputRegisters_336__6,inputRegisters_336__5,
           inputRegisters_336__4,inputRegisters_336__3,inputRegisters_336__2,
           inputRegisters_336__1,inputRegisters_336__0}), .en (
           enableRegister_336), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_336__15,registerOutputs_336__14,
           registerOutputs_336__13,registerOutputs_336__12,
           registerOutputs_336__11,registerOutputs_336__10,
           registerOutputs_336__9,registerOutputs_336__8,registerOutputs_336__7,
           registerOutputs_336__6,registerOutputs_336__5,registerOutputs_336__4,
           registerOutputs_336__3,registerOutputs_336__2,registerOutputs_336__1,
           registerOutputs_336__0})) ;
    Mux2_16 loop1_337_y (.A ({nx35981,nx36123,nx36265,nx36407,nx36549,nx36691,
            nx36833,nx36975,nx37117,nx37259,nx37401,nx37543,nx37685,nx37827,
            nx37969,nx38111}), .B ({nx33737,nx33875,nx34013,nx34151,nx34289,
            nx34427,nx34567,nx34707,nx34849,nx34991,nx35133,nx35275,nx35417,
            nx35559,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35701), .C ({inputRegisters_337__15,inputRegisters_337__14,
            inputRegisters_337__13,inputRegisters_337__12,inputRegisters_337__11
            ,inputRegisters_337__10,inputRegisters_337__9,inputRegisters_337__8,
            inputRegisters_337__7,inputRegisters_337__6,inputRegisters_337__5,
            inputRegisters_337__4,inputRegisters_337__3,inputRegisters_337__2,
            inputRegisters_337__1,inputRegisters_337__0})) ;
    Reg_16 loop1_337_x (.D ({inputRegisters_337__15,inputRegisters_337__14,
           inputRegisters_337__13,inputRegisters_337__12,inputRegisters_337__11,
           inputRegisters_337__10,inputRegisters_337__9,inputRegisters_337__8,
           inputRegisters_337__7,inputRegisters_337__6,inputRegisters_337__5,
           inputRegisters_337__4,inputRegisters_337__3,inputRegisters_337__2,
           inputRegisters_337__1,inputRegisters_337__0}), .en (
           enableRegister_337), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_337__15,registerOutputs_337__14,
           registerOutputs_337__13,registerOutputs_337__12,
           registerOutputs_337__11,registerOutputs_337__10,
           registerOutputs_337__9,registerOutputs_337__8,registerOutputs_337__7,
           registerOutputs_337__6,registerOutputs_337__5,registerOutputs_337__4,
           registerOutputs_337__3,registerOutputs_337__2,registerOutputs_337__1,
           registerOutputs_337__0})) ;
    Mux2_16 loop1_338_y (.A ({nx35981,nx36123,nx36265,nx36407,nx36549,nx36691,
            nx36833,nx36975,nx37117,nx37259,nx37401,nx37543,nx37685,nx37827,
            nx37969,nx38111}), .B ({nx33737,nx33875,nx34013,nx34151,nx34289,
            nx34429,nx34567,nx34707,nx34849,nx34991,nx35133,nx35275,nx35417,
            nx35559,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35701), .C ({inputRegisters_338__15,inputRegisters_338__14,
            inputRegisters_338__13,inputRegisters_338__12,inputRegisters_338__11
            ,inputRegisters_338__10,inputRegisters_338__9,inputRegisters_338__8,
            inputRegisters_338__7,inputRegisters_338__6,inputRegisters_338__5,
            inputRegisters_338__4,inputRegisters_338__3,inputRegisters_338__2,
            inputRegisters_338__1,inputRegisters_338__0})) ;
    Reg_16 loop1_338_x (.D ({inputRegisters_338__15,inputRegisters_338__14,
           inputRegisters_338__13,inputRegisters_338__12,inputRegisters_338__11,
           inputRegisters_338__10,inputRegisters_338__9,inputRegisters_338__8,
           inputRegisters_338__7,inputRegisters_338__6,inputRegisters_338__5,
           inputRegisters_338__4,inputRegisters_338__3,inputRegisters_338__2,
           inputRegisters_338__1,inputRegisters_338__0}), .en (
           enableRegister_338), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_338__15,registerOutputs_338__14,
           registerOutputs_338__13,registerOutputs_338__12,
           registerOutputs_338__11,registerOutputs_338__10,
           registerOutputs_338__9,registerOutputs_338__8,registerOutputs_338__7,
           registerOutputs_338__6,registerOutputs_338__5,registerOutputs_338__4,
           registerOutputs_338__3,registerOutputs_338__2,registerOutputs_338__1,
           registerOutputs_338__0})) ;
    Mux2_16 loop1_339_y (.A ({nx35981,nx36123,nx36265,nx36407,nx36549,nx36691,
            nx36833,nx36975,nx37117,nx37259,nx37401,nx37543,nx37685,nx37827,
            nx37969,nx38111}), .B ({nx33737,nx33875,nx34013,nx34151,nx34291,
            nx34429,nx34567,nx34707,nx34849,nx34991,nx35133,nx35275,nx35417,
            nx35559,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35701), .C ({inputRegisters_339__15,inputRegisters_339__14,
            inputRegisters_339__13,inputRegisters_339__12,inputRegisters_339__11
            ,inputRegisters_339__10,inputRegisters_339__9,inputRegisters_339__8,
            inputRegisters_339__7,inputRegisters_339__6,inputRegisters_339__5,
            inputRegisters_339__4,inputRegisters_339__3,inputRegisters_339__2,
            inputRegisters_339__1,inputRegisters_339__0})) ;
    Reg_16 loop1_339_x (.D ({inputRegisters_339__15,inputRegisters_339__14,
           inputRegisters_339__13,inputRegisters_339__12,inputRegisters_339__11,
           inputRegisters_339__10,inputRegisters_339__9,inputRegisters_339__8,
           inputRegisters_339__7,inputRegisters_339__6,inputRegisters_339__5,
           inputRegisters_339__4,inputRegisters_339__3,inputRegisters_339__2,
           inputRegisters_339__1,inputRegisters_339__0}), .en (
           enableRegister_339), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_339__15,registerOutputs_339__14,
           registerOutputs_339__13,registerOutputs_339__12,
           registerOutputs_339__11,registerOutputs_339__10,
           registerOutputs_339__9,registerOutputs_339__8,registerOutputs_339__7,
           registerOutputs_339__6,registerOutputs_339__5,registerOutputs_339__4,
           registerOutputs_339__3,registerOutputs_339__2,registerOutputs_339__1,
           registerOutputs_339__0})) ;
    Mux2_16 loop1_340_y (.A ({nx35981,nx36123,nx36265,nx36407,nx36549,nx36691,
            nx36833,nx36975,nx37117,nx37259,nx37401,nx37543,nx37685,nx37827,
            nx37969,nx38111}), .B ({nx33737,nx33875,nx34013,nx34153,nx34291,
            nx34429,nx34567,nx34707,nx34849,nx34991,nx35133,nx35275,nx35417,
            nx35559,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35701), .C ({inputRegisters_340__15,inputRegisters_340__14,
            inputRegisters_340__13,inputRegisters_340__12,inputRegisters_340__11
            ,inputRegisters_340__10,inputRegisters_340__9,inputRegisters_340__8,
            inputRegisters_340__7,inputRegisters_340__6,inputRegisters_340__5,
            inputRegisters_340__4,inputRegisters_340__3,inputRegisters_340__2,
            inputRegisters_340__1,inputRegisters_340__0})) ;
    Reg_16 loop1_340_x (.D ({inputRegisters_340__15,inputRegisters_340__14,
           inputRegisters_340__13,inputRegisters_340__12,inputRegisters_340__11,
           inputRegisters_340__10,inputRegisters_340__9,inputRegisters_340__8,
           inputRegisters_340__7,inputRegisters_340__6,inputRegisters_340__5,
           inputRegisters_340__4,inputRegisters_340__3,inputRegisters_340__2,
           inputRegisters_340__1,inputRegisters_340__0}), .en (
           enableRegister_340), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_340__15,registerOutputs_340__14,
           registerOutputs_340__13,registerOutputs_340__12,
           registerOutputs_340__11,registerOutputs_340__10,
           registerOutputs_340__9,registerOutputs_340__8,registerOutputs_340__7,
           registerOutputs_340__6,registerOutputs_340__5,registerOutputs_340__4,
           registerOutputs_340__3,registerOutputs_340__2,registerOutputs_340__1,
           registerOutputs_340__0})) ;
    Mux2_16 loop1_341_y (.A ({nx35981,nx36123,nx36265,nx36407,nx36549,nx36691,
            nx36833,nx36975,nx37117,nx37259,nx37401,nx37543,nx37685,nx37827,
            nx37969,nx38111}), .B ({nx33737,nx33875,nx34015,nx34153,nx34291,
            nx34429,nx34567,nx34707,nx34849,nx34991,nx35133,nx35275,nx35417,
            nx35559,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35701), .C ({inputRegisters_341__15,inputRegisters_341__14,
            inputRegisters_341__13,inputRegisters_341__12,inputRegisters_341__11
            ,inputRegisters_341__10,inputRegisters_341__9,inputRegisters_341__8,
            inputRegisters_341__7,inputRegisters_341__6,inputRegisters_341__5,
            inputRegisters_341__4,inputRegisters_341__3,inputRegisters_341__2,
            inputRegisters_341__1,inputRegisters_341__0})) ;
    Reg_16 loop1_341_x (.D ({inputRegisters_341__15,inputRegisters_341__14,
           inputRegisters_341__13,inputRegisters_341__12,inputRegisters_341__11,
           inputRegisters_341__10,inputRegisters_341__9,inputRegisters_341__8,
           inputRegisters_341__7,inputRegisters_341__6,inputRegisters_341__5,
           inputRegisters_341__4,inputRegisters_341__3,inputRegisters_341__2,
           inputRegisters_341__1,inputRegisters_341__0}), .en (
           enableRegister_341), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_341__15,registerOutputs_341__14,
           registerOutputs_341__13,registerOutputs_341__12,
           registerOutputs_341__11,registerOutputs_341__10,
           registerOutputs_341__9,registerOutputs_341__8,registerOutputs_341__7,
           registerOutputs_341__6,registerOutputs_341__5,registerOutputs_341__4,
           registerOutputs_341__3,registerOutputs_341__2,registerOutputs_341__1,
           registerOutputs_341__0})) ;
    Mux2_16 loop1_342_y (.A ({nx35981,nx36123,nx36265,nx36407,nx36549,nx36691,
            nx36833,nx36975,nx37117,nx37259,nx37401,nx37543,nx37685,nx37827,
            nx37969,nx38111}), .B ({nx33737,nx33877,nx34015,nx34153,nx34291,
            nx34429,nx34567,nx34707,nx34849,nx34991,nx35133,nx35275,nx35417,
            nx35559,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35701), .C ({inputRegisters_342__15,inputRegisters_342__14,
            inputRegisters_342__13,inputRegisters_342__12,inputRegisters_342__11
            ,inputRegisters_342__10,inputRegisters_342__9,inputRegisters_342__8,
            inputRegisters_342__7,inputRegisters_342__6,inputRegisters_342__5,
            inputRegisters_342__4,inputRegisters_342__3,inputRegisters_342__2,
            inputRegisters_342__1,inputRegisters_342__0})) ;
    Reg_16 loop1_342_x (.D ({inputRegisters_342__15,inputRegisters_342__14,
           inputRegisters_342__13,inputRegisters_342__12,inputRegisters_342__11,
           inputRegisters_342__10,inputRegisters_342__9,inputRegisters_342__8,
           inputRegisters_342__7,inputRegisters_342__6,inputRegisters_342__5,
           inputRegisters_342__4,inputRegisters_342__3,inputRegisters_342__2,
           inputRegisters_342__1,inputRegisters_342__0}), .en (
           enableRegister_342), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_342__15,registerOutputs_342__14,
           registerOutputs_342__13,registerOutputs_342__12,
           registerOutputs_342__11,registerOutputs_342__10,
           registerOutputs_342__9,registerOutputs_342__8,registerOutputs_342__7,
           registerOutputs_342__6,registerOutputs_342__5,registerOutputs_342__4,
           registerOutputs_342__3,registerOutputs_342__2,registerOutputs_342__1,
           registerOutputs_342__0})) ;
    Mux2_16 loop1_343_y (.A ({nx35983,nx36125,nx36267,nx36409,nx36551,nx36693,
            nx36835,nx36977,nx37119,nx37261,nx37403,nx37545,nx37687,nx37829,
            nx37971,nx38113}), .B ({nx33739,nx33877,nx34015,nx34153,nx34291,
            nx34429,nx34567,nx34709,nx34851,nx34993,nx35135,nx35277,nx35419,
            nx35561,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35703), .C ({inputRegisters_343__15,inputRegisters_343__14,
            inputRegisters_343__13,inputRegisters_343__12,inputRegisters_343__11
            ,inputRegisters_343__10,inputRegisters_343__9,inputRegisters_343__8,
            inputRegisters_343__7,inputRegisters_343__6,inputRegisters_343__5,
            inputRegisters_343__4,inputRegisters_343__3,inputRegisters_343__2,
            inputRegisters_343__1,inputRegisters_343__0})) ;
    Reg_16 loop1_343_x (.D ({inputRegisters_343__15,inputRegisters_343__14,
           inputRegisters_343__13,inputRegisters_343__12,inputRegisters_343__11,
           inputRegisters_343__10,inputRegisters_343__9,inputRegisters_343__8,
           inputRegisters_343__7,inputRegisters_343__6,inputRegisters_343__5,
           inputRegisters_343__4,inputRegisters_343__3,inputRegisters_343__2,
           inputRegisters_343__1,inputRegisters_343__0}), .en (
           enableRegister_343), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_343__15,registerOutputs_343__14,
           registerOutputs_343__13,registerOutputs_343__12,
           registerOutputs_343__11,registerOutputs_343__10,
           registerOutputs_343__9,registerOutputs_343__8,registerOutputs_343__7,
           registerOutputs_343__6,registerOutputs_343__5,registerOutputs_343__4,
           registerOutputs_343__3,registerOutputs_343__2,registerOutputs_343__1,
           registerOutputs_343__0})) ;
    Mux2_16 loop1_344_y (.A ({nx35983,nx36125,nx36267,nx36409,nx36551,nx36693,
            nx36835,nx36977,nx37119,nx37261,nx37403,nx37545,nx37687,nx37829,
            nx37971,nx38113}), .B ({nx33739,nx33877,nx34015,nx34153,nx34291,
            nx34429,nx34569,nx34709,nx34851,nx34993,nx35135,nx35277,nx35419,
            nx35561,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35703), .C ({inputRegisters_344__15,inputRegisters_344__14,
            inputRegisters_344__13,inputRegisters_344__12,inputRegisters_344__11
            ,inputRegisters_344__10,inputRegisters_344__9,inputRegisters_344__8,
            inputRegisters_344__7,inputRegisters_344__6,inputRegisters_344__5,
            inputRegisters_344__4,inputRegisters_344__3,inputRegisters_344__2,
            inputRegisters_344__1,inputRegisters_344__0})) ;
    Reg_16 loop1_344_x (.D ({inputRegisters_344__15,inputRegisters_344__14,
           inputRegisters_344__13,inputRegisters_344__12,inputRegisters_344__11,
           inputRegisters_344__10,inputRegisters_344__9,inputRegisters_344__8,
           inputRegisters_344__7,inputRegisters_344__6,inputRegisters_344__5,
           inputRegisters_344__4,inputRegisters_344__3,inputRegisters_344__2,
           inputRegisters_344__1,inputRegisters_344__0}), .en (
           enableRegister_344), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_344__15,registerOutputs_344__14,
           registerOutputs_344__13,registerOutputs_344__12,
           registerOutputs_344__11,registerOutputs_344__10,
           registerOutputs_344__9,registerOutputs_344__8,registerOutputs_344__7,
           registerOutputs_344__6,registerOutputs_344__5,registerOutputs_344__4,
           registerOutputs_344__3,registerOutputs_344__2,registerOutputs_344__1,
           registerOutputs_344__0})) ;
    Mux2_16 loop1_345_y (.A ({nx35983,nx36125,nx36267,nx36409,nx36551,nx36693,
            nx36835,nx36977,nx37119,nx37261,nx37403,nx37545,nx37687,nx37829,
            nx37971,nx38113}), .B ({nx33739,nx33877,nx34015,nx34153,nx34291,
            nx34431,nx34569,nx34709,nx34851,nx34993,nx35135,nx35277,nx35419,
            nx35561,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35703), .C ({inputRegisters_345__15,inputRegisters_345__14,
            inputRegisters_345__13,inputRegisters_345__12,inputRegisters_345__11
            ,inputRegisters_345__10,inputRegisters_345__9,inputRegisters_345__8,
            inputRegisters_345__7,inputRegisters_345__6,inputRegisters_345__5,
            inputRegisters_345__4,inputRegisters_345__3,inputRegisters_345__2,
            inputRegisters_345__1,inputRegisters_345__0})) ;
    Reg_16 loop1_345_x (.D ({inputRegisters_345__15,inputRegisters_345__14,
           inputRegisters_345__13,inputRegisters_345__12,inputRegisters_345__11,
           inputRegisters_345__10,inputRegisters_345__9,inputRegisters_345__8,
           inputRegisters_345__7,inputRegisters_345__6,inputRegisters_345__5,
           inputRegisters_345__4,inputRegisters_345__3,inputRegisters_345__2,
           inputRegisters_345__1,inputRegisters_345__0}), .en (
           enableRegister_345), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_345__15,registerOutputs_345__14,
           registerOutputs_345__13,registerOutputs_345__12,
           registerOutputs_345__11,registerOutputs_345__10,
           registerOutputs_345__9,registerOutputs_345__8,registerOutputs_345__7,
           registerOutputs_345__6,registerOutputs_345__5,registerOutputs_345__4,
           registerOutputs_345__3,registerOutputs_345__2,registerOutputs_345__1,
           registerOutputs_345__0})) ;
    Mux2_16 loop1_346_y (.A ({nx35983,nx36125,nx36267,nx36409,nx36551,nx36693,
            nx36835,nx36977,nx37119,nx37261,nx37403,nx37545,nx37687,nx37829,
            nx37971,nx38113}), .B ({nx33739,nx33877,nx34015,nx34153,nx34293,
            nx34431,nx34569,nx34709,nx34851,nx34993,nx35135,nx35277,nx35419,
            nx35561,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35703), .C ({inputRegisters_346__15,inputRegisters_346__14,
            inputRegisters_346__13,inputRegisters_346__12,inputRegisters_346__11
            ,inputRegisters_346__10,inputRegisters_346__9,inputRegisters_346__8,
            inputRegisters_346__7,inputRegisters_346__6,inputRegisters_346__5,
            inputRegisters_346__4,inputRegisters_346__3,inputRegisters_346__2,
            inputRegisters_346__1,inputRegisters_346__0})) ;
    Reg_16 loop1_346_x (.D ({inputRegisters_346__15,inputRegisters_346__14,
           inputRegisters_346__13,inputRegisters_346__12,inputRegisters_346__11,
           inputRegisters_346__10,inputRegisters_346__9,inputRegisters_346__8,
           inputRegisters_346__7,inputRegisters_346__6,inputRegisters_346__5,
           inputRegisters_346__4,inputRegisters_346__3,inputRegisters_346__2,
           inputRegisters_346__1,inputRegisters_346__0}), .en (
           enableRegister_346), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_346__15,registerOutputs_346__14,
           registerOutputs_346__13,registerOutputs_346__12,
           registerOutputs_346__11,registerOutputs_346__10,
           registerOutputs_346__9,registerOutputs_346__8,registerOutputs_346__7,
           registerOutputs_346__6,registerOutputs_346__5,registerOutputs_346__4,
           registerOutputs_346__3,registerOutputs_346__2,registerOutputs_346__1,
           registerOutputs_346__0})) ;
    Mux2_16 loop1_347_y (.A ({nx35983,nx36125,nx36267,nx36409,nx36551,nx36693,
            nx36835,nx36977,nx37119,nx37261,nx37403,nx37545,nx37687,nx37829,
            nx37971,nx38113}), .B ({nx33739,nx33877,nx34015,nx34155,nx34293,
            nx34431,nx34569,nx34709,nx34851,nx34993,nx35135,nx35277,nx35419,
            nx35561,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35703), .C ({inputRegisters_347__15,inputRegisters_347__14,
            inputRegisters_347__13,inputRegisters_347__12,inputRegisters_347__11
            ,inputRegisters_347__10,inputRegisters_347__9,inputRegisters_347__8,
            inputRegisters_347__7,inputRegisters_347__6,inputRegisters_347__5,
            inputRegisters_347__4,inputRegisters_347__3,inputRegisters_347__2,
            inputRegisters_347__1,inputRegisters_347__0})) ;
    Reg_16 loop1_347_x (.D ({inputRegisters_347__15,inputRegisters_347__14,
           inputRegisters_347__13,inputRegisters_347__12,inputRegisters_347__11,
           inputRegisters_347__10,inputRegisters_347__9,inputRegisters_347__8,
           inputRegisters_347__7,inputRegisters_347__6,inputRegisters_347__5,
           inputRegisters_347__4,inputRegisters_347__3,inputRegisters_347__2,
           inputRegisters_347__1,inputRegisters_347__0}), .en (
           enableRegister_347), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_347__15,registerOutputs_347__14,
           registerOutputs_347__13,registerOutputs_347__12,
           registerOutputs_347__11,registerOutputs_347__10,
           registerOutputs_347__9,registerOutputs_347__8,registerOutputs_347__7,
           registerOutputs_347__6,registerOutputs_347__5,registerOutputs_347__4,
           registerOutputs_347__3,registerOutputs_347__2,registerOutputs_347__1,
           registerOutputs_347__0})) ;
    Mux2_16 loop1_348_y (.A ({nx35983,nx36125,nx36267,nx36409,nx36551,nx36693,
            nx36835,nx36977,nx37119,nx37261,nx37403,nx37545,nx37687,nx37829,
            nx37971,nx38113}), .B ({nx33739,nx33877,nx34017,nx34155,nx34293,
            nx34431,nx34569,nx34709,nx34851,nx34993,nx35135,nx35277,nx35419,
            nx35561,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35703), .C ({inputRegisters_348__15,inputRegisters_348__14,
            inputRegisters_348__13,inputRegisters_348__12,inputRegisters_348__11
            ,inputRegisters_348__10,inputRegisters_348__9,inputRegisters_348__8,
            inputRegisters_348__7,inputRegisters_348__6,inputRegisters_348__5,
            inputRegisters_348__4,inputRegisters_348__3,inputRegisters_348__2,
            inputRegisters_348__1,inputRegisters_348__0})) ;
    Reg_16 loop1_348_x (.D ({inputRegisters_348__15,inputRegisters_348__14,
           inputRegisters_348__13,inputRegisters_348__12,inputRegisters_348__11,
           inputRegisters_348__10,inputRegisters_348__9,inputRegisters_348__8,
           inputRegisters_348__7,inputRegisters_348__6,inputRegisters_348__5,
           inputRegisters_348__4,inputRegisters_348__3,inputRegisters_348__2,
           inputRegisters_348__1,inputRegisters_348__0}), .en (
           enableRegister_348), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_348__15,registerOutputs_348__14,
           registerOutputs_348__13,registerOutputs_348__12,
           registerOutputs_348__11,registerOutputs_348__10,
           registerOutputs_348__9,registerOutputs_348__8,registerOutputs_348__7,
           registerOutputs_348__6,registerOutputs_348__5,registerOutputs_348__4,
           registerOutputs_348__3,registerOutputs_348__2,registerOutputs_348__1,
           registerOutputs_348__0})) ;
    Mux2_16 loop1_349_y (.A ({nx35983,nx36125,nx36267,nx36409,nx36551,nx36693,
            nx36835,nx36977,nx37119,nx37261,nx37403,nx37545,nx37687,nx37829,
            nx37971,nx38113}), .B ({nx33739,nx33879,nx34017,nx34155,nx34293,
            nx34431,nx34569,nx34709,nx34851,nx34993,nx35135,nx35277,nx35419,
            nx35561,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35703), .C ({inputRegisters_349__15,inputRegisters_349__14,
            inputRegisters_349__13,inputRegisters_349__12,inputRegisters_349__11
            ,inputRegisters_349__10,inputRegisters_349__9,inputRegisters_349__8,
            inputRegisters_349__7,inputRegisters_349__6,inputRegisters_349__5,
            inputRegisters_349__4,inputRegisters_349__3,inputRegisters_349__2,
            inputRegisters_349__1,inputRegisters_349__0})) ;
    Reg_16 loop1_349_x (.D ({inputRegisters_349__15,inputRegisters_349__14,
           inputRegisters_349__13,inputRegisters_349__12,inputRegisters_349__11,
           inputRegisters_349__10,inputRegisters_349__9,inputRegisters_349__8,
           inputRegisters_349__7,inputRegisters_349__6,inputRegisters_349__5,
           inputRegisters_349__4,inputRegisters_349__3,inputRegisters_349__2,
           inputRegisters_349__1,inputRegisters_349__0}), .en (
           enableRegister_349), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_349__15,registerOutputs_349__14,
           registerOutputs_349__13,registerOutputs_349__12,
           registerOutputs_349__11,registerOutputs_349__10,
           registerOutputs_349__9,registerOutputs_349__8,registerOutputs_349__7,
           registerOutputs_349__6,registerOutputs_349__5,registerOutputs_349__4,
           registerOutputs_349__3,registerOutputs_349__2,registerOutputs_349__1,
           registerOutputs_349__0})) ;
    Mux2_16 loop1_350_y (.A ({nx35985,nx36127,nx36269,nx36411,nx36553,nx36695,
            nx36837,nx36979,nx37121,nx37263,nx37405,nx37547,nx37689,nx37831,
            nx37973,nx38115}), .B ({nx33741,nx33879,nx34017,nx34155,nx34293,
            nx34431,nx34569,nx34711,nx34853,nx34995,nx35137,nx35279,nx35421,
            nx35563,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35705), .C ({inputRegisters_350__15,inputRegisters_350__14,
            inputRegisters_350__13,inputRegisters_350__12,inputRegisters_350__11
            ,inputRegisters_350__10,inputRegisters_350__9,inputRegisters_350__8,
            inputRegisters_350__7,inputRegisters_350__6,inputRegisters_350__5,
            inputRegisters_350__4,inputRegisters_350__3,inputRegisters_350__2,
            inputRegisters_350__1,inputRegisters_350__0})) ;
    Reg_16 loop1_350_x (.D ({inputRegisters_350__15,inputRegisters_350__14,
           inputRegisters_350__13,inputRegisters_350__12,inputRegisters_350__11,
           inputRegisters_350__10,inputRegisters_350__9,inputRegisters_350__8,
           inputRegisters_350__7,inputRegisters_350__6,inputRegisters_350__5,
           inputRegisters_350__4,inputRegisters_350__3,inputRegisters_350__2,
           inputRegisters_350__1,inputRegisters_350__0}), .en (
           enableRegister_350), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_350__15,registerOutputs_350__14,
           registerOutputs_350__13,registerOutputs_350__12,
           registerOutputs_350__11,registerOutputs_350__10,
           registerOutputs_350__9,registerOutputs_350__8,registerOutputs_350__7,
           registerOutputs_350__6,registerOutputs_350__5,registerOutputs_350__4,
           registerOutputs_350__3,registerOutputs_350__2,registerOutputs_350__1,
           registerOutputs_350__0})) ;
    Mux2_16 loop1_351_y (.A ({nx35985,nx36127,nx36269,nx36411,nx36553,nx36695,
            nx36837,nx36979,nx37121,nx37263,nx37405,nx37547,nx37689,nx37831,
            nx37973,nx38115}), .B ({nx33741,nx33879,nx34017,nx34155,nx34293,
            nx34431,nx34571,nx34711,nx34853,nx34995,nx35137,nx35279,nx35421,
            nx35563,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35705), .C ({inputRegisters_351__15,inputRegisters_351__14,
            inputRegisters_351__13,inputRegisters_351__12,inputRegisters_351__11
            ,inputRegisters_351__10,inputRegisters_351__9,inputRegisters_351__8,
            inputRegisters_351__7,inputRegisters_351__6,inputRegisters_351__5,
            inputRegisters_351__4,inputRegisters_351__3,inputRegisters_351__2,
            inputRegisters_351__1,inputRegisters_351__0})) ;
    Reg_16 loop1_351_x (.D ({inputRegisters_351__15,inputRegisters_351__14,
           inputRegisters_351__13,inputRegisters_351__12,inputRegisters_351__11,
           inputRegisters_351__10,inputRegisters_351__9,inputRegisters_351__8,
           inputRegisters_351__7,inputRegisters_351__6,inputRegisters_351__5,
           inputRegisters_351__4,inputRegisters_351__3,inputRegisters_351__2,
           inputRegisters_351__1,inputRegisters_351__0}), .en (
           enableRegister_351), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_351__15,registerOutputs_351__14,
           registerOutputs_351__13,registerOutputs_351__12,
           registerOutputs_351__11,registerOutputs_351__10,
           registerOutputs_351__9,registerOutputs_351__8,registerOutputs_351__7,
           registerOutputs_351__6,registerOutputs_351__5,registerOutputs_351__4,
           registerOutputs_351__3,registerOutputs_351__2,registerOutputs_351__1,
           registerOutputs_351__0})) ;
    Mux2_16 loop1_352_y (.A ({nx35985,nx36127,nx36269,nx36411,nx36553,nx36695,
            nx36837,nx36979,nx37121,nx37263,nx37405,nx37547,nx37689,nx37831,
            nx37973,nx38115}), .B ({nx33741,nx33879,nx34017,nx34155,nx34293,
            nx34433,nx34571,nx34711,nx34853,nx34995,nx35137,nx35279,nx35421,
            nx35563,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35705), .C ({inputRegisters_352__15,inputRegisters_352__14,
            inputRegisters_352__13,inputRegisters_352__12,inputRegisters_352__11
            ,inputRegisters_352__10,inputRegisters_352__9,inputRegisters_352__8,
            inputRegisters_352__7,inputRegisters_352__6,inputRegisters_352__5,
            inputRegisters_352__4,inputRegisters_352__3,inputRegisters_352__2,
            inputRegisters_352__1,inputRegisters_352__0})) ;
    Reg_16 loop1_352_x (.D ({inputRegisters_352__15,inputRegisters_352__14,
           inputRegisters_352__13,inputRegisters_352__12,inputRegisters_352__11,
           inputRegisters_352__10,inputRegisters_352__9,inputRegisters_352__8,
           inputRegisters_352__7,inputRegisters_352__6,inputRegisters_352__5,
           inputRegisters_352__4,inputRegisters_352__3,inputRegisters_352__2,
           inputRegisters_352__1,inputRegisters_352__0}), .en (
           enableRegister_352), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_352__15,registerOutputs_352__14,
           registerOutputs_352__13,registerOutputs_352__12,
           registerOutputs_352__11,registerOutputs_352__10,
           registerOutputs_352__9,registerOutputs_352__8,registerOutputs_352__7,
           registerOutputs_352__6,registerOutputs_352__5,registerOutputs_352__4,
           registerOutputs_352__3,registerOutputs_352__2,registerOutputs_352__1,
           registerOutputs_352__0})) ;
    Mux2_16 loop1_353_y (.A ({nx35985,nx36127,nx36269,nx36411,nx36553,nx36695,
            nx36837,nx36979,nx37121,nx37263,nx37405,nx37547,nx37689,nx37831,
            nx37973,nx38115}), .B ({nx33741,nx33879,nx34017,nx34155,nx34295,
            nx34433,nx34571,nx34711,nx34853,nx34995,nx35137,nx35279,nx35421,
            nx35563,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35705), .C ({inputRegisters_353__15,inputRegisters_353__14,
            inputRegisters_353__13,inputRegisters_353__12,inputRegisters_353__11
            ,inputRegisters_353__10,inputRegisters_353__9,inputRegisters_353__8,
            inputRegisters_353__7,inputRegisters_353__6,inputRegisters_353__5,
            inputRegisters_353__4,inputRegisters_353__3,inputRegisters_353__2,
            inputRegisters_353__1,inputRegisters_353__0})) ;
    Reg_16 loop1_353_x (.D ({inputRegisters_353__15,inputRegisters_353__14,
           inputRegisters_353__13,inputRegisters_353__12,inputRegisters_353__11,
           inputRegisters_353__10,inputRegisters_353__9,inputRegisters_353__8,
           inputRegisters_353__7,inputRegisters_353__6,inputRegisters_353__5,
           inputRegisters_353__4,inputRegisters_353__3,inputRegisters_353__2,
           inputRegisters_353__1,inputRegisters_353__0}), .en (
           enableRegister_353), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_353__15,registerOutputs_353__14,
           registerOutputs_353__13,registerOutputs_353__12,
           registerOutputs_353__11,registerOutputs_353__10,
           registerOutputs_353__9,registerOutputs_353__8,registerOutputs_353__7,
           registerOutputs_353__6,registerOutputs_353__5,registerOutputs_353__4,
           registerOutputs_353__3,registerOutputs_353__2,registerOutputs_353__1,
           registerOutputs_353__0})) ;
    Mux2_16 loop1_354_y (.A ({nx35985,nx36127,nx36269,nx36411,nx36553,nx36695,
            nx36837,nx36979,nx37121,nx37263,nx37405,nx37547,nx37689,nx37831,
            nx37973,nx38115}), .B ({nx33741,nx33879,nx34017,nx34157,nx34295,
            nx34433,nx34571,nx34711,nx34853,nx34995,nx35137,nx35279,nx35421,
            nx35563,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35705), .C ({inputRegisters_354__15,inputRegisters_354__14,
            inputRegisters_354__13,inputRegisters_354__12,inputRegisters_354__11
            ,inputRegisters_354__10,inputRegisters_354__9,inputRegisters_354__8,
            inputRegisters_354__7,inputRegisters_354__6,inputRegisters_354__5,
            inputRegisters_354__4,inputRegisters_354__3,inputRegisters_354__2,
            inputRegisters_354__1,inputRegisters_354__0})) ;
    Reg_16 loop1_354_x (.D ({inputRegisters_354__15,inputRegisters_354__14,
           inputRegisters_354__13,inputRegisters_354__12,inputRegisters_354__11,
           inputRegisters_354__10,inputRegisters_354__9,inputRegisters_354__8,
           inputRegisters_354__7,inputRegisters_354__6,inputRegisters_354__5,
           inputRegisters_354__4,inputRegisters_354__3,inputRegisters_354__2,
           inputRegisters_354__1,inputRegisters_354__0}), .en (
           enableRegister_354), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_354__15,registerOutputs_354__14,
           registerOutputs_354__13,registerOutputs_354__12,
           registerOutputs_354__11,registerOutputs_354__10,
           registerOutputs_354__9,registerOutputs_354__8,registerOutputs_354__7,
           registerOutputs_354__6,registerOutputs_354__5,registerOutputs_354__4,
           registerOutputs_354__3,registerOutputs_354__2,registerOutputs_354__1,
           registerOutputs_354__0})) ;
    Mux2_16 loop1_355_y (.A ({nx35985,nx36127,nx36269,nx36411,nx36553,nx36695,
            nx36837,nx36979,nx37121,nx37263,nx37405,nx37547,nx37689,nx37831,
            nx37973,nx38115}), .B ({nx33741,nx33879,nx34019,nx34157,nx34295,
            nx34433,nx34571,nx34711,nx34853,nx34995,nx35137,nx35279,nx35421,
            nx35563,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35705), .C ({inputRegisters_355__15,inputRegisters_355__14,
            inputRegisters_355__13,inputRegisters_355__12,inputRegisters_355__11
            ,inputRegisters_355__10,inputRegisters_355__9,inputRegisters_355__8,
            inputRegisters_355__7,inputRegisters_355__6,inputRegisters_355__5,
            inputRegisters_355__4,inputRegisters_355__3,inputRegisters_355__2,
            inputRegisters_355__1,inputRegisters_355__0})) ;
    Reg_16 loop1_355_x (.D ({inputRegisters_355__15,inputRegisters_355__14,
           inputRegisters_355__13,inputRegisters_355__12,inputRegisters_355__11,
           inputRegisters_355__10,inputRegisters_355__9,inputRegisters_355__8,
           inputRegisters_355__7,inputRegisters_355__6,inputRegisters_355__5,
           inputRegisters_355__4,inputRegisters_355__3,inputRegisters_355__2,
           inputRegisters_355__1,inputRegisters_355__0}), .en (
           enableRegister_355), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_355__15,registerOutputs_355__14,
           registerOutputs_355__13,registerOutputs_355__12,
           registerOutputs_355__11,registerOutputs_355__10,
           registerOutputs_355__9,registerOutputs_355__8,registerOutputs_355__7,
           registerOutputs_355__6,registerOutputs_355__5,registerOutputs_355__4,
           registerOutputs_355__3,registerOutputs_355__2,registerOutputs_355__1,
           registerOutputs_355__0})) ;
    Mux2_16 loop1_356_y (.A ({nx35985,nx36127,nx36269,nx36411,nx36553,nx36695,
            nx36837,nx36979,nx37121,nx37263,nx37405,nx37547,nx37689,nx37831,
            nx37973,nx38115}), .B ({nx33741,nx33881,nx34019,nx34157,nx34295,
            nx34433,nx34571,nx34711,nx34853,nx34995,nx35137,nx35279,nx35421,
            nx35563,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35705), .C ({inputRegisters_356__15,inputRegisters_356__14,
            inputRegisters_356__13,inputRegisters_356__12,inputRegisters_356__11
            ,inputRegisters_356__10,inputRegisters_356__9,inputRegisters_356__8,
            inputRegisters_356__7,inputRegisters_356__6,inputRegisters_356__5,
            inputRegisters_356__4,inputRegisters_356__3,inputRegisters_356__2,
            inputRegisters_356__1,inputRegisters_356__0})) ;
    Reg_16 loop1_356_x (.D ({inputRegisters_356__15,inputRegisters_356__14,
           inputRegisters_356__13,inputRegisters_356__12,inputRegisters_356__11,
           inputRegisters_356__10,inputRegisters_356__9,inputRegisters_356__8,
           inputRegisters_356__7,inputRegisters_356__6,inputRegisters_356__5,
           inputRegisters_356__4,inputRegisters_356__3,inputRegisters_356__2,
           inputRegisters_356__1,inputRegisters_356__0}), .en (
           enableRegister_356), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_356__15,registerOutputs_356__14,
           registerOutputs_356__13,registerOutputs_356__12,
           registerOutputs_356__11,registerOutputs_356__10,
           registerOutputs_356__9,registerOutputs_356__8,registerOutputs_356__7,
           registerOutputs_356__6,registerOutputs_356__5,registerOutputs_356__4,
           registerOutputs_356__3,registerOutputs_356__2,registerOutputs_356__1,
           registerOutputs_356__0})) ;
    Mux2_16 loop1_357_y (.A ({nx35987,nx36129,nx36271,nx36413,nx36555,nx36697,
            nx36839,nx36981,nx37123,nx37265,nx37407,nx37549,nx37691,nx37833,
            nx37975,nx38117}), .B ({nx33743,nx33881,nx34019,nx34157,nx34295,
            nx34433,nx34571,nx34713,nx34855,nx34997,nx35139,nx35281,nx35423,
            nx35565,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35707), .C ({inputRegisters_357__15,inputRegisters_357__14,
            inputRegisters_357__13,inputRegisters_357__12,inputRegisters_357__11
            ,inputRegisters_357__10,inputRegisters_357__9,inputRegisters_357__8,
            inputRegisters_357__7,inputRegisters_357__6,inputRegisters_357__5,
            inputRegisters_357__4,inputRegisters_357__3,inputRegisters_357__2,
            inputRegisters_357__1,inputRegisters_357__0})) ;
    Reg_16 loop1_357_x (.D ({inputRegisters_357__15,inputRegisters_357__14,
           inputRegisters_357__13,inputRegisters_357__12,inputRegisters_357__11,
           inputRegisters_357__10,inputRegisters_357__9,inputRegisters_357__8,
           inputRegisters_357__7,inputRegisters_357__6,inputRegisters_357__5,
           inputRegisters_357__4,inputRegisters_357__3,inputRegisters_357__2,
           inputRegisters_357__1,inputRegisters_357__0}), .en (
           enableRegister_357), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_357__15,registerOutputs_357__14,
           registerOutputs_357__13,registerOutputs_357__12,
           registerOutputs_357__11,registerOutputs_357__10,
           registerOutputs_357__9,registerOutputs_357__8,registerOutputs_357__7,
           registerOutputs_357__6,registerOutputs_357__5,registerOutputs_357__4,
           registerOutputs_357__3,registerOutputs_357__2,registerOutputs_357__1,
           registerOutputs_357__0})) ;
    Mux2_16 loop1_358_y (.A ({nx35987,nx36129,nx36271,nx36413,nx36555,nx36697,
            nx36839,nx36981,nx37123,nx37265,nx37407,nx37549,nx37691,nx37833,
            nx37975,nx38117}), .B ({nx33743,nx33881,nx34019,nx34157,nx34295,
            nx34433,nx34573,nx34713,nx34855,nx34997,nx35139,nx35281,nx35423,
            nx35565,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35707), .C ({inputRegisters_358__15,inputRegisters_358__14,
            inputRegisters_358__13,inputRegisters_358__12,inputRegisters_358__11
            ,inputRegisters_358__10,inputRegisters_358__9,inputRegisters_358__8,
            inputRegisters_358__7,inputRegisters_358__6,inputRegisters_358__5,
            inputRegisters_358__4,inputRegisters_358__3,inputRegisters_358__2,
            inputRegisters_358__1,inputRegisters_358__0})) ;
    Reg_16 loop1_358_x (.D ({inputRegisters_358__15,inputRegisters_358__14,
           inputRegisters_358__13,inputRegisters_358__12,inputRegisters_358__11,
           inputRegisters_358__10,inputRegisters_358__9,inputRegisters_358__8,
           inputRegisters_358__7,inputRegisters_358__6,inputRegisters_358__5,
           inputRegisters_358__4,inputRegisters_358__3,inputRegisters_358__2,
           inputRegisters_358__1,inputRegisters_358__0}), .en (
           enableRegister_358), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_358__15,registerOutputs_358__14,
           registerOutputs_358__13,registerOutputs_358__12,
           registerOutputs_358__11,registerOutputs_358__10,
           registerOutputs_358__9,registerOutputs_358__8,registerOutputs_358__7,
           registerOutputs_358__6,registerOutputs_358__5,registerOutputs_358__4,
           registerOutputs_358__3,registerOutputs_358__2,registerOutputs_358__1,
           registerOutputs_358__0})) ;
    Mux2_16 loop1_359_y (.A ({nx35987,nx36129,nx36271,nx36413,nx36555,nx36697,
            nx36839,nx36981,nx37123,nx37265,nx37407,nx37549,nx37691,nx37833,
            nx37975,nx38117}), .B ({nx33743,nx33881,nx34019,nx34157,nx34295,
            nx34435,nx34573,nx34713,nx34855,nx34997,nx35139,nx35281,nx35423,
            nx35565,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35707), .C ({inputRegisters_359__15,inputRegisters_359__14,
            inputRegisters_359__13,inputRegisters_359__12,inputRegisters_359__11
            ,inputRegisters_359__10,inputRegisters_359__9,inputRegisters_359__8,
            inputRegisters_359__7,inputRegisters_359__6,inputRegisters_359__5,
            inputRegisters_359__4,inputRegisters_359__3,inputRegisters_359__2,
            inputRegisters_359__1,inputRegisters_359__0})) ;
    Reg_16 loop1_359_x (.D ({inputRegisters_359__15,inputRegisters_359__14,
           inputRegisters_359__13,inputRegisters_359__12,inputRegisters_359__11,
           inputRegisters_359__10,inputRegisters_359__9,inputRegisters_359__8,
           inputRegisters_359__7,inputRegisters_359__6,inputRegisters_359__5,
           inputRegisters_359__4,inputRegisters_359__3,inputRegisters_359__2,
           inputRegisters_359__1,inputRegisters_359__0}), .en (
           enableRegister_359), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_359__15,registerOutputs_359__14,
           registerOutputs_359__13,registerOutputs_359__12,
           registerOutputs_359__11,registerOutputs_359__10,
           registerOutputs_359__9,registerOutputs_359__8,registerOutputs_359__7,
           registerOutputs_359__6,registerOutputs_359__5,registerOutputs_359__4,
           registerOutputs_359__3,registerOutputs_359__2,registerOutputs_359__1,
           registerOutputs_359__0})) ;
    Mux2_16 loop1_360_y (.A ({nx35987,nx36129,nx36271,nx36413,nx36555,nx36697,
            nx36839,nx36981,nx37123,nx37265,nx37407,nx37549,nx37691,nx37833,
            nx37975,nx38117}), .B ({nx33743,nx33881,nx34019,nx34157,nx34297,
            nx34435,nx34573,nx34713,nx34855,nx34997,nx35139,nx35281,nx35423,
            nx35565,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35707), .C ({inputRegisters_360__15,inputRegisters_360__14,
            inputRegisters_360__13,inputRegisters_360__12,inputRegisters_360__11
            ,inputRegisters_360__10,inputRegisters_360__9,inputRegisters_360__8,
            inputRegisters_360__7,inputRegisters_360__6,inputRegisters_360__5,
            inputRegisters_360__4,inputRegisters_360__3,inputRegisters_360__2,
            inputRegisters_360__1,inputRegisters_360__0})) ;
    Reg_16 loop1_360_x (.D ({inputRegisters_360__15,inputRegisters_360__14,
           inputRegisters_360__13,inputRegisters_360__12,inputRegisters_360__11,
           inputRegisters_360__10,inputRegisters_360__9,inputRegisters_360__8,
           inputRegisters_360__7,inputRegisters_360__6,inputRegisters_360__5,
           inputRegisters_360__4,inputRegisters_360__3,inputRegisters_360__2,
           inputRegisters_360__1,inputRegisters_360__0}), .en (
           enableRegister_360), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_360__15,registerOutputs_360__14,
           registerOutputs_360__13,registerOutputs_360__12,
           registerOutputs_360__11,registerOutputs_360__10,
           registerOutputs_360__9,registerOutputs_360__8,registerOutputs_360__7,
           registerOutputs_360__6,registerOutputs_360__5,registerOutputs_360__4,
           registerOutputs_360__3,registerOutputs_360__2,registerOutputs_360__1,
           registerOutputs_360__0})) ;
    Mux2_16 loop1_361_y (.A ({nx35987,nx36129,nx36271,nx36413,nx36555,nx36697,
            nx36839,nx36981,nx37123,nx37265,nx37407,nx37549,nx37691,nx37833,
            nx37975,nx38117}), .B ({nx33743,nx33881,nx34019,nx34159,nx34297,
            nx34435,nx34573,nx34713,nx34855,nx34997,nx35139,nx35281,nx35423,
            nx35565,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35707), .C ({inputRegisters_361__15,inputRegisters_361__14,
            inputRegisters_361__13,inputRegisters_361__12,inputRegisters_361__11
            ,inputRegisters_361__10,inputRegisters_361__9,inputRegisters_361__8,
            inputRegisters_361__7,inputRegisters_361__6,inputRegisters_361__5,
            inputRegisters_361__4,inputRegisters_361__3,inputRegisters_361__2,
            inputRegisters_361__1,inputRegisters_361__0})) ;
    Reg_16 loop1_361_x (.D ({inputRegisters_361__15,inputRegisters_361__14,
           inputRegisters_361__13,inputRegisters_361__12,inputRegisters_361__11,
           inputRegisters_361__10,inputRegisters_361__9,inputRegisters_361__8,
           inputRegisters_361__7,inputRegisters_361__6,inputRegisters_361__5,
           inputRegisters_361__4,inputRegisters_361__3,inputRegisters_361__2,
           inputRegisters_361__1,inputRegisters_361__0}), .en (
           enableRegister_361), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_361__15,registerOutputs_361__14,
           registerOutputs_361__13,registerOutputs_361__12,
           registerOutputs_361__11,registerOutputs_361__10,
           registerOutputs_361__9,registerOutputs_361__8,registerOutputs_361__7,
           registerOutputs_361__6,registerOutputs_361__5,registerOutputs_361__4,
           registerOutputs_361__3,registerOutputs_361__2,registerOutputs_361__1,
           registerOutputs_361__0})) ;
    Mux2_16 loop1_362_y (.A ({nx35987,nx36129,nx36271,nx36413,nx36555,nx36697,
            nx36839,nx36981,nx37123,nx37265,nx37407,nx37549,nx37691,nx37833,
            nx37975,nx38117}), .B ({nx33743,nx33881,nx34021,nx34159,nx34297,
            nx34435,nx34573,nx34713,nx34855,nx34997,nx35139,nx35281,nx35423,
            nx35565,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35707), .C ({inputRegisters_362__15,inputRegisters_362__14,
            inputRegisters_362__13,inputRegisters_362__12,inputRegisters_362__11
            ,inputRegisters_362__10,inputRegisters_362__9,inputRegisters_362__8,
            inputRegisters_362__7,inputRegisters_362__6,inputRegisters_362__5,
            inputRegisters_362__4,inputRegisters_362__3,inputRegisters_362__2,
            inputRegisters_362__1,inputRegisters_362__0})) ;
    Reg_16 loop1_362_x (.D ({inputRegisters_362__15,inputRegisters_362__14,
           inputRegisters_362__13,inputRegisters_362__12,inputRegisters_362__11,
           inputRegisters_362__10,inputRegisters_362__9,inputRegisters_362__8,
           inputRegisters_362__7,inputRegisters_362__6,inputRegisters_362__5,
           inputRegisters_362__4,inputRegisters_362__3,inputRegisters_362__2,
           inputRegisters_362__1,inputRegisters_362__0}), .en (
           enableRegister_362), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_362__15,registerOutputs_362__14,
           registerOutputs_362__13,registerOutputs_362__12,
           registerOutputs_362__11,registerOutputs_362__10,
           registerOutputs_362__9,registerOutputs_362__8,registerOutputs_362__7,
           registerOutputs_362__6,registerOutputs_362__5,registerOutputs_362__4,
           registerOutputs_362__3,registerOutputs_362__2,registerOutputs_362__1,
           registerOutputs_362__0})) ;
    Mux2_16 loop1_363_y (.A ({nx35987,nx36129,nx36271,nx36413,nx36555,nx36697,
            nx36839,nx36981,nx37123,nx37265,nx37407,nx37549,nx37691,nx37833,
            nx37975,nx38117}), .B ({nx33743,nx33883,nx34021,nx34159,nx34297,
            nx34435,nx34573,nx34713,nx34855,nx34997,nx35139,nx35281,nx35423,
            nx35565,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35707), .C ({inputRegisters_363__15,inputRegisters_363__14,
            inputRegisters_363__13,inputRegisters_363__12,inputRegisters_363__11
            ,inputRegisters_363__10,inputRegisters_363__9,inputRegisters_363__8,
            inputRegisters_363__7,inputRegisters_363__6,inputRegisters_363__5,
            inputRegisters_363__4,inputRegisters_363__3,inputRegisters_363__2,
            inputRegisters_363__1,inputRegisters_363__0})) ;
    Reg_16 loop1_363_x (.D ({inputRegisters_363__15,inputRegisters_363__14,
           inputRegisters_363__13,inputRegisters_363__12,inputRegisters_363__11,
           inputRegisters_363__10,inputRegisters_363__9,inputRegisters_363__8,
           inputRegisters_363__7,inputRegisters_363__6,inputRegisters_363__5,
           inputRegisters_363__4,inputRegisters_363__3,inputRegisters_363__2,
           inputRegisters_363__1,inputRegisters_363__0}), .en (
           enableRegister_363), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_363__15,registerOutputs_363__14,
           registerOutputs_363__13,registerOutputs_363__12,
           registerOutputs_363__11,registerOutputs_363__10,
           registerOutputs_363__9,registerOutputs_363__8,registerOutputs_363__7,
           registerOutputs_363__6,registerOutputs_363__5,registerOutputs_363__4,
           registerOutputs_363__3,registerOutputs_363__2,registerOutputs_363__1,
           registerOutputs_363__0})) ;
    Mux2_16 loop1_364_y (.A ({nx35989,nx36131,nx36273,nx36415,nx36557,nx36699,
            nx36841,nx36983,nx37125,nx37267,nx37409,nx37551,nx37693,nx37835,
            nx37977,nx38119}), .B ({nx33745,nx33883,nx34021,nx34159,nx34297,
            nx34435,nx34573,nx34715,nx34857,nx34999,nx35141,nx35283,nx35425,
            nx35567,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35709), .C ({inputRegisters_364__15,inputRegisters_364__14,
            inputRegisters_364__13,inputRegisters_364__12,inputRegisters_364__11
            ,inputRegisters_364__10,inputRegisters_364__9,inputRegisters_364__8,
            inputRegisters_364__7,inputRegisters_364__6,inputRegisters_364__5,
            inputRegisters_364__4,inputRegisters_364__3,inputRegisters_364__2,
            inputRegisters_364__1,inputRegisters_364__0})) ;
    Reg_16 loop1_364_x (.D ({inputRegisters_364__15,inputRegisters_364__14,
           inputRegisters_364__13,inputRegisters_364__12,inputRegisters_364__11,
           inputRegisters_364__10,inputRegisters_364__9,inputRegisters_364__8,
           inputRegisters_364__7,inputRegisters_364__6,inputRegisters_364__5,
           inputRegisters_364__4,inputRegisters_364__3,inputRegisters_364__2,
           inputRegisters_364__1,inputRegisters_364__0}), .en (
           enableRegister_364), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_364__15,registerOutputs_364__14,
           registerOutputs_364__13,registerOutputs_364__12,
           registerOutputs_364__11,registerOutputs_364__10,
           registerOutputs_364__9,registerOutputs_364__8,registerOutputs_364__7,
           registerOutputs_364__6,registerOutputs_364__5,registerOutputs_364__4,
           registerOutputs_364__3,registerOutputs_364__2,registerOutputs_364__1,
           registerOutputs_364__0})) ;
    Mux2_16 loop1_365_y (.A ({nx35989,nx36131,nx36273,nx36415,nx36557,nx36699,
            nx36841,nx36983,nx37125,nx37267,nx37409,nx37551,nx37693,nx37835,
            nx37977,nx38119}), .B ({nx33745,nx33883,nx34021,nx34159,nx34297,
            nx34435,nx34575,nx34715,nx34857,nx34999,nx35141,nx35283,nx35425,
            nx35567,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35709), .C ({inputRegisters_365__15,inputRegisters_365__14,
            inputRegisters_365__13,inputRegisters_365__12,inputRegisters_365__11
            ,inputRegisters_365__10,inputRegisters_365__9,inputRegisters_365__8,
            inputRegisters_365__7,inputRegisters_365__6,inputRegisters_365__5,
            inputRegisters_365__4,inputRegisters_365__3,inputRegisters_365__2,
            inputRegisters_365__1,inputRegisters_365__0})) ;
    Reg_16 loop1_365_x (.D ({inputRegisters_365__15,inputRegisters_365__14,
           inputRegisters_365__13,inputRegisters_365__12,inputRegisters_365__11,
           inputRegisters_365__10,inputRegisters_365__9,inputRegisters_365__8,
           inputRegisters_365__7,inputRegisters_365__6,inputRegisters_365__5,
           inputRegisters_365__4,inputRegisters_365__3,inputRegisters_365__2,
           inputRegisters_365__1,inputRegisters_365__0}), .en (
           enableRegister_365), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_365__15,registerOutputs_365__14,
           registerOutputs_365__13,registerOutputs_365__12,
           registerOutputs_365__11,registerOutputs_365__10,
           registerOutputs_365__9,registerOutputs_365__8,registerOutputs_365__7,
           registerOutputs_365__6,registerOutputs_365__5,registerOutputs_365__4,
           registerOutputs_365__3,registerOutputs_365__2,registerOutputs_365__1,
           registerOutputs_365__0})) ;
    Mux2_16 loop1_366_y (.A ({nx35989,nx36131,nx36273,nx36415,nx36557,nx36699,
            nx36841,nx36983,nx37125,nx37267,nx37409,nx37551,nx37693,nx37835,
            nx37977,nx38119}), .B ({nx33745,nx33883,nx34021,nx34159,nx34297,
            nx34437,nx34575,nx34715,nx34857,nx34999,nx35141,nx35283,nx35425,
            nx35567,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35709), .C ({inputRegisters_366__15,inputRegisters_366__14,
            inputRegisters_366__13,inputRegisters_366__12,inputRegisters_366__11
            ,inputRegisters_366__10,inputRegisters_366__9,inputRegisters_366__8,
            inputRegisters_366__7,inputRegisters_366__6,inputRegisters_366__5,
            inputRegisters_366__4,inputRegisters_366__3,inputRegisters_366__2,
            inputRegisters_366__1,inputRegisters_366__0})) ;
    Reg_16 loop1_366_x (.D ({inputRegisters_366__15,inputRegisters_366__14,
           inputRegisters_366__13,inputRegisters_366__12,inputRegisters_366__11,
           inputRegisters_366__10,inputRegisters_366__9,inputRegisters_366__8,
           inputRegisters_366__7,inputRegisters_366__6,inputRegisters_366__5,
           inputRegisters_366__4,inputRegisters_366__3,inputRegisters_366__2,
           inputRegisters_366__1,inputRegisters_366__0}), .en (
           enableRegister_366), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_366__15,registerOutputs_366__14,
           registerOutputs_366__13,registerOutputs_366__12,
           registerOutputs_366__11,registerOutputs_366__10,
           registerOutputs_366__9,registerOutputs_366__8,registerOutputs_366__7,
           registerOutputs_366__6,registerOutputs_366__5,registerOutputs_366__4,
           registerOutputs_366__3,registerOutputs_366__2,registerOutputs_366__1,
           registerOutputs_366__0})) ;
    Mux2_16 loop1_367_y (.A ({nx35989,nx36131,nx36273,nx36415,nx36557,nx36699,
            nx36841,nx36983,nx37125,nx37267,nx37409,nx37551,nx37693,nx37835,
            nx37977,nx38119}), .B ({nx33745,nx33883,nx34021,nx34159,nx34299,
            nx34437,nx34575,nx34715,nx34857,nx34999,nx35141,nx35283,nx35425,
            nx35567,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35709), .C ({inputRegisters_367__15,inputRegisters_367__14,
            inputRegisters_367__13,inputRegisters_367__12,inputRegisters_367__11
            ,inputRegisters_367__10,inputRegisters_367__9,inputRegisters_367__8,
            inputRegisters_367__7,inputRegisters_367__6,inputRegisters_367__5,
            inputRegisters_367__4,inputRegisters_367__3,inputRegisters_367__2,
            inputRegisters_367__1,inputRegisters_367__0})) ;
    Reg_16 loop1_367_x (.D ({inputRegisters_367__15,inputRegisters_367__14,
           inputRegisters_367__13,inputRegisters_367__12,inputRegisters_367__11,
           inputRegisters_367__10,inputRegisters_367__9,inputRegisters_367__8,
           inputRegisters_367__7,inputRegisters_367__6,inputRegisters_367__5,
           inputRegisters_367__4,inputRegisters_367__3,inputRegisters_367__2,
           inputRegisters_367__1,inputRegisters_367__0}), .en (
           enableRegister_367), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_367__15,registerOutputs_367__14,
           registerOutputs_367__13,registerOutputs_367__12,
           registerOutputs_367__11,registerOutputs_367__10,
           registerOutputs_367__9,registerOutputs_367__8,registerOutputs_367__7,
           registerOutputs_367__6,registerOutputs_367__5,registerOutputs_367__4,
           registerOutputs_367__3,registerOutputs_367__2,registerOutputs_367__1,
           registerOutputs_367__0})) ;
    Mux2_16 loop1_368_y (.A ({nx35989,nx36131,nx36273,nx36415,nx36557,nx36699,
            nx36841,nx36983,nx37125,nx37267,nx37409,nx37551,nx37693,nx37835,
            nx37977,nx38119}), .B ({nx33745,nx33883,nx34021,nx34161,nx34299,
            nx34437,nx34575,nx34715,nx34857,nx34999,nx35141,nx35283,nx35425,
            nx35567,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35709), .C ({inputRegisters_368__15,inputRegisters_368__14,
            inputRegisters_368__13,inputRegisters_368__12,inputRegisters_368__11
            ,inputRegisters_368__10,inputRegisters_368__9,inputRegisters_368__8,
            inputRegisters_368__7,inputRegisters_368__6,inputRegisters_368__5,
            inputRegisters_368__4,inputRegisters_368__3,inputRegisters_368__2,
            inputRegisters_368__1,inputRegisters_368__0})) ;
    Reg_16 loop1_368_x (.D ({inputRegisters_368__15,inputRegisters_368__14,
           inputRegisters_368__13,inputRegisters_368__12,inputRegisters_368__11,
           inputRegisters_368__10,inputRegisters_368__9,inputRegisters_368__8,
           inputRegisters_368__7,inputRegisters_368__6,inputRegisters_368__5,
           inputRegisters_368__4,inputRegisters_368__3,inputRegisters_368__2,
           inputRegisters_368__1,inputRegisters_368__0}), .en (
           enableRegister_368), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_368__15,registerOutputs_368__14,
           registerOutputs_368__13,registerOutputs_368__12,
           registerOutputs_368__11,registerOutputs_368__10,
           registerOutputs_368__9,registerOutputs_368__8,registerOutputs_368__7,
           registerOutputs_368__6,registerOutputs_368__5,registerOutputs_368__4,
           registerOutputs_368__3,registerOutputs_368__2,registerOutputs_368__1,
           registerOutputs_368__0})) ;
    Mux2_16 loop1_369_y (.A ({nx35989,nx36131,nx36273,nx36415,nx36557,nx36699,
            nx36841,nx36983,nx37125,nx37267,nx37409,nx37551,nx37693,nx37835,
            nx37977,nx38119}), .B ({nx33745,nx33883,nx34023,nx34161,nx34299,
            nx34437,nx34575,nx34715,nx34857,nx34999,nx35141,nx35283,nx35425,
            nx35567,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35709), .C ({inputRegisters_369__15,inputRegisters_369__14,
            inputRegisters_369__13,inputRegisters_369__12,inputRegisters_369__11
            ,inputRegisters_369__10,inputRegisters_369__9,inputRegisters_369__8,
            inputRegisters_369__7,inputRegisters_369__6,inputRegisters_369__5,
            inputRegisters_369__4,inputRegisters_369__3,inputRegisters_369__2,
            inputRegisters_369__1,inputRegisters_369__0})) ;
    Reg_16 loop1_369_x (.D ({inputRegisters_369__15,inputRegisters_369__14,
           inputRegisters_369__13,inputRegisters_369__12,inputRegisters_369__11,
           inputRegisters_369__10,inputRegisters_369__9,inputRegisters_369__8,
           inputRegisters_369__7,inputRegisters_369__6,inputRegisters_369__5,
           inputRegisters_369__4,inputRegisters_369__3,inputRegisters_369__2,
           inputRegisters_369__1,inputRegisters_369__0}), .en (
           enableRegister_369), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_369__15,registerOutputs_369__14,
           registerOutputs_369__13,registerOutputs_369__12,
           registerOutputs_369__11,registerOutputs_369__10,
           registerOutputs_369__9,registerOutputs_369__8,registerOutputs_369__7,
           registerOutputs_369__6,registerOutputs_369__5,registerOutputs_369__4,
           registerOutputs_369__3,registerOutputs_369__2,registerOutputs_369__1,
           registerOutputs_369__0})) ;
    Mux2_16 loop1_370_y (.A ({nx35989,nx36131,nx36273,nx36415,nx36557,nx36699,
            nx36841,nx36983,nx37125,nx37267,nx37409,nx37551,nx37693,nx37835,
            nx37977,nx38119}), .B ({nx33745,nx33885,nx34023,nx34161,nx34299,
            nx34437,nx34575,nx34715,nx34857,nx34999,nx35141,nx35283,nx35425,
            nx35567,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35709), .C ({inputRegisters_370__15,inputRegisters_370__14,
            inputRegisters_370__13,inputRegisters_370__12,inputRegisters_370__11
            ,inputRegisters_370__10,inputRegisters_370__9,inputRegisters_370__8,
            inputRegisters_370__7,inputRegisters_370__6,inputRegisters_370__5,
            inputRegisters_370__4,inputRegisters_370__3,inputRegisters_370__2,
            inputRegisters_370__1,inputRegisters_370__0})) ;
    Reg_16 loop1_370_x (.D ({inputRegisters_370__15,inputRegisters_370__14,
           inputRegisters_370__13,inputRegisters_370__12,inputRegisters_370__11,
           inputRegisters_370__10,inputRegisters_370__9,inputRegisters_370__8,
           inputRegisters_370__7,inputRegisters_370__6,inputRegisters_370__5,
           inputRegisters_370__4,inputRegisters_370__3,inputRegisters_370__2,
           inputRegisters_370__1,inputRegisters_370__0}), .en (
           enableRegister_370), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_370__15,registerOutputs_370__14,
           registerOutputs_370__13,registerOutputs_370__12,
           registerOutputs_370__11,registerOutputs_370__10,
           registerOutputs_370__9,registerOutputs_370__8,registerOutputs_370__7,
           registerOutputs_370__6,registerOutputs_370__5,registerOutputs_370__4,
           registerOutputs_370__3,registerOutputs_370__2,registerOutputs_370__1,
           registerOutputs_370__0})) ;
    Mux2_16 loop1_371_y (.A ({nx35991,nx36133,nx36275,nx36417,nx36559,nx36701,
            nx36843,nx36985,nx37127,nx37269,nx37411,nx37553,nx37695,nx37837,
            nx37979,nx38121}), .B ({nx33747,nx33885,nx34023,nx34161,nx34299,
            nx34437,nx34575,nx34717,nx34859,nx35001,nx35143,nx35285,nx35427,
            nx35569,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35711), .C ({inputRegisters_371__15,inputRegisters_371__14,
            inputRegisters_371__13,inputRegisters_371__12,inputRegisters_371__11
            ,inputRegisters_371__10,inputRegisters_371__9,inputRegisters_371__8,
            inputRegisters_371__7,inputRegisters_371__6,inputRegisters_371__5,
            inputRegisters_371__4,inputRegisters_371__3,inputRegisters_371__2,
            inputRegisters_371__1,inputRegisters_371__0})) ;
    Reg_16 loop1_371_x (.D ({inputRegisters_371__15,inputRegisters_371__14,
           inputRegisters_371__13,inputRegisters_371__12,inputRegisters_371__11,
           inputRegisters_371__10,inputRegisters_371__9,inputRegisters_371__8,
           inputRegisters_371__7,inputRegisters_371__6,inputRegisters_371__5,
           inputRegisters_371__4,inputRegisters_371__3,inputRegisters_371__2,
           inputRegisters_371__1,inputRegisters_371__0}), .en (
           enableRegister_371), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_371__15,registerOutputs_371__14,
           registerOutputs_371__13,registerOutputs_371__12,
           registerOutputs_371__11,registerOutputs_371__10,
           registerOutputs_371__9,registerOutputs_371__8,registerOutputs_371__7,
           registerOutputs_371__6,registerOutputs_371__5,registerOutputs_371__4,
           registerOutputs_371__3,registerOutputs_371__2,registerOutputs_371__1,
           registerOutputs_371__0})) ;
    Mux2_16 loop1_372_y (.A ({nx35991,nx36133,nx36275,nx36417,nx36559,nx36701,
            nx36843,nx36985,nx37127,nx37269,nx37411,nx37553,nx37695,nx37837,
            nx37979,nx38121}), .B ({nx33747,nx33885,nx34023,nx34161,nx34299,
            nx34437,nx34577,nx34717,nx34859,nx35001,nx35143,nx35285,nx35427,
            nx35569,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35711), .C ({inputRegisters_372__15,inputRegisters_372__14,
            inputRegisters_372__13,inputRegisters_372__12,inputRegisters_372__11
            ,inputRegisters_372__10,inputRegisters_372__9,inputRegisters_372__8,
            inputRegisters_372__7,inputRegisters_372__6,inputRegisters_372__5,
            inputRegisters_372__4,inputRegisters_372__3,inputRegisters_372__2,
            inputRegisters_372__1,inputRegisters_372__0})) ;
    Reg_16 loop1_372_x (.D ({inputRegisters_372__15,inputRegisters_372__14,
           inputRegisters_372__13,inputRegisters_372__12,inputRegisters_372__11,
           inputRegisters_372__10,inputRegisters_372__9,inputRegisters_372__8,
           inputRegisters_372__7,inputRegisters_372__6,inputRegisters_372__5,
           inputRegisters_372__4,inputRegisters_372__3,inputRegisters_372__2,
           inputRegisters_372__1,inputRegisters_372__0}), .en (
           enableRegister_372), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_372__15,registerOutputs_372__14,
           registerOutputs_372__13,registerOutputs_372__12,
           registerOutputs_372__11,registerOutputs_372__10,
           registerOutputs_372__9,registerOutputs_372__8,registerOutputs_372__7,
           registerOutputs_372__6,registerOutputs_372__5,registerOutputs_372__4,
           registerOutputs_372__3,registerOutputs_372__2,registerOutputs_372__1,
           registerOutputs_372__0})) ;
    Mux2_16 loop1_373_y (.A ({nx35991,nx36133,nx36275,nx36417,nx36559,nx36701,
            nx36843,nx36985,nx37127,nx37269,nx37411,nx37553,nx37695,nx37837,
            nx37979,nx38121}), .B ({nx33747,nx33885,nx34023,nx34161,nx34299,
            nx34439,nx34577,nx34717,nx34859,nx35001,nx35143,nx35285,nx35427,
            nx35569,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35711), .C ({inputRegisters_373__15,inputRegisters_373__14,
            inputRegisters_373__13,inputRegisters_373__12,inputRegisters_373__11
            ,inputRegisters_373__10,inputRegisters_373__9,inputRegisters_373__8,
            inputRegisters_373__7,inputRegisters_373__6,inputRegisters_373__5,
            inputRegisters_373__4,inputRegisters_373__3,inputRegisters_373__2,
            inputRegisters_373__1,inputRegisters_373__0})) ;
    Reg_16 loop1_373_x (.D ({inputRegisters_373__15,inputRegisters_373__14,
           inputRegisters_373__13,inputRegisters_373__12,inputRegisters_373__11,
           inputRegisters_373__10,inputRegisters_373__9,inputRegisters_373__8,
           inputRegisters_373__7,inputRegisters_373__6,inputRegisters_373__5,
           inputRegisters_373__4,inputRegisters_373__3,inputRegisters_373__2,
           inputRegisters_373__1,inputRegisters_373__0}), .en (
           enableRegister_373), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_373__15,registerOutputs_373__14,
           registerOutputs_373__13,registerOutputs_373__12,
           registerOutputs_373__11,registerOutputs_373__10,
           registerOutputs_373__9,registerOutputs_373__8,registerOutputs_373__7,
           registerOutputs_373__6,registerOutputs_373__5,registerOutputs_373__4,
           registerOutputs_373__3,registerOutputs_373__2,registerOutputs_373__1,
           registerOutputs_373__0})) ;
    Mux2_16 loop1_374_y (.A ({nx35991,nx36133,nx36275,nx36417,nx36559,nx36701,
            nx36843,nx36985,nx37127,nx37269,nx37411,nx37553,nx37695,nx37837,
            nx37979,nx38121}), .B ({nx33747,nx33885,nx34023,nx34161,nx34301,
            nx34439,nx34577,nx34717,nx34859,nx35001,nx35143,nx35285,nx35427,
            nx35569,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35711), .C ({inputRegisters_374__15,inputRegisters_374__14,
            inputRegisters_374__13,inputRegisters_374__12,inputRegisters_374__11
            ,inputRegisters_374__10,inputRegisters_374__9,inputRegisters_374__8,
            inputRegisters_374__7,inputRegisters_374__6,inputRegisters_374__5,
            inputRegisters_374__4,inputRegisters_374__3,inputRegisters_374__2,
            inputRegisters_374__1,inputRegisters_374__0})) ;
    Reg_16 loop1_374_x (.D ({inputRegisters_374__15,inputRegisters_374__14,
           inputRegisters_374__13,inputRegisters_374__12,inputRegisters_374__11,
           inputRegisters_374__10,inputRegisters_374__9,inputRegisters_374__8,
           inputRegisters_374__7,inputRegisters_374__6,inputRegisters_374__5,
           inputRegisters_374__4,inputRegisters_374__3,inputRegisters_374__2,
           inputRegisters_374__1,inputRegisters_374__0}), .en (
           enableRegister_374), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_374__15,registerOutputs_374__14,
           registerOutputs_374__13,registerOutputs_374__12,
           registerOutputs_374__11,registerOutputs_374__10,
           registerOutputs_374__9,registerOutputs_374__8,registerOutputs_374__7,
           registerOutputs_374__6,registerOutputs_374__5,registerOutputs_374__4,
           registerOutputs_374__3,registerOutputs_374__2,registerOutputs_374__1,
           registerOutputs_374__0})) ;
    Mux2_16 loop1_375_y (.A ({nx35991,nx36133,nx36275,nx36417,nx36559,nx36701,
            nx36843,nx36985,nx37127,nx37269,nx37411,nx37553,nx37695,nx37837,
            nx37979,nx38121}), .B ({nx33747,nx33885,nx34023,nx34163,nx34301,
            nx34439,nx34577,nx34717,nx34859,nx35001,nx35143,nx35285,nx35427,
            nx35569,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35711), .C ({inputRegisters_375__15,inputRegisters_375__14,
            inputRegisters_375__13,inputRegisters_375__12,inputRegisters_375__11
            ,inputRegisters_375__10,inputRegisters_375__9,inputRegisters_375__8,
            inputRegisters_375__7,inputRegisters_375__6,inputRegisters_375__5,
            inputRegisters_375__4,inputRegisters_375__3,inputRegisters_375__2,
            inputRegisters_375__1,inputRegisters_375__0})) ;
    Reg_16 loop1_375_x (.D ({inputRegisters_375__15,inputRegisters_375__14,
           inputRegisters_375__13,inputRegisters_375__12,inputRegisters_375__11,
           inputRegisters_375__10,inputRegisters_375__9,inputRegisters_375__8,
           inputRegisters_375__7,inputRegisters_375__6,inputRegisters_375__5,
           inputRegisters_375__4,inputRegisters_375__3,inputRegisters_375__2,
           inputRegisters_375__1,inputRegisters_375__0}), .en (
           enableRegister_375), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_375__15,registerOutputs_375__14,
           registerOutputs_375__13,registerOutputs_375__12,
           registerOutputs_375__11,registerOutputs_375__10,
           registerOutputs_375__9,registerOutputs_375__8,registerOutputs_375__7,
           registerOutputs_375__6,registerOutputs_375__5,registerOutputs_375__4,
           registerOutputs_375__3,registerOutputs_375__2,registerOutputs_375__1,
           registerOutputs_375__0})) ;
    Mux2_16 loop1_376_y (.A ({nx35991,nx36133,nx36275,nx36417,nx36559,nx36701,
            nx36843,nx36985,nx37127,nx37269,nx37411,nx37553,nx37695,nx37837,
            nx37979,nx38121}), .B ({nx33747,nx33885,nx34025,nx34163,nx34301,
            nx34439,nx34577,nx34717,nx34859,nx35001,nx35143,nx35285,nx35427,
            nx35569,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35711), .C ({inputRegisters_376__15,inputRegisters_376__14,
            inputRegisters_376__13,inputRegisters_376__12,inputRegisters_376__11
            ,inputRegisters_376__10,inputRegisters_376__9,inputRegisters_376__8,
            inputRegisters_376__7,inputRegisters_376__6,inputRegisters_376__5,
            inputRegisters_376__4,inputRegisters_376__3,inputRegisters_376__2,
            inputRegisters_376__1,inputRegisters_376__0})) ;
    Reg_16 loop1_376_x (.D ({inputRegisters_376__15,inputRegisters_376__14,
           inputRegisters_376__13,inputRegisters_376__12,inputRegisters_376__11,
           inputRegisters_376__10,inputRegisters_376__9,inputRegisters_376__8,
           inputRegisters_376__7,inputRegisters_376__6,inputRegisters_376__5,
           inputRegisters_376__4,inputRegisters_376__3,inputRegisters_376__2,
           inputRegisters_376__1,inputRegisters_376__0}), .en (
           enableRegister_376), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_376__15,registerOutputs_376__14,
           registerOutputs_376__13,registerOutputs_376__12,
           registerOutputs_376__11,registerOutputs_376__10,
           registerOutputs_376__9,registerOutputs_376__8,registerOutputs_376__7,
           registerOutputs_376__6,registerOutputs_376__5,registerOutputs_376__4,
           registerOutputs_376__3,registerOutputs_376__2,registerOutputs_376__1,
           registerOutputs_376__0})) ;
    Mux2_16 loop1_377_y (.A ({nx35991,nx36133,nx36275,nx36417,nx36559,nx36701,
            nx36843,nx36985,nx37127,nx37269,nx37411,nx37553,nx37695,nx37837,
            nx37979,nx38121}), .B ({nx33747,nx33887,nx34025,nx34163,nx34301,
            nx34439,nx34577,nx34717,nx34859,nx35001,nx35143,nx35285,nx35427,
            nx35569,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35711), .C ({inputRegisters_377__15,inputRegisters_377__14,
            inputRegisters_377__13,inputRegisters_377__12,inputRegisters_377__11
            ,inputRegisters_377__10,inputRegisters_377__9,inputRegisters_377__8,
            inputRegisters_377__7,inputRegisters_377__6,inputRegisters_377__5,
            inputRegisters_377__4,inputRegisters_377__3,inputRegisters_377__2,
            inputRegisters_377__1,inputRegisters_377__0})) ;
    Reg_16 loop1_377_x (.D ({inputRegisters_377__15,inputRegisters_377__14,
           inputRegisters_377__13,inputRegisters_377__12,inputRegisters_377__11,
           inputRegisters_377__10,inputRegisters_377__9,inputRegisters_377__8,
           inputRegisters_377__7,inputRegisters_377__6,inputRegisters_377__5,
           inputRegisters_377__4,inputRegisters_377__3,inputRegisters_377__2,
           inputRegisters_377__1,inputRegisters_377__0}), .en (
           enableRegister_377), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_377__15,registerOutputs_377__14,
           registerOutputs_377__13,registerOutputs_377__12,
           registerOutputs_377__11,registerOutputs_377__10,
           registerOutputs_377__9,registerOutputs_377__8,registerOutputs_377__7,
           registerOutputs_377__6,registerOutputs_377__5,registerOutputs_377__4,
           registerOutputs_377__3,registerOutputs_377__2,registerOutputs_377__1,
           registerOutputs_377__0})) ;
    Mux2_16 loop1_378_y (.A ({nx35993,nx36135,nx36277,nx36419,nx36561,nx36703,
            nx36845,nx36987,nx37129,nx37271,nx37413,nx37555,nx37697,nx37839,
            nx37981,nx38123}), .B ({nx33749,nx33887,nx34025,nx34163,nx34301,
            nx34439,nx34577,nx34719,nx34861,nx35003,nx35145,nx35287,nx35429,
            nx35571,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35713), .C ({inputRegisters_378__15,inputRegisters_378__14,
            inputRegisters_378__13,inputRegisters_378__12,inputRegisters_378__11
            ,inputRegisters_378__10,inputRegisters_378__9,inputRegisters_378__8,
            inputRegisters_378__7,inputRegisters_378__6,inputRegisters_378__5,
            inputRegisters_378__4,inputRegisters_378__3,inputRegisters_378__2,
            inputRegisters_378__1,inputRegisters_378__0})) ;
    Reg_16 loop1_378_x (.D ({inputRegisters_378__15,inputRegisters_378__14,
           inputRegisters_378__13,inputRegisters_378__12,inputRegisters_378__11,
           inputRegisters_378__10,inputRegisters_378__9,inputRegisters_378__8,
           inputRegisters_378__7,inputRegisters_378__6,inputRegisters_378__5,
           inputRegisters_378__4,inputRegisters_378__3,inputRegisters_378__2,
           inputRegisters_378__1,inputRegisters_378__0}), .en (
           enableRegister_378), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_378__15,registerOutputs_378__14,
           registerOutputs_378__13,registerOutputs_378__12,
           registerOutputs_378__11,registerOutputs_378__10,
           registerOutputs_378__9,registerOutputs_378__8,registerOutputs_378__7,
           registerOutputs_378__6,registerOutputs_378__5,registerOutputs_378__4,
           registerOutputs_378__3,registerOutputs_378__2,registerOutputs_378__1,
           registerOutputs_378__0})) ;
    Mux2_16 loop1_379_y (.A ({nx35993,nx36135,nx36277,nx36419,nx36561,nx36703,
            nx36845,nx36987,nx37129,nx37271,nx37413,nx37555,nx37697,nx37839,
            nx37981,nx38123}), .B ({nx33749,nx33887,nx34025,nx34163,nx34301,
            nx34439,nx34579,nx34719,nx34861,nx35003,nx35145,nx35287,nx35429,
            nx35571,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35713), .C ({inputRegisters_379__15,inputRegisters_379__14,
            inputRegisters_379__13,inputRegisters_379__12,inputRegisters_379__11
            ,inputRegisters_379__10,inputRegisters_379__9,inputRegisters_379__8,
            inputRegisters_379__7,inputRegisters_379__6,inputRegisters_379__5,
            inputRegisters_379__4,inputRegisters_379__3,inputRegisters_379__2,
            inputRegisters_379__1,inputRegisters_379__0})) ;
    Reg_16 loop1_379_x (.D ({inputRegisters_379__15,inputRegisters_379__14,
           inputRegisters_379__13,inputRegisters_379__12,inputRegisters_379__11,
           inputRegisters_379__10,inputRegisters_379__9,inputRegisters_379__8,
           inputRegisters_379__7,inputRegisters_379__6,inputRegisters_379__5,
           inputRegisters_379__4,inputRegisters_379__3,inputRegisters_379__2,
           inputRegisters_379__1,inputRegisters_379__0}), .en (
           enableRegister_379), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_379__15,registerOutputs_379__14,
           registerOutputs_379__13,registerOutputs_379__12,
           registerOutputs_379__11,registerOutputs_379__10,
           registerOutputs_379__9,registerOutputs_379__8,registerOutputs_379__7,
           registerOutputs_379__6,registerOutputs_379__5,registerOutputs_379__4,
           registerOutputs_379__3,registerOutputs_379__2,registerOutputs_379__1,
           registerOutputs_379__0})) ;
    Mux2_16 loop1_380_y (.A ({nx35993,nx36135,nx36277,nx36419,nx36561,nx36703,
            nx36845,nx36987,nx37129,nx37271,nx37413,nx37555,nx37697,nx37839,
            nx37981,nx38123}), .B ({nx33749,nx33887,nx34025,nx34163,nx34301,
            nx34441,nx34579,nx34719,nx34861,nx35003,nx35145,nx35287,nx35429,
            nx35571,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35713), .C ({inputRegisters_380__15,inputRegisters_380__14,
            inputRegisters_380__13,inputRegisters_380__12,inputRegisters_380__11
            ,inputRegisters_380__10,inputRegisters_380__9,inputRegisters_380__8,
            inputRegisters_380__7,inputRegisters_380__6,inputRegisters_380__5,
            inputRegisters_380__4,inputRegisters_380__3,inputRegisters_380__2,
            inputRegisters_380__1,inputRegisters_380__0})) ;
    Reg_16 loop1_380_x (.D ({inputRegisters_380__15,inputRegisters_380__14,
           inputRegisters_380__13,inputRegisters_380__12,inputRegisters_380__11,
           inputRegisters_380__10,inputRegisters_380__9,inputRegisters_380__8,
           inputRegisters_380__7,inputRegisters_380__6,inputRegisters_380__5,
           inputRegisters_380__4,inputRegisters_380__3,inputRegisters_380__2,
           inputRegisters_380__1,inputRegisters_380__0}), .en (
           enableRegister_380), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_380__15,registerOutputs_380__14,
           registerOutputs_380__13,registerOutputs_380__12,
           registerOutputs_380__11,registerOutputs_380__10,
           registerOutputs_380__9,registerOutputs_380__8,registerOutputs_380__7,
           registerOutputs_380__6,registerOutputs_380__5,registerOutputs_380__4,
           registerOutputs_380__3,registerOutputs_380__2,registerOutputs_380__1,
           registerOutputs_380__0})) ;
    Mux2_16 loop1_381_y (.A ({nx35993,nx36135,nx36277,nx36419,nx36561,nx36703,
            nx36845,nx36987,nx37129,nx37271,nx37413,nx37555,nx37697,nx37839,
            nx37981,nx38123}), .B ({nx33749,nx33887,nx34025,nx34163,nx34303,
            nx34441,nx34579,nx34719,nx34861,nx35003,nx35145,nx35287,nx35429,
            nx35571,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35713), .C ({inputRegisters_381__15,inputRegisters_381__14,
            inputRegisters_381__13,inputRegisters_381__12,inputRegisters_381__11
            ,inputRegisters_381__10,inputRegisters_381__9,inputRegisters_381__8,
            inputRegisters_381__7,inputRegisters_381__6,inputRegisters_381__5,
            inputRegisters_381__4,inputRegisters_381__3,inputRegisters_381__2,
            inputRegisters_381__1,inputRegisters_381__0})) ;
    Reg_16 loop1_381_x (.D ({inputRegisters_381__15,inputRegisters_381__14,
           inputRegisters_381__13,inputRegisters_381__12,inputRegisters_381__11,
           inputRegisters_381__10,inputRegisters_381__9,inputRegisters_381__8,
           inputRegisters_381__7,inputRegisters_381__6,inputRegisters_381__5,
           inputRegisters_381__4,inputRegisters_381__3,inputRegisters_381__2,
           inputRegisters_381__1,inputRegisters_381__0}), .en (
           enableRegister_381), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_381__15,registerOutputs_381__14,
           registerOutputs_381__13,registerOutputs_381__12,
           registerOutputs_381__11,registerOutputs_381__10,
           registerOutputs_381__9,registerOutputs_381__8,registerOutputs_381__7,
           registerOutputs_381__6,registerOutputs_381__5,registerOutputs_381__4,
           registerOutputs_381__3,registerOutputs_381__2,registerOutputs_381__1,
           registerOutputs_381__0})) ;
    Mux2_16 loop1_382_y (.A ({nx35993,nx36135,nx36277,nx36419,nx36561,nx36703,
            nx36845,nx36987,nx37129,nx37271,nx37413,nx37555,nx37697,nx37839,
            nx37981,nx38123}), .B ({nx33749,nx33887,nx34025,nx34165,nx34303,
            nx34441,nx34579,nx34719,nx34861,nx35003,nx35145,nx35287,nx35429,
            nx35571,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35713), .C ({inputRegisters_382__15,inputRegisters_382__14,
            inputRegisters_382__13,inputRegisters_382__12,inputRegisters_382__11
            ,inputRegisters_382__10,inputRegisters_382__9,inputRegisters_382__8,
            inputRegisters_382__7,inputRegisters_382__6,inputRegisters_382__5,
            inputRegisters_382__4,inputRegisters_382__3,inputRegisters_382__2,
            inputRegisters_382__1,inputRegisters_382__0})) ;
    Reg_16 loop1_382_x (.D ({inputRegisters_382__15,inputRegisters_382__14,
           inputRegisters_382__13,inputRegisters_382__12,inputRegisters_382__11,
           inputRegisters_382__10,inputRegisters_382__9,inputRegisters_382__8,
           inputRegisters_382__7,inputRegisters_382__6,inputRegisters_382__5,
           inputRegisters_382__4,inputRegisters_382__3,inputRegisters_382__2,
           inputRegisters_382__1,inputRegisters_382__0}), .en (
           enableRegister_382), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_382__15,registerOutputs_382__14,
           registerOutputs_382__13,registerOutputs_382__12,
           registerOutputs_382__11,registerOutputs_382__10,
           registerOutputs_382__9,registerOutputs_382__8,registerOutputs_382__7,
           registerOutputs_382__6,registerOutputs_382__5,registerOutputs_382__4,
           registerOutputs_382__3,registerOutputs_382__2,registerOutputs_382__1,
           registerOutputs_382__0})) ;
    Mux2_16 loop1_383_y (.A ({nx35993,nx36135,nx36277,nx36419,nx36561,nx36703,
            nx36845,nx36987,nx37129,nx37271,nx37413,nx37555,nx37697,nx37839,
            nx37981,nx38123}), .B ({nx33749,nx33887,nx34027,nx34165,nx34303,
            nx34441,nx34579,nx34719,nx34861,nx35003,nx35145,nx35287,nx35429,
            nx35571,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35713), .C ({inputRegisters_383__15,inputRegisters_383__14,
            inputRegisters_383__13,inputRegisters_383__12,inputRegisters_383__11
            ,inputRegisters_383__10,inputRegisters_383__9,inputRegisters_383__8,
            inputRegisters_383__7,inputRegisters_383__6,inputRegisters_383__5,
            inputRegisters_383__4,inputRegisters_383__3,inputRegisters_383__2,
            inputRegisters_383__1,inputRegisters_383__0})) ;
    Reg_16 loop1_383_x (.D ({inputRegisters_383__15,inputRegisters_383__14,
           inputRegisters_383__13,inputRegisters_383__12,inputRegisters_383__11,
           inputRegisters_383__10,inputRegisters_383__9,inputRegisters_383__8,
           inputRegisters_383__7,inputRegisters_383__6,inputRegisters_383__5,
           inputRegisters_383__4,inputRegisters_383__3,inputRegisters_383__2,
           inputRegisters_383__1,inputRegisters_383__0}), .en (
           enableRegister_383), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_383__15,registerOutputs_383__14,
           registerOutputs_383__13,registerOutputs_383__12,
           registerOutputs_383__11,registerOutputs_383__10,
           registerOutputs_383__9,registerOutputs_383__8,registerOutputs_383__7,
           registerOutputs_383__6,registerOutputs_383__5,registerOutputs_383__4,
           registerOutputs_383__3,registerOutputs_383__2,registerOutputs_383__1,
           registerOutputs_383__0})) ;
    Mux2_16 loop1_384_y (.A ({nx35993,nx36135,nx36277,nx36419,nx36561,nx36703,
            nx36845,nx36987,nx37129,nx37271,nx37413,nx37555,nx37697,nx37839,
            nx37981,nx38123}), .B ({nx33749,nx33889,nx34027,nx34165,nx34303,
            nx34441,nx34579,nx34719,nx34861,nx35003,nx35145,nx35287,nx35429,
            nx35571,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35713), .C ({inputRegisters_384__15,inputRegisters_384__14,
            inputRegisters_384__13,inputRegisters_384__12,inputRegisters_384__11
            ,inputRegisters_384__10,inputRegisters_384__9,inputRegisters_384__8,
            inputRegisters_384__7,inputRegisters_384__6,inputRegisters_384__5,
            inputRegisters_384__4,inputRegisters_384__3,inputRegisters_384__2,
            inputRegisters_384__1,inputRegisters_384__0})) ;
    Reg_16 loop1_384_x (.D ({inputRegisters_384__15,inputRegisters_384__14,
           inputRegisters_384__13,inputRegisters_384__12,inputRegisters_384__11,
           inputRegisters_384__10,inputRegisters_384__9,inputRegisters_384__8,
           inputRegisters_384__7,inputRegisters_384__6,inputRegisters_384__5,
           inputRegisters_384__4,inputRegisters_384__3,inputRegisters_384__2,
           inputRegisters_384__1,inputRegisters_384__0}), .en (
           enableRegister_384), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_384__15,registerOutputs_384__14,
           registerOutputs_384__13,registerOutputs_384__12,
           registerOutputs_384__11,registerOutputs_384__10,
           registerOutputs_384__9,registerOutputs_384__8,registerOutputs_384__7,
           registerOutputs_384__6,registerOutputs_384__5,registerOutputs_384__4,
           registerOutputs_384__3,registerOutputs_384__2,registerOutputs_384__1,
           registerOutputs_384__0})) ;
    Mux2_16 loop1_385_y (.A ({nx35995,nx36137,nx36279,nx36421,nx36563,nx36705,
            nx36847,nx36989,nx37131,nx37273,nx37415,nx37557,nx37699,nx37841,
            nx37983,nx38125}), .B ({nx33751,nx33889,nx34027,nx34165,nx34303,
            nx34441,nx34579,nx34721,nx34863,nx35005,nx35147,nx35289,nx35431,
            nx35573,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35715), .C ({inputRegisters_385__15,inputRegisters_385__14,
            inputRegisters_385__13,inputRegisters_385__12,inputRegisters_385__11
            ,inputRegisters_385__10,inputRegisters_385__9,inputRegisters_385__8,
            inputRegisters_385__7,inputRegisters_385__6,inputRegisters_385__5,
            inputRegisters_385__4,inputRegisters_385__3,inputRegisters_385__2,
            inputRegisters_385__1,inputRegisters_385__0})) ;
    Reg_16 loop1_385_x (.D ({inputRegisters_385__15,inputRegisters_385__14,
           inputRegisters_385__13,inputRegisters_385__12,inputRegisters_385__11,
           inputRegisters_385__10,inputRegisters_385__9,inputRegisters_385__8,
           inputRegisters_385__7,inputRegisters_385__6,inputRegisters_385__5,
           inputRegisters_385__4,inputRegisters_385__3,inputRegisters_385__2,
           inputRegisters_385__1,inputRegisters_385__0}), .en (
           enableRegister_385), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_385__15,registerOutputs_385__14,
           registerOutputs_385__13,registerOutputs_385__12,
           registerOutputs_385__11,registerOutputs_385__10,
           registerOutputs_385__9,registerOutputs_385__8,registerOutputs_385__7,
           registerOutputs_385__6,registerOutputs_385__5,registerOutputs_385__4,
           registerOutputs_385__3,registerOutputs_385__2,registerOutputs_385__1,
           registerOutputs_385__0})) ;
    Mux2_16 loop1_386_y (.A ({nx35995,nx36137,nx36279,nx36421,nx36563,nx36705,
            nx36847,nx36989,nx37131,nx37273,nx37415,nx37557,nx37699,nx37841,
            nx37983,nx38125}), .B ({nx33751,nx33889,nx34027,nx34165,nx34303,
            nx34441,nx34581,nx34721,nx34863,nx35005,nx35147,nx35289,nx35431,
            nx35573,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35715), .C ({inputRegisters_386__15,inputRegisters_386__14,
            inputRegisters_386__13,inputRegisters_386__12,inputRegisters_386__11
            ,inputRegisters_386__10,inputRegisters_386__9,inputRegisters_386__8,
            inputRegisters_386__7,inputRegisters_386__6,inputRegisters_386__5,
            inputRegisters_386__4,inputRegisters_386__3,inputRegisters_386__2,
            inputRegisters_386__1,inputRegisters_386__0})) ;
    Reg_16 loop1_386_x (.D ({inputRegisters_386__15,inputRegisters_386__14,
           inputRegisters_386__13,inputRegisters_386__12,inputRegisters_386__11,
           inputRegisters_386__10,inputRegisters_386__9,inputRegisters_386__8,
           inputRegisters_386__7,inputRegisters_386__6,inputRegisters_386__5,
           inputRegisters_386__4,inputRegisters_386__3,inputRegisters_386__2,
           inputRegisters_386__1,inputRegisters_386__0}), .en (
           enableRegister_386), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_386__15,registerOutputs_386__14,
           registerOutputs_386__13,registerOutputs_386__12,
           registerOutputs_386__11,registerOutputs_386__10,
           registerOutputs_386__9,registerOutputs_386__8,registerOutputs_386__7,
           registerOutputs_386__6,registerOutputs_386__5,registerOutputs_386__4,
           registerOutputs_386__3,registerOutputs_386__2,registerOutputs_386__1,
           registerOutputs_386__0})) ;
    Mux2_16 loop1_387_y (.A ({nx35995,nx36137,nx36279,nx36421,nx36563,nx36705,
            nx36847,nx36989,nx37131,nx37273,nx37415,nx37557,nx37699,nx37841,
            nx37983,nx38125}), .B ({nx33751,nx33889,nx34027,nx34165,nx34303,
            nx34443,nx34581,nx34721,nx34863,nx35005,nx35147,nx35289,nx35431,
            nx35573,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35715), .C ({inputRegisters_387__15,inputRegisters_387__14,
            inputRegisters_387__13,inputRegisters_387__12,inputRegisters_387__11
            ,inputRegisters_387__10,inputRegisters_387__9,inputRegisters_387__8,
            inputRegisters_387__7,inputRegisters_387__6,inputRegisters_387__5,
            inputRegisters_387__4,inputRegisters_387__3,inputRegisters_387__2,
            inputRegisters_387__1,inputRegisters_387__0})) ;
    Reg_16 loop1_387_x (.D ({inputRegisters_387__15,inputRegisters_387__14,
           inputRegisters_387__13,inputRegisters_387__12,inputRegisters_387__11,
           inputRegisters_387__10,inputRegisters_387__9,inputRegisters_387__8,
           inputRegisters_387__7,inputRegisters_387__6,inputRegisters_387__5,
           inputRegisters_387__4,inputRegisters_387__3,inputRegisters_387__2,
           inputRegisters_387__1,inputRegisters_387__0}), .en (
           enableRegister_387), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_387__15,registerOutputs_387__14,
           registerOutputs_387__13,registerOutputs_387__12,
           registerOutputs_387__11,registerOutputs_387__10,
           registerOutputs_387__9,registerOutputs_387__8,registerOutputs_387__7,
           registerOutputs_387__6,registerOutputs_387__5,registerOutputs_387__4,
           registerOutputs_387__3,registerOutputs_387__2,registerOutputs_387__1,
           registerOutputs_387__0})) ;
    Mux2_16 loop1_388_y (.A ({nx35995,nx36137,nx36279,nx36421,nx36563,nx36705,
            nx36847,nx36989,nx37131,nx37273,nx37415,nx37557,nx37699,nx37841,
            nx37983,nx38125}), .B ({nx33751,nx33889,nx34027,nx34165,nx34305,
            nx34443,nx34581,nx34721,nx34863,nx35005,nx35147,nx35289,nx35431,
            nx35573,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35715), .C ({inputRegisters_388__15,inputRegisters_388__14,
            inputRegisters_388__13,inputRegisters_388__12,inputRegisters_388__11
            ,inputRegisters_388__10,inputRegisters_388__9,inputRegisters_388__8,
            inputRegisters_388__7,inputRegisters_388__6,inputRegisters_388__5,
            inputRegisters_388__4,inputRegisters_388__3,inputRegisters_388__2,
            inputRegisters_388__1,inputRegisters_388__0})) ;
    Reg_16 loop1_388_x (.D ({inputRegisters_388__15,inputRegisters_388__14,
           inputRegisters_388__13,inputRegisters_388__12,inputRegisters_388__11,
           inputRegisters_388__10,inputRegisters_388__9,inputRegisters_388__8,
           inputRegisters_388__7,inputRegisters_388__6,inputRegisters_388__5,
           inputRegisters_388__4,inputRegisters_388__3,inputRegisters_388__2,
           inputRegisters_388__1,inputRegisters_388__0}), .en (
           enableRegister_388), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_388__15,registerOutputs_388__14,
           registerOutputs_388__13,registerOutputs_388__12,
           registerOutputs_388__11,registerOutputs_388__10,
           registerOutputs_388__9,registerOutputs_388__8,registerOutputs_388__7,
           registerOutputs_388__6,registerOutputs_388__5,registerOutputs_388__4,
           registerOutputs_388__3,registerOutputs_388__2,registerOutputs_388__1,
           registerOutputs_388__0})) ;
    Mux2_16 loop1_389_y (.A ({nx35995,nx36137,nx36279,nx36421,nx36563,nx36705,
            nx36847,nx36989,nx37131,nx37273,nx37415,nx37557,nx37699,nx37841,
            nx37983,nx38125}), .B ({nx33751,nx33889,nx34027,nx34167,nx34305,
            nx34443,nx34581,nx34721,nx34863,nx35005,nx35147,nx35289,nx35431,
            nx35573,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35715), .C ({inputRegisters_389__15,inputRegisters_389__14,
            inputRegisters_389__13,inputRegisters_389__12,inputRegisters_389__11
            ,inputRegisters_389__10,inputRegisters_389__9,inputRegisters_389__8,
            inputRegisters_389__7,inputRegisters_389__6,inputRegisters_389__5,
            inputRegisters_389__4,inputRegisters_389__3,inputRegisters_389__2,
            inputRegisters_389__1,inputRegisters_389__0})) ;
    Reg_16 loop1_389_x (.D ({inputRegisters_389__15,inputRegisters_389__14,
           inputRegisters_389__13,inputRegisters_389__12,inputRegisters_389__11,
           inputRegisters_389__10,inputRegisters_389__9,inputRegisters_389__8,
           inputRegisters_389__7,inputRegisters_389__6,inputRegisters_389__5,
           inputRegisters_389__4,inputRegisters_389__3,inputRegisters_389__2,
           inputRegisters_389__1,inputRegisters_389__0}), .en (
           enableRegister_389), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_389__15,registerOutputs_389__14,
           registerOutputs_389__13,registerOutputs_389__12,
           registerOutputs_389__11,registerOutputs_389__10,
           registerOutputs_389__9,registerOutputs_389__8,registerOutputs_389__7,
           registerOutputs_389__6,registerOutputs_389__5,registerOutputs_389__4,
           registerOutputs_389__3,registerOutputs_389__2,registerOutputs_389__1,
           registerOutputs_389__0})) ;
    Mux2_16 loop1_390_y (.A ({nx35995,nx36137,nx36279,nx36421,nx36563,nx36705,
            nx36847,nx36989,nx37131,nx37273,nx37415,nx37557,nx37699,nx37841,
            nx37983,nx38125}), .B ({nx33751,nx33889,nx34029,nx34167,nx34305,
            nx34443,nx34581,nx34721,nx34863,nx35005,nx35147,nx35289,nx35431,
            nx35573,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35715), .C ({inputRegisters_390__15,inputRegisters_390__14,
            inputRegisters_390__13,inputRegisters_390__12,inputRegisters_390__11
            ,inputRegisters_390__10,inputRegisters_390__9,inputRegisters_390__8,
            inputRegisters_390__7,inputRegisters_390__6,inputRegisters_390__5,
            inputRegisters_390__4,inputRegisters_390__3,inputRegisters_390__2,
            inputRegisters_390__1,inputRegisters_390__0})) ;
    Reg_16 loop1_390_x (.D ({inputRegisters_390__15,inputRegisters_390__14,
           inputRegisters_390__13,inputRegisters_390__12,inputRegisters_390__11,
           inputRegisters_390__10,inputRegisters_390__9,inputRegisters_390__8,
           inputRegisters_390__7,inputRegisters_390__6,inputRegisters_390__5,
           inputRegisters_390__4,inputRegisters_390__3,inputRegisters_390__2,
           inputRegisters_390__1,inputRegisters_390__0}), .en (
           enableRegister_390), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_390__15,registerOutputs_390__14,
           registerOutputs_390__13,registerOutputs_390__12,
           registerOutputs_390__11,registerOutputs_390__10,
           registerOutputs_390__9,registerOutputs_390__8,registerOutputs_390__7,
           registerOutputs_390__6,registerOutputs_390__5,registerOutputs_390__4,
           registerOutputs_390__3,registerOutputs_390__2,registerOutputs_390__1,
           registerOutputs_390__0})) ;
    Mux2_16 loop1_391_y (.A ({nx35995,nx36137,nx36279,nx36421,nx36563,nx36705,
            nx36847,nx36989,nx37131,nx37273,nx37415,nx37557,nx37699,nx37841,
            nx37983,nx38125}), .B ({nx33751,nx33891,nx34029,nx34167,nx34305,
            nx34443,nx34581,nx34721,nx34863,nx35005,nx35147,nx35289,nx35431,
            nx35573,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35715), .C ({inputRegisters_391__15,inputRegisters_391__14,
            inputRegisters_391__13,inputRegisters_391__12,inputRegisters_391__11
            ,inputRegisters_391__10,inputRegisters_391__9,inputRegisters_391__8,
            inputRegisters_391__7,inputRegisters_391__6,inputRegisters_391__5,
            inputRegisters_391__4,inputRegisters_391__3,inputRegisters_391__2,
            inputRegisters_391__1,inputRegisters_391__0})) ;
    Reg_16 loop1_391_x (.D ({inputRegisters_391__15,inputRegisters_391__14,
           inputRegisters_391__13,inputRegisters_391__12,inputRegisters_391__11,
           inputRegisters_391__10,inputRegisters_391__9,inputRegisters_391__8,
           inputRegisters_391__7,inputRegisters_391__6,inputRegisters_391__5,
           inputRegisters_391__4,inputRegisters_391__3,inputRegisters_391__2,
           inputRegisters_391__1,inputRegisters_391__0}), .en (
           enableRegister_391), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_391__15,registerOutputs_391__14,
           registerOutputs_391__13,registerOutputs_391__12,
           registerOutputs_391__11,registerOutputs_391__10,
           registerOutputs_391__9,registerOutputs_391__8,registerOutputs_391__7,
           registerOutputs_391__6,registerOutputs_391__5,registerOutputs_391__4,
           registerOutputs_391__3,registerOutputs_391__2,registerOutputs_391__1,
           registerOutputs_391__0})) ;
    Mux2_16 loop1_392_y (.A ({nx35997,nx36139,nx36281,nx36423,nx36565,nx36707,
            nx36849,nx36991,nx37133,nx37275,nx37417,nx37559,nx37701,nx37843,
            nx37985,nx38127}), .B ({nx33753,nx33891,nx34029,nx34167,nx34305,
            nx34443,nx34581,nx34723,nx34865,nx35007,nx35149,nx35291,nx35433,
            nx35575,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35717), .C ({inputRegisters_392__15,inputRegisters_392__14,
            inputRegisters_392__13,inputRegisters_392__12,inputRegisters_392__11
            ,inputRegisters_392__10,inputRegisters_392__9,inputRegisters_392__8,
            inputRegisters_392__7,inputRegisters_392__6,inputRegisters_392__5,
            inputRegisters_392__4,inputRegisters_392__3,inputRegisters_392__2,
            inputRegisters_392__1,inputRegisters_392__0})) ;
    Reg_16 loop1_392_x (.D ({inputRegisters_392__15,inputRegisters_392__14,
           inputRegisters_392__13,inputRegisters_392__12,inputRegisters_392__11,
           inputRegisters_392__10,inputRegisters_392__9,inputRegisters_392__8,
           inputRegisters_392__7,inputRegisters_392__6,inputRegisters_392__5,
           inputRegisters_392__4,inputRegisters_392__3,inputRegisters_392__2,
           inputRegisters_392__1,inputRegisters_392__0}), .en (
           enableRegister_392), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_392__15,registerOutputs_392__14,
           registerOutputs_392__13,registerOutputs_392__12,
           registerOutputs_392__11,registerOutputs_392__10,
           registerOutputs_392__9,registerOutputs_392__8,registerOutputs_392__7,
           registerOutputs_392__6,registerOutputs_392__5,registerOutputs_392__4,
           registerOutputs_392__3,registerOutputs_392__2,registerOutputs_392__1,
           registerOutputs_392__0})) ;
    Mux2_16 loop1_393_y (.A ({nx35997,nx36139,nx36281,nx36423,nx36565,nx36707,
            nx36849,nx36991,nx37133,nx37275,nx37417,nx37559,nx37701,nx37843,
            nx37985,nx38127}), .B ({nx33753,nx33891,nx34029,nx34167,nx34305,
            nx34443,nx34583,nx34723,nx34865,nx35007,nx35149,nx35291,nx35433,
            nx35575,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35717), .C ({inputRegisters_393__15,inputRegisters_393__14,
            inputRegisters_393__13,inputRegisters_393__12,inputRegisters_393__11
            ,inputRegisters_393__10,inputRegisters_393__9,inputRegisters_393__8,
            inputRegisters_393__7,inputRegisters_393__6,inputRegisters_393__5,
            inputRegisters_393__4,inputRegisters_393__3,inputRegisters_393__2,
            inputRegisters_393__1,inputRegisters_393__0})) ;
    Reg_16 loop1_393_x (.D ({inputRegisters_393__15,inputRegisters_393__14,
           inputRegisters_393__13,inputRegisters_393__12,inputRegisters_393__11,
           inputRegisters_393__10,inputRegisters_393__9,inputRegisters_393__8,
           inputRegisters_393__7,inputRegisters_393__6,inputRegisters_393__5,
           inputRegisters_393__4,inputRegisters_393__3,inputRegisters_393__2,
           inputRegisters_393__1,inputRegisters_393__0}), .en (
           enableRegister_393), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_393__15,registerOutputs_393__14,
           registerOutputs_393__13,registerOutputs_393__12,
           registerOutputs_393__11,registerOutputs_393__10,
           registerOutputs_393__9,registerOutputs_393__8,registerOutputs_393__7,
           registerOutputs_393__6,registerOutputs_393__5,registerOutputs_393__4,
           registerOutputs_393__3,registerOutputs_393__2,registerOutputs_393__1,
           registerOutputs_393__0})) ;
    Mux2_16 loop1_394_y (.A ({nx35997,nx36139,nx36281,nx36423,nx36565,nx36707,
            nx36849,nx36991,nx37133,nx37275,nx37417,nx37559,nx37701,nx37843,
            nx37985,nx38127}), .B ({nx33753,nx33891,nx34029,nx34167,nx34305,
            nx34445,nx34583,nx34723,nx34865,nx35007,nx35149,nx35291,nx35433,
            nx35575,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35717), .C ({inputRegisters_394__15,inputRegisters_394__14,
            inputRegisters_394__13,inputRegisters_394__12,inputRegisters_394__11
            ,inputRegisters_394__10,inputRegisters_394__9,inputRegisters_394__8,
            inputRegisters_394__7,inputRegisters_394__6,inputRegisters_394__5,
            inputRegisters_394__4,inputRegisters_394__3,inputRegisters_394__2,
            inputRegisters_394__1,inputRegisters_394__0})) ;
    Reg_16 loop1_394_x (.D ({inputRegisters_394__15,inputRegisters_394__14,
           inputRegisters_394__13,inputRegisters_394__12,inputRegisters_394__11,
           inputRegisters_394__10,inputRegisters_394__9,inputRegisters_394__8,
           inputRegisters_394__7,inputRegisters_394__6,inputRegisters_394__5,
           inputRegisters_394__4,inputRegisters_394__3,inputRegisters_394__2,
           inputRegisters_394__1,inputRegisters_394__0}), .en (
           enableRegister_394), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_394__15,registerOutputs_394__14,
           registerOutputs_394__13,registerOutputs_394__12,
           registerOutputs_394__11,registerOutputs_394__10,
           registerOutputs_394__9,registerOutputs_394__8,registerOutputs_394__7,
           registerOutputs_394__6,registerOutputs_394__5,registerOutputs_394__4,
           registerOutputs_394__3,registerOutputs_394__2,registerOutputs_394__1,
           registerOutputs_394__0})) ;
    Mux2_16 loop1_395_y (.A ({nx35997,nx36139,nx36281,nx36423,nx36565,nx36707,
            nx36849,nx36991,nx37133,nx37275,nx37417,nx37559,nx37701,nx37843,
            nx37985,nx38127}), .B ({nx33753,nx33891,nx34029,nx34167,nx34307,
            nx34445,nx34583,nx34723,nx34865,nx35007,nx35149,nx35291,nx35433,
            nx35575,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35717), .C ({inputRegisters_395__15,inputRegisters_395__14,
            inputRegisters_395__13,inputRegisters_395__12,inputRegisters_395__11
            ,inputRegisters_395__10,inputRegisters_395__9,inputRegisters_395__8,
            inputRegisters_395__7,inputRegisters_395__6,inputRegisters_395__5,
            inputRegisters_395__4,inputRegisters_395__3,inputRegisters_395__2,
            inputRegisters_395__1,inputRegisters_395__0})) ;
    Reg_16 loop1_395_x (.D ({inputRegisters_395__15,inputRegisters_395__14,
           inputRegisters_395__13,inputRegisters_395__12,inputRegisters_395__11,
           inputRegisters_395__10,inputRegisters_395__9,inputRegisters_395__8,
           inputRegisters_395__7,inputRegisters_395__6,inputRegisters_395__5,
           inputRegisters_395__4,inputRegisters_395__3,inputRegisters_395__2,
           inputRegisters_395__1,inputRegisters_395__0}), .en (
           enableRegister_395), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_395__15,registerOutputs_395__14,
           registerOutputs_395__13,registerOutputs_395__12,
           registerOutputs_395__11,registerOutputs_395__10,
           registerOutputs_395__9,registerOutputs_395__8,registerOutputs_395__7,
           registerOutputs_395__6,registerOutputs_395__5,registerOutputs_395__4,
           registerOutputs_395__3,registerOutputs_395__2,registerOutputs_395__1,
           registerOutputs_395__0})) ;
    Mux2_16 loop1_396_y (.A ({nx35997,nx36139,nx36281,nx36423,nx36565,nx36707,
            nx36849,nx36991,nx37133,nx37275,nx37417,nx37559,nx37701,nx37843,
            nx37985,nx38127}), .B ({nx33753,nx33891,nx34029,nx34169,nx34307,
            nx34445,nx34583,nx34723,nx34865,nx35007,nx35149,nx35291,nx35433,
            nx35575,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35717), .C ({inputRegisters_396__15,inputRegisters_396__14,
            inputRegisters_396__13,inputRegisters_396__12,inputRegisters_396__11
            ,inputRegisters_396__10,inputRegisters_396__9,inputRegisters_396__8,
            inputRegisters_396__7,inputRegisters_396__6,inputRegisters_396__5,
            inputRegisters_396__4,inputRegisters_396__3,inputRegisters_396__2,
            inputRegisters_396__1,inputRegisters_396__0})) ;
    Reg_16 loop1_396_x (.D ({inputRegisters_396__15,inputRegisters_396__14,
           inputRegisters_396__13,inputRegisters_396__12,inputRegisters_396__11,
           inputRegisters_396__10,inputRegisters_396__9,inputRegisters_396__8,
           inputRegisters_396__7,inputRegisters_396__6,inputRegisters_396__5,
           inputRegisters_396__4,inputRegisters_396__3,inputRegisters_396__2,
           inputRegisters_396__1,inputRegisters_396__0}), .en (
           enableRegister_396), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_396__15,registerOutputs_396__14,
           registerOutputs_396__13,registerOutputs_396__12,
           registerOutputs_396__11,registerOutputs_396__10,
           registerOutputs_396__9,registerOutputs_396__8,registerOutputs_396__7,
           registerOutputs_396__6,registerOutputs_396__5,registerOutputs_396__4,
           registerOutputs_396__3,registerOutputs_396__2,registerOutputs_396__1,
           registerOutputs_396__0})) ;
    Mux2_16 loop1_397_y (.A ({nx35997,nx36139,nx36281,nx36423,nx36565,nx36707,
            nx36849,nx36991,nx37133,nx37275,nx37417,nx37559,nx37701,nx37843,
            nx37985,nx38127}), .B ({nx33753,nx33891,nx34031,nx34169,nx34307,
            nx34445,nx34583,nx34723,nx34865,nx35007,nx35149,nx35291,nx35433,
            nx35575,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35717), .C ({inputRegisters_397__15,inputRegisters_397__14,
            inputRegisters_397__13,inputRegisters_397__12,inputRegisters_397__11
            ,inputRegisters_397__10,inputRegisters_397__9,inputRegisters_397__8,
            inputRegisters_397__7,inputRegisters_397__6,inputRegisters_397__5,
            inputRegisters_397__4,inputRegisters_397__3,inputRegisters_397__2,
            inputRegisters_397__1,inputRegisters_397__0})) ;
    Reg_16 loop1_397_x (.D ({inputRegisters_397__15,inputRegisters_397__14,
           inputRegisters_397__13,inputRegisters_397__12,inputRegisters_397__11,
           inputRegisters_397__10,inputRegisters_397__9,inputRegisters_397__8,
           inputRegisters_397__7,inputRegisters_397__6,inputRegisters_397__5,
           inputRegisters_397__4,inputRegisters_397__3,inputRegisters_397__2,
           inputRegisters_397__1,inputRegisters_397__0}), .en (
           enableRegister_397), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_397__15,registerOutputs_397__14,
           registerOutputs_397__13,registerOutputs_397__12,
           registerOutputs_397__11,registerOutputs_397__10,
           registerOutputs_397__9,registerOutputs_397__8,registerOutputs_397__7,
           registerOutputs_397__6,registerOutputs_397__5,registerOutputs_397__4,
           registerOutputs_397__3,registerOutputs_397__2,registerOutputs_397__1,
           registerOutputs_397__0})) ;
    Mux2_16 loop1_398_y (.A ({nx35997,nx36139,nx36281,nx36423,nx36565,nx36707,
            nx36849,nx36991,nx37133,nx37275,nx37417,nx37559,nx37701,nx37843,
            nx37985,nx38127}), .B ({nx33753,nx33893,nx34031,nx34169,nx34307,
            nx34445,nx34583,nx34723,nx34865,nx35007,nx35149,nx35291,nx35433,
            nx35575,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35717), .C ({inputRegisters_398__15,inputRegisters_398__14,
            inputRegisters_398__13,inputRegisters_398__12,inputRegisters_398__11
            ,inputRegisters_398__10,inputRegisters_398__9,inputRegisters_398__8,
            inputRegisters_398__7,inputRegisters_398__6,inputRegisters_398__5,
            inputRegisters_398__4,inputRegisters_398__3,inputRegisters_398__2,
            inputRegisters_398__1,inputRegisters_398__0})) ;
    Reg_16 loop1_398_x (.D ({inputRegisters_398__15,inputRegisters_398__14,
           inputRegisters_398__13,inputRegisters_398__12,inputRegisters_398__11,
           inputRegisters_398__10,inputRegisters_398__9,inputRegisters_398__8,
           inputRegisters_398__7,inputRegisters_398__6,inputRegisters_398__5,
           inputRegisters_398__4,inputRegisters_398__3,inputRegisters_398__2,
           inputRegisters_398__1,inputRegisters_398__0}), .en (
           enableRegister_398), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_398__15,registerOutputs_398__14,
           registerOutputs_398__13,registerOutputs_398__12,
           registerOutputs_398__11,registerOutputs_398__10,
           registerOutputs_398__9,registerOutputs_398__8,registerOutputs_398__7,
           registerOutputs_398__6,registerOutputs_398__5,registerOutputs_398__4,
           registerOutputs_398__3,registerOutputs_398__2,registerOutputs_398__1,
           registerOutputs_398__0})) ;
    Mux2_16 loop1_399_y (.A ({nx35999,nx36141,nx36283,nx36425,nx36567,nx36709,
            nx36851,nx36993,nx37135,nx37277,nx37419,nx37561,nx37703,nx37845,
            nx37987,nx38129}), .B ({nx33755,nx33893,nx34031,nx34169,nx34307,
            nx34445,nx34583,nx34725,nx34867,nx35009,nx35151,nx35293,nx35435,
            nx35577,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35719), .C ({inputRegisters_399__15,inputRegisters_399__14,
            inputRegisters_399__13,inputRegisters_399__12,inputRegisters_399__11
            ,inputRegisters_399__10,inputRegisters_399__9,inputRegisters_399__8,
            inputRegisters_399__7,inputRegisters_399__6,inputRegisters_399__5,
            inputRegisters_399__4,inputRegisters_399__3,inputRegisters_399__2,
            inputRegisters_399__1,inputRegisters_399__0})) ;
    Reg_16 loop1_399_x (.D ({inputRegisters_399__15,inputRegisters_399__14,
           inputRegisters_399__13,inputRegisters_399__12,inputRegisters_399__11,
           inputRegisters_399__10,inputRegisters_399__9,inputRegisters_399__8,
           inputRegisters_399__7,inputRegisters_399__6,inputRegisters_399__5,
           inputRegisters_399__4,inputRegisters_399__3,inputRegisters_399__2,
           inputRegisters_399__1,inputRegisters_399__0}), .en (
           enableRegister_399), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_399__15,registerOutputs_399__14,
           registerOutputs_399__13,registerOutputs_399__12,
           registerOutputs_399__11,registerOutputs_399__10,
           registerOutputs_399__9,registerOutputs_399__8,registerOutputs_399__7,
           registerOutputs_399__6,registerOutputs_399__5,registerOutputs_399__4,
           registerOutputs_399__3,registerOutputs_399__2,registerOutputs_399__1,
           registerOutputs_399__0})) ;
    Mux2_16 loop1_400_y (.A ({nx35999,nx36141,nx36283,nx36425,nx36567,nx36709,
            nx36851,nx36993,nx37135,nx37277,nx37419,nx37561,nx37703,nx37845,
            nx37987,nx38129}), .B ({nx33755,nx33893,nx34031,nx34169,nx34307,
            nx34445,nx34585,nx34725,nx34867,nx35009,nx35151,nx35293,nx35435,
            nx35577,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35719), .C ({inputRegisters_400__15,inputRegisters_400__14,
            inputRegisters_400__13,inputRegisters_400__12,inputRegisters_400__11
            ,inputRegisters_400__10,inputRegisters_400__9,inputRegisters_400__8,
            inputRegisters_400__7,inputRegisters_400__6,inputRegisters_400__5,
            inputRegisters_400__4,inputRegisters_400__3,inputRegisters_400__2,
            inputRegisters_400__1,inputRegisters_400__0})) ;
    Reg_16 loop1_400_x (.D ({inputRegisters_400__15,inputRegisters_400__14,
           inputRegisters_400__13,inputRegisters_400__12,inputRegisters_400__11,
           inputRegisters_400__10,inputRegisters_400__9,inputRegisters_400__8,
           inputRegisters_400__7,inputRegisters_400__6,inputRegisters_400__5,
           inputRegisters_400__4,inputRegisters_400__3,inputRegisters_400__2,
           inputRegisters_400__1,inputRegisters_400__0}), .en (
           enableRegister_400), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_400__15,registerOutputs_400__14,
           registerOutputs_400__13,registerOutputs_400__12,
           registerOutputs_400__11,registerOutputs_400__10,
           registerOutputs_400__9,registerOutputs_400__8,registerOutputs_400__7,
           registerOutputs_400__6,registerOutputs_400__5,registerOutputs_400__4,
           registerOutputs_400__3,registerOutputs_400__2,registerOutputs_400__1,
           registerOutputs_400__0})) ;
    Mux2_16 loop1_401_y (.A ({nx35999,nx36141,nx36283,nx36425,nx36567,nx36709,
            nx36851,nx36993,nx37135,nx37277,nx37419,nx37561,nx37703,nx37845,
            nx37987,nx38129}), .B ({nx33755,nx33893,nx34031,nx34169,nx34307,
            nx34447,nx34585,nx34725,nx34867,nx35009,nx35151,nx35293,nx35435,
            nx35577,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35719), .C ({inputRegisters_401__15,inputRegisters_401__14,
            inputRegisters_401__13,inputRegisters_401__12,inputRegisters_401__11
            ,inputRegisters_401__10,inputRegisters_401__9,inputRegisters_401__8,
            inputRegisters_401__7,inputRegisters_401__6,inputRegisters_401__5,
            inputRegisters_401__4,inputRegisters_401__3,inputRegisters_401__2,
            inputRegisters_401__1,inputRegisters_401__0})) ;
    Reg_16 loop1_401_x (.D ({inputRegisters_401__15,inputRegisters_401__14,
           inputRegisters_401__13,inputRegisters_401__12,inputRegisters_401__11,
           inputRegisters_401__10,inputRegisters_401__9,inputRegisters_401__8,
           inputRegisters_401__7,inputRegisters_401__6,inputRegisters_401__5,
           inputRegisters_401__4,inputRegisters_401__3,inputRegisters_401__2,
           inputRegisters_401__1,inputRegisters_401__0}), .en (
           enableRegister_401), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_401__15,registerOutputs_401__14,
           registerOutputs_401__13,registerOutputs_401__12,
           registerOutputs_401__11,registerOutputs_401__10,
           registerOutputs_401__9,registerOutputs_401__8,registerOutputs_401__7,
           registerOutputs_401__6,registerOutputs_401__5,registerOutputs_401__4,
           registerOutputs_401__3,registerOutputs_401__2,registerOutputs_401__1,
           registerOutputs_401__0})) ;
    Mux2_16 loop1_402_y (.A ({nx35999,nx36141,nx36283,nx36425,nx36567,nx36709,
            nx36851,nx36993,nx37135,nx37277,nx37419,nx37561,nx37703,nx37845,
            nx37987,nx38129}), .B ({nx33755,nx33893,nx34031,nx34169,nx34309,
            nx34447,nx34585,nx34725,nx34867,nx35009,nx35151,nx35293,nx35435,
            nx35577,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35719), .C ({inputRegisters_402__15,inputRegisters_402__14,
            inputRegisters_402__13,inputRegisters_402__12,inputRegisters_402__11
            ,inputRegisters_402__10,inputRegisters_402__9,inputRegisters_402__8,
            inputRegisters_402__7,inputRegisters_402__6,inputRegisters_402__5,
            inputRegisters_402__4,inputRegisters_402__3,inputRegisters_402__2,
            inputRegisters_402__1,inputRegisters_402__0})) ;
    Reg_16 loop1_402_x (.D ({inputRegisters_402__15,inputRegisters_402__14,
           inputRegisters_402__13,inputRegisters_402__12,inputRegisters_402__11,
           inputRegisters_402__10,inputRegisters_402__9,inputRegisters_402__8,
           inputRegisters_402__7,inputRegisters_402__6,inputRegisters_402__5,
           inputRegisters_402__4,inputRegisters_402__3,inputRegisters_402__2,
           inputRegisters_402__1,inputRegisters_402__0}), .en (
           enableRegister_402), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_402__15,registerOutputs_402__14,
           registerOutputs_402__13,registerOutputs_402__12,
           registerOutputs_402__11,registerOutputs_402__10,
           registerOutputs_402__9,registerOutputs_402__8,registerOutputs_402__7,
           registerOutputs_402__6,registerOutputs_402__5,registerOutputs_402__4,
           registerOutputs_402__3,registerOutputs_402__2,registerOutputs_402__1,
           registerOutputs_402__0})) ;
    Mux2_16 loop1_403_y (.A ({nx35999,nx36141,nx36283,nx36425,nx36567,nx36709,
            nx36851,nx36993,nx37135,nx37277,nx37419,nx37561,nx37703,nx37845,
            nx37987,nx38129}), .B ({nx33755,nx33893,nx34031,nx34171,nx34309,
            nx34447,nx34585,nx34725,nx34867,nx35009,nx35151,nx35293,nx35435,
            nx35577,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35719), .C ({inputRegisters_403__15,inputRegisters_403__14,
            inputRegisters_403__13,inputRegisters_403__12,inputRegisters_403__11
            ,inputRegisters_403__10,inputRegisters_403__9,inputRegisters_403__8,
            inputRegisters_403__7,inputRegisters_403__6,inputRegisters_403__5,
            inputRegisters_403__4,inputRegisters_403__3,inputRegisters_403__2,
            inputRegisters_403__1,inputRegisters_403__0})) ;
    Reg_16 loop1_403_x (.D ({inputRegisters_403__15,inputRegisters_403__14,
           inputRegisters_403__13,inputRegisters_403__12,inputRegisters_403__11,
           inputRegisters_403__10,inputRegisters_403__9,inputRegisters_403__8,
           inputRegisters_403__7,inputRegisters_403__6,inputRegisters_403__5,
           inputRegisters_403__4,inputRegisters_403__3,inputRegisters_403__2,
           inputRegisters_403__1,inputRegisters_403__0}), .en (
           enableRegister_403), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_403__15,registerOutputs_403__14,
           registerOutputs_403__13,registerOutputs_403__12,
           registerOutputs_403__11,registerOutputs_403__10,
           registerOutputs_403__9,registerOutputs_403__8,registerOutputs_403__7,
           registerOutputs_403__6,registerOutputs_403__5,registerOutputs_403__4,
           registerOutputs_403__3,registerOutputs_403__2,registerOutputs_403__1,
           registerOutputs_403__0})) ;
    Mux2_16 loop1_404_y (.A ({nx35999,nx36141,nx36283,nx36425,nx36567,nx36709,
            nx36851,nx36993,nx37135,nx37277,nx37419,nx37561,nx37703,nx37845,
            nx37987,nx38129}), .B ({nx33755,nx33893,nx34033,nx34171,nx34309,
            nx34447,nx34585,nx34725,nx34867,nx35009,nx35151,nx35293,nx35435,
            nx35577,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35719), .C ({inputRegisters_404__15,inputRegisters_404__14,
            inputRegisters_404__13,inputRegisters_404__12,inputRegisters_404__11
            ,inputRegisters_404__10,inputRegisters_404__9,inputRegisters_404__8,
            inputRegisters_404__7,inputRegisters_404__6,inputRegisters_404__5,
            inputRegisters_404__4,inputRegisters_404__3,inputRegisters_404__2,
            inputRegisters_404__1,inputRegisters_404__0})) ;
    Reg_16 loop1_404_x (.D ({inputRegisters_404__15,inputRegisters_404__14,
           inputRegisters_404__13,inputRegisters_404__12,inputRegisters_404__11,
           inputRegisters_404__10,inputRegisters_404__9,inputRegisters_404__8,
           inputRegisters_404__7,inputRegisters_404__6,inputRegisters_404__5,
           inputRegisters_404__4,inputRegisters_404__3,inputRegisters_404__2,
           inputRegisters_404__1,inputRegisters_404__0}), .en (
           enableRegister_404), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_404__15,registerOutputs_404__14,
           registerOutputs_404__13,registerOutputs_404__12,
           registerOutputs_404__11,registerOutputs_404__10,
           registerOutputs_404__9,registerOutputs_404__8,registerOutputs_404__7,
           registerOutputs_404__6,registerOutputs_404__5,registerOutputs_404__4,
           registerOutputs_404__3,registerOutputs_404__2,registerOutputs_404__1,
           registerOutputs_404__0})) ;
    Mux2_16 loop1_405_y (.A ({nx35999,nx36141,nx36283,nx36425,nx36567,nx36709,
            nx36851,nx36993,nx37135,nx37277,nx37419,nx37561,nx37703,nx37845,
            nx37987,nx38129}), .B ({nx33755,nx33895,nx34033,nx34171,nx34309,
            nx34447,nx34585,nx34725,nx34867,nx35009,nx35151,nx35293,nx35435,
            nx35577,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35719), .C ({inputRegisters_405__15,inputRegisters_405__14,
            inputRegisters_405__13,inputRegisters_405__12,inputRegisters_405__11
            ,inputRegisters_405__10,inputRegisters_405__9,inputRegisters_405__8,
            inputRegisters_405__7,inputRegisters_405__6,inputRegisters_405__5,
            inputRegisters_405__4,inputRegisters_405__3,inputRegisters_405__2,
            inputRegisters_405__1,inputRegisters_405__0})) ;
    Reg_16 loop1_405_x (.D ({inputRegisters_405__15,inputRegisters_405__14,
           inputRegisters_405__13,inputRegisters_405__12,inputRegisters_405__11,
           inputRegisters_405__10,inputRegisters_405__9,inputRegisters_405__8,
           inputRegisters_405__7,inputRegisters_405__6,inputRegisters_405__5,
           inputRegisters_405__4,inputRegisters_405__3,inputRegisters_405__2,
           inputRegisters_405__1,inputRegisters_405__0}), .en (
           enableRegister_405), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_405__15,registerOutputs_405__14,
           registerOutputs_405__13,registerOutputs_405__12,
           registerOutputs_405__11,registerOutputs_405__10,
           registerOutputs_405__9,registerOutputs_405__8,registerOutputs_405__7,
           registerOutputs_405__6,registerOutputs_405__5,registerOutputs_405__4,
           registerOutputs_405__3,registerOutputs_405__2,registerOutputs_405__1,
           registerOutputs_405__0})) ;
    Mux2_16 loop1_406_y (.A ({nx36001,nx36143,nx36285,nx36427,nx36569,nx36711,
            nx36853,nx36995,nx37137,nx37279,nx37421,nx37563,nx37705,nx37847,
            nx37989,nx38131}), .B ({nx33757,nx33895,nx34033,nx34171,nx34309,
            nx34447,nx34585,nx34727,nx34869,nx35011,nx35153,nx35295,nx35437,
            nx35579,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35721), .C ({inputRegisters_406__15,inputRegisters_406__14,
            inputRegisters_406__13,inputRegisters_406__12,inputRegisters_406__11
            ,inputRegisters_406__10,inputRegisters_406__9,inputRegisters_406__8,
            inputRegisters_406__7,inputRegisters_406__6,inputRegisters_406__5,
            inputRegisters_406__4,inputRegisters_406__3,inputRegisters_406__2,
            inputRegisters_406__1,inputRegisters_406__0})) ;
    Reg_16 loop1_406_x (.D ({inputRegisters_406__15,inputRegisters_406__14,
           inputRegisters_406__13,inputRegisters_406__12,inputRegisters_406__11,
           inputRegisters_406__10,inputRegisters_406__9,inputRegisters_406__8,
           inputRegisters_406__7,inputRegisters_406__6,inputRegisters_406__5,
           inputRegisters_406__4,inputRegisters_406__3,inputRegisters_406__2,
           inputRegisters_406__1,inputRegisters_406__0}), .en (
           enableRegister_406), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_406__15,registerOutputs_406__14,
           registerOutputs_406__13,registerOutputs_406__12,
           registerOutputs_406__11,registerOutputs_406__10,
           registerOutputs_406__9,registerOutputs_406__8,registerOutputs_406__7,
           registerOutputs_406__6,registerOutputs_406__5,registerOutputs_406__4,
           registerOutputs_406__3,registerOutputs_406__2,registerOutputs_406__1,
           registerOutputs_406__0})) ;
    Mux2_16 loop1_407_y (.A ({nx36001,nx36143,nx36285,nx36427,nx36569,nx36711,
            nx36853,nx36995,nx37137,nx37279,nx37421,nx37563,nx37705,nx37847,
            nx37989,nx38131}), .B ({nx33757,nx33895,nx34033,nx34171,nx34309,
            nx34447,nx34587,nx34727,nx34869,nx35011,nx35153,nx35295,nx35437,
            nx35579,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35721), .C ({inputRegisters_407__15,inputRegisters_407__14,
            inputRegisters_407__13,inputRegisters_407__12,inputRegisters_407__11
            ,inputRegisters_407__10,inputRegisters_407__9,inputRegisters_407__8,
            inputRegisters_407__7,inputRegisters_407__6,inputRegisters_407__5,
            inputRegisters_407__4,inputRegisters_407__3,inputRegisters_407__2,
            inputRegisters_407__1,inputRegisters_407__0})) ;
    Reg_16 loop1_407_x (.D ({inputRegisters_407__15,inputRegisters_407__14,
           inputRegisters_407__13,inputRegisters_407__12,inputRegisters_407__11,
           inputRegisters_407__10,inputRegisters_407__9,inputRegisters_407__8,
           inputRegisters_407__7,inputRegisters_407__6,inputRegisters_407__5,
           inputRegisters_407__4,inputRegisters_407__3,inputRegisters_407__2,
           inputRegisters_407__1,inputRegisters_407__0}), .en (
           enableRegister_407), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_407__15,registerOutputs_407__14,
           registerOutputs_407__13,registerOutputs_407__12,
           registerOutputs_407__11,registerOutputs_407__10,
           registerOutputs_407__9,registerOutputs_407__8,registerOutputs_407__7,
           registerOutputs_407__6,registerOutputs_407__5,registerOutputs_407__4,
           registerOutputs_407__3,registerOutputs_407__2,registerOutputs_407__1,
           registerOutputs_407__0})) ;
    Mux2_16 loop1_408_y (.A ({nx36001,nx36143,nx36285,nx36427,nx36569,nx36711,
            nx36853,nx36995,nx37137,nx37279,nx37421,nx37563,nx37705,nx37847,
            nx37989,nx38131}), .B ({nx33757,nx33895,nx34033,nx34171,nx34309,
            nx34449,nx34587,nx34727,nx34869,nx35011,nx35153,nx35295,nx35437,
            nx35579,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35721), .C ({inputRegisters_408__15,inputRegisters_408__14,
            inputRegisters_408__13,inputRegisters_408__12,inputRegisters_408__11
            ,inputRegisters_408__10,inputRegisters_408__9,inputRegisters_408__8,
            inputRegisters_408__7,inputRegisters_408__6,inputRegisters_408__5,
            inputRegisters_408__4,inputRegisters_408__3,inputRegisters_408__2,
            inputRegisters_408__1,inputRegisters_408__0})) ;
    Reg_16 loop1_408_x (.D ({inputRegisters_408__15,inputRegisters_408__14,
           inputRegisters_408__13,inputRegisters_408__12,inputRegisters_408__11,
           inputRegisters_408__10,inputRegisters_408__9,inputRegisters_408__8,
           inputRegisters_408__7,inputRegisters_408__6,inputRegisters_408__5,
           inputRegisters_408__4,inputRegisters_408__3,inputRegisters_408__2,
           inputRegisters_408__1,inputRegisters_408__0}), .en (
           enableRegister_408), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_408__15,registerOutputs_408__14,
           registerOutputs_408__13,registerOutputs_408__12,
           registerOutputs_408__11,registerOutputs_408__10,
           registerOutputs_408__9,registerOutputs_408__8,registerOutputs_408__7,
           registerOutputs_408__6,registerOutputs_408__5,registerOutputs_408__4,
           registerOutputs_408__3,registerOutputs_408__2,registerOutputs_408__1,
           registerOutputs_408__0})) ;
    Mux2_16 loop1_409_y (.A ({nx36001,nx36143,nx36285,nx36427,nx36569,nx36711,
            nx36853,nx36995,nx37137,nx37279,nx37421,nx37563,nx37705,nx37847,
            nx37989,nx38131}), .B ({nx33757,nx33895,nx34033,nx34171,nx34311,
            nx34449,nx34587,nx34727,nx34869,nx35011,nx35153,nx35295,nx35437,
            nx35579,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35721), .C ({inputRegisters_409__15,inputRegisters_409__14,
            inputRegisters_409__13,inputRegisters_409__12,inputRegisters_409__11
            ,inputRegisters_409__10,inputRegisters_409__9,inputRegisters_409__8,
            inputRegisters_409__7,inputRegisters_409__6,inputRegisters_409__5,
            inputRegisters_409__4,inputRegisters_409__3,inputRegisters_409__2,
            inputRegisters_409__1,inputRegisters_409__0})) ;
    Reg_16 loop1_409_x (.D ({inputRegisters_409__15,inputRegisters_409__14,
           inputRegisters_409__13,inputRegisters_409__12,inputRegisters_409__11,
           inputRegisters_409__10,inputRegisters_409__9,inputRegisters_409__8,
           inputRegisters_409__7,inputRegisters_409__6,inputRegisters_409__5,
           inputRegisters_409__4,inputRegisters_409__3,inputRegisters_409__2,
           inputRegisters_409__1,inputRegisters_409__0}), .en (
           enableRegister_409), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_409__15,registerOutputs_409__14,
           registerOutputs_409__13,registerOutputs_409__12,
           registerOutputs_409__11,registerOutputs_409__10,
           registerOutputs_409__9,registerOutputs_409__8,registerOutputs_409__7,
           registerOutputs_409__6,registerOutputs_409__5,registerOutputs_409__4,
           registerOutputs_409__3,registerOutputs_409__2,registerOutputs_409__1,
           registerOutputs_409__0})) ;
    Mux2_16 loop1_410_y (.A ({nx36001,nx36143,nx36285,nx36427,nx36569,nx36711,
            nx36853,nx36995,nx37137,nx37279,nx37421,nx37563,nx37705,nx37847,
            nx37989,nx38131}), .B ({nx33757,nx33895,nx34033,nx34173,nx34311,
            nx34449,nx34587,nx34727,nx34869,nx35011,nx35153,nx35295,nx35437,
            nx35579,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35721), .C ({inputRegisters_410__15,inputRegisters_410__14,
            inputRegisters_410__13,inputRegisters_410__12,inputRegisters_410__11
            ,inputRegisters_410__10,inputRegisters_410__9,inputRegisters_410__8,
            inputRegisters_410__7,inputRegisters_410__6,inputRegisters_410__5,
            inputRegisters_410__4,inputRegisters_410__3,inputRegisters_410__2,
            inputRegisters_410__1,inputRegisters_410__0})) ;
    Reg_16 loop1_410_x (.D ({inputRegisters_410__15,inputRegisters_410__14,
           inputRegisters_410__13,inputRegisters_410__12,inputRegisters_410__11,
           inputRegisters_410__10,inputRegisters_410__9,inputRegisters_410__8,
           inputRegisters_410__7,inputRegisters_410__6,inputRegisters_410__5,
           inputRegisters_410__4,inputRegisters_410__3,inputRegisters_410__2,
           inputRegisters_410__1,inputRegisters_410__0}), .en (
           enableRegister_410), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_410__15,registerOutputs_410__14,
           registerOutputs_410__13,registerOutputs_410__12,
           registerOutputs_410__11,registerOutputs_410__10,
           registerOutputs_410__9,registerOutputs_410__8,registerOutputs_410__7,
           registerOutputs_410__6,registerOutputs_410__5,registerOutputs_410__4,
           registerOutputs_410__3,registerOutputs_410__2,registerOutputs_410__1,
           registerOutputs_410__0})) ;
    Mux2_16 loop1_411_y (.A ({nx36001,nx36143,nx36285,nx36427,nx36569,nx36711,
            nx36853,nx36995,nx37137,nx37279,nx37421,nx37563,nx37705,nx37847,
            nx37989,nx38131}), .B ({nx33757,nx33895,nx34035,nx34173,nx34311,
            nx34449,nx34587,nx34727,nx34869,nx35011,nx35153,nx35295,nx35437,
            nx35579,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35721), .C ({inputRegisters_411__15,inputRegisters_411__14,
            inputRegisters_411__13,inputRegisters_411__12,inputRegisters_411__11
            ,inputRegisters_411__10,inputRegisters_411__9,inputRegisters_411__8,
            inputRegisters_411__7,inputRegisters_411__6,inputRegisters_411__5,
            inputRegisters_411__4,inputRegisters_411__3,inputRegisters_411__2,
            inputRegisters_411__1,inputRegisters_411__0})) ;
    Reg_16 loop1_411_x (.D ({inputRegisters_411__15,inputRegisters_411__14,
           inputRegisters_411__13,inputRegisters_411__12,inputRegisters_411__11,
           inputRegisters_411__10,inputRegisters_411__9,inputRegisters_411__8,
           inputRegisters_411__7,inputRegisters_411__6,inputRegisters_411__5,
           inputRegisters_411__4,inputRegisters_411__3,inputRegisters_411__2,
           inputRegisters_411__1,inputRegisters_411__0}), .en (
           enableRegister_411), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_411__15,registerOutputs_411__14,
           registerOutputs_411__13,registerOutputs_411__12,
           registerOutputs_411__11,registerOutputs_411__10,
           registerOutputs_411__9,registerOutputs_411__8,registerOutputs_411__7,
           registerOutputs_411__6,registerOutputs_411__5,registerOutputs_411__4,
           registerOutputs_411__3,registerOutputs_411__2,registerOutputs_411__1,
           registerOutputs_411__0})) ;
    Mux2_16 loop1_412_y (.A ({nx36001,nx36143,nx36285,nx36427,nx36569,nx36711,
            nx36853,nx36995,nx37137,nx37279,nx37421,nx37563,nx37705,nx37847,
            nx37989,nx38131}), .B ({nx33757,nx33897,nx34035,nx34173,nx34311,
            nx34449,nx34587,nx34727,nx34869,nx35011,nx35153,nx35295,nx35437,
            nx35579,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35721), .C ({inputRegisters_412__15,inputRegisters_412__14,
            inputRegisters_412__13,inputRegisters_412__12,inputRegisters_412__11
            ,inputRegisters_412__10,inputRegisters_412__9,inputRegisters_412__8,
            inputRegisters_412__7,inputRegisters_412__6,inputRegisters_412__5,
            inputRegisters_412__4,inputRegisters_412__3,inputRegisters_412__2,
            inputRegisters_412__1,inputRegisters_412__0})) ;
    Reg_16 loop1_412_x (.D ({inputRegisters_412__15,inputRegisters_412__14,
           inputRegisters_412__13,inputRegisters_412__12,inputRegisters_412__11,
           inputRegisters_412__10,inputRegisters_412__9,inputRegisters_412__8,
           inputRegisters_412__7,inputRegisters_412__6,inputRegisters_412__5,
           inputRegisters_412__4,inputRegisters_412__3,inputRegisters_412__2,
           inputRegisters_412__1,inputRegisters_412__0}), .en (
           enableRegister_412), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_412__15,registerOutputs_412__14,
           registerOutputs_412__13,registerOutputs_412__12,
           registerOutputs_412__11,registerOutputs_412__10,
           registerOutputs_412__9,registerOutputs_412__8,registerOutputs_412__7,
           registerOutputs_412__6,registerOutputs_412__5,registerOutputs_412__4,
           registerOutputs_412__3,registerOutputs_412__2,registerOutputs_412__1,
           registerOutputs_412__0})) ;
    Mux2_16 loop1_413_y (.A ({nx36003,nx36145,nx36287,nx36429,nx36571,nx36713,
            nx36855,nx36997,nx37139,nx37281,nx37423,nx37565,nx37707,nx37849,
            nx37991,nx38133}), .B ({nx33759,nx33897,nx34035,nx34173,nx34311,
            nx34449,nx34587,nx34729,nx34871,nx35013,nx35155,nx35297,nx35439,
            nx35581,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35723), .C ({inputRegisters_413__15,inputRegisters_413__14,
            inputRegisters_413__13,inputRegisters_413__12,inputRegisters_413__11
            ,inputRegisters_413__10,inputRegisters_413__9,inputRegisters_413__8,
            inputRegisters_413__7,inputRegisters_413__6,inputRegisters_413__5,
            inputRegisters_413__4,inputRegisters_413__3,inputRegisters_413__2,
            inputRegisters_413__1,inputRegisters_413__0})) ;
    Reg_16 loop1_413_x (.D ({inputRegisters_413__15,inputRegisters_413__14,
           inputRegisters_413__13,inputRegisters_413__12,inputRegisters_413__11,
           inputRegisters_413__10,inputRegisters_413__9,inputRegisters_413__8,
           inputRegisters_413__7,inputRegisters_413__6,inputRegisters_413__5,
           inputRegisters_413__4,inputRegisters_413__3,inputRegisters_413__2,
           inputRegisters_413__1,inputRegisters_413__0}), .en (
           enableRegister_413), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_413__15,registerOutputs_413__14,
           registerOutputs_413__13,registerOutputs_413__12,
           registerOutputs_413__11,registerOutputs_413__10,
           registerOutputs_413__9,registerOutputs_413__8,registerOutputs_413__7,
           registerOutputs_413__6,registerOutputs_413__5,registerOutputs_413__4,
           registerOutputs_413__3,registerOutputs_413__2,registerOutputs_413__1,
           registerOutputs_413__0})) ;
    Mux2_16 loop1_414_y (.A ({nx36003,nx36145,nx36287,nx36429,nx36571,nx36713,
            nx36855,nx36997,nx37139,nx37281,nx37423,nx37565,nx37707,nx37849,
            nx37991,nx38133}), .B ({nx33759,nx33897,nx34035,nx34173,nx34311,
            nx34449,nx34589,nx34729,nx34871,nx35013,nx35155,nx35297,nx35439,
            nx35581,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35723), .C ({inputRegisters_414__15,inputRegisters_414__14,
            inputRegisters_414__13,inputRegisters_414__12,inputRegisters_414__11
            ,inputRegisters_414__10,inputRegisters_414__9,inputRegisters_414__8,
            inputRegisters_414__7,inputRegisters_414__6,inputRegisters_414__5,
            inputRegisters_414__4,inputRegisters_414__3,inputRegisters_414__2,
            inputRegisters_414__1,inputRegisters_414__0})) ;
    Reg_16 loop1_414_x (.D ({inputRegisters_414__15,inputRegisters_414__14,
           inputRegisters_414__13,inputRegisters_414__12,inputRegisters_414__11,
           inputRegisters_414__10,inputRegisters_414__9,inputRegisters_414__8,
           inputRegisters_414__7,inputRegisters_414__6,inputRegisters_414__5,
           inputRegisters_414__4,inputRegisters_414__3,inputRegisters_414__2,
           inputRegisters_414__1,inputRegisters_414__0}), .en (
           enableRegister_414), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_414__15,registerOutputs_414__14,
           registerOutputs_414__13,registerOutputs_414__12,
           registerOutputs_414__11,registerOutputs_414__10,
           registerOutputs_414__9,registerOutputs_414__8,registerOutputs_414__7,
           registerOutputs_414__6,registerOutputs_414__5,registerOutputs_414__4,
           registerOutputs_414__3,registerOutputs_414__2,registerOutputs_414__1,
           registerOutputs_414__0})) ;
    Mux2_16 loop1_415_y (.A ({nx36003,nx36145,nx36287,nx36429,nx36571,nx36713,
            nx36855,nx36997,nx37139,nx37281,nx37423,nx37565,nx37707,nx37849,
            nx37991,nx38133}), .B ({nx33759,nx33897,nx34035,nx34173,nx34311,
            nx34451,nx34589,nx34729,nx34871,nx35013,nx35155,nx35297,nx35439,
            nx35581,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35723), .C ({inputRegisters_415__15,inputRegisters_415__14,
            inputRegisters_415__13,inputRegisters_415__12,inputRegisters_415__11
            ,inputRegisters_415__10,inputRegisters_415__9,inputRegisters_415__8,
            inputRegisters_415__7,inputRegisters_415__6,inputRegisters_415__5,
            inputRegisters_415__4,inputRegisters_415__3,inputRegisters_415__2,
            inputRegisters_415__1,inputRegisters_415__0})) ;
    Reg_16 loop1_415_x (.D ({inputRegisters_415__15,inputRegisters_415__14,
           inputRegisters_415__13,inputRegisters_415__12,inputRegisters_415__11,
           inputRegisters_415__10,inputRegisters_415__9,inputRegisters_415__8,
           inputRegisters_415__7,inputRegisters_415__6,inputRegisters_415__5,
           inputRegisters_415__4,inputRegisters_415__3,inputRegisters_415__2,
           inputRegisters_415__1,inputRegisters_415__0}), .en (
           enableRegister_415), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_415__15,registerOutputs_415__14,
           registerOutputs_415__13,registerOutputs_415__12,
           registerOutputs_415__11,registerOutputs_415__10,
           registerOutputs_415__9,registerOutputs_415__8,registerOutputs_415__7,
           registerOutputs_415__6,registerOutputs_415__5,registerOutputs_415__4,
           registerOutputs_415__3,registerOutputs_415__2,registerOutputs_415__1,
           registerOutputs_415__0})) ;
    Mux2_16 loop1_416_y (.A ({nx36003,nx36145,nx36287,nx36429,nx36571,nx36713,
            nx36855,nx36997,nx37139,nx37281,nx37423,nx37565,nx37707,nx37849,
            nx37991,nx38133}), .B ({nx33759,nx33897,nx34035,nx34173,nx34313,
            nx34451,nx34589,nx34729,nx34871,nx35013,nx35155,nx35297,nx35439,
            nx35581,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35723), .C ({inputRegisters_416__15,inputRegisters_416__14,
            inputRegisters_416__13,inputRegisters_416__12,inputRegisters_416__11
            ,inputRegisters_416__10,inputRegisters_416__9,inputRegisters_416__8,
            inputRegisters_416__7,inputRegisters_416__6,inputRegisters_416__5,
            inputRegisters_416__4,inputRegisters_416__3,inputRegisters_416__2,
            inputRegisters_416__1,inputRegisters_416__0})) ;
    Reg_16 loop1_416_x (.D ({inputRegisters_416__15,inputRegisters_416__14,
           inputRegisters_416__13,inputRegisters_416__12,inputRegisters_416__11,
           inputRegisters_416__10,inputRegisters_416__9,inputRegisters_416__8,
           inputRegisters_416__7,inputRegisters_416__6,inputRegisters_416__5,
           inputRegisters_416__4,inputRegisters_416__3,inputRegisters_416__2,
           inputRegisters_416__1,inputRegisters_416__0}), .en (
           enableRegister_416), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_416__15,registerOutputs_416__14,
           registerOutputs_416__13,registerOutputs_416__12,
           registerOutputs_416__11,registerOutputs_416__10,
           registerOutputs_416__9,registerOutputs_416__8,registerOutputs_416__7,
           registerOutputs_416__6,registerOutputs_416__5,registerOutputs_416__4,
           registerOutputs_416__3,registerOutputs_416__2,registerOutputs_416__1,
           registerOutputs_416__0})) ;
    Mux2_16 loop1_417_y (.A ({nx36003,nx36145,nx36287,nx36429,nx36571,nx36713,
            nx36855,nx36997,nx37139,nx37281,nx37423,nx37565,nx37707,nx37849,
            nx37991,nx38133}), .B ({nx33759,nx33897,nx34035,nx34175,nx34313,
            nx34451,nx34589,nx34729,nx34871,nx35013,nx35155,nx35297,nx35439,
            nx35581,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35723), .C ({inputRegisters_417__15,inputRegisters_417__14,
            inputRegisters_417__13,inputRegisters_417__12,inputRegisters_417__11
            ,inputRegisters_417__10,inputRegisters_417__9,inputRegisters_417__8,
            inputRegisters_417__7,inputRegisters_417__6,inputRegisters_417__5,
            inputRegisters_417__4,inputRegisters_417__3,inputRegisters_417__2,
            inputRegisters_417__1,inputRegisters_417__0})) ;
    Reg_16 loop1_417_x (.D ({inputRegisters_417__15,inputRegisters_417__14,
           inputRegisters_417__13,inputRegisters_417__12,inputRegisters_417__11,
           inputRegisters_417__10,inputRegisters_417__9,inputRegisters_417__8,
           inputRegisters_417__7,inputRegisters_417__6,inputRegisters_417__5,
           inputRegisters_417__4,inputRegisters_417__3,inputRegisters_417__2,
           inputRegisters_417__1,inputRegisters_417__0}), .en (
           enableRegister_417), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_417__15,registerOutputs_417__14,
           registerOutputs_417__13,registerOutputs_417__12,
           registerOutputs_417__11,registerOutputs_417__10,
           registerOutputs_417__9,registerOutputs_417__8,registerOutputs_417__7,
           registerOutputs_417__6,registerOutputs_417__5,registerOutputs_417__4,
           registerOutputs_417__3,registerOutputs_417__2,registerOutputs_417__1,
           registerOutputs_417__0})) ;
    Mux2_16 loop1_418_y (.A ({nx36003,nx36145,nx36287,nx36429,nx36571,nx36713,
            nx36855,nx36997,nx37139,nx37281,nx37423,nx37565,nx37707,nx37849,
            nx37991,nx38133}), .B ({nx33759,nx33897,nx34037,nx34175,nx34313,
            nx34451,nx34589,nx34729,nx34871,nx35013,nx35155,nx35297,nx35439,
            nx35581,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35723), .C ({inputRegisters_418__15,inputRegisters_418__14,
            inputRegisters_418__13,inputRegisters_418__12,inputRegisters_418__11
            ,inputRegisters_418__10,inputRegisters_418__9,inputRegisters_418__8,
            inputRegisters_418__7,inputRegisters_418__6,inputRegisters_418__5,
            inputRegisters_418__4,inputRegisters_418__3,inputRegisters_418__2,
            inputRegisters_418__1,inputRegisters_418__0})) ;
    Reg_16 loop1_418_x (.D ({inputRegisters_418__15,inputRegisters_418__14,
           inputRegisters_418__13,inputRegisters_418__12,inputRegisters_418__11,
           inputRegisters_418__10,inputRegisters_418__9,inputRegisters_418__8,
           inputRegisters_418__7,inputRegisters_418__6,inputRegisters_418__5,
           inputRegisters_418__4,inputRegisters_418__3,inputRegisters_418__2,
           inputRegisters_418__1,inputRegisters_418__0}), .en (
           enableRegister_418), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_418__15,registerOutputs_418__14,
           registerOutputs_418__13,registerOutputs_418__12,
           registerOutputs_418__11,registerOutputs_418__10,
           registerOutputs_418__9,registerOutputs_418__8,registerOutputs_418__7,
           registerOutputs_418__6,registerOutputs_418__5,registerOutputs_418__4,
           registerOutputs_418__3,registerOutputs_418__2,registerOutputs_418__1,
           registerOutputs_418__0})) ;
    Mux2_16 loop1_419_y (.A ({nx36003,nx36145,nx36287,nx36429,nx36571,nx36713,
            nx36855,nx36997,nx37139,nx37281,nx37423,nx37565,nx37707,nx37849,
            nx37991,nx38133}), .B ({nx33759,nx33899,nx34037,nx34175,nx34313,
            nx34451,nx34589,nx34729,nx34871,nx35013,nx35155,nx35297,nx35439,
            nx35581,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35723), .C ({inputRegisters_419__15,inputRegisters_419__14,
            inputRegisters_419__13,inputRegisters_419__12,inputRegisters_419__11
            ,inputRegisters_419__10,inputRegisters_419__9,inputRegisters_419__8,
            inputRegisters_419__7,inputRegisters_419__6,inputRegisters_419__5,
            inputRegisters_419__4,inputRegisters_419__3,inputRegisters_419__2,
            inputRegisters_419__1,inputRegisters_419__0})) ;
    Reg_16 loop1_419_x (.D ({inputRegisters_419__15,inputRegisters_419__14,
           inputRegisters_419__13,inputRegisters_419__12,inputRegisters_419__11,
           inputRegisters_419__10,inputRegisters_419__9,inputRegisters_419__8,
           inputRegisters_419__7,inputRegisters_419__6,inputRegisters_419__5,
           inputRegisters_419__4,inputRegisters_419__3,inputRegisters_419__2,
           inputRegisters_419__1,inputRegisters_419__0}), .en (
           enableRegister_419), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_419__15,registerOutputs_419__14,
           registerOutputs_419__13,registerOutputs_419__12,
           registerOutputs_419__11,registerOutputs_419__10,
           registerOutputs_419__9,registerOutputs_419__8,registerOutputs_419__7,
           registerOutputs_419__6,registerOutputs_419__5,registerOutputs_419__4,
           registerOutputs_419__3,registerOutputs_419__2,registerOutputs_419__1,
           registerOutputs_419__0})) ;
    Mux2_16 loop1_420_y (.A ({nx36005,nx36147,nx36289,nx36431,nx36573,nx36715,
            nx36857,nx36999,nx37141,nx37283,nx37425,nx37567,nx37709,nx37851,
            nx37993,nx38135}), .B ({nx33761,nx33899,nx34037,nx34175,nx34313,
            nx34451,nx34589,nx34731,nx34873,nx35015,nx35157,nx35299,nx35441,
            nx35583,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35725), .C ({inputRegisters_420__15,inputRegisters_420__14,
            inputRegisters_420__13,inputRegisters_420__12,inputRegisters_420__11
            ,inputRegisters_420__10,inputRegisters_420__9,inputRegisters_420__8,
            inputRegisters_420__7,inputRegisters_420__6,inputRegisters_420__5,
            inputRegisters_420__4,inputRegisters_420__3,inputRegisters_420__2,
            inputRegisters_420__1,inputRegisters_420__0})) ;
    Reg_16 loop1_420_x (.D ({inputRegisters_420__15,inputRegisters_420__14,
           inputRegisters_420__13,inputRegisters_420__12,inputRegisters_420__11,
           inputRegisters_420__10,inputRegisters_420__9,inputRegisters_420__8,
           inputRegisters_420__7,inputRegisters_420__6,inputRegisters_420__5,
           inputRegisters_420__4,inputRegisters_420__3,inputRegisters_420__2,
           inputRegisters_420__1,inputRegisters_420__0}), .en (
           enableRegister_420), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_420__15,registerOutputs_420__14,
           registerOutputs_420__13,registerOutputs_420__12,
           registerOutputs_420__11,registerOutputs_420__10,
           registerOutputs_420__9,registerOutputs_420__8,registerOutputs_420__7,
           registerOutputs_420__6,registerOutputs_420__5,registerOutputs_420__4,
           registerOutputs_420__3,registerOutputs_420__2,registerOutputs_420__1,
           registerOutputs_420__0})) ;
    Mux2_16 loop1_421_y (.A ({nx36005,nx36147,nx36289,nx36431,nx36573,nx36715,
            nx36857,nx36999,nx37141,nx37283,nx37425,nx37567,nx37709,nx37851,
            nx37993,nx38135}), .B ({nx33761,nx33899,nx34037,nx34175,nx34313,
            nx34451,nx34591,nx34731,nx34873,nx35015,nx35157,nx35299,nx35441,
            nx35583,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35725), .C ({inputRegisters_421__15,inputRegisters_421__14,
            inputRegisters_421__13,inputRegisters_421__12,inputRegisters_421__11
            ,inputRegisters_421__10,inputRegisters_421__9,inputRegisters_421__8,
            inputRegisters_421__7,inputRegisters_421__6,inputRegisters_421__5,
            inputRegisters_421__4,inputRegisters_421__3,inputRegisters_421__2,
            inputRegisters_421__1,inputRegisters_421__0})) ;
    Reg_16 loop1_421_x (.D ({inputRegisters_421__15,inputRegisters_421__14,
           inputRegisters_421__13,inputRegisters_421__12,inputRegisters_421__11,
           inputRegisters_421__10,inputRegisters_421__9,inputRegisters_421__8,
           inputRegisters_421__7,inputRegisters_421__6,inputRegisters_421__5,
           inputRegisters_421__4,inputRegisters_421__3,inputRegisters_421__2,
           inputRegisters_421__1,inputRegisters_421__0}), .en (
           enableRegister_421), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_421__15,registerOutputs_421__14,
           registerOutputs_421__13,registerOutputs_421__12,
           registerOutputs_421__11,registerOutputs_421__10,
           registerOutputs_421__9,registerOutputs_421__8,registerOutputs_421__7,
           registerOutputs_421__6,registerOutputs_421__5,registerOutputs_421__4,
           registerOutputs_421__3,registerOutputs_421__2,registerOutputs_421__1,
           registerOutputs_421__0})) ;
    Mux2_16 loop1_422_y (.A ({nx36005,nx36147,nx36289,nx36431,nx36573,nx36715,
            nx36857,nx36999,nx37141,nx37283,nx37425,nx37567,nx37709,nx37851,
            nx37993,nx38135}), .B ({nx33761,nx33899,nx34037,nx34175,nx34313,
            nx34453,nx34591,nx34731,nx34873,nx35015,nx35157,nx35299,nx35441,
            nx35583,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35725), .C ({inputRegisters_422__15,inputRegisters_422__14,
            inputRegisters_422__13,inputRegisters_422__12,inputRegisters_422__11
            ,inputRegisters_422__10,inputRegisters_422__9,inputRegisters_422__8,
            inputRegisters_422__7,inputRegisters_422__6,inputRegisters_422__5,
            inputRegisters_422__4,inputRegisters_422__3,inputRegisters_422__2,
            inputRegisters_422__1,inputRegisters_422__0})) ;
    Reg_16 loop1_422_x (.D ({inputRegisters_422__15,inputRegisters_422__14,
           inputRegisters_422__13,inputRegisters_422__12,inputRegisters_422__11,
           inputRegisters_422__10,inputRegisters_422__9,inputRegisters_422__8,
           inputRegisters_422__7,inputRegisters_422__6,inputRegisters_422__5,
           inputRegisters_422__4,inputRegisters_422__3,inputRegisters_422__2,
           inputRegisters_422__1,inputRegisters_422__0}), .en (
           enableRegister_422), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_422__15,registerOutputs_422__14,
           registerOutputs_422__13,registerOutputs_422__12,
           registerOutputs_422__11,registerOutputs_422__10,
           registerOutputs_422__9,registerOutputs_422__8,registerOutputs_422__7,
           registerOutputs_422__6,registerOutputs_422__5,registerOutputs_422__4,
           registerOutputs_422__3,registerOutputs_422__2,registerOutputs_422__1,
           registerOutputs_422__0})) ;
    Mux2_16 loop1_423_y (.A ({nx36005,nx36147,nx36289,nx36431,nx36573,nx36715,
            nx36857,nx36999,nx37141,nx37283,nx37425,nx37567,nx37709,nx37851,
            nx37993,nx38135}), .B ({nx33761,nx33899,nx34037,nx34175,nx34315,
            nx34453,nx34591,nx34731,nx34873,nx35015,nx35157,nx35299,nx35441,
            nx35583,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35725), .C ({inputRegisters_423__15,inputRegisters_423__14,
            inputRegisters_423__13,inputRegisters_423__12,inputRegisters_423__11
            ,inputRegisters_423__10,inputRegisters_423__9,inputRegisters_423__8,
            inputRegisters_423__7,inputRegisters_423__6,inputRegisters_423__5,
            inputRegisters_423__4,inputRegisters_423__3,inputRegisters_423__2,
            inputRegisters_423__1,inputRegisters_423__0})) ;
    Reg_16 loop1_423_x (.D ({inputRegisters_423__15,inputRegisters_423__14,
           inputRegisters_423__13,inputRegisters_423__12,inputRegisters_423__11,
           inputRegisters_423__10,inputRegisters_423__9,inputRegisters_423__8,
           inputRegisters_423__7,inputRegisters_423__6,inputRegisters_423__5,
           inputRegisters_423__4,inputRegisters_423__3,inputRegisters_423__2,
           inputRegisters_423__1,inputRegisters_423__0}), .en (
           enableRegister_423), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_423__15,registerOutputs_423__14,
           registerOutputs_423__13,registerOutputs_423__12,
           registerOutputs_423__11,registerOutputs_423__10,
           registerOutputs_423__9,registerOutputs_423__8,registerOutputs_423__7,
           registerOutputs_423__6,registerOutputs_423__5,registerOutputs_423__4,
           registerOutputs_423__3,registerOutputs_423__2,registerOutputs_423__1,
           registerOutputs_423__0})) ;
    Mux2_16 loop1_424_y (.A ({nx36005,nx36147,nx36289,nx36431,nx36573,nx36715,
            nx36857,nx36999,nx37141,nx37283,nx37425,nx37567,nx37709,nx37851,
            nx37993,nx38135}), .B ({nx33761,nx33899,nx34037,nx34177,nx34315,
            nx34453,nx34591,nx34731,nx34873,nx35015,nx35157,nx35299,nx35441,
            nx35583,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35725), .C ({inputRegisters_424__15,inputRegisters_424__14,
            inputRegisters_424__13,inputRegisters_424__12,inputRegisters_424__11
            ,inputRegisters_424__10,inputRegisters_424__9,inputRegisters_424__8,
            inputRegisters_424__7,inputRegisters_424__6,inputRegisters_424__5,
            inputRegisters_424__4,inputRegisters_424__3,inputRegisters_424__2,
            inputRegisters_424__1,inputRegisters_424__0})) ;
    Reg_16 loop1_424_x (.D ({inputRegisters_424__15,inputRegisters_424__14,
           inputRegisters_424__13,inputRegisters_424__12,inputRegisters_424__11,
           inputRegisters_424__10,inputRegisters_424__9,inputRegisters_424__8,
           inputRegisters_424__7,inputRegisters_424__6,inputRegisters_424__5,
           inputRegisters_424__4,inputRegisters_424__3,inputRegisters_424__2,
           inputRegisters_424__1,inputRegisters_424__0}), .en (
           enableRegister_424), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_424__15,registerOutputs_424__14,
           registerOutputs_424__13,registerOutputs_424__12,
           registerOutputs_424__11,registerOutputs_424__10,
           registerOutputs_424__9,registerOutputs_424__8,registerOutputs_424__7,
           registerOutputs_424__6,registerOutputs_424__5,registerOutputs_424__4,
           registerOutputs_424__3,registerOutputs_424__2,registerOutputs_424__1,
           registerOutputs_424__0})) ;
    Mux2_16 loop1_425_y (.A ({nx36005,nx36147,nx36289,nx36431,nx36573,nx36715,
            nx36857,nx36999,nx37141,nx37283,nx37425,nx37567,nx37709,nx37851,
            nx37993,nx38135}), .B ({nx33761,nx33899,nx34039,nx34177,nx34315,
            nx34453,nx34591,nx34731,nx34873,nx35015,nx35157,nx35299,nx35441,
            nx35583,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35725), .C ({inputRegisters_425__15,inputRegisters_425__14,
            inputRegisters_425__13,inputRegisters_425__12,inputRegisters_425__11
            ,inputRegisters_425__10,inputRegisters_425__9,inputRegisters_425__8,
            inputRegisters_425__7,inputRegisters_425__6,inputRegisters_425__5,
            inputRegisters_425__4,inputRegisters_425__3,inputRegisters_425__2,
            inputRegisters_425__1,inputRegisters_425__0})) ;
    Reg_16 loop1_425_x (.D ({inputRegisters_425__15,inputRegisters_425__14,
           inputRegisters_425__13,inputRegisters_425__12,inputRegisters_425__11,
           inputRegisters_425__10,inputRegisters_425__9,inputRegisters_425__8,
           inputRegisters_425__7,inputRegisters_425__6,inputRegisters_425__5,
           inputRegisters_425__4,inputRegisters_425__3,inputRegisters_425__2,
           inputRegisters_425__1,inputRegisters_425__0}), .en (
           enableRegister_425), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_425__15,registerOutputs_425__14,
           registerOutputs_425__13,registerOutputs_425__12,
           registerOutputs_425__11,registerOutputs_425__10,
           registerOutputs_425__9,registerOutputs_425__8,registerOutputs_425__7,
           registerOutputs_425__6,registerOutputs_425__5,registerOutputs_425__4,
           registerOutputs_425__3,registerOutputs_425__2,registerOutputs_425__1,
           registerOutputs_425__0})) ;
    Mux2_16 loop1_426_y (.A ({nx36005,nx36147,nx36289,nx36431,nx36573,nx36715,
            nx36857,nx36999,nx37141,nx37283,nx37425,nx37567,nx37709,nx37851,
            nx37993,nx38135}), .B ({nx33761,nx33901,nx34039,nx34177,nx34315,
            nx34453,nx34591,nx34731,nx34873,nx35015,nx35157,nx35299,nx35441,
            nx35583,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35725), .C ({inputRegisters_426__15,inputRegisters_426__14,
            inputRegisters_426__13,inputRegisters_426__12,inputRegisters_426__11
            ,inputRegisters_426__10,inputRegisters_426__9,inputRegisters_426__8,
            inputRegisters_426__7,inputRegisters_426__6,inputRegisters_426__5,
            inputRegisters_426__4,inputRegisters_426__3,inputRegisters_426__2,
            inputRegisters_426__1,inputRegisters_426__0})) ;
    Reg_16 loop1_426_x (.D ({inputRegisters_426__15,inputRegisters_426__14,
           inputRegisters_426__13,inputRegisters_426__12,inputRegisters_426__11,
           inputRegisters_426__10,inputRegisters_426__9,inputRegisters_426__8,
           inputRegisters_426__7,inputRegisters_426__6,inputRegisters_426__5,
           inputRegisters_426__4,inputRegisters_426__3,inputRegisters_426__2,
           inputRegisters_426__1,inputRegisters_426__0}), .en (
           enableRegister_426), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_426__15,registerOutputs_426__14,
           registerOutputs_426__13,registerOutputs_426__12,
           registerOutputs_426__11,registerOutputs_426__10,
           registerOutputs_426__9,registerOutputs_426__8,registerOutputs_426__7,
           registerOutputs_426__6,registerOutputs_426__5,registerOutputs_426__4,
           registerOutputs_426__3,registerOutputs_426__2,registerOutputs_426__1,
           registerOutputs_426__0})) ;
    Mux2_16 loop1_427_y (.A ({nx36007,nx36149,nx36291,nx36433,nx36575,nx36717,
            nx36859,nx37001,nx37143,nx37285,nx37427,nx37569,nx37711,nx37853,
            nx37995,nx38137}), .B ({nx33763,nx33901,nx34039,nx34177,nx34315,
            nx34453,nx34591,nx34733,nx34875,nx35017,nx35159,nx35301,nx35443,
            nx35585,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35727), .C ({inputRegisters_427__15,inputRegisters_427__14,
            inputRegisters_427__13,inputRegisters_427__12,inputRegisters_427__11
            ,inputRegisters_427__10,inputRegisters_427__9,inputRegisters_427__8,
            inputRegisters_427__7,inputRegisters_427__6,inputRegisters_427__5,
            inputRegisters_427__4,inputRegisters_427__3,inputRegisters_427__2,
            inputRegisters_427__1,inputRegisters_427__0})) ;
    Reg_16 loop1_427_x (.D ({inputRegisters_427__15,inputRegisters_427__14,
           inputRegisters_427__13,inputRegisters_427__12,inputRegisters_427__11,
           inputRegisters_427__10,inputRegisters_427__9,inputRegisters_427__8,
           inputRegisters_427__7,inputRegisters_427__6,inputRegisters_427__5,
           inputRegisters_427__4,inputRegisters_427__3,inputRegisters_427__2,
           inputRegisters_427__1,inputRegisters_427__0}), .en (
           enableRegister_427), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_427__15,registerOutputs_427__14,
           registerOutputs_427__13,registerOutputs_427__12,
           registerOutputs_427__11,registerOutputs_427__10,
           registerOutputs_427__9,registerOutputs_427__8,registerOutputs_427__7,
           registerOutputs_427__6,registerOutputs_427__5,registerOutputs_427__4,
           registerOutputs_427__3,registerOutputs_427__2,registerOutputs_427__1,
           registerOutputs_427__0})) ;
    Mux2_16 loop1_428_y (.A ({nx36007,nx36149,nx36291,nx36433,nx36575,nx36717,
            nx36859,nx37001,nx37143,nx37285,nx37427,nx37569,nx37711,nx37853,
            nx37995,nx38137}), .B ({nx33763,nx33901,nx34039,nx34177,nx34315,
            nx34453,nx34593,nx34733,nx34875,nx35017,nx35159,nx35301,nx35443,
            nx35585,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35727), .C ({inputRegisters_428__15,inputRegisters_428__14,
            inputRegisters_428__13,inputRegisters_428__12,inputRegisters_428__11
            ,inputRegisters_428__10,inputRegisters_428__9,inputRegisters_428__8,
            inputRegisters_428__7,inputRegisters_428__6,inputRegisters_428__5,
            inputRegisters_428__4,inputRegisters_428__3,inputRegisters_428__2,
            inputRegisters_428__1,inputRegisters_428__0})) ;
    Reg_16 loop1_428_x (.D ({inputRegisters_428__15,inputRegisters_428__14,
           inputRegisters_428__13,inputRegisters_428__12,inputRegisters_428__11,
           inputRegisters_428__10,inputRegisters_428__9,inputRegisters_428__8,
           inputRegisters_428__7,inputRegisters_428__6,inputRegisters_428__5,
           inputRegisters_428__4,inputRegisters_428__3,inputRegisters_428__2,
           inputRegisters_428__1,inputRegisters_428__0}), .en (
           enableRegister_428), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_428__15,registerOutputs_428__14,
           registerOutputs_428__13,registerOutputs_428__12,
           registerOutputs_428__11,registerOutputs_428__10,
           registerOutputs_428__9,registerOutputs_428__8,registerOutputs_428__7,
           registerOutputs_428__6,registerOutputs_428__5,registerOutputs_428__4,
           registerOutputs_428__3,registerOutputs_428__2,registerOutputs_428__1,
           registerOutputs_428__0})) ;
    Mux2_16 loop1_429_y (.A ({nx36007,nx36149,nx36291,nx36433,nx36575,nx36717,
            nx36859,nx37001,nx37143,nx37285,nx37427,nx37569,nx37711,nx37853,
            nx37995,nx38137}), .B ({nx33763,nx33901,nx34039,nx34177,nx34315,
            nx34455,nx34593,nx34733,nx34875,nx35017,nx35159,nx35301,nx35443,
            nx35585,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35727), .C ({inputRegisters_429__15,inputRegisters_429__14,
            inputRegisters_429__13,inputRegisters_429__12,inputRegisters_429__11
            ,inputRegisters_429__10,inputRegisters_429__9,inputRegisters_429__8,
            inputRegisters_429__7,inputRegisters_429__6,inputRegisters_429__5,
            inputRegisters_429__4,inputRegisters_429__3,inputRegisters_429__2,
            inputRegisters_429__1,inputRegisters_429__0})) ;
    Reg_16 loop1_429_x (.D ({inputRegisters_429__15,inputRegisters_429__14,
           inputRegisters_429__13,inputRegisters_429__12,inputRegisters_429__11,
           inputRegisters_429__10,inputRegisters_429__9,inputRegisters_429__8,
           inputRegisters_429__7,inputRegisters_429__6,inputRegisters_429__5,
           inputRegisters_429__4,inputRegisters_429__3,inputRegisters_429__2,
           inputRegisters_429__1,inputRegisters_429__0}), .en (
           enableRegister_429), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_429__15,registerOutputs_429__14,
           registerOutputs_429__13,registerOutputs_429__12,
           registerOutputs_429__11,registerOutputs_429__10,
           registerOutputs_429__9,registerOutputs_429__8,registerOutputs_429__7,
           registerOutputs_429__6,registerOutputs_429__5,registerOutputs_429__4,
           registerOutputs_429__3,registerOutputs_429__2,registerOutputs_429__1,
           registerOutputs_429__0})) ;
    Mux2_16 loop1_430_y (.A ({nx36007,nx36149,nx36291,nx36433,nx36575,nx36717,
            nx36859,nx37001,nx37143,nx37285,nx37427,nx37569,nx37711,nx37853,
            nx37995,nx38137}), .B ({nx33763,nx33901,nx34039,nx34177,nx34317,
            nx34455,nx34593,nx34733,nx34875,nx35017,nx35159,nx35301,nx35443,
            nx35585,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35727), .C ({inputRegisters_430__15,inputRegisters_430__14,
            inputRegisters_430__13,inputRegisters_430__12,inputRegisters_430__11
            ,inputRegisters_430__10,inputRegisters_430__9,inputRegisters_430__8,
            inputRegisters_430__7,inputRegisters_430__6,inputRegisters_430__5,
            inputRegisters_430__4,inputRegisters_430__3,inputRegisters_430__2,
            inputRegisters_430__1,inputRegisters_430__0})) ;
    Reg_16 loop1_430_x (.D ({inputRegisters_430__15,inputRegisters_430__14,
           inputRegisters_430__13,inputRegisters_430__12,inputRegisters_430__11,
           inputRegisters_430__10,inputRegisters_430__9,inputRegisters_430__8,
           inputRegisters_430__7,inputRegisters_430__6,inputRegisters_430__5,
           inputRegisters_430__4,inputRegisters_430__3,inputRegisters_430__2,
           inputRegisters_430__1,inputRegisters_430__0}), .en (
           enableRegister_430), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_430__15,registerOutputs_430__14,
           registerOutputs_430__13,registerOutputs_430__12,
           registerOutputs_430__11,registerOutputs_430__10,
           registerOutputs_430__9,registerOutputs_430__8,registerOutputs_430__7,
           registerOutputs_430__6,registerOutputs_430__5,registerOutputs_430__4,
           registerOutputs_430__3,registerOutputs_430__2,registerOutputs_430__1,
           registerOutputs_430__0})) ;
    Mux2_16 loop1_431_y (.A ({nx36007,nx36149,nx36291,nx36433,nx36575,nx36717,
            nx36859,nx37001,nx37143,nx37285,nx37427,nx37569,nx37711,nx37853,
            nx37995,nx38137}), .B ({nx33763,nx33901,nx34039,nx34179,nx34317,
            nx34455,nx34593,nx34733,nx34875,nx35017,nx35159,nx35301,nx35443,
            nx35585,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35727), .C ({inputRegisters_431__15,inputRegisters_431__14,
            inputRegisters_431__13,inputRegisters_431__12,inputRegisters_431__11
            ,inputRegisters_431__10,inputRegisters_431__9,inputRegisters_431__8,
            inputRegisters_431__7,inputRegisters_431__6,inputRegisters_431__5,
            inputRegisters_431__4,inputRegisters_431__3,inputRegisters_431__2,
            inputRegisters_431__1,inputRegisters_431__0})) ;
    Reg_16 loop1_431_x (.D ({inputRegisters_431__15,inputRegisters_431__14,
           inputRegisters_431__13,inputRegisters_431__12,inputRegisters_431__11,
           inputRegisters_431__10,inputRegisters_431__9,inputRegisters_431__8,
           inputRegisters_431__7,inputRegisters_431__6,inputRegisters_431__5,
           inputRegisters_431__4,inputRegisters_431__3,inputRegisters_431__2,
           inputRegisters_431__1,inputRegisters_431__0}), .en (
           enableRegister_431), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_431__15,registerOutputs_431__14,
           registerOutputs_431__13,registerOutputs_431__12,
           registerOutputs_431__11,registerOutputs_431__10,
           registerOutputs_431__9,registerOutputs_431__8,registerOutputs_431__7,
           registerOutputs_431__6,registerOutputs_431__5,registerOutputs_431__4,
           registerOutputs_431__3,registerOutputs_431__2,registerOutputs_431__1,
           registerOutputs_431__0})) ;
    Mux2_16 loop1_432_y (.A ({nx36007,nx36149,nx36291,nx36433,nx36575,nx36717,
            nx36859,nx37001,nx37143,nx37285,nx37427,nx37569,nx37711,nx37853,
            nx37995,nx38137}), .B ({nx33763,nx33901,nx34041,nx34179,nx34317,
            nx34455,nx34593,nx34733,nx34875,nx35017,nx35159,nx35301,nx35443,
            nx35585,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35727), .C ({inputRegisters_432__15,inputRegisters_432__14,
            inputRegisters_432__13,inputRegisters_432__12,inputRegisters_432__11
            ,inputRegisters_432__10,inputRegisters_432__9,inputRegisters_432__8,
            inputRegisters_432__7,inputRegisters_432__6,inputRegisters_432__5,
            inputRegisters_432__4,inputRegisters_432__3,inputRegisters_432__2,
            inputRegisters_432__1,inputRegisters_432__0})) ;
    Reg_16 loop1_432_x (.D ({inputRegisters_432__15,inputRegisters_432__14,
           inputRegisters_432__13,inputRegisters_432__12,inputRegisters_432__11,
           inputRegisters_432__10,inputRegisters_432__9,inputRegisters_432__8,
           inputRegisters_432__7,inputRegisters_432__6,inputRegisters_432__5,
           inputRegisters_432__4,inputRegisters_432__3,inputRegisters_432__2,
           inputRegisters_432__1,inputRegisters_432__0}), .en (
           enableRegister_432), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_432__15,registerOutputs_432__14,
           registerOutputs_432__13,registerOutputs_432__12,
           registerOutputs_432__11,registerOutputs_432__10,
           registerOutputs_432__9,registerOutputs_432__8,registerOutputs_432__7,
           registerOutputs_432__6,registerOutputs_432__5,registerOutputs_432__4,
           registerOutputs_432__3,registerOutputs_432__2,registerOutputs_432__1,
           registerOutputs_432__0})) ;
    Mux2_16 loop1_433_y (.A ({nx36007,nx36149,nx36291,nx36433,nx36575,nx36717,
            nx36859,nx37001,nx37143,nx37285,nx37427,nx37569,nx37711,nx37853,
            nx37995,nx38137}), .B ({nx33763,nx33903,nx34041,nx34179,nx34317,
            nx34455,nx34593,nx34733,nx34875,nx35017,nx35159,nx35301,nx35443,
            nx35585,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35727), .C ({inputRegisters_433__15,inputRegisters_433__14,
            inputRegisters_433__13,inputRegisters_433__12,inputRegisters_433__11
            ,inputRegisters_433__10,inputRegisters_433__9,inputRegisters_433__8,
            inputRegisters_433__7,inputRegisters_433__6,inputRegisters_433__5,
            inputRegisters_433__4,inputRegisters_433__3,inputRegisters_433__2,
            inputRegisters_433__1,inputRegisters_433__0})) ;
    Reg_16 loop1_433_x (.D ({inputRegisters_433__15,inputRegisters_433__14,
           inputRegisters_433__13,inputRegisters_433__12,inputRegisters_433__11,
           inputRegisters_433__10,inputRegisters_433__9,inputRegisters_433__8,
           inputRegisters_433__7,inputRegisters_433__6,inputRegisters_433__5,
           inputRegisters_433__4,inputRegisters_433__3,inputRegisters_433__2,
           inputRegisters_433__1,inputRegisters_433__0}), .en (
           enableRegister_433), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_433__15,registerOutputs_433__14,
           registerOutputs_433__13,registerOutputs_433__12,
           registerOutputs_433__11,registerOutputs_433__10,
           registerOutputs_433__9,registerOutputs_433__8,registerOutputs_433__7,
           registerOutputs_433__6,registerOutputs_433__5,registerOutputs_433__4,
           registerOutputs_433__3,registerOutputs_433__2,registerOutputs_433__1,
           registerOutputs_433__0})) ;
    Mux2_16 loop1_434_y (.A ({nx36009,nx36151,nx36293,nx36435,nx36577,nx36719,
            nx36861,nx37003,nx37145,nx37287,nx37429,nx37571,nx37713,nx37855,
            nx37997,nx38139}), .B ({nx33765,nx33903,nx34041,nx34179,nx34317,
            nx34455,nx34593,nx34735,nx34877,nx35019,nx35161,nx35303,nx35445,
            nx35587,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35729), .C ({inputRegisters_434__15,inputRegisters_434__14,
            inputRegisters_434__13,inputRegisters_434__12,inputRegisters_434__11
            ,inputRegisters_434__10,inputRegisters_434__9,inputRegisters_434__8,
            inputRegisters_434__7,inputRegisters_434__6,inputRegisters_434__5,
            inputRegisters_434__4,inputRegisters_434__3,inputRegisters_434__2,
            inputRegisters_434__1,inputRegisters_434__0})) ;
    Reg_16 loop1_434_x (.D ({inputRegisters_434__15,inputRegisters_434__14,
           inputRegisters_434__13,inputRegisters_434__12,inputRegisters_434__11,
           inputRegisters_434__10,inputRegisters_434__9,inputRegisters_434__8,
           inputRegisters_434__7,inputRegisters_434__6,inputRegisters_434__5,
           inputRegisters_434__4,inputRegisters_434__3,inputRegisters_434__2,
           inputRegisters_434__1,inputRegisters_434__0}), .en (
           enableRegister_434), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_434__15,registerOutputs_434__14,
           registerOutputs_434__13,registerOutputs_434__12,
           registerOutputs_434__11,registerOutputs_434__10,
           registerOutputs_434__9,registerOutputs_434__8,registerOutputs_434__7,
           registerOutputs_434__6,registerOutputs_434__5,registerOutputs_434__4,
           registerOutputs_434__3,registerOutputs_434__2,registerOutputs_434__1,
           registerOutputs_434__0})) ;
    Mux2_16 loop1_435_y (.A ({nx36009,nx36151,nx36293,nx36435,nx36577,nx36719,
            nx36861,nx37003,nx37145,nx37287,nx37429,nx37571,nx37713,nx37855,
            nx37997,nx38139}), .B ({nx33765,nx33903,nx34041,nx34179,nx34317,
            nx34455,nx34595,nx34735,nx34877,nx35019,nx35161,nx35303,nx35445,
            nx35587,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35729), .C ({inputRegisters_435__15,inputRegisters_435__14,
            inputRegisters_435__13,inputRegisters_435__12,inputRegisters_435__11
            ,inputRegisters_435__10,inputRegisters_435__9,inputRegisters_435__8,
            inputRegisters_435__7,inputRegisters_435__6,inputRegisters_435__5,
            inputRegisters_435__4,inputRegisters_435__3,inputRegisters_435__2,
            inputRegisters_435__1,inputRegisters_435__0})) ;
    Reg_16 loop1_435_x (.D ({inputRegisters_435__15,inputRegisters_435__14,
           inputRegisters_435__13,inputRegisters_435__12,inputRegisters_435__11,
           inputRegisters_435__10,inputRegisters_435__9,inputRegisters_435__8,
           inputRegisters_435__7,inputRegisters_435__6,inputRegisters_435__5,
           inputRegisters_435__4,inputRegisters_435__3,inputRegisters_435__2,
           inputRegisters_435__1,inputRegisters_435__0}), .en (
           enableRegister_435), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_435__15,registerOutputs_435__14,
           registerOutputs_435__13,registerOutputs_435__12,
           registerOutputs_435__11,registerOutputs_435__10,
           registerOutputs_435__9,registerOutputs_435__8,registerOutputs_435__7,
           registerOutputs_435__6,registerOutputs_435__5,registerOutputs_435__4,
           registerOutputs_435__3,registerOutputs_435__2,registerOutputs_435__1,
           registerOutputs_435__0})) ;
    Mux2_16 loop1_436_y (.A ({nx36009,nx36151,nx36293,nx36435,nx36577,nx36719,
            nx36861,nx37003,nx37145,nx37287,nx37429,nx37571,nx37713,nx37855,
            nx37997,nx38139}), .B ({nx33765,nx33903,nx34041,nx34179,nx34317,
            nx34457,nx34595,nx34735,nx34877,nx35019,nx35161,nx35303,nx35445,
            nx35587,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35729), .C ({inputRegisters_436__15,inputRegisters_436__14,
            inputRegisters_436__13,inputRegisters_436__12,inputRegisters_436__11
            ,inputRegisters_436__10,inputRegisters_436__9,inputRegisters_436__8,
            inputRegisters_436__7,inputRegisters_436__6,inputRegisters_436__5,
            inputRegisters_436__4,inputRegisters_436__3,inputRegisters_436__2,
            inputRegisters_436__1,inputRegisters_436__0})) ;
    Reg_16 loop1_436_x (.D ({inputRegisters_436__15,inputRegisters_436__14,
           inputRegisters_436__13,inputRegisters_436__12,inputRegisters_436__11,
           inputRegisters_436__10,inputRegisters_436__9,inputRegisters_436__8,
           inputRegisters_436__7,inputRegisters_436__6,inputRegisters_436__5,
           inputRegisters_436__4,inputRegisters_436__3,inputRegisters_436__2,
           inputRegisters_436__1,inputRegisters_436__0}), .en (
           enableRegister_436), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_436__15,registerOutputs_436__14,
           registerOutputs_436__13,registerOutputs_436__12,
           registerOutputs_436__11,registerOutputs_436__10,
           registerOutputs_436__9,registerOutputs_436__8,registerOutputs_436__7,
           registerOutputs_436__6,registerOutputs_436__5,registerOutputs_436__4,
           registerOutputs_436__3,registerOutputs_436__2,registerOutputs_436__1,
           registerOutputs_436__0})) ;
    Mux2_16 loop1_437_y (.A ({nx36009,nx36151,nx36293,nx36435,nx36577,nx36719,
            nx36861,nx37003,nx37145,nx37287,nx37429,nx37571,nx37713,nx37855,
            nx37997,nx38139}), .B ({nx33765,nx33903,nx34041,nx34179,nx34319,
            nx34457,nx34595,nx34735,nx34877,nx35019,nx35161,nx35303,nx35445,
            nx35587,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35729), .C ({inputRegisters_437__15,inputRegisters_437__14,
            inputRegisters_437__13,inputRegisters_437__12,inputRegisters_437__11
            ,inputRegisters_437__10,inputRegisters_437__9,inputRegisters_437__8,
            inputRegisters_437__7,inputRegisters_437__6,inputRegisters_437__5,
            inputRegisters_437__4,inputRegisters_437__3,inputRegisters_437__2,
            inputRegisters_437__1,inputRegisters_437__0})) ;
    Reg_16 loop1_437_x (.D ({inputRegisters_437__15,inputRegisters_437__14,
           inputRegisters_437__13,inputRegisters_437__12,inputRegisters_437__11,
           inputRegisters_437__10,inputRegisters_437__9,inputRegisters_437__8,
           inputRegisters_437__7,inputRegisters_437__6,inputRegisters_437__5,
           inputRegisters_437__4,inputRegisters_437__3,inputRegisters_437__2,
           inputRegisters_437__1,inputRegisters_437__0}), .en (
           enableRegister_437), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_437__15,registerOutputs_437__14,
           registerOutputs_437__13,registerOutputs_437__12,
           registerOutputs_437__11,registerOutputs_437__10,
           registerOutputs_437__9,registerOutputs_437__8,registerOutputs_437__7,
           registerOutputs_437__6,registerOutputs_437__5,registerOutputs_437__4,
           registerOutputs_437__3,registerOutputs_437__2,registerOutputs_437__1,
           registerOutputs_437__0})) ;
    Mux2_16 loop1_438_y (.A ({nx36009,nx36151,nx36293,nx36435,nx36577,nx36719,
            nx36861,nx37003,nx37145,nx37287,nx37429,nx37571,nx37713,nx37855,
            nx37997,nx38139}), .B ({nx33765,nx33903,nx34041,nx34181,nx34319,
            nx34457,nx34595,nx34735,nx34877,nx35019,nx35161,nx35303,nx35445,
            nx35587,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35729), .C ({inputRegisters_438__15,inputRegisters_438__14,
            inputRegisters_438__13,inputRegisters_438__12,inputRegisters_438__11
            ,inputRegisters_438__10,inputRegisters_438__9,inputRegisters_438__8,
            inputRegisters_438__7,inputRegisters_438__6,inputRegisters_438__5,
            inputRegisters_438__4,inputRegisters_438__3,inputRegisters_438__2,
            inputRegisters_438__1,inputRegisters_438__0})) ;
    Reg_16 loop1_438_x (.D ({inputRegisters_438__15,inputRegisters_438__14,
           inputRegisters_438__13,inputRegisters_438__12,inputRegisters_438__11,
           inputRegisters_438__10,inputRegisters_438__9,inputRegisters_438__8,
           inputRegisters_438__7,inputRegisters_438__6,inputRegisters_438__5,
           inputRegisters_438__4,inputRegisters_438__3,inputRegisters_438__2,
           inputRegisters_438__1,inputRegisters_438__0}), .en (
           enableRegister_438), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_438__15,registerOutputs_438__14,
           registerOutputs_438__13,registerOutputs_438__12,
           registerOutputs_438__11,registerOutputs_438__10,
           registerOutputs_438__9,registerOutputs_438__8,registerOutputs_438__7,
           registerOutputs_438__6,registerOutputs_438__5,registerOutputs_438__4,
           registerOutputs_438__3,registerOutputs_438__2,registerOutputs_438__1,
           registerOutputs_438__0})) ;
    Mux2_16 loop1_439_y (.A ({nx36009,nx36151,nx36293,nx36435,nx36577,nx36719,
            nx36861,nx37003,nx37145,nx37287,nx37429,nx37571,nx37713,nx37855,
            nx37997,nx38139}), .B ({nx33765,nx33903,nx34043,nx34181,nx34319,
            nx34457,nx34595,nx34735,nx34877,nx35019,nx35161,nx35303,nx35445,
            nx35587,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35729), .C ({inputRegisters_439__15,inputRegisters_439__14,
            inputRegisters_439__13,inputRegisters_439__12,inputRegisters_439__11
            ,inputRegisters_439__10,inputRegisters_439__9,inputRegisters_439__8,
            inputRegisters_439__7,inputRegisters_439__6,inputRegisters_439__5,
            inputRegisters_439__4,inputRegisters_439__3,inputRegisters_439__2,
            inputRegisters_439__1,inputRegisters_439__0})) ;
    Reg_16 loop1_439_x (.D ({inputRegisters_439__15,inputRegisters_439__14,
           inputRegisters_439__13,inputRegisters_439__12,inputRegisters_439__11,
           inputRegisters_439__10,inputRegisters_439__9,inputRegisters_439__8,
           inputRegisters_439__7,inputRegisters_439__6,inputRegisters_439__5,
           inputRegisters_439__4,inputRegisters_439__3,inputRegisters_439__2,
           inputRegisters_439__1,inputRegisters_439__0}), .en (
           enableRegister_439), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_439__15,registerOutputs_439__14,
           registerOutputs_439__13,registerOutputs_439__12,
           registerOutputs_439__11,registerOutputs_439__10,
           registerOutputs_439__9,registerOutputs_439__8,registerOutputs_439__7,
           registerOutputs_439__6,registerOutputs_439__5,registerOutputs_439__4,
           registerOutputs_439__3,registerOutputs_439__2,registerOutputs_439__1,
           registerOutputs_439__0})) ;
    Mux2_16 loop1_440_y (.A ({nx36009,nx36151,nx36293,nx36435,nx36577,nx36719,
            nx36861,nx37003,nx37145,nx37287,nx37429,nx37571,nx37713,nx37855,
            nx37997,nx38139}), .B ({nx33765,nx33905,nx34043,nx34181,nx34319,
            nx34457,nx34595,nx34735,nx34877,nx35019,nx35161,nx35303,nx35445,
            nx35587,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35729), .C ({inputRegisters_440__15,inputRegisters_440__14,
            inputRegisters_440__13,inputRegisters_440__12,inputRegisters_440__11
            ,inputRegisters_440__10,inputRegisters_440__9,inputRegisters_440__8,
            inputRegisters_440__7,inputRegisters_440__6,inputRegisters_440__5,
            inputRegisters_440__4,inputRegisters_440__3,inputRegisters_440__2,
            inputRegisters_440__1,inputRegisters_440__0})) ;
    Reg_16 loop1_440_x (.D ({inputRegisters_440__15,inputRegisters_440__14,
           inputRegisters_440__13,inputRegisters_440__12,inputRegisters_440__11,
           inputRegisters_440__10,inputRegisters_440__9,inputRegisters_440__8,
           inputRegisters_440__7,inputRegisters_440__6,inputRegisters_440__5,
           inputRegisters_440__4,inputRegisters_440__3,inputRegisters_440__2,
           inputRegisters_440__1,inputRegisters_440__0}), .en (
           enableRegister_440), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_440__15,registerOutputs_440__14,
           registerOutputs_440__13,registerOutputs_440__12,
           registerOutputs_440__11,registerOutputs_440__10,
           registerOutputs_440__9,registerOutputs_440__8,registerOutputs_440__7,
           registerOutputs_440__6,registerOutputs_440__5,registerOutputs_440__4,
           registerOutputs_440__3,registerOutputs_440__2,registerOutputs_440__1,
           registerOutputs_440__0})) ;
    Mux2_16 loop1_441_y (.A ({nx36011,nx36153,nx36295,nx36437,nx36579,nx36721,
            nx36863,nx37005,nx37147,nx37289,nx37431,nx37573,nx37715,nx37857,
            nx37999,nx38141}), .B ({nx33767,nx33905,nx34043,nx34181,nx34319,
            nx34457,nx34595,nx34737,nx34879,nx35021,nx35163,nx35305,nx35447,
            nx35589,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35731), .C ({inputRegisters_441__15,inputRegisters_441__14,
            inputRegisters_441__13,inputRegisters_441__12,inputRegisters_441__11
            ,inputRegisters_441__10,inputRegisters_441__9,inputRegisters_441__8,
            inputRegisters_441__7,inputRegisters_441__6,inputRegisters_441__5,
            inputRegisters_441__4,inputRegisters_441__3,inputRegisters_441__2,
            inputRegisters_441__1,inputRegisters_441__0})) ;
    Reg_16 loop1_441_x (.D ({inputRegisters_441__15,inputRegisters_441__14,
           inputRegisters_441__13,inputRegisters_441__12,inputRegisters_441__11,
           inputRegisters_441__10,inputRegisters_441__9,inputRegisters_441__8,
           inputRegisters_441__7,inputRegisters_441__6,inputRegisters_441__5,
           inputRegisters_441__4,inputRegisters_441__3,inputRegisters_441__2,
           inputRegisters_441__1,inputRegisters_441__0}), .en (
           enableRegister_441), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_441__15,registerOutputs_441__14,
           registerOutputs_441__13,registerOutputs_441__12,
           registerOutputs_441__11,registerOutputs_441__10,
           registerOutputs_441__9,registerOutputs_441__8,registerOutputs_441__7,
           registerOutputs_441__6,registerOutputs_441__5,registerOutputs_441__4,
           registerOutputs_441__3,registerOutputs_441__2,registerOutputs_441__1,
           registerOutputs_441__0})) ;
    Mux2_16 loop1_442_y (.A ({nx36011,nx36153,nx36295,nx36437,nx36579,nx36721,
            nx36863,nx37005,nx37147,nx37289,nx37431,nx37573,nx37715,nx37857,
            nx37999,nx38141}), .B ({nx33767,nx33905,nx34043,nx34181,nx34319,
            nx34457,nx34597,nx34737,nx34879,nx35021,nx35163,nx35305,nx35447,
            nx35589,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35731), .C ({inputRegisters_442__15,inputRegisters_442__14,
            inputRegisters_442__13,inputRegisters_442__12,inputRegisters_442__11
            ,inputRegisters_442__10,inputRegisters_442__9,inputRegisters_442__8,
            inputRegisters_442__7,inputRegisters_442__6,inputRegisters_442__5,
            inputRegisters_442__4,inputRegisters_442__3,inputRegisters_442__2,
            inputRegisters_442__1,inputRegisters_442__0})) ;
    Reg_16 loop1_442_x (.D ({inputRegisters_442__15,inputRegisters_442__14,
           inputRegisters_442__13,inputRegisters_442__12,inputRegisters_442__11,
           inputRegisters_442__10,inputRegisters_442__9,inputRegisters_442__8,
           inputRegisters_442__7,inputRegisters_442__6,inputRegisters_442__5,
           inputRegisters_442__4,inputRegisters_442__3,inputRegisters_442__2,
           inputRegisters_442__1,inputRegisters_442__0}), .en (
           enableRegister_442), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_442__15,registerOutputs_442__14,
           registerOutputs_442__13,registerOutputs_442__12,
           registerOutputs_442__11,registerOutputs_442__10,
           registerOutputs_442__9,registerOutputs_442__8,registerOutputs_442__7,
           registerOutputs_442__6,registerOutputs_442__5,registerOutputs_442__4,
           registerOutputs_442__3,registerOutputs_442__2,registerOutputs_442__1,
           registerOutputs_442__0})) ;
    Mux2_16 loop1_443_y (.A ({nx36011,nx36153,nx36295,nx36437,nx36579,nx36721,
            nx36863,nx37005,nx37147,nx37289,nx37431,nx37573,nx37715,nx37857,
            nx37999,nx38141}), .B ({nx33767,nx33905,nx34043,nx34181,nx34319,
            nx34459,nx34597,nx34737,nx34879,nx35021,nx35163,nx35305,nx35447,
            nx35589,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35731), .C ({inputRegisters_443__15,inputRegisters_443__14,
            inputRegisters_443__13,inputRegisters_443__12,inputRegisters_443__11
            ,inputRegisters_443__10,inputRegisters_443__9,inputRegisters_443__8,
            inputRegisters_443__7,inputRegisters_443__6,inputRegisters_443__5,
            inputRegisters_443__4,inputRegisters_443__3,inputRegisters_443__2,
            inputRegisters_443__1,inputRegisters_443__0})) ;
    Reg_16 loop1_443_x (.D ({inputRegisters_443__15,inputRegisters_443__14,
           inputRegisters_443__13,inputRegisters_443__12,inputRegisters_443__11,
           inputRegisters_443__10,inputRegisters_443__9,inputRegisters_443__8,
           inputRegisters_443__7,inputRegisters_443__6,inputRegisters_443__5,
           inputRegisters_443__4,inputRegisters_443__3,inputRegisters_443__2,
           inputRegisters_443__1,inputRegisters_443__0}), .en (
           enableRegister_443), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_443__15,registerOutputs_443__14,
           registerOutputs_443__13,registerOutputs_443__12,
           registerOutputs_443__11,registerOutputs_443__10,
           registerOutputs_443__9,registerOutputs_443__8,registerOutputs_443__7,
           registerOutputs_443__6,registerOutputs_443__5,registerOutputs_443__4,
           registerOutputs_443__3,registerOutputs_443__2,registerOutputs_443__1,
           registerOutputs_443__0})) ;
    Mux2_16 loop1_444_y (.A ({nx36011,nx36153,nx36295,nx36437,nx36579,nx36721,
            nx36863,nx37005,nx37147,nx37289,nx37431,nx37573,nx37715,nx37857,
            nx37999,nx38141}), .B ({nx33767,nx33905,nx34043,nx34181,nx34321,
            nx34459,nx34597,nx34737,nx34879,nx35021,nx35163,nx35305,nx35447,
            nx35589,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35731), .C ({inputRegisters_444__15,inputRegisters_444__14,
            inputRegisters_444__13,inputRegisters_444__12,inputRegisters_444__11
            ,inputRegisters_444__10,inputRegisters_444__9,inputRegisters_444__8,
            inputRegisters_444__7,inputRegisters_444__6,inputRegisters_444__5,
            inputRegisters_444__4,inputRegisters_444__3,inputRegisters_444__2,
            inputRegisters_444__1,inputRegisters_444__0})) ;
    Reg_16 loop1_444_x (.D ({inputRegisters_444__15,inputRegisters_444__14,
           inputRegisters_444__13,inputRegisters_444__12,inputRegisters_444__11,
           inputRegisters_444__10,inputRegisters_444__9,inputRegisters_444__8,
           inputRegisters_444__7,inputRegisters_444__6,inputRegisters_444__5,
           inputRegisters_444__4,inputRegisters_444__3,inputRegisters_444__2,
           inputRegisters_444__1,inputRegisters_444__0}), .en (
           enableRegister_444), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_444__15,registerOutputs_444__14,
           registerOutputs_444__13,registerOutputs_444__12,
           registerOutputs_444__11,registerOutputs_444__10,
           registerOutputs_444__9,registerOutputs_444__8,registerOutputs_444__7,
           registerOutputs_444__6,registerOutputs_444__5,registerOutputs_444__4,
           registerOutputs_444__3,registerOutputs_444__2,registerOutputs_444__1,
           registerOutputs_444__0})) ;
    Mux2_16 loop1_445_y (.A ({nx36011,nx36153,nx36295,nx36437,nx36579,nx36721,
            nx36863,nx37005,nx37147,nx37289,nx37431,nx37573,nx37715,nx37857,
            nx37999,nx38141}), .B ({nx33767,nx33905,nx34043,nx34183,nx34321,
            nx34459,nx34597,nx34737,nx34879,nx35021,nx35163,nx35305,nx35447,
            nx35589,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35731), .C ({inputRegisters_445__15,inputRegisters_445__14,
            inputRegisters_445__13,inputRegisters_445__12,inputRegisters_445__11
            ,inputRegisters_445__10,inputRegisters_445__9,inputRegisters_445__8,
            inputRegisters_445__7,inputRegisters_445__6,inputRegisters_445__5,
            inputRegisters_445__4,inputRegisters_445__3,inputRegisters_445__2,
            inputRegisters_445__1,inputRegisters_445__0})) ;
    Reg_16 loop1_445_x (.D ({inputRegisters_445__15,inputRegisters_445__14,
           inputRegisters_445__13,inputRegisters_445__12,inputRegisters_445__11,
           inputRegisters_445__10,inputRegisters_445__9,inputRegisters_445__8,
           inputRegisters_445__7,inputRegisters_445__6,inputRegisters_445__5,
           inputRegisters_445__4,inputRegisters_445__3,inputRegisters_445__2,
           inputRegisters_445__1,inputRegisters_445__0}), .en (
           enableRegister_445), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_445__15,registerOutputs_445__14,
           registerOutputs_445__13,registerOutputs_445__12,
           registerOutputs_445__11,registerOutputs_445__10,
           registerOutputs_445__9,registerOutputs_445__8,registerOutputs_445__7,
           registerOutputs_445__6,registerOutputs_445__5,registerOutputs_445__4,
           registerOutputs_445__3,registerOutputs_445__2,registerOutputs_445__1,
           registerOutputs_445__0})) ;
    Mux2_16 loop1_446_y (.A ({nx36011,nx36153,nx36295,nx36437,nx36579,nx36721,
            nx36863,nx37005,nx37147,nx37289,nx37431,nx37573,nx37715,nx37857,
            nx37999,nx38141}), .B ({nx33767,nx33905,nx34045,nx34183,nx34321,
            nx34459,nx34597,nx34737,nx34879,nx35021,nx35163,nx35305,nx35447,
            nx35589,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35731), .C ({inputRegisters_446__15,inputRegisters_446__14,
            inputRegisters_446__13,inputRegisters_446__12,inputRegisters_446__11
            ,inputRegisters_446__10,inputRegisters_446__9,inputRegisters_446__8,
            inputRegisters_446__7,inputRegisters_446__6,inputRegisters_446__5,
            inputRegisters_446__4,inputRegisters_446__3,inputRegisters_446__2,
            inputRegisters_446__1,inputRegisters_446__0})) ;
    Reg_16 loop1_446_x (.D ({inputRegisters_446__15,inputRegisters_446__14,
           inputRegisters_446__13,inputRegisters_446__12,inputRegisters_446__11,
           inputRegisters_446__10,inputRegisters_446__9,inputRegisters_446__8,
           inputRegisters_446__7,inputRegisters_446__6,inputRegisters_446__5,
           inputRegisters_446__4,inputRegisters_446__3,inputRegisters_446__2,
           inputRegisters_446__1,inputRegisters_446__0}), .en (
           enableRegister_446), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_446__15,registerOutputs_446__14,
           registerOutputs_446__13,registerOutputs_446__12,
           registerOutputs_446__11,registerOutputs_446__10,
           registerOutputs_446__9,registerOutputs_446__8,registerOutputs_446__7,
           registerOutputs_446__6,registerOutputs_446__5,registerOutputs_446__4,
           registerOutputs_446__3,registerOutputs_446__2,registerOutputs_446__1,
           registerOutputs_446__0})) ;
    Mux2_16 loop1_447_y (.A ({nx36011,nx36153,nx36295,nx36437,nx36579,nx36721,
            nx36863,nx37005,nx37147,nx37289,nx37431,nx37573,nx37715,nx37857,
            nx37999,nx38141}), .B ({nx33767,nx33907,nx34045,nx34183,nx34321,
            nx34459,nx34597,nx34737,nx34879,nx35021,nx35163,nx35305,nx35447,
            nx35589,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35731), .C ({inputRegisters_447__15,inputRegisters_447__14,
            inputRegisters_447__13,inputRegisters_447__12,inputRegisters_447__11
            ,inputRegisters_447__10,inputRegisters_447__9,inputRegisters_447__8,
            inputRegisters_447__7,inputRegisters_447__6,inputRegisters_447__5,
            inputRegisters_447__4,inputRegisters_447__3,inputRegisters_447__2,
            inputRegisters_447__1,inputRegisters_447__0})) ;
    Reg_16 loop1_447_x (.D ({inputRegisters_447__15,inputRegisters_447__14,
           inputRegisters_447__13,inputRegisters_447__12,inputRegisters_447__11,
           inputRegisters_447__10,inputRegisters_447__9,inputRegisters_447__8,
           inputRegisters_447__7,inputRegisters_447__6,inputRegisters_447__5,
           inputRegisters_447__4,inputRegisters_447__3,inputRegisters_447__2,
           inputRegisters_447__1,inputRegisters_447__0}), .en (
           enableRegister_447), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_447__15,registerOutputs_447__14,
           registerOutputs_447__13,registerOutputs_447__12,
           registerOutputs_447__11,registerOutputs_447__10,
           registerOutputs_447__9,registerOutputs_447__8,registerOutputs_447__7,
           registerOutputs_447__6,registerOutputs_447__5,registerOutputs_447__4,
           registerOutputs_447__3,registerOutputs_447__2,registerOutputs_447__1,
           registerOutputs_447__0})) ;
    Mux2_16 loop1_448_y (.A ({nx36013,nx36155,nx36297,nx36439,nx36581,nx36723,
            nx36865,nx37007,nx37149,nx37291,nx37433,nx37575,nx37717,nx37859,
            nx38001,nx38143}), .B ({nx33769,nx33907,nx34045,nx34183,nx34321,
            nx34459,nx34597,nx34739,nx34881,nx35023,nx35165,nx35307,nx35449,
            nx35591,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35733), .C ({inputRegisters_448__15,inputRegisters_448__14,
            inputRegisters_448__13,inputRegisters_448__12,inputRegisters_448__11
            ,inputRegisters_448__10,inputRegisters_448__9,inputRegisters_448__8,
            inputRegisters_448__7,inputRegisters_448__6,inputRegisters_448__5,
            inputRegisters_448__4,inputRegisters_448__3,inputRegisters_448__2,
            inputRegisters_448__1,inputRegisters_448__0})) ;
    Reg_16 loop1_448_x (.D ({inputRegisters_448__15,inputRegisters_448__14,
           inputRegisters_448__13,inputRegisters_448__12,inputRegisters_448__11,
           inputRegisters_448__10,inputRegisters_448__9,inputRegisters_448__8,
           inputRegisters_448__7,inputRegisters_448__6,inputRegisters_448__5,
           inputRegisters_448__4,inputRegisters_448__3,inputRegisters_448__2,
           inputRegisters_448__1,inputRegisters_448__0}), .en (
           enableRegister_448), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_448__15,registerOutputs_448__14,
           registerOutputs_448__13,registerOutputs_448__12,
           registerOutputs_448__11,registerOutputs_448__10,
           registerOutputs_448__9,registerOutputs_448__8,registerOutputs_448__7,
           registerOutputs_448__6,registerOutputs_448__5,registerOutputs_448__4,
           registerOutputs_448__3,registerOutputs_448__2,registerOutputs_448__1,
           registerOutputs_448__0})) ;
    Mux2_16 loop1_449_y (.A ({nx36013,nx36155,nx36297,nx36439,nx36581,nx36723,
            nx36865,nx37007,nx37149,nx37291,nx37433,nx37575,nx37717,nx37859,
            nx38001,nx38143}), .B ({nx33769,nx33907,nx34045,nx34183,nx34321,
            nx34459,nx34599,nx34739,nx34881,nx35023,nx35165,nx35307,nx35449,
            nx35591,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35733), .C ({inputRegisters_449__15,inputRegisters_449__14,
            inputRegisters_449__13,inputRegisters_449__12,inputRegisters_449__11
            ,inputRegisters_449__10,inputRegisters_449__9,inputRegisters_449__8,
            inputRegisters_449__7,inputRegisters_449__6,inputRegisters_449__5,
            inputRegisters_449__4,inputRegisters_449__3,inputRegisters_449__2,
            inputRegisters_449__1,inputRegisters_449__0})) ;
    Reg_16 loop1_449_x (.D ({inputRegisters_449__15,inputRegisters_449__14,
           inputRegisters_449__13,inputRegisters_449__12,inputRegisters_449__11,
           inputRegisters_449__10,inputRegisters_449__9,inputRegisters_449__8,
           inputRegisters_449__7,inputRegisters_449__6,inputRegisters_449__5,
           inputRegisters_449__4,inputRegisters_449__3,inputRegisters_449__2,
           inputRegisters_449__1,inputRegisters_449__0}), .en (
           enableRegister_449), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_449__15,registerOutputs_449__14,
           registerOutputs_449__13,registerOutputs_449__12,
           registerOutputs_449__11,registerOutputs_449__10,
           registerOutputs_449__9,registerOutputs_449__8,registerOutputs_449__7,
           registerOutputs_449__6,registerOutputs_449__5,registerOutputs_449__4,
           registerOutputs_449__3,registerOutputs_449__2,registerOutputs_449__1,
           registerOutputs_449__0})) ;
    Mux2_16 loop1_450_y (.A ({nx36013,nx36155,nx36297,nx36439,nx36581,nx36723,
            nx36865,nx37007,nx37149,nx37291,nx37433,nx37575,nx37717,nx37859,
            nx38001,nx38143}), .B ({nx33769,nx33907,nx34045,nx34183,nx34321,
            nx34461,nx34599,nx34739,nx34881,nx35023,nx35165,nx35307,nx35449,
            nx35591,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35733), .C ({inputRegisters_450__15,inputRegisters_450__14,
            inputRegisters_450__13,inputRegisters_450__12,inputRegisters_450__11
            ,inputRegisters_450__10,inputRegisters_450__9,inputRegisters_450__8,
            inputRegisters_450__7,inputRegisters_450__6,inputRegisters_450__5,
            inputRegisters_450__4,inputRegisters_450__3,inputRegisters_450__2,
            inputRegisters_450__1,inputRegisters_450__0})) ;
    Reg_16 loop1_450_x (.D ({inputRegisters_450__15,inputRegisters_450__14,
           inputRegisters_450__13,inputRegisters_450__12,inputRegisters_450__11,
           inputRegisters_450__10,inputRegisters_450__9,inputRegisters_450__8,
           inputRegisters_450__7,inputRegisters_450__6,inputRegisters_450__5,
           inputRegisters_450__4,inputRegisters_450__3,inputRegisters_450__2,
           inputRegisters_450__1,inputRegisters_450__0}), .en (
           enableRegister_450), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_450__15,registerOutputs_450__14,
           registerOutputs_450__13,registerOutputs_450__12,
           registerOutputs_450__11,registerOutputs_450__10,
           registerOutputs_450__9,registerOutputs_450__8,registerOutputs_450__7,
           registerOutputs_450__6,registerOutputs_450__5,registerOutputs_450__4,
           registerOutputs_450__3,registerOutputs_450__2,registerOutputs_450__1,
           registerOutputs_450__0})) ;
    Mux2_16 loop1_451_y (.A ({nx36013,nx36155,nx36297,nx36439,nx36581,nx36723,
            nx36865,nx37007,nx37149,nx37291,nx37433,nx37575,nx37717,nx37859,
            nx38001,nx38143}), .B ({nx33769,nx33907,nx34045,nx34183,nx34323,
            nx34461,nx34599,nx34739,nx34881,nx35023,nx35165,nx35307,nx35449,
            nx35591,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35733), .C ({inputRegisters_451__15,inputRegisters_451__14,
            inputRegisters_451__13,inputRegisters_451__12,inputRegisters_451__11
            ,inputRegisters_451__10,inputRegisters_451__9,inputRegisters_451__8,
            inputRegisters_451__7,inputRegisters_451__6,inputRegisters_451__5,
            inputRegisters_451__4,inputRegisters_451__3,inputRegisters_451__2,
            inputRegisters_451__1,inputRegisters_451__0})) ;
    Reg_16 loop1_451_x (.D ({inputRegisters_451__15,inputRegisters_451__14,
           inputRegisters_451__13,inputRegisters_451__12,inputRegisters_451__11,
           inputRegisters_451__10,inputRegisters_451__9,inputRegisters_451__8,
           inputRegisters_451__7,inputRegisters_451__6,inputRegisters_451__5,
           inputRegisters_451__4,inputRegisters_451__3,inputRegisters_451__2,
           inputRegisters_451__1,inputRegisters_451__0}), .en (
           enableRegister_451), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_451__15,registerOutputs_451__14,
           registerOutputs_451__13,registerOutputs_451__12,
           registerOutputs_451__11,registerOutputs_451__10,
           registerOutputs_451__9,registerOutputs_451__8,registerOutputs_451__7,
           registerOutputs_451__6,registerOutputs_451__5,registerOutputs_451__4,
           registerOutputs_451__3,registerOutputs_451__2,registerOutputs_451__1,
           registerOutputs_451__0})) ;
    Mux2_16 loop1_452_y (.A ({nx36013,nx36155,nx36297,nx36439,nx36581,nx36723,
            nx36865,nx37007,nx37149,nx37291,nx37433,nx37575,nx37717,nx37859,
            nx38001,nx38143}), .B ({nx33769,nx33907,nx34045,nx34185,nx34323,
            nx34461,nx34599,nx34739,nx34881,nx35023,nx35165,nx35307,nx35449,
            nx35591,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35733), .C ({inputRegisters_452__15,inputRegisters_452__14,
            inputRegisters_452__13,inputRegisters_452__12,inputRegisters_452__11
            ,inputRegisters_452__10,inputRegisters_452__9,inputRegisters_452__8,
            inputRegisters_452__7,inputRegisters_452__6,inputRegisters_452__5,
            inputRegisters_452__4,inputRegisters_452__3,inputRegisters_452__2,
            inputRegisters_452__1,inputRegisters_452__0})) ;
    Reg_16 loop1_452_x (.D ({inputRegisters_452__15,inputRegisters_452__14,
           inputRegisters_452__13,inputRegisters_452__12,inputRegisters_452__11,
           inputRegisters_452__10,inputRegisters_452__9,inputRegisters_452__8,
           inputRegisters_452__7,inputRegisters_452__6,inputRegisters_452__5,
           inputRegisters_452__4,inputRegisters_452__3,inputRegisters_452__2,
           inputRegisters_452__1,inputRegisters_452__0}), .en (
           enableRegister_452), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_452__15,registerOutputs_452__14,
           registerOutputs_452__13,registerOutputs_452__12,
           registerOutputs_452__11,registerOutputs_452__10,
           registerOutputs_452__9,registerOutputs_452__8,registerOutputs_452__7,
           registerOutputs_452__6,registerOutputs_452__5,registerOutputs_452__4,
           registerOutputs_452__3,registerOutputs_452__2,registerOutputs_452__1,
           registerOutputs_452__0})) ;
    Mux2_16 loop1_453_y (.A ({nx36013,nx36155,nx36297,nx36439,nx36581,nx36723,
            nx36865,nx37007,nx37149,nx37291,nx37433,nx37575,nx37717,nx37859,
            nx38001,nx38143}), .B ({nx33769,nx33907,nx34047,nx34185,nx34323,
            nx34461,nx34599,nx34739,nx34881,nx35023,nx35165,nx35307,nx35449,
            nx35591,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35733), .C ({inputRegisters_453__15,inputRegisters_453__14,
            inputRegisters_453__13,inputRegisters_453__12,inputRegisters_453__11
            ,inputRegisters_453__10,inputRegisters_453__9,inputRegisters_453__8,
            inputRegisters_453__7,inputRegisters_453__6,inputRegisters_453__5,
            inputRegisters_453__4,inputRegisters_453__3,inputRegisters_453__2,
            inputRegisters_453__1,inputRegisters_453__0})) ;
    Reg_16 loop1_453_x (.D ({inputRegisters_453__15,inputRegisters_453__14,
           inputRegisters_453__13,inputRegisters_453__12,inputRegisters_453__11,
           inputRegisters_453__10,inputRegisters_453__9,inputRegisters_453__8,
           inputRegisters_453__7,inputRegisters_453__6,inputRegisters_453__5,
           inputRegisters_453__4,inputRegisters_453__3,inputRegisters_453__2,
           inputRegisters_453__1,inputRegisters_453__0}), .en (
           enableRegister_453), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_453__15,registerOutputs_453__14,
           registerOutputs_453__13,registerOutputs_453__12,
           registerOutputs_453__11,registerOutputs_453__10,
           registerOutputs_453__9,registerOutputs_453__8,registerOutputs_453__7,
           registerOutputs_453__6,registerOutputs_453__5,registerOutputs_453__4,
           registerOutputs_453__3,registerOutputs_453__2,registerOutputs_453__1,
           registerOutputs_453__0})) ;
    Mux2_16 loop1_454_y (.A ({nx36013,nx36155,nx36297,nx36439,nx36581,nx36723,
            nx36865,nx37007,nx37149,nx37291,nx37433,nx37575,nx37717,nx37859,
            nx38001,nx38143}), .B ({nx33769,nx33909,nx34047,nx34185,nx34323,
            nx34461,nx34599,nx34739,nx34881,nx35023,nx35165,nx35307,nx35449,
            nx35591,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35733), .C ({inputRegisters_454__15,inputRegisters_454__14,
            inputRegisters_454__13,inputRegisters_454__12,inputRegisters_454__11
            ,inputRegisters_454__10,inputRegisters_454__9,inputRegisters_454__8,
            inputRegisters_454__7,inputRegisters_454__6,inputRegisters_454__5,
            inputRegisters_454__4,inputRegisters_454__3,inputRegisters_454__2,
            inputRegisters_454__1,inputRegisters_454__0})) ;
    Reg_16 loop1_454_x (.D ({inputRegisters_454__15,inputRegisters_454__14,
           inputRegisters_454__13,inputRegisters_454__12,inputRegisters_454__11,
           inputRegisters_454__10,inputRegisters_454__9,inputRegisters_454__8,
           inputRegisters_454__7,inputRegisters_454__6,inputRegisters_454__5,
           inputRegisters_454__4,inputRegisters_454__3,inputRegisters_454__2,
           inputRegisters_454__1,inputRegisters_454__0}), .en (
           enableRegister_454), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_454__15,registerOutputs_454__14,
           registerOutputs_454__13,registerOutputs_454__12,
           registerOutputs_454__11,registerOutputs_454__10,
           registerOutputs_454__9,registerOutputs_454__8,registerOutputs_454__7,
           registerOutputs_454__6,registerOutputs_454__5,registerOutputs_454__4,
           registerOutputs_454__3,registerOutputs_454__2,registerOutputs_454__1,
           registerOutputs_454__0})) ;
    Mux2_16 loop1_455_y (.A ({nx36015,nx36157,nx36299,nx36441,nx36583,nx36725,
            nx36867,nx37009,nx37151,nx37293,nx37435,nx37577,nx37719,nx37861,
            nx38003,nx38145}), .B ({nx33771,nx33909,nx34047,nx34185,nx34323,
            nx34461,nx34599,nx34741,nx34883,nx35025,nx35167,nx35309,nx35451,
            nx35593,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35735), .C ({inputRegisters_455__15,inputRegisters_455__14,
            inputRegisters_455__13,inputRegisters_455__12,inputRegisters_455__11
            ,inputRegisters_455__10,inputRegisters_455__9,inputRegisters_455__8,
            inputRegisters_455__7,inputRegisters_455__6,inputRegisters_455__5,
            inputRegisters_455__4,inputRegisters_455__3,inputRegisters_455__2,
            inputRegisters_455__1,inputRegisters_455__0})) ;
    Reg_16 loop1_455_x (.D ({inputRegisters_455__15,inputRegisters_455__14,
           inputRegisters_455__13,inputRegisters_455__12,inputRegisters_455__11,
           inputRegisters_455__10,inputRegisters_455__9,inputRegisters_455__8,
           inputRegisters_455__7,inputRegisters_455__6,inputRegisters_455__5,
           inputRegisters_455__4,inputRegisters_455__3,inputRegisters_455__2,
           inputRegisters_455__1,inputRegisters_455__0}), .en (
           enableRegister_455), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_455__15,registerOutputs_455__14,
           registerOutputs_455__13,registerOutputs_455__12,
           registerOutputs_455__11,registerOutputs_455__10,
           registerOutputs_455__9,registerOutputs_455__8,registerOutputs_455__7,
           registerOutputs_455__6,registerOutputs_455__5,registerOutputs_455__4,
           registerOutputs_455__3,registerOutputs_455__2,registerOutputs_455__1,
           registerOutputs_455__0})) ;
    Mux2_16 loop1_456_y (.A ({nx36015,nx36157,nx36299,nx36441,nx36583,nx36725,
            nx36867,nx37009,nx37151,nx37293,nx37435,nx37577,nx37719,nx37861,
            nx38003,nx38145}), .B ({nx33771,nx33909,nx34047,nx34185,nx34323,
            nx34461,nx34601,nx34741,nx34883,nx35025,nx35167,nx35309,nx35451,
            nx35593,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35735), .C ({inputRegisters_456__15,inputRegisters_456__14,
            inputRegisters_456__13,inputRegisters_456__12,inputRegisters_456__11
            ,inputRegisters_456__10,inputRegisters_456__9,inputRegisters_456__8,
            inputRegisters_456__7,inputRegisters_456__6,inputRegisters_456__5,
            inputRegisters_456__4,inputRegisters_456__3,inputRegisters_456__2,
            inputRegisters_456__1,inputRegisters_456__0})) ;
    Reg_16 loop1_456_x (.D ({inputRegisters_456__15,inputRegisters_456__14,
           inputRegisters_456__13,inputRegisters_456__12,inputRegisters_456__11,
           inputRegisters_456__10,inputRegisters_456__9,inputRegisters_456__8,
           inputRegisters_456__7,inputRegisters_456__6,inputRegisters_456__5,
           inputRegisters_456__4,inputRegisters_456__3,inputRegisters_456__2,
           inputRegisters_456__1,inputRegisters_456__0}), .en (
           enableRegister_456), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_456__15,registerOutputs_456__14,
           registerOutputs_456__13,registerOutputs_456__12,
           registerOutputs_456__11,registerOutputs_456__10,
           registerOutputs_456__9,registerOutputs_456__8,registerOutputs_456__7,
           registerOutputs_456__6,registerOutputs_456__5,registerOutputs_456__4,
           registerOutputs_456__3,registerOutputs_456__2,registerOutputs_456__1,
           registerOutputs_456__0})) ;
    Mux2_16 loop1_457_y (.A ({nx36015,nx36157,nx36299,nx36441,nx36583,nx36725,
            nx36867,nx37009,nx37151,nx37293,nx37435,nx37577,nx37719,nx37861,
            nx38003,nx38145}), .B ({nx33771,nx33909,nx34047,nx34185,nx34323,
            nx34463,nx34601,nx34741,nx34883,nx35025,nx35167,nx35309,nx35451,
            nx35593,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35735), .C ({inputRegisters_457__15,inputRegisters_457__14,
            inputRegisters_457__13,inputRegisters_457__12,inputRegisters_457__11
            ,inputRegisters_457__10,inputRegisters_457__9,inputRegisters_457__8,
            inputRegisters_457__7,inputRegisters_457__6,inputRegisters_457__5,
            inputRegisters_457__4,inputRegisters_457__3,inputRegisters_457__2,
            inputRegisters_457__1,inputRegisters_457__0})) ;
    Reg_16 loop1_457_x (.D ({inputRegisters_457__15,inputRegisters_457__14,
           inputRegisters_457__13,inputRegisters_457__12,inputRegisters_457__11,
           inputRegisters_457__10,inputRegisters_457__9,inputRegisters_457__8,
           inputRegisters_457__7,inputRegisters_457__6,inputRegisters_457__5,
           inputRegisters_457__4,inputRegisters_457__3,inputRegisters_457__2,
           inputRegisters_457__1,inputRegisters_457__0}), .en (
           enableRegister_457), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_457__15,registerOutputs_457__14,
           registerOutputs_457__13,registerOutputs_457__12,
           registerOutputs_457__11,registerOutputs_457__10,
           registerOutputs_457__9,registerOutputs_457__8,registerOutputs_457__7,
           registerOutputs_457__6,registerOutputs_457__5,registerOutputs_457__4,
           registerOutputs_457__3,registerOutputs_457__2,registerOutputs_457__1,
           registerOutputs_457__0})) ;
    Mux2_16 loop1_458_y (.A ({nx36015,nx36157,nx36299,nx36441,nx36583,nx36725,
            nx36867,nx37009,nx37151,nx37293,nx37435,nx37577,nx37719,nx37861,
            nx38003,nx38145}), .B ({nx33771,nx33909,nx34047,nx34185,nx34325,
            nx34463,nx34601,nx34741,nx34883,nx35025,nx35167,nx35309,nx35451,
            nx35593,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35735), .C ({inputRegisters_458__15,inputRegisters_458__14,
            inputRegisters_458__13,inputRegisters_458__12,inputRegisters_458__11
            ,inputRegisters_458__10,inputRegisters_458__9,inputRegisters_458__8,
            inputRegisters_458__7,inputRegisters_458__6,inputRegisters_458__5,
            inputRegisters_458__4,inputRegisters_458__3,inputRegisters_458__2,
            inputRegisters_458__1,inputRegisters_458__0})) ;
    Reg_16 loop1_458_x (.D ({inputRegisters_458__15,inputRegisters_458__14,
           inputRegisters_458__13,inputRegisters_458__12,inputRegisters_458__11,
           inputRegisters_458__10,inputRegisters_458__9,inputRegisters_458__8,
           inputRegisters_458__7,inputRegisters_458__6,inputRegisters_458__5,
           inputRegisters_458__4,inputRegisters_458__3,inputRegisters_458__2,
           inputRegisters_458__1,inputRegisters_458__0}), .en (
           enableRegister_458), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_458__15,registerOutputs_458__14,
           registerOutputs_458__13,registerOutputs_458__12,
           registerOutputs_458__11,registerOutputs_458__10,
           registerOutputs_458__9,registerOutputs_458__8,registerOutputs_458__7,
           registerOutputs_458__6,registerOutputs_458__5,registerOutputs_458__4,
           registerOutputs_458__3,registerOutputs_458__2,registerOutputs_458__1,
           registerOutputs_458__0})) ;
    Mux2_16 loop1_459_y (.A ({nx36015,nx36157,nx36299,nx36441,nx36583,nx36725,
            nx36867,nx37009,nx37151,nx37293,nx37435,nx37577,nx37719,nx37861,
            nx38003,nx38145}), .B ({nx33771,nx33909,nx34047,nx34187,nx34325,
            nx34463,nx34601,nx34741,nx34883,nx35025,nx35167,nx35309,nx35451,
            nx35593,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35735), .C ({inputRegisters_459__15,inputRegisters_459__14,
            inputRegisters_459__13,inputRegisters_459__12,inputRegisters_459__11
            ,inputRegisters_459__10,inputRegisters_459__9,inputRegisters_459__8,
            inputRegisters_459__7,inputRegisters_459__6,inputRegisters_459__5,
            inputRegisters_459__4,inputRegisters_459__3,inputRegisters_459__2,
            inputRegisters_459__1,inputRegisters_459__0})) ;
    Reg_16 loop1_459_x (.D ({inputRegisters_459__15,inputRegisters_459__14,
           inputRegisters_459__13,inputRegisters_459__12,inputRegisters_459__11,
           inputRegisters_459__10,inputRegisters_459__9,inputRegisters_459__8,
           inputRegisters_459__7,inputRegisters_459__6,inputRegisters_459__5,
           inputRegisters_459__4,inputRegisters_459__3,inputRegisters_459__2,
           inputRegisters_459__1,inputRegisters_459__0}), .en (
           enableRegister_459), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_459__15,registerOutputs_459__14,
           registerOutputs_459__13,registerOutputs_459__12,
           registerOutputs_459__11,registerOutputs_459__10,
           registerOutputs_459__9,registerOutputs_459__8,registerOutputs_459__7,
           registerOutputs_459__6,registerOutputs_459__5,registerOutputs_459__4,
           registerOutputs_459__3,registerOutputs_459__2,registerOutputs_459__1,
           registerOutputs_459__0})) ;
    Mux2_16 loop1_460_y (.A ({nx36015,nx36157,nx36299,nx36441,nx36583,nx36725,
            nx36867,nx37009,nx37151,nx37293,nx37435,nx37577,nx37719,nx37861,
            nx38003,nx38145}), .B ({nx33771,nx33909,nx34049,nx34187,nx34325,
            nx34463,nx34601,nx34741,nx34883,nx35025,nx35167,nx35309,nx35451,
            nx35593,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35735), .C ({inputRegisters_460__15,inputRegisters_460__14,
            inputRegisters_460__13,inputRegisters_460__12,inputRegisters_460__11
            ,inputRegisters_460__10,inputRegisters_460__9,inputRegisters_460__8,
            inputRegisters_460__7,inputRegisters_460__6,inputRegisters_460__5,
            inputRegisters_460__4,inputRegisters_460__3,inputRegisters_460__2,
            inputRegisters_460__1,inputRegisters_460__0})) ;
    Reg_16 loop1_460_x (.D ({inputRegisters_460__15,inputRegisters_460__14,
           inputRegisters_460__13,inputRegisters_460__12,inputRegisters_460__11,
           inputRegisters_460__10,inputRegisters_460__9,inputRegisters_460__8,
           inputRegisters_460__7,inputRegisters_460__6,inputRegisters_460__5,
           inputRegisters_460__4,inputRegisters_460__3,inputRegisters_460__2,
           inputRegisters_460__1,inputRegisters_460__0}), .en (
           enableRegister_460), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_460__15,registerOutputs_460__14,
           registerOutputs_460__13,registerOutputs_460__12,
           registerOutputs_460__11,registerOutputs_460__10,
           registerOutputs_460__9,registerOutputs_460__8,registerOutputs_460__7,
           registerOutputs_460__6,registerOutputs_460__5,registerOutputs_460__4,
           registerOutputs_460__3,registerOutputs_460__2,registerOutputs_460__1,
           registerOutputs_460__0})) ;
    Mux2_16 loop1_461_y (.A ({nx36015,nx36157,nx36299,nx36441,nx36583,nx36725,
            nx36867,nx37009,nx37151,nx37293,nx37435,nx37577,nx37719,nx37861,
            nx38003,nx38145}), .B ({nx33771,nx33911,nx34049,nx34187,nx34325,
            nx34463,nx34601,nx34741,nx34883,nx35025,nx35167,nx35309,nx35451,
            nx35593,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35735), .C ({inputRegisters_461__15,inputRegisters_461__14,
            inputRegisters_461__13,inputRegisters_461__12,inputRegisters_461__11
            ,inputRegisters_461__10,inputRegisters_461__9,inputRegisters_461__8,
            inputRegisters_461__7,inputRegisters_461__6,inputRegisters_461__5,
            inputRegisters_461__4,inputRegisters_461__3,inputRegisters_461__2,
            inputRegisters_461__1,inputRegisters_461__0})) ;
    Reg_16 loop1_461_x (.D ({inputRegisters_461__15,inputRegisters_461__14,
           inputRegisters_461__13,inputRegisters_461__12,inputRegisters_461__11,
           inputRegisters_461__10,inputRegisters_461__9,inputRegisters_461__8,
           inputRegisters_461__7,inputRegisters_461__6,inputRegisters_461__5,
           inputRegisters_461__4,inputRegisters_461__3,inputRegisters_461__2,
           inputRegisters_461__1,inputRegisters_461__0}), .en (
           enableRegister_461), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_461__15,registerOutputs_461__14,
           registerOutputs_461__13,registerOutputs_461__12,
           registerOutputs_461__11,registerOutputs_461__10,
           registerOutputs_461__9,registerOutputs_461__8,registerOutputs_461__7,
           registerOutputs_461__6,registerOutputs_461__5,registerOutputs_461__4,
           registerOutputs_461__3,registerOutputs_461__2,registerOutputs_461__1,
           registerOutputs_461__0})) ;
    Mux2_16 loop1_462_y (.A ({nx36017,nx36159,nx36301,nx36443,nx36585,nx36727,
            nx36869,nx37011,nx37153,nx37295,nx37437,nx37579,nx37721,nx37863,
            nx38005,nx38147}), .B ({nx33773,nx33911,nx34049,nx34187,nx34325,
            nx34463,nx34601,nx34743,nx34885,nx35027,nx35169,nx35311,nx35453,
            nx35595,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35737), .C ({inputRegisters_462__15,inputRegisters_462__14,
            inputRegisters_462__13,inputRegisters_462__12,inputRegisters_462__11
            ,inputRegisters_462__10,inputRegisters_462__9,inputRegisters_462__8,
            inputRegisters_462__7,inputRegisters_462__6,inputRegisters_462__5,
            inputRegisters_462__4,inputRegisters_462__3,inputRegisters_462__2,
            inputRegisters_462__1,inputRegisters_462__0})) ;
    Reg_16 loop1_462_x (.D ({inputRegisters_462__15,inputRegisters_462__14,
           inputRegisters_462__13,inputRegisters_462__12,inputRegisters_462__11,
           inputRegisters_462__10,inputRegisters_462__9,inputRegisters_462__8,
           inputRegisters_462__7,inputRegisters_462__6,inputRegisters_462__5,
           inputRegisters_462__4,inputRegisters_462__3,inputRegisters_462__2,
           inputRegisters_462__1,inputRegisters_462__0}), .en (
           enableRegister_462), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_462__15,registerOutputs_462__14,
           registerOutputs_462__13,registerOutputs_462__12,
           registerOutputs_462__11,registerOutputs_462__10,
           registerOutputs_462__9,registerOutputs_462__8,registerOutputs_462__7,
           registerOutputs_462__6,registerOutputs_462__5,registerOutputs_462__4,
           registerOutputs_462__3,registerOutputs_462__2,registerOutputs_462__1,
           registerOutputs_462__0})) ;
    Mux2_16 loop1_463_y (.A ({nx36017,nx36159,nx36301,nx36443,nx36585,nx36727,
            nx36869,nx37011,nx37153,nx37295,nx37437,nx37579,nx37721,nx37863,
            nx38005,nx38147}), .B ({nx33773,nx33911,nx34049,nx34187,nx34325,
            nx34463,nx34603,nx34743,nx34885,nx35027,nx35169,nx35311,nx35453,
            nx35595,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35737), .C ({inputRegisters_463__15,inputRegisters_463__14,
            inputRegisters_463__13,inputRegisters_463__12,inputRegisters_463__11
            ,inputRegisters_463__10,inputRegisters_463__9,inputRegisters_463__8,
            inputRegisters_463__7,inputRegisters_463__6,inputRegisters_463__5,
            inputRegisters_463__4,inputRegisters_463__3,inputRegisters_463__2,
            inputRegisters_463__1,inputRegisters_463__0})) ;
    Reg_16 loop1_463_x (.D ({inputRegisters_463__15,inputRegisters_463__14,
           inputRegisters_463__13,inputRegisters_463__12,inputRegisters_463__11,
           inputRegisters_463__10,inputRegisters_463__9,inputRegisters_463__8,
           inputRegisters_463__7,inputRegisters_463__6,inputRegisters_463__5,
           inputRegisters_463__4,inputRegisters_463__3,inputRegisters_463__2,
           inputRegisters_463__1,inputRegisters_463__0}), .en (
           enableRegister_463), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_463__15,registerOutputs_463__14,
           registerOutputs_463__13,registerOutputs_463__12,
           registerOutputs_463__11,registerOutputs_463__10,
           registerOutputs_463__9,registerOutputs_463__8,registerOutputs_463__7,
           registerOutputs_463__6,registerOutputs_463__5,registerOutputs_463__4,
           registerOutputs_463__3,registerOutputs_463__2,registerOutputs_463__1,
           registerOutputs_463__0})) ;
    Mux2_16 loop1_464_y (.A ({nx36017,nx36159,nx36301,nx36443,nx36585,nx36727,
            nx36869,nx37011,nx37153,nx37295,nx37437,nx37579,nx37721,nx37863,
            nx38005,nx38147}), .B ({nx33773,nx33911,nx34049,nx34187,nx34325,
            nx34465,nx34603,nx34743,nx34885,nx35027,nx35169,nx35311,nx35453,
            nx35595,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35737), .C ({inputRegisters_464__15,inputRegisters_464__14,
            inputRegisters_464__13,inputRegisters_464__12,inputRegisters_464__11
            ,inputRegisters_464__10,inputRegisters_464__9,inputRegisters_464__8,
            inputRegisters_464__7,inputRegisters_464__6,inputRegisters_464__5,
            inputRegisters_464__4,inputRegisters_464__3,inputRegisters_464__2,
            inputRegisters_464__1,inputRegisters_464__0})) ;
    Reg_16 loop1_464_x (.D ({inputRegisters_464__15,inputRegisters_464__14,
           inputRegisters_464__13,inputRegisters_464__12,inputRegisters_464__11,
           inputRegisters_464__10,inputRegisters_464__9,inputRegisters_464__8,
           inputRegisters_464__7,inputRegisters_464__6,inputRegisters_464__5,
           inputRegisters_464__4,inputRegisters_464__3,inputRegisters_464__2,
           inputRegisters_464__1,inputRegisters_464__0}), .en (
           enableRegister_464), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_464__15,registerOutputs_464__14,
           registerOutputs_464__13,registerOutputs_464__12,
           registerOutputs_464__11,registerOutputs_464__10,
           registerOutputs_464__9,registerOutputs_464__8,registerOutputs_464__7,
           registerOutputs_464__6,registerOutputs_464__5,registerOutputs_464__4,
           registerOutputs_464__3,registerOutputs_464__2,registerOutputs_464__1,
           registerOutputs_464__0})) ;
    Mux2_16 loop1_465_y (.A ({nx36017,nx36159,nx36301,nx36443,nx36585,nx36727,
            nx36869,nx37011,nx37153,nx37295,nx37437,nx37579,nx37721,nx37863,
            nx38005,nx38147}), .B ({nx33773,nx33911,nx34049,nx34187,nx34327,
            nx34465,nx34603,nx34743,nx34885,nx35027,nx35169,nx35311,nx35453,
            nx35595,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35737), .C ({inputRegisters_465__15,inputRegisters_465__14,
            inputRegisters_465__13,inputRegisters_465__12,inputRegisters_465__11
            ,inputRegisters_465__10,inputRegisters_465__9,inputRegisters_465__8,
            inputRegisters_465__7,inputRegisters_465__6,inputRegisters_465__5,
            inputRegisters_465__4,inputRegisters_465__3,inputRegisters_465__2,
            inputRegisters_465__1,inputRegisters_465__0})) ;
    Reg_16 loop1_465_x (.D ({inputRegisters_465__15,inputRegisters_465__14,
           inputRegisters_465__13,inputRegisters_465__12,inputRegisters_465__11,
           inputRegisters_465__10,inputRegisters_465__9,inputRegisters_465__8,
           inputRegisters_465__7,inputRegisters_465__6,inputRegisters_465__5,
           inputRegisters_465__4,inputRegisters_465__3,inputRegisters_465__2,
           inputRegisters_465__1,inputRegisters_465__0}), .en (
           enableRegister_465), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_465__15,registerOutputs_465__14,
           registerOutputs_465__13,registerOutputs_465__12,
           registerOutputs_465__11,registerOutputs_465__10,
           registerOutputs_465__9,registerOutputs_465__8,registerOutputs_465__7,
           registerOutputs_465__6,registerOutputs_465__5,registerOutputs_465__4,
           registerOutputs_465__3,registerOutputs_465__2,registerOutputs_465__1,
           registerOutputs_465__0})) ;
    Mux2_16 loop1_466_y (.A ({nx36017,nx36159,nx36301,nx36443,nx36585,nx36727,
            nx36869,nx37011,nx37153,nx37295,nx37437,nx37579,nx37721,nx37863,
            nx38005,nx38147}), .B ({nx33773,nx33911,nx34049,nx34189,nx34327,
            nx34465,nx34603,nx34743,nx34885,nx35027,nx35169,nx35311,nx35453,
            nx35595,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35737), .C ({inputRegisters_466__15,inputRegisters_466__14,
            inputRegisters_466__13,inputRegisters_466__12,inputRegisters_466__11
            ,inputRegisters_466__10,inputRegisters_466__9,inputRegisters_466__8,
            inputRegisters_466__7,inputRegisters_466__6,inputRegisters_466__5,
            inputRegisters_466__4,inputRegisters_466__3,inputRegisters_466__2,
            inputRegisters_466__1,inputRegisters_466__0})) ;
    Reg_16 loop1_466_x (.D ({inputRegisters_466__15,inputRegisters_466__14,
           inputRegisters_466__13,inputRegisters_466__12,inputRegisters_466__11,
           inputRegisters_466__10,inputRegisters_466__9,inputRegisters_466__8,
           inputRegisters_466__7,inputRegisters_466__6,inputRegisters_466__5,
           inputRegisters_466__4,inputRegisters_466__3,inputRegisters_466__2,
           inputRegisters_466__1,inputRegisters_466__0}), .en (
           enableRegister_466), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_466__15,registerOutputs_466__14,
           registerOutputs_466__13,registerOutputs_466__12,
           registerOutputs_466__11,registerOutputs_466__10,
           registerOutputs_466__9,registerOutputs_466__8,registerOutputs_466__7,
           registerOutputs_466__6,registerOutputs_466__5,registerOutputs_466__4,
           registerOutputs_466__3,registerOutputs_466__2,registerOutputs_466__1,
           registerOutputs_466__0})) ;
    Mux2_16 loop1_467_y (.A ({nx36017,nx36159,nx36301,nx36443,nx36585,nx36727,
            nx36869,nx37011,nx37153,nx37295,nx37437,nx37579,nx37721,nx37863,
            nx38005,nx38147}), .B ({nx33773,nx33911,nx34051,nx34189,nx34327,
            nx34465,nx34603,nx34743,nx34885,nx35027,nx35169,nx35311,nx35453,
            nx35595,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35737), .C ({inputRegisters_467__15,inputRegisters_467__14,
            inputRegisters_467__13,inputRegisters_467__12,inputRegisters_467__11
            ,inputRegisters_467__10,inputRegisters_467__9,inputRegisters_467__8,
            inputRegisters_467__7,inputRegisters_467__6,inputRegisters_467__5,
            inputRegisters_467__4,inputRegisters_467__3,inputRegisters_467__2,
            inputRegisters_467__1,inputRegisters_467__0})) ;
    Reg_16 loop1_467_x (.D ({inputRegisters_467__15,inputRegisters_467__14,
           inputRegisters_467__13,inputRegisters_467__12,inputRegisters_467__11,
           inputRegisters_467__10,inputRegisters_467__9,inputRegisters_467__8,
           inputRegisters_467__7,inputRegisters_467__6,inputRegisters_467__5,
           inputRegisters_467__4,inputRegisters_467__3,inputRegisters_467__2,
           inputRegisters_467__1,inputRegisters_467__0}), .en (
           enableRegister_467), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_467__15,registerOutputs_467__14,
           registerOutputs_467__13,registerOutputs_467__12,
           registerOutputs_467__11,registerOutputs_467__10,
           registerOutputs_467__9,registerOutputs_467__8,registerOutputs_467__7,
           registerOutputs_467__6,registerOutputs_467__5,registerOutputs_467__4,
           registerOutputs_467__3,registerOutputs_467__2,registerOutputs_467__1,
           registerOutputs_467__0})) ;
    Mux2_16 loop1_468_y (.A ({nx36017,nx36159,nx36301,nx36443,nx36585,nx36727,
            nx36869,nx37011,nx37153,nx37295,nx37437,nx37579,nx37721,nx37863,
            nx38005,nx38147}), .B ({nx33773,nx33913,nx34051,nx34189,nx34327,
            nx34465,nx34603,nx34743,nx34885,nx35027,nx35169,nx35311,nx35453,
            nx35595,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35737), .C ({inputRegisters_468__15,inputRegisters_468__14,
            inputRegisters_468__13,inputRegisters_468__12,inputRegisters_468__11
            ,inputRegisters_468__10,inputRegisters_468__9,inputRegisters_468__8,
            inputRegisters_468__7,inputRegisters_468__6,inputRegisters_468__5,
            inputRegisters_468__4,inputRegisters_468__3,inputRegisters_468__2,
            inputRegisters_468__1,inputRegisters_468__0})) ;
    Reg_16 loop1_468_x (.D ({inputRegisters_468__15,inputRegisters_468__14,
           inputRegisters_468__13,inputRegisters_468__12,inputRegisters_468__11,
           inputRegisters_468__10,inputRegisters_468__9,inputRegisters_468__8,
           inputRegisters_468__7,inputRegisters_468__6,inputRegisters_468__5,
           inputRegisters_468__4,inputRegisters_468__3,inputRegisters_468__2,
           inputRegisters_468__1,inputRegisters_468__0}), .en (
           enableRegister_468), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_468__15,registerOutputs_468__14,
           registerOutputs_468__13,registerOutputs_468__12,
           registerOutputs_468__11,registerOutputs_468__10,
           registerOutputs_468__9,registerOutputs_468__8,registerOutputs_468__7,
           registerOutputs_468__6,registerOutputs_468__5,registerOutputs_468__4,
           registerOutputs_468__3,registerOutputs_468__2,registerOutputs_468__1,
           registerOutputs_468__0})) ;
    Mux2_16 loop1_469_y (.A ({nx36019,nx36161,nx36303,nx36445,nx36587,nx36729,
            nx36871,nx37013,nx37155,nx37297,nx37439,nx37581,nx37723,nx37865,
            nx38007,nx38149}), .B ({nx33775,nx33913,nx34051,nx34189,nx34327,
            nx34465,nx34603,nx34745,nx34887,nx35029,nx35171,nx35313,nx35455,
            nx35597,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35739), .C ({inputRegisters_469__15,inputRegisters_469__14,
            inputRegisters_469__13,inputRegisters_469__12,inputRegisters_469__11
            ,inputRegisters_469__10,inputRegisters_469__9,inputRegisters_469__8,
            inputRegisters_469__7,inputRegisters_469__6,inputRegisters_469__5,
            inputRegisters_469__4,inputRegisters_469__3,inputRegisters_469__2,
            inputRegisters_469__1,inputRegisters_469__0})) ;
    Reg_16 loop1_469_x (.D ({inputRegisters_469__15,inputRegisters_469__14,
           inputRegisters_469__13,inputRegisters_469__12,inputRegisters_469__11,
           inputRegisters_469__10,inputRegisters_469__9,inputRegisters_469__8,
           inputRegisters_469__7,inputRegisters_469__6,inputRegisters_469__5,
           inputRegisters_469__4,inputRegisters_469__3,inputRegisters_469__2,
           inputRegisters_469__1,inputRegisters_469__0}), .en (
           enableRegister_469), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_469__15,registerOutputs_469__14,
           registerOutputs_469__13,registerOutputs_469__12,
           registerOutputs_469__11,registerOutputs_469__10,
           registerOutputs_469__9,registerOutputs_469__8,registerOutputs_469__7,
           registerOutputs_469__6,registerOutputs_469__5,registerOutputs_469__4,
           registerOutputs_469__3,registerOutputs_469__2,registerOutputs_469__1,
           registerOutputs_469__0})) ;
    Mux2_16 loop1_470_y (.A ({nx36019,nx36161,nx36303,nx36445,nx36587,nx36729,
            nx36871,nx37013,nx37155,nx37297,nx37439,nx37581,nx37723,nx37865,
            nx38007,nx38149}), .B ({nx33775,nx33913,nx34051,nx34189,nx34327,
            nx34465,nx34605,nx34745,nx34887,nx35029,nx35171,nx35313,nx35455,
            nx35597,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35739), .C ({inputRegisters_470__15,inputRegisters_470__14,
            inputRegisters_470__13,inputRegisters_470__12,inputRegisters_470__11
            ,inputRegisters_470__10,inputRegisters_470__9,inputRegisters_470__8,
            inputRegisters_470__7,inputRegisters_470__6,inputRegisters_470__5,
            inputRegisters_470__4,inputRegisters_470__3,inputRegisters_470__2,
            inputRegisters_470__1,inputRegisters_470__0})) ;
    Reg_16 loop1_470_x (.D ({inputRegisters_470__15,inputRegisters_470__14,
           inputRegisters_470__13,inputRegisters_470__12,inputRegisters_470__11,
           inputRegisters_470__10,inputRegisters_470__9,inputRegisters_470__8,
           inputRegisters_470__7,inputRegisters_470__6,inputRegisters_470__5,
           inputRegisters_470__4,inputRegisters_470__3,inputRegisters_470__2,
           inputRegisters_470__1,inputRegisters_470__0}), .en (
           enableRegister_470), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_470__15,registerOutputs_470__14,
           registerOutputs_470__13,registerOutputs_470__12,
           registerOutputs_470__11,registerOutputs_470__10,
           registerOutputs_470__9,registerOutputs_470__8,registerOutputs_470__7,
           registerOutputs_470__6,registerOutputs_470__5,registerOutputs_470__4,
           registerOutputs_470__3,registerOutputs_470__2,registerOutputs_470__1,
           registerOutputs_470__0})) ;
    Mux2_16 loop1_471_y (.A ({nx36019,nx36161,nx36303,nx36445,nx36587,nx36729,
            nx36871,nx37013,nx37155,nx37297,nx37439,nx37581,nx37723,nx37865,
            nx38007,nx38149}), .B ({nx33775,nx33913,nx34051,nx34189,nx34327,
            nx34467,nx34605,nx34745,nx34887,nx35029,nx35171,nx35313,nx35455,
            nx35597,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35739), .C ({inputRegisters_471__15,inputRegisters_471__14,
            inputRegisters_471__13,inputRegisters_471__12,inputRegisters_471__11
            ,inputRegisters_471__10,inputRegisters_471__9,inputRegisters_471__8,
            inputRegisters_471__7,inputRegisters_471__6,inputRegisters_471__5,
            inputRegisters_471__4,inputRegisters_471__3,inputRegisters_471__2,
            inputRegisters_471__1,inputRegisters_471__0})) ;
    Reg_16 loop1_471_x (.D ({inputRegisters_471__15,inputRegisters_471__14,
           inputRegisters_471__13,inputRegisters_471__12,inputRegisters_471__11,
           inputRegisters_471__10,inputRegisters_471__9,inputRegisters_471__8,
           inputRegisters_471__7,inputRegisters_471__6,inputRegisters_471__5,
           inputRegisters_471__4,inputRegisters_471__3,inputRegisters_471__2,
           inputRegisters_471__1,inputRegisters_471__0}), .en (
           enableRegister_471), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_471__15,registerOutputs_471__14,
           registerOutputs_471__13,registerOutputs_471__12,
           registerOutputs_471__11,registerOutputs_471__10,
           registerOutputs_471__9,registerOutputs_471__8,registerOutputs_471__7,
           registerOutputs_471__6,registerOutputs_471__5,registerOutputs_471__4,
           registerOutputs_471__3,registerOutputs_471__2,registerOutputs_471__1,
           registerOutputs_471__0})) ;
    Mux2_16 loop1_472_y (.A ({nx36019,nx36161,nx36303,nx36445,nx36587,nx36729,
            nx36871,nx37013,nx37155,nx37297,nx37439,nx37581,nx37723,nx37865,
            nx38007,nx38149}), .B ({nx33775,nx33913,nx34051,nx34189,nx34329,
            nx34467,nx34605,nx34745,nx34887,nx35029,nx35171,nx35313,nx35455,
            nx35597,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35739), .C ({inputRegisters_472__15,inputRegisters_472__14,
            inputRegisters_472__13,inputRegisters_472__12,inputRegisters_472__11
            ,inputRegisters_472__10,inputRegisters_472__9,inputRegisters_472__8,
            inputRegisters_472__7,inputRegisters_472__6,inputRegisters_472__5,
            inputRegisters_472__4,inputRegisters_472__3,inputRegisters_472__2,
            inputRegisters_472__1,inputRegisters_472__0})) ;
    Reg_16 loop1_472_x (.D ({inputRegisters_472__15,inputRegisters_472__14,
           inputRegisters_472__13,inputRegisters_472__12,inputRegisters_472__11,
           inputRegisters_472__10,inputRegisters_472__9,inputRegisters_472__8,
           inputRegisters_472__7,inputRegisters_472__6,inputRegisters_472__5,
           inputRegisters_472__4,inputRegisters_472__3,inputRegisters_472__2,
           inputRegisters_472__1,inputRegisters_472__0}), .en (
           enableRegister_472), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_472__15,registerOutputs_472__14,
           registerOutputs_472__13,registerOutputs_472__12,
           registerOutputs_472__11,registerOutputs_472__10,
           registerOutputs_472__9,registerOutputs_472__8,registerOutputs_472__7,
           registerOutputs_472__6,registerOutputs_472__5,registerOutputs_472__4,
           registerOutputs_472__3,registerOutputs_472__2,registerOutputs_472__1,
           registerOutputs_472__0})) ;
    Mux2_16 loop1_473_y (.A ({nx36019,nx36161,nx36303,nx36445,nx36587,nx36729,
            nx36871,nx37013,nx37155,nx37297,nx37439,nx37581,nx37723,nx37865,
            nx38007,nx38149}), .B ({nx33775,nx33913,nx34051,nx34191,nx34329,
            nx34467,nx34605,nx34745,nx34887,nx35029,nx35171,nx35313,nx35455,
            nx35597,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35739), .C ({inputRegisters_473__15,inputRegisters_473__14,
            inputRegisters_473__13,inputRegisters_473__12,inputRegisters_473__11
            ,inputRegisters_473__10,inputRegisters_473__9,inputRegisters_473__8,
            inputRegisters_473__7,inputRegisters_473__6,inputRegisters_473__5,
            inputRegisters_473__4,inputRegisters_473__3,inputRegisters_473__2,
            inputRegisters_473__1,inputRegisters_473__0})) ;
    Reg_16 loop1_473_x (.D ({inputRegisters_473__15,inputRegisters_473__14,
           inputRegisters_473__13,inputRegisters_473__12,inputRegisters_473__11,
           inputRegisters_473__10,inputRegisters_473__9,inputRegisters_473__8,
           inputRegisters_473__7,inputRegisters_473__6,inputRegisters_473__5,
           inputRegisters_473__4,inputRegisters_473__3,inputRegisters_473__2,
           inputRegisters_473__1,inputRegisters_473__0}), .en (
           enableRegister_473), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_473__15,registerOutputs_473__14,
           registerOutputs_473__13,registerOutputs_473__12,
           registerOutputs_473__11,registerOutputs_473__10,
           registerOutputs_473__9,registerOutputs_473__8,registerOutputs_473__7,
           registerOutputs_473__6,registerOutputs_473__5,registerOutputs_473__4,
           registerOutputs_473__3,registerOutputs_473__2,registerOutputs_473__1,
           registerOutputs_473__0})) ;
    Mux2_16 loop1_474_y (.A ({nx36019,nx36161,nx36303,nx36445,nx36587,nx36729,
            nx36871,nx37013,nx37155,nx37297,nx37439,nx37581,nx37723,nx37865,
            nx38007,nx38149}), .B ({nx33775,nx33913,nx34053,nx34191,nx34329,
            nx34467,nx34605,nx34745,nx34887,nx35029,nx35171,nx35313,nx35455,
            nx35597,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35739), .C ({inputRegisters_474__15,inputRegisters_474__14,
            inputRegisters_474__13,inputRegisters_474__12,inputRegisters_474__11
            ,inputRegisters_474__10,inputRegisters_474__9,inputRegisters_474__8,
            inputRegisters_474__7,inputRegisters_474__6,inputRegisters_474__5,
            inputRegisters_474__4,inputRegisters_474__3,inputRegisters_474__2,
            inputRegisters_474__1,inputRegisters_474__0})) ;
    Reg_16 loop1_474_x (.D ({inputRegisters_474__15,inputRegisters_474__14,
           inputRegisters_474__13,inputRegisters_474__12,inputRegisters_474__11,
           inputRegisters_474__10,inputRegisters_474__9,inputRegisters_474__8,
           inputRegisters_474__7,inputRegisters_474__6,inputRegisters_474__5,
           inputRegisters_474__4,inputRegisters_474__3,inputRegisters_474__2,
           inputRegisters_474__1,inputRegisters_474__0}), .en (
           enableRegister_474), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_474__15,registerOutputs_474__14,
           registerOutputs_474__13,registerOutputs_474__12,
           registerOutputs_474__11,registerOutputs_474__10,
           registerOutputs_474__9,registerOutputs_474__8,registerOutputs_474__7,
           registerOutputs_474__6,registerOutputs_474__5,registerOutputs_474__4,
           registerOutputs_474__3,registerOutputs_474__2,registerOutputs_474__1,
           registerOutputs_474__0})) ;
    Mux2_16 loop1_475_y (.A ({nx36019,nx36161,nx36303,nx36445,nx36587,nx36729,
            nx36871,nx37013,nx37155,nx37297,nx37439,nx37581,nx37723,nx37865,
            nx38007,nx38149}), .B ({nx33775,nx33915,nx34053,nx34191,nx34329,
            nx34467,nx34605,nx34745,nx34887,nx35029,nx35171,nx35313,nx35455,
            nx35597,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35739), .C ({inputRegisters_475__15,inputRegisters_475__14,
            inputRegisters_475__13,inputRegisters_475__12,inputRegisters_475__11
            ,inputRegisters_475__10,inputRegisters_475__9,inputRegisters_475__8,
            inputRegisters_475__7,inputRegisters_475__6,inputRegisters_475__5,
            inputRegisters_475__4,inputRegisters_475__3,inputRegisters_475__2,
            inputRegisters_475__1,inputRegisters_475__0})) ;
    Reg_16 loop1_475_x (.D ({inputRegisters_475__15,inputRegisters_475__14,
           inputRegisters_475__13,inputRegisters_475__12,inputRegisters_475__11,
           inputRegisters_475__10,inputRegisters_475__9,inputRegisters_475__8,
           inputRegisters_475__7,inputRegisters_475__6,inputRegisters_475__5,
           inputRegisters_475__4,inputRegisters_475__3,inputRegisters_475__2,
           inputRegisters_475__1,inputRegisters_475__0}), .en (
           enableRegister_475), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_475__15,registerOutputs_475__14,
           registerOutputs_475__13,registerOutputs_475__12,
           registerOutputs_475__11,registerOutputs_475__10,
           registerOutputs_475__9,registerOutputs_475__8,registerOutputs_475__7,
           registerOutputs_475__6,registerOutputs_475__5,registerOutputs_475__4,
           registerOutputs_475__3,registerOutputs_475__2,registerOutputs_475__1,
           registerOutputs_475__0})) ;
    Mux2_16 loop1_476_y (.A ({nx36021,nx36163,nx36305,nx36447,nx36589,nx36731,
            nx36873,nx37015,nx37157,nx37299,nx37441,nx37583,nx37725,nx37867,
            nx38009,nx38151}), .B ({nx33777,nx33915,nx34053,nx34191,nx34329,
            nx34467,nx34605,nx34747,nx34889,nx35031,nx35173,nx35315,nx35457,
            nx35599,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35741), .C ({inputRegisters_476__15,inputRegisters_476__14,
            inputRegisters_476__13,inputRegisters_476__12,inputRegisters_476__11
            ,inputRegisters_476__10,inputRegisters_476__9,inputRegisters_476__8,
            inputRegisters_476__7,inputRegisters_476__6,inputRegisters_476__5,
            inputRegisters_476__4,inputRegisters_476__3,inputRegisters_476__2,
            inputRegisters_476__1,inputRegisters_476__0})) ;
    Reg_16 loop1_476_x (.D ({inputRegisters_476__15,inputRegisters_476__14,
           inputRegisters_476__13,inputRegisters_476__12,inputRegisters_476__11,
           inputRegisters_476__10,inputRegisters_476__9,inputRegisters_476__8,
           inputRegisters_476__7,inputRegisters_476__6,inputRegisters_476__5,
           inputRegisters_476__4,inputRegisters_476__3,inputRegisters_476__2,
           inputRegisters_476__1,inputRegisters_476__0}), .en (
           enableRegister_476), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_476__15,registerOutputs_476__14,
           registerOutputs_476__13,registerOutputs_476__12,
           registerOutputs_476__11,registerOutputs_476__10,
           registerOutputs_476__9,registerOutputs_476__8,registerOutputs_476__7,
           registerOutputs_476__6,registerOutputs_476__5,registerOutputs_476__4,
           registerOutputs_476__3,registerOutputs_476__2,registerOutputs_476__1,
           registerOutputs_476__0})) ;
    Mux2_16 loop1_477_y (.A ({nx36021,nx36163,nx36305,nx36447,nx36589,nx36731,
            nx36873,nx37015,nx37157,nx37299,nx37441,nx37583,nx37725,nx37867,
            nx38009,nx38151}), .B ({nx33777,nx33915,nx34053,nx34191,nx34329,
            nx34467,nx34607,nx34747,nx34889,nx35031,nx35173,nx35315,nx35457,
            nx35599,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35741), .C ({inputRegisters_477__15,inputRegisters_477__14,
            inputRegisters_477__13,inputRegisters_477__12,inputRegisters_477__11
            ,inputRegisters_477__10,inputRegisters_477__9,inputRegisters_477__8,
            inputRegisters_477__7,inputRegisters_477__6,inputRegisters_477__5,
            inputRegisters_477__4,inputRegisters_477__3,inputRegisters_477__2,
            inputRegisters_477__1,inputRegisters_477__0})) ;
    Reg_16 loop1_477_x (.D ({inputRegisters_477__15,inputRegisters_477__14,
           inputRegisters_477__13,inputRegisters_477__12,inputRegisters_477__11,
           inputRegisters_477__10,inputRegisters_477__9,inputRegisters_477__8,
           inputRegisters_477__7,inputRegisters_477__6,inputRegisters_477__5,
           inputRegisters_477__4,inputRegisters_477__3,inputRegisters_477__2,
           inputRegisters_477__1,inputRegisters_477__0}), .en (
           enableRegister_477), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_477__15,registerOutputs_477__14,
           registerOutputs_477__13,registerOutputs_477__12,
           registerOutputs_477__11,registerOutputs_477__10,
           registerOutputs_477__9,registerOutputs_477__8,registerOutputs_477__7,
           registerOutputs_477__6,registerOutputs_477__5,registerOutputs_477__4,
           registerOutputs_477__3,registerOutputs_477__2,registerOutputs_477__1,
           registerOutputs_477__0})) ;
    Mux2_16 loop1_478_y (.A ({nx36021,nx36163,nx36305,nx36447,nx36589,nx36731,
            nx36873,nx37015,nx37157,nx37299,nx37441,nx37583,nx37725,nx37867,
            nx38009,nx38151}), .B ({nx33777,nx33915,nx34053,nx34191,nx34329,
            nx34469,nx34607,nx34747,nx34889,nx35031,nx35173,nx35315,nx35457,
            nx35599,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35741), .C ({inputRegisters_478__15,inputRegisters_478__14,
            inputRegisters_478__13,inputRegisters_478__12,inputRegisters_478__11
            ,inputRegisters_478__10,inputRegisters_478__9,inputRegisters_478__8,
            inputRegisters_478__7,inputRegisters_478__6,inputRegisters_478__5,
            inputRegisters_478__4,inputRegisters_478__3,inputRegisters_478__2,
            inputRegisters_478__1,inputRegisters_478__0})) ;
    Reg_16 loop1_478_x (.D ({inputRegisters_478__15,inputRegisters_478__14,
           inputRegisters_478__13,inputRegisters_478__12,inputRegisters_478__11,
           inputRegisters_478__10,inputRegisters_478__9,inputRegisters_478__8,
           inputRegisters_478__7,inputRegisters_478__6,inputRegisters_478__5,
           inputRegisters_478__4,inputRegisters_478__3,inputRegisters_478__2,
           inputRegisters_478__1,inputRegisters_478__0}), .en (
           enableRegister_478), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_478__15,registerOutputs_478__14,
           registerOutputs_478__13,registerOutputs_478__12,
           registerOutputs_478__11,registerOutputs_478__10,
           registerOutputs_478__9,registerOutputs_478__8,registerOutputs_478__7,
           registerOutputs_478__6,registerOutputs_478__5,registerOutputs_478__4,
           registerOutputs_478__3,registerOutputs_478__2,registerOutputs_478__1,
           registerOutputs_478__0})) ;
    Mux2_16 loop1_479_y (.A ({nx36021,nx36163,nx36305,nx36447,nx36589,nx36731,
            nx36873,nx37015,nx37157,nx37299,nx37441,nx37583,nx37725,nx37867,
            nx38009,nx38151}), .B ({nx33777,nx33915,nx34053,nx34191,nx34331,
            nx34469,nx34607,nx34747,nx34889,nx35031,nx35173,nx35315,nx35457,
            nx35599,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35741), .C ({inputRegisters_479__15,inputRegisters_479__14,
            inputRegisters_479__13,inputRegisters_479__12,inputRegisters_479__11
            ,inputRegisters_479__10,inputRegisters_479__9,inputRegisters_479__8,
            inputRegisters_479__7,inputRegisters_479__6,inputRegisters_479__5,
            inputRegisters_479__4,inputRegisters_479__3,inputRegisters_479__2,
            inputRegisters_479__1,inputRegisters_479__0})) ;
    Reg_16 loop1_479_x (.D ({inputRegisters_479__15,inputRegisters_479__14,
           inputRegisters_479__13,inputRegisters_479__12,inputRegisters_479__11,
           inputRegisters_479__10,inputRegisters_479__9,inputRegisters_479__8,
           inputRegisters_479__7,inputRegisters_479__6,inputRegisters_479__5,
           inputRegisters_479__4,inputRegisters_479__3,inputRegisters_479__2,
           inputRegisters_479__1,inputRegisters_479__0}), .en (
           enableRegister_479), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_479__15,registerOutputs_479__14,
           registerOutputs_479__13,registerOutputs_479__12,
           registerOutputs_479__11,registerOutputs_479__10,
           registerOutputs_479__9,registerOutputs_479__8,registerOutputs_479__7,
           registerOutputs_479__6,registerOutputs_479__5,registerOutputs_479__4,
           registerOutputs_479__3,registerOutputs_479__2,registerOutputs_479__1,
           registerOutputs_479__0})) ;
    Mux2_16 loop1_480_y (.A ({nx36021,nx36163,nx36305,nx36447,nx36589,nx36731,
            nx36873,nx37015,nx37157,nx37299,nx37441,nx37583,nx37725,nx37867,
            nx38009,nx38151}), .B ({nx33777,nx33915,nx34053,nx34193,nx34331,
            nx34469,nx34607,nx34747,nx34889,nx35031,nx35173,nx35315,nx35457,
            nx35599,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35741), .C ({inputRegisters_480__15,inputRegisters_480__14,
            inputRegisters_480__13,inputRegisters_480__12,inputRegisters_480__11
            ,inputRegisters_480__10,inputRegisters_480__9,inputRegisters_480__8,
            inputRegisters_480__7,inputRegisters_480__6,inputRegisters_480__5,
            inputRegisters_480__4,inputRegisters_480__3,inputRegisters_480__2,
            inputRegisters_480__1,inputRegisters_480__0})) ;
    Reg_16 loop1_480_x (.D ({inputRegisters_480__15,inputRegisters_480__14,
           inputRegisters_480__13,inputRegisters_480__12,inputRegisters_480__11,
           inputRegisters_480__10,inputRegisters_480__9,inputRegisters_480__8,
           inputRegisters_480__7,inputRegisters_480__6,inputRegisters_480__5,
           inputRegisters_480__4,inputRegisters_480__3,inputRegisters_480__2,
           inputRegisters_480__1,inputRegisters_480__0}), .en (
           enableRegister_480), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_480__15,registerOutputs_480__14,
           registerOutputs_480__13,registerOutputs_480__12,
           registerOutputs_480__11,registerOutputs_480__10,
           registerOutputs_480__9,registerOutputs_480__8,registerOutputs_480__7,
           registerOutputs_480__6,registerOutputs_480__5,registerOutputs_480__4,
           registerOutputs_480__3,registerOutputs_480__2,registerOutputs_480__1,
           registerOutputs_480__0})) ;
    Mux2_16 loop1_481_y (.A ({nx36021,nx36163,nx36305,nx36447,nx36589,nx36731,
            nx36873,nx37015,nx37157,nx37299,nx37441,nx37583,nx37725,nx37867,
            nx38009,nx38151}), .B ({nx33777,nx33915,nx34055,nx34193,nx34331,
            nx34469,nx34607,nx34747,nx34889,nx35031,nx35173,nx35315,nx35457,
            nx35599,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35741), .C ({inputRegisters_481__15,inputRegisters_481__14,
            inputRegisters_481__13,inputRegisters_481__12,inputRegisters_481__11
            ,inputRegisters_481__10,inputRegisters_481__9,inputRegisters_481__8,
            inputRegisters_481__7,inputRegisters_481__6,inputRegisters_481__5,
            inputRegisters_481__4,inputRegisters_481__3,inputRegisters_481__2,
            inputRegisters_481__1,inputRegisters_481__0})) ;
    Reg_16 loop1_481_x (.D ({inputRegisters_481__15,inputRegisters_481__14,
           inputRegisters_481__13,inputRegisters_481__12,inputRegisters_481__11,
           inputRegisters_481__10,inputRegisters_481__9,inputRegisters_481__8,
           inputRegisters_481__7,inputRegisters_481__6,inputRegisters_481__5,
           inputRegisters_481__4,inputRegisters_481__3,inputRegisters_481__2,
           inputRegisters_481__1,inputRegisters_481__0}), .en (
           enableRegister_481), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_481__15,registerOutputs_481__14,
           registerOutputs_481__13,registerOutputs_481__12,
           registerOutputs_481__11,registerOutputs_481__10,
           registerOutputs_481__9,registerOutputs_481__8,registerOutputs_481__7,
           registerOutputs_481__6,registerOutputs_481__5,registerOutputs_481__4,
           registerOutputs_481__3,registerOutputs_481__2,registerOutputs_481__1,
           registerOutputs_481__0})) ;
    Mux2_16 loop1_482_y (.A ({nx36021,nx36163,nx36305,nx36447,nx36589,nx36731,
            nx36873,nx37015,nx37157,nx37299,nx37441,nx37583,nx37725,nx37867,
            nx38009,nx38151}), .B ({nx33777,nx33917,nx34055,nx34193,nx34331,
            nx34469,nx34607,nx34747,nx34889,nx35031,nx35173,nx35315,nx35457,
            nx35599,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35741), .C ({inputRegisters_482__15,inputRegisters_482__14,
            inputRegisters_482__13,inputRegisters_482__12,inputRegisters_482__11
            ,inputRegisters_482__10,inputRegisters_482__9,inputRegisters_482__8,
            inputRegisters_482__7,inputRegisters_482__6,inputRegisters_482__5,
            inputRegisters_482__4,inputRegisters_482__3,inputRegisters_482__2,
            inputRegisters_482__1,inputRegisters_482__0})) ;
    Reg_16 loop1_482_x (.D ({inputRegisters_482__15,inputRegisters_482__14,
           inputRegisters_482__13,inputRegisters_482__12,inputRegisters_482__11,
           inputRegisters_482__10,inputRegisters_482__9,inputRegisters_482__8,
           inputRegisters_482__7,inputRegisters_482__6,inputRegisters_482__5,
           inputRegisters_482__4,inputRegisters_482__3,inputRegisters_482__2,
           inputRegisters_482__1,inputRegisters_482__0}), .en (
           enableRegister_482), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_482__15,registerOutputs_482__14,
           registerOutputs_482__13,registerOutputs_482__12,
           registerOutputs_482__11,registerOutputs_482__10,
           registerOutputs_482__9,registerOutputs_482__8,registerOutputs_482__7,
           registerOutputs_482__6,registerOutputs_482__5,registerOutputs_482__4,
           registerOutputs_482__3,registerOutputs_482__2,registerOutputs_482__1,
           registerOutputs_482__0})) ;
    Mux2_16 loop1_483_y (.A ({nx36023,nx36165,nx36307,nx36449,nx36591,nx36733,
            nx36875,nx37017,nx37159,nx37301,nx37443,nx37585,nx37727,nx37869,
            nx38011,nx38153}), .B ({nx33779,nx33917,nx34055,nx34193,nx34331,
            nx34469,nx34607,nx34749,nx34891,nx35033,nx35175,nx35317,nx35459,
            nx35601,registerOutputs_484__15,registerOutputs_484__15}), .S (
            nx35743), .C ({inputRegisters_483__15,inputRegisters_483__14,
            inputRegisters_483__13,inputRegisters_483__12,inputRegisters_483__11
            ,inputRegisters_483__10,inputRegisters_483__9,inputRegisters_483__8,
            inputRegisters_483__7,inputRegisters_483__6,inputRegisters_483__5,
            inputRegisters_483__4,inputRegisters_483__3,inputRegisters_483__2,
            inputRegisters_483__1,inputRegisters_483__0})) ;
    Reg_16 loop1_483_x (.D ({inputRegisters_483__15,inputRegisters_483__14,
           inputRegisters_483__13,inputRegisters_483__12,inputRegisters_483__11,
           inputRegisters_483__10,inputRegisters_483__9,inputRegisters_483__8,
           inputRegisters_483__7,inputRegisters_483__6,inputRegisters_483__5,
           inputRegisters_483__4,inputRegisters_483__3,inputRegisters_483__2,
           inputRegisters_483__1,inputRegisters_483__0}), .en (
           enableRegister_483), .clk (clk), .rst (resetRegisters), .Q ({
           registerOutputs_483__15,registerOutputs_483__14,
           registerOutputs_483__13,registerOutputs_483__12,
           registerOutputs_483__11,registerOutputs_483__10,
           registerOutputs_483__9,registerOutputs_483__8,registerOutputs_483__7,
           registerOutputs_483__6,registerOutputs_483__5,registerOutputs_483__4,
           registerOutputs_483__3,registerOutputs_483__2,registerOutputs_483__1,
           registerOutputs_483__0})) ;
    Mux_512 selectedRegisterMUX (.inputs_0__15 (registerOutputs_0__15), .inputs_0__14 (
            registerOutputs_0__14), .inputs_0__13 (registerOutputs_0__13), .inputs_0__12 (
            registerOutputs_0__12), .inputs_0__11 (registerOutputs_0__11), .inputs_0__10 (
            registerOutputs_0__10), .inputs_0__9 (registerOutputs_0__9), .inputs_0__8 (
            registerOutputs_0__8), .inputs_0__7 (registerOutputs_0__7), .inputs_0__6 (
            registerOutputs_0__6), .inputs_0__5 (registerOutputs_0__5), .inputs_0__4 (
            registerOutputs_0__4), .inputs_0__3 (registerOutputs_0__3), .inputs_0__2 (
            registerOutputs_0__2), .inputs_0__1 (registerOutputs_0__1), .inputs_0__0 (
            registerOutputs_0__0), .inputs_1__15 (registerOutputs_1__15), .inputs_1__14 (
            registerOutputs_1__14), .inputs_1__13 (registerOutputs_1__13), .inputs_1__12 (
            registerOutputs_1__12), .inputs_1__11 (registerOutputs_1__11), .inputs_1__10 (
            registerOutputs_1__10), .inputs_1__9 (registerOutputs_1__9), .inputs_1__8 (
            registerOutputs_1__8), .inputs_1__7 (registerOutputs_1__7), .inputs_1__6 (
            registerOutputs_1__6), .inputs_1__5 (registerOutputs_1__5), .inputs_1__4 (
            registerOutputs_1__4), .inputs_1__3 (registerOutputs_1__3), .inputs_1__2 (
            registerOutputs_1__2), .inputs_1__1 (registerOutputs_1__1), .inputs_1__0 (
            registerOutputs_1__0), .inputs_2__15 (registerOutputs_2__15), .inputs_2__14 (
            registerOutputs_2__14), .inputs_2__13 (registerOutputs_2__13), .inputs_2__12 (
            registerOutputs_2__12), .inputs_2__11 (registerOutputs_2__11), .inputs_2__10 (
            registerOutputs_2__10), .inputs_2__9 (registerOutputs_2__9), .inputs_2__8 (
            registerOutputs_2__8), .inputs_2__7 (registerOutputs_2__7), .inputs_2__6 (
            registerOutputs_2__6), .inputs_2__5 (registerOutputs_2__5), .inputs_2__4 (
            registerOutputs_2__4), .inputs_2__3 (registerOutputs_2__3), .inputs_2__2 (
            registerOutputs_2__2), .inputs_2__1 (registerOutputs_2__1), .inputs_2__0 (
            registerOutputs_2__0), .inputs_3__15 (registerOutputs_3__15), .inputs_3__14 (
            registerOutputs_3__14), .inputs_3__13 (registerOutputs_3__13), .inputs_3__12 (
            registerOutputs_3__12), .inputs_3__11 (registerOutputs_3__11), .inputs_3__10 (
            registerOutputs_3__10), .inputs_3__9 (registerOutputs_3__9), .inputs_3__8 (
            registerOutputs_3__8), .inputs_3__7 (registerOutputs_3__7), .inputs_3__6 (
            registerOutputs_3__6), .inputs_3__5 (registerOutputs_3__5), .inputs_3__4 (
            registerOutputs_3__4), .inputs_3__3 (registerOutputs_3__3), .inputs_3__2 (
            registerOutputs_3__2), .inputs_3__1 (registerOutputs_3__1), .inputs_3__0 (
            registerOutputs_3__0), .inputs_4__15 (registerOutputs_4__15), .inputs_4__14 (
            registerOutputs_4__14), .inputs_4__13 (registerOutputs_4__13), .inputs_4__12 (
            registerOutputs_4__12), .inputs_4__11 (registerOutputs_4__11), .inputs_4__10 (
            registerOutputs_4__10), .inputs_4__9 (registerOutputs_4__9), .inputs_4__8 (
            registerOutputs_4__8), .inputs_4__7 (registerOutputs_4__7), .inputs_4__6 (
            registerOutputs_4__6), .inputs_4__5 (registerOutputs_4__5), .inputs_4__4 (
            registerOutputs_4__4), .inputs_4__3 (registerOutputs_4__3), .inputs_4__2 (
            registerOutputs_4__2), .inputs_4__1 (registerOutputs_4__1), .inputs_4__0 (
            registerOutputs_4__0), .inputs_5__15 (registerOutputs_5__15), .inputs_5__14 (
            registerOutputs_5__14), .inputs_5__13 (registerOutputs_5__13), .inputs_5__12 (
            registerOutputs_5__12), .inputs_5__11 (registerOutputs_5__11), .inputs_5__10 (
            registerOutputs_5__10), .inputs_5__9 (registerOutputs_5__9), .inputs_5__8 (
            registerOutputs_5__8), .inputs_5__7 (registerOutputs_5__7), .inputs_5__6 (
            registerOutputs_5__6), .inputs_5__5 (registerOutputs_5__5), .inputs_5__4 (
            registerOutputs_5__4), .inputs_5__3 (registerOutputs_5__3), .inputs_5__2 (
            registerOutputs_5__2), .inputs_5__1 (registerOutputs_5__1), .inputs_5__0 (
            registerOutputs_5__0), .inputs_6__15 (registerOutputs_6__15), .inputs_6__14 (
            registerOutputs_6__14), .inputs_6__13 (registerOutputs_6__13), .inputs_6__12 (
            registerOutputs_6__12), .inputs_6__11 (registerOutputs_6__11), .inputs_6__10 (
            registerOutputs_6__10), .inputs_6__9 (registerOutputs_6__9), .inputs_6__8 (
            registerOutputs_6__8), .inputs_6__7 (registerOutputs_6__7), .inputs_6__6 (
            registerOutputs_6__6), .inputs_6__5 (registerOutputs_6__5), .inputs_6__4 (
            registerOutputs_6__4), .inputs_6__3 (registerOutputs_6__3), .inputs_6__2 (
            registerOutputs_6__2), .inputs_6__1 (registerOutputs_6__1), .inputs_6__0 (
            registerOutputs_6__0), .inputs_7__15 (registerOutputs_7__15), .inputs_7__14 (
            registerOutputs_7__14), .inputs_7__13 (registerOutputs_7__13), .inputs_7__12 (
            registerOutputs_7__12), .inputs_7__11 (registerOutputs_7__11), .inputs_7__10 (
            registerOutputs_7__10), .inputs_7__9 (registerOutputs_7__9), .inputs_7__8 (
            registerOutputs_7__8), .inputs_7__7 (registerOutputs_7__7), .inputs_7__6 (
            registerOutputs_7__6), .inputs_7__5 (registerOutputs_7__5), .inputs_7__4 (
            registerOutputs_7__4), .inputs_7__3 (registerOutputs_7__3), .inputs_7__2 (
            registerOutputs_7__2), .inputs_7__1 (registerOutputs_7__1), .inputs_7__0 (
            registerOutputs_7__0), .inputs_8__15 (registerOutputs_8__15), .inputs_8__14 (
            registerOutputs_8__14), .inputs_8__13 (registerOutputs_8__13), .inputs_8__12 (
            registerOutputs_8__12), .inputs_8__11 (registerOutputs_8__11), .inputs_8__10 (
            registerOutputs_8__10), .inputs_8__9 (registerOutputs_8__9), .inputs_8__8 (
            registerOutputs_8__8), .inputs_8__7 (registerOutputs_8__7), .inputs_8__6 (
            registerOutputs_8__6), .inputs_8__5 (registerOutputs_8__5), .inputs_8__4 (
            registerOutputs_8__4), .inputs_8__3 (registerOutputs_8__3), .inputs_8__2 (
            registerOutputs_8__2), .inputs_8__1 (registerOutputs_8__1), .inputs_8__0 (
            registerOutputs_8__0), .inputs_9__15 (registerOutputs_9__15), .inputs_9__14 (
            registerOutputs_9__14), .inputs_9__13 (registerOutputs_9__13), .inputs_9__12 (
            registerOutputs_9__12), .inputs_9__11 (registerOutputs_9__11), .inputs_9__10 (
            registerOutputs_9__10), .inputs_9__9 (registerOutputs_9__9), .inputs_9__8 (
            registerOutputs_9__8), .inputs_9__7 (registerOutputs_9__7), .inputs_9__6 (
            registerOutputs_9__6), .inputs_9__5 (registerOutputs_9__5), .inputs_9__4 (
            registerOutputs_9__4), .inputs_9__3 (registerOutputs_9__3), .inputs_9__2 (
            registerOutputs_9__2), .inputs_9__1 (registerOutputs_9__1), .inputs_9__0 (
            registerOutputs_9__0), .inputs_10__15 (registerOutputs_10__15), .inputs_10__14 (
            registerOutputs_10__14), .inputs_10__13 (registerOutputs_10__13), .inputs_10__12 (
            registerOutputs_10__12), .inputs_10__11 (registerOutputs_10__11), .inputs_10__10 (
            registerOutputs_10__10), .inputs_10__9 (registerOutputs_10__9), .inputs_10__8 (
            registerOutputs_10__8), .inputs_10__7 (registerOutputs_10__7), .inputs_10__6 (
            registerOutputs_10__6), .inputs_10__5 (registerOutputs_10__5), .inputs_10__4 (
            registerOutputs_10__4), .inputs_10__3 (registerOutputs_10__3), .inputs_10__2 (
            registerOutputs_10__2), .inputs_10__1 (registerOutputs_10__1), .inputs_10__0 (
            registerOutputs_10__0), .inputs_11__15 (registerOutputs_11__15), .inputs_11__14 (
            registerOutputs_11__14), .inputs_11__13 (registerOutputs_11__13), .inputs_11__12 (
            registerOutputs_11__12), .inputs_11__11 (registerOutputs_11__11), .inputs_11__10 (
            registerOutputs_11__10), .inputs_11__9 (registerOutputs_11__9), .inputs_11__8 (
            registerOutputs_11__8), .inputs_11__7 (registerOutputs_11__7), .inputs_11__6 (
            registerOutputs_11__6), .inputs_11__5 (registerOutputs_11__5), .inputs_11__4 (
            registerOutputs_11__4), .inputs_11__3 (registerOutputs_11__3), .inputs_11__2 (
            registerOutputs_11__2), .inputs_11__1 (registerOutputs_11__1), .inputs_11__0 (
            registerOutputs_11__0), .inputs_12__15 (registerOutputs_12__15), .inputs_12__14 (
            registerOutputs_12__14), .inputs_12__13 (registerOutputs_12__13), .inputs_12__12 (
            registerOutputs_12__12), .inputs_12__11 (registerOutputs_12__11), .inputs_12__10 (
            registerOutputs_12__10), .inputs_12__9 (registerOutputs_12__9), .inputs_12__8 (
            registerOutputs_12__8), .inputs_12__7 (registerOutputs_12__7), .inputs_12__6 (
            registerOutputs_12__6), .inputs_12__5 (registerOutputs_12__5), .inputs_12__4 (
            registerOutputs_12__4), .inputs_12__3 (registerOutputs_12__3), .inputs_12__2 (
            registerOutputs_12__2), .inputs_12__1 (registerOutputs_12__1), .inputs_12__0 (
            registerOutputs_12__0), .inputs_13__15 (registerOutputs_13__15), .inputs_13__14 (
            registerOutputs_13__14), .inputs_13__13 (registerOutputs_13__13), .inputs_13__12 (
            registerOutputs_13__12), .inputs_13__11 (registerOutputs_13__11), .inputs_13__10 (
            registerOutputs_13__10), .inputs_13__9 (registerOutputs_13__9), .inputs_13__8 (
            registerOutputs_13__8), .inputs_13__7 (registerOutputs_13__7), .inputs_13__6 (
            registerOutputs_13__6), .inputs_13__5 (registerOutputs_13__5), .inputs_13__4 (
            registerOutputs_13__4), .inputs_13__3 (registerOutputs_13__3), .inputs_13__2 (
            registerOutputs_13__2), .inputs_13__1 (registerOutputs_13__1), .inputs_13__0 (
            registerOutputs_13__0), .inputs_14__15 (registerOutputs_14__15), .inputs_14__14 (
            registerOutputs_14__14), .inputs_14__13 (registerOutputs_14__13), .inputs_14__12 (
            registerOutputs_14__12), .inputs_14__11 (registerOutputs_14__11), .inputs_14__10 (
            registerOutputs_14__10), .inputs_14__9 (registerOutputs_14__9), .inputs_14__8 (
            registerOutputs_14__8), .inputs_14__7 (registerOutputs_14__7), .inputs_14__6 (
            registerOutputs_14__6), .inputs_14__5 (registerOutputs_14__5), .inputs_14__4 (
            registerOutputs_14__4), .inputs_14__3 (registerOutputs_14__3), .inputs_14__2 (
            registerOutputs_14__2), .inputs_14__1 (registerOutputs_14__1), .inputs_14__0 (
            registerOutputs_14__0), .inputs_15__15 (registerOutputs_15__15), .inputs_15__14 (
            registerOutputs_15__14), .inputs_15__13 (registerOutputs_15__13), .inputs_15__12 (
            registerOutputs_15__12), .inputs_15__11 (registerOutputs_15__11), .inputs_15__10 (
            registerOutputs_15__10), .inputs_15__9 (registerOutputs_15__9), .inputs_15__8 (
            registerOutputs_15__8), .inputs_15__7 (registerOutputs_15__7), .inputs_15__6 (
            registerOutputs_15__6), .inputs_15__5 (registerOutputs_15__5), .inputs_15__4 (
            registerOutputs_15__4), .inputs_15__3 (registerOutputs_15__3), .inputs_15__2 (
            registerOutputs_15__2), .inputs_15__1 (registerOutputs_15__1), .inputs_15__0 (
            registerOutputs_15__0), .inputs_16__15 (registerOutputs_16__15), .inputs_16__14 (
            registerOutputs_16__14), .inputs_16__13 (registerOutputs_16__13), .inputs_16__12 (
            registerOutputs_16__12), .inputs_16__11 (registerOutputs_16__11), .inputs_16__10 (
            registerOutputs_16__10), .inputs_16__9 (registerOutputs_16__9), .inputs_16__8 (
            registerOutputs_16__8), .inputs_16__7 (registerOutputs_16__7), .inputs_16__6 (
            registerOutputs_16__6), .inputs_16__5 (registerOutputs_16__5), .inputs_16__4 (
            registerOutputs_16__4), .inputs_16__3 (registerOutputs_16__3), .inputs_16__2 (
            registerOutputs_16__2), .inputs_16__1 (registerOutputs_16__1), .inputs_16__0 (
            registerOutputs_16__0), .inputs_17__15 (registerOutputs_17__15), .inputs_17__14 (
            registerOutputs_17__14), .inputs_17__13 (registerOutputs_17__13), .inputs_17__12 (
            registerOutputs_17__12), .inputs_17__11 (registerOutputs_17__11), .inputs_17__10 (
            registerOutputs_17__10), .inputs_17__9 (registerOutputs_17__9), .inputs_17__8 (
            registerOutputs_17__8), .inputs_17__7 (registerOutputs_17__7), .inputs_17__6 (
            registerOutputs_17__6), .inputs_17__5 (registerOutputs_17__5), .inputs_17__4 (
            registerOutputs_17__4), .inputs_17__3 (registerOutputs_17__3), .inputs_17__2 (
            registerOutputs_17__2), .inputs_17__1 (registerOutputs_17__1), .inputs_17__0 (
            registerOutputs_17__0), .inputs_18__15 (registerOutputs_18__15), .inputs_18__14 (
            registerOutputs_18__14), .inputs_18__13 (registerOutputs_18__13), .inputs_18__12 (
            registerOutputs_18__12), .inputs_18__11 (registerOutputs_18__11), .inputs_18__10 (
            registerOutputs_18__10), .inputs_18__9 (registerOutputs_18__9), .inputs_18__8 (
            registerOutputs_18__8), .inputs_18__7 (registerOutputs_18__7), .inputs_18__6 (
            registerOutputs_18__6), .inputs_18__5 (registerOutputs_18__5), .inputs_18__4 (
            registerOutputs_18__4), .inputs_18__3 (registerOutputs_18__3), .inputs_18__2 (
            registerOutputs_18__2), .inputs_18__1 (registerOutputs_18__1), .inputs_18__0 (
            registerOutputs_18__0), .inputs_19__15 (registerOutputs_19__15), .inputs_19__14 (
            registerOutputs_19__14), .inputs_19__13 (registerOutputs_19__13), .inputs_19__12 (
            registerOutputs_19__12), .inputs_19__11 (registerOutputs_19__11), .inputs_19__10 (
            registerOutputs_19__10), .inputs_19__9 (registerOutputs_19__9), .inputs_19__8 (
            registerOutputs_19__8), .inputs_19__7 (registerOutputs_19__7), .inputs_19__6 (
            registerOutputs_19__6), .inputs_19__5 (registerOutputs_19__5), .inputs_19__4 (
            registerOutputs_19__4), .inputs_19__3 (registerOutputs_19__3), .inputs_19__2 (
            registerOutputs_19__2), .inputs_19__1 (registerOutputs_19__1), .inputs_19__0 (
            registerOutputs_19__0), .inputs_20__15 (registerOutputs_20__15), .inputs_20__14 (
            registerOutputs_20__14), .inputs_20__13 (registerOutputs_20__13), .inputs_20__12 (
            registerOutputs_20__12), .inputs_20__11 (registerOutputs_20__11), .inputs_20__10 (
            registerOutputs_20__10), .inputs_20__9 (registerOutputs_20__9), .inputs_20__8 (
            registerOutputs_20__8), .inputs_20__7 (registerOutputs_20__7), .inputs_20__6 (
            registerOutputs_20__6), .inputs_20__5 (registerOutputs_20__5), .inputs_20__4 (
            registerOutputs_20__4), .inputs_20__3 (registerOutputs_20__3), .inputs_20__2 (
            registerOutputs_20__2), .inputs_20__1 (registerOutputs_20__1), .inputs_20__0 (
            registerOutputs_20__0), .inputs_21__15 (registerOutputs_21__15), .inputs_21__14 (
            registerOutputs_21__14), .inputs_21__13 (registerOutputs_21__13), .inputs_21__12 (
            registerOutputs_21__12), .inputs_21__11 (registerOutputs_21__11), .inputs_21__10 (
            registerOutputs_21__10), .inputs_21__9 (registerOutputs_21__9), .inputs_21__8 (
            registerOutputs_21__8), .inputs_21__7 (registerOutputs_21__7), .inputs_21__6 (
            registerOutputs_21__6), .inputs_21__5 (registerOutputs_21__5), .inputs_21__4 (
            registerOutputs_21__4), .inputs_21__3 (registerOutputs_21__3), .inputs_21__2 (
            registerOutputs_21__2), .inputs_21__1 (registerOutputs_21__1), .inputs_21__0 (
            registerOutputs_21__0), .inputs_22__15 (registerOutputs_22__15), .inputs_22__14 (
            registerOutputs_22__14), .inputs_22__13 (registerOutputs_22__13), .inputs_22__12 (
            registerOutputs_22__12), .inputs_22__11 (registerOutputs_22__11), .inputs_22__10 (
            registerOutputs_22__10), .inputs_22__9 (registerOutputs_22__9), .inputs_22__8 (
            registerOutputs_22__8), .inputs_22__7 (registerOutputs_22__7), .inputs_22__6 (
            registerOutputs_22__6), .inputs_22__5 (registerOutputs_22__5), .inputs_22__4 (
            registerOutputs_22__4), .inputs_22__3 (registerOutputs_22__3), .inputs_22__2 (
            registerOutputs_22__2), .inputs_22__1 (registerOutputs_22__1), .inputs_22__0 (
            registerOutputs_22__0), .inputs_23__15 (registerOutputs_23__15), .inputs_23__14 (
            registerOutputs_23__14), .inputs_23__13 (registerOutputs_23__13), .inputs_23__12 (
            registerOutputs_23__12), .inputs_23__11 (registerOutputs_23__11), .inputs_23__10 (
            registerOutputs_23__10), .inputs_23__9 (registerOutputs_23__9), .inputs_23__8 (
            registerOutputs_23__8), .inputs_23__7 (registerOutputs_23__7), .inputs_23__6 (
            registerOutputs_23__6), .inputs_23__5 (registerOutputs_23__5), .inputs_23__4 (
            registerOutputs_23__4), .inputs_23__3 (registerOutputs_23__3), .inputs_23__2 (
            registerOutputs_23__2), .inputs_23__1 (registerOutputs_23__1), .inputs_23__0 (
            registerOutputs_23__0), .inputs_24__15 (registerOutputs_24__15), .inputs_24__14 (
            registerOutputs_24__14), .inputs_24__13 (registerOutputs_24__13), .inputs_24__12 (
            registerOutputs_24__12), .inputs_24__11 (registerOutputs_24__11), .inputs_24__10 (
            registerOutputs_24__10), .inputs_24__9 (registerOutputs_24__9), .inputs_24__8 (
            registerOutputs_24__8), .inputs_24__7 (registerOutputs_24__7), .inputs_24__6 (
            registerOutputs_24__6), .inputs_24__5 (registerOutputs_24__5), .inputs_24__4 (
            registerOutputs_24__4), .inputs_24__3 (registerOutputs_24__3), .inputs_24__2 (
            registerOutputs_24__2), .inputs_24__1 (registerOutputs_24__1), .inputs_24__0 (
            registerOutputs_24__0), .inputs_25__15 (registerOutputs_25__15), .inputs_25__14 (
            registerOutputs_25__14), .inputs_25__13 (registerOutputs_25__13), .inputs_25__12 (
            registerOutputs_25__12), .inputs_25__11 (registerOutputs_25__11), .inputs_25__10 (
            registerOutputs_25__10), .inputs_25__9 (registerOutputs_25__9), .inputs_25__8 (
            registerOutputs_25__8), .inputs_25__7 (registerOutputs_25__7), .inputs_25__6 (
            registerOutputs_25__6), .inputs_25__5 (registerOutputs_25__5), .inputs_25__4 (
            registerOutputs_25__4), .inputs_25__3 (registerOutputs_25__3), .inputs_25__2 (
            registerOutputs_25__2), .inputs_25__1 (registerOutputs_25__1), .inputs_25__0 (
            registerOutputs_25__0), .inputs_26__15 (registerOutputs_26__15), .inputs_26__14 (
            registerOutputs_26__14), .inputs_26__13 (registerOutputs_26__13), .inputs_26__12 (
            registerOutputs_26__12), .inputs_26__11 (registerOutputs_26__11), .inputs_26__10 (
            registerOutputs_26__10), .inputs_26__9 (registerOutputs_26__9), .inputs_26__8 (
            registerOutputs_26__8), .inputs_26__7 (registerOutputs_26__7), .inputs_26__6 (
            registerOutputs_26__6), .inputs_26__5 (registerOutputs_26__5), .inputs_26__4 (
            registerOutputs_26__4), .inputs_26__3 (registerOutputs_26__3), .inputs_26__2 (
            registerOutputs_26__2), .inputs_26__1 (registerOutputs_26__1), .inputs_26__0 (
            registerOutputs_26__0), .inputs_27__15 (registerOutputs_27__15), .inputs_27__14 (
            registerOutputs_27__14), .inputs_27__13 (registerOutputs_27__13), .inputs_27__12 (
            registerOutputs_27__12), .inputs_27__11 (registerOutputs_27__11), .inputs_27__10 (
            registerOutputs_27__10), .inputs_27__9 (registerOutputs_27__9), .inputs_27__8 (
            registerOutputs_27__8), .inputs_27__7 (registerOutputs_27__7), .inputs_27__6 (
            registerOutputs_27__6), .inputs_27__5 (registerOutputs_27__5), .inputs_27__4 (
            registerOutputs_27__4), .inputs_27__3 (registerOutputs_27__3), .inputs_27__2 (
            registerOutputs_27__2), .inputs_27__1 (registerOutputs_27__1), .inputs_27__0 (
            registerOutputs_27__0), .inputs_28__15 (registerOutputs_28__15), .inputs_28__14 (
            registerOutputs_28__14), .inputs_28__13 (registerOutputs_28__13), .inputs_28__12 (
            registerOutputs_28__12), .inputs_28__11 (registerOutputs_28__11), .inputs_28__10 (
            registerOutputs_28__10), .inputs_28__9 (registerOutputs_28__9), .inputs_28__8 (
            registerOutputs_28__8), .inputs_28__7 (registerOutputs_28__7), .inputs_28__6 (
            registerOutputs_28__6), .inputs_28__5 (registerOutputs_28__5), .inputs_28__4 (
            registerOutputs_28__4), .inputs_28__3 (registerOutputs_28__3), .inputs_28__2 (
            registerOutputs_28__2), .inputs_28__1 (registerOutputs_28__1), .inputs_28__0 (
            registerOutputs_28__0), .inputs_29__15 (registerOutputs_29__15), .inputs_29__14 (
            registerOutputs_29__14), .inputs_29__13 (registerOutputs_29__13), .inputs_29__12 (
            registerOutputs_29__12), .inputs_29__11 (registerOutputs_29__11), .inputs_29__10 (
            registerOutputs_29__10), .inputs_29__9 (registerOutputs_29__9), .inputs_29__8 (
            registerOutputs_29__8), .inputs_29__7 (registerOutputs_29__7), .inputs_29__6 (
            registerOutputs_29__6), .inputs_29__5 (registerOutputs_29__5), .inputs_29__4 (
            registerOutputs_29__4), .inputs_29__3 (registerOutputs_29__3), .inputs_29__2 (
            registerOutputs_29__2), .inputs_29__1 (registerOutputs_29__1), .inputs_29__0 (
            registerOutputs_29__0), .inputs_30__15 (registerOutputs_30__15), .inputs_30__14 (
            registerOutputs_30__14), .inputs_30__13 (registerOutputs_30__13), .inputs_30__12 (
            registerOutputs_30__12), .inputs_30__11 (registerOutputs_30__11), .inputs_30__10 (
            registerOutputs_30__10), .inputs_30__9 (registerOutputs_30__9), .inputs_30__8 (
            registerOutputs_30__8), .inputs_30__7 (registerOutputs_30__7), .inputs_30__6 (
            registerOutputs_30__6), .inputs_30__5 (registerOutputs_30__5), .inputs_30__4 (
            registerOutputs_30__4), .inputs_30__3 (registerOutputs_30__3), .inputs_30__2 (
            registerOutputs_30__2), .inputs_30__1 (registerOutputs_30__1), .inputs_30__0 (
            registerOutputs_30__0), .inputs_31__15 (registerOutputs_31__15), .inputs_31__14 (
            registerOutputs_31__14), .inputs_31__13 (registerOutputs_31__13), .inputs_31__12 (
            registerOutputs_31__12), .inputs_31__11 (registerOutputs_31__11), .inputs_31__10 (
            registerOutputs_31__10), .inputs_31__9 (registerOutputs_31__9), .inputs_31__8 (
            registerOutputs_31__8), .inputs_31__7 (registerOutputs_31__7), .inputs_31__6 (
            registerOutputs_31__6), .inputs_31__5 (registerOutputs_31__5), .inputs_31__4 (
            registerOutputs_31__4), .inputs_31__3 (registerOutputs_31__3), .inputs_31__2 (
            registerOutputs_31__2), .inputs_31__1 (registerOutputs_31__1), .inputs_31__0 (
            registerOutputs_31__0), .inputs_32__15 (registerOutputs_32__15), .inputs_32__14 (
            registerOutputs_32__14), .inputs_32__13 (registerOutputs_32__13), .inputs_32__12 (
            registerOutputs_32__12), .inputs_32__11 (registerOutputs_32__11), .inputs_32__10 (
            registerOutputs_32__10), .inputs_32__9 (registerOutputs_32__9), .inputs_32__8 (
            registerOutputs_32__8), .inputs_32__7 (registerOutputs_32__7), .inputs_32__6 (
            registerOutputs_32__6), .inputs_32__5 (registerOutputs_32__5), .inputs_32__4 (
            registerOutputs_32__4), .inputs_32__3 (registerOutputs_32__3), .inputs_32__2 (
            registerOutputs_32__2), .inputs_32__1 (registerOutputs_32__1), .inputs_32__0 (
            registerOutputs_32__0), .inputs_33__15 (registerOutputs_33__15), .inputs_33__14 (
            registerOutputs_33__14), .inputs_33__13 (registerOutputs_33__13), .inputs_33__12 (
            registerOutputs_33__12), .inputs_33__11 (registerOutputs_33__11), .inputs_33__10 (
            registerOutputs_33__10), .inputs_33__9 (registerOutputs_33__9), .inputs_33__8 (
            registerOutputs_33__8), .inputs_33__7 (registerOutputs_33__7), .inputs_33__6 (
            registerOutputs_33__6), .inputs_33__5 (registerOutputs_33__5), .inputs_33__4 (
            registerOutputs_33__4), .inputs_33__3 (registerOutputs_33__3), .inputs_33__2 (
            registerOutputs_33__2), .inputs_33__1 (registerOutputs_33__1), .inputs_33__0 (
            registerOutputs_33__0), .inputs_34__15 (registerOutputs_34__15), .inputs_34__14 (
            registerOutputs_34__14), .inputs_34__13 (registerOutputs_34__13), .inputs_34__12 (
            registerOutputs_34__12), .inputs_34__11 (registerOutputs_34__11), .inputs_34__10 (
            registerOutputs_34__10), .inputs_34__9 (registerOutputs_34__9), .inputs_34__8 (
            registerOutputs_34__8), .inputs_34__7 (registerOutputs_34__7), .inputs_34__6 (
            registerOutputs_34__6), .inputs_34__5 (registerOutputs_34__5), .inputs_34__4 (
            registerOutputs_34__4), .inputs_34__3 (registerOutputs_34__3), .inputs_34__2 (
            registerOutputs_34__2), .inputs_34__1 (registerOutputs_34__1), .inputs_34__0 (
            registerOutputs_34__0), .inputs_35__15 (registerOutputs_35__15), .inputs_35__14 (
            registerOutputs_35__14), .inputs_35__13 (registerOutputs_35__13), .inputs_35__12 (
            registerOutputs_35__12), .inputs_35__11 (registerOutputs_35__11), .inputs_35__10 (
            registerOutputs_35__10), .inputs_35__9 (registerOutputs_35__9), .inputs_35__8 (
            registerOutputs_35__8), .inputs_35__7 (registerOutputs_35__7), .inputs_35__6 (
            registerOutputs_35__6), .inputs_35__5 (registerOutputs_35__5), .inputs_35__4 (
            registerOutputs_35__4), .inputs_35__3 (registerOutputs_35__3), .inputs_35__2 (
            registerOutputs_35__2), .inputs_35__1 (registerOutputs_35__1), .inputs_35__0 (
            registerOutputs_35__0), .inputs_36__15 (registerOutputs_36__15), .inputs_36__14 (
            registerOutputs_36__14), .inputs_36__13 (registerOutputs_36__13), .inputs_36__12 (
            registerOutputs_36__12), .inputs_36__11 (registerOutputs_36__11), .inputs_36__10 (
            registerOutputs_36__10), .inputs_36__9 (registerOutputs_36__9), .inputs_36__8 (
            registerOutputs_36__8), .inputs_36__7 (registerOutputs_36__7), .inputs_36__6 (
            registerOutputs_36__6), .inputs_36__5 (registerOutputs_36__5), .inputs_36__4 (
            registerOutputs_36__4), .inputs_36__3 (registerOutputs_36__3), .inputs_36__2 (
            registerOutputs_36__2), .inputs_36__1 (registerOutputs_36__1), .inputs_36__0 (
            registerOutputs_36__0), .inputs_37__15 (registerOutputs_37__15), .inputs_37__14 (
            registerOutputs_37__14), .inputs_37__13 (registerOutputs_37__13), .inputs_37__12 (
            registerOutputs_37__12), .inputs_37__11 (registerOutputs_37__11), .inputs_37__10 (
            registerOutputs_37__10), .inputs_37__9 (registerOutputs_37__9), .inputs_37__8 (
            registerOutputs_37__8), .inputs_37__7 (registerOutputs_37__7), .inputs_37__6 (
            registerOutputs_37__6), .inputs_37__5 (registerOutputs_37__5), .inputs_37__4 (
            registerOutputs_37__4), .inputs_37__3 (registerOutputs_37__3), .inputs_37__2 (
            registerOutputs_37__2), .inputs_37__1 (registerOutputs_37__1), .inputs_37__0 (
            registerOutputs_37__0), .inputs_38__15 (registerOutputs_38__15), .inputs_38__14 (
            registerOutputs_38__14), .inputs_38__13 (registerOutputs_38__13), .inputs_38__12 (
            registerOutputs_38__12), .inputs_38__11 (registerOutputs_38__11), .inputs_38__10 (
            registerOutputs_38__10), .inputs_38__9 (registerOutputs_38__9), .inputs_38__8 (
            registerOutputs_38__8), .inputs_38__7 (registerOutputs_38__7), .inputs_38__6 (
            registerOutputs_38__6), .inputs_38__5 (registerOutputs_38__5), .inputs_38__4 (
            registerOutputs_38__4), .inputs_38__3 (registerOutputs_38__3), .inputs_38__2 (
            registerOutputs_38__2), .inputs_38__1 (registerOutputs_38__1), .inputs_38__0 (
            registerOutputs_38__0), .inputs_39__15 (registerOutputs_39__15), .inputs_39__14 (
            registerOutputs_39__14), .inputs_39__13 (registerOutputs_39__13), .inputs_39__12 (
            registerOutputs_39__12), .inputs_39__11 (registerOutputs_39__11), .inputs_39__10 (
            registerOutputs_39__10), .inputs_39__9 (registerOutputs_39__9), .inputs_39__8 (
            registerOutputs_39__8), .inputs_39__7 (registerOutputs_39__7), .inputs_39__6 (
            registerOutputs_39__6), .inputs_39__5 (registerOutputs_39__5), .inputs_39__4 (
            registerOutputs_39__4), .inputs_39__3 (registerOutputs_39__3), .inputs_39__2 (
            registerOutputs_39__2), .inputs_39__1 (registerOutputs_39__1), .inputs_39__0 (
            registerOutputs_39__0), .inputs_40__15 (registerOutputs_40__15), .inputs_40__14 (
            registerOutputs_40__14), .inputs_40__13 (registerOutputs_40__13), .inputs_40__12 (
            registerOutputs_40__12), .inputs_40__11 (registerOutputs_40__11), .inputs_40__10 (
            registerOutputs_40__10), .inputs_40__9 (registerOutputs_40__9), .inputs_40__8 (
            registerOutputs_40__8), .inputs_40__7 (registerOutputs_40__7), .inputs_40__6 (
            registerOutputs_40__6), .inputs_40__5 (registerOutputs_40__5), .inputs_40__4 (
            registerOutputs_40__4), .inputs_40__3 (registerOutputs_40__3), .inputs_40__2 (
            registerOutputs_40__2), .inputs_40__1 (registerOutputs_40__1), .inputs_40__0 (
            registerOutputs_40__0), .inputs_41__15 (registerOutputs_41__15), .inputs_41__14 (
            registerOutputs_41__14), .inputs_41__13 (registerOutputs_41__13), .inputs_41__12 (
            registerOutputs_41__12), .inputs_41__11 (registerOutputs_41__11), .inputs_41__10 (
            registerOutputs_41__10), .inputs_41__9 (registerOutputs_41__9), .inputs_41__8 (
            registerOutputs_41__8), .inputs_41__7 (registerOutputs_41__7), .inputs_41__6 (
            registerOutputs_41__6), .inputs_41__5 (registerOutputs_41__5), .inputs_41__4 (
            registerOutputs_41__4), .inputs_41__3 (registerOutputs_41__3), .inputs_41__2 (
            registerOutputs_41__2), .inputs_41__1 (registerOutputs_41__1), .inputs_41__0 (
            registerOutputs_41__0), .inputs_42__15 (registerOutputs_42__15), .inputs_42__14 (
            registerOutputs_42__14), .inputs_42__13 (registerOutputs_42__13), .inputs_42__12 (
            registerOutputs_42__12), .inputs_42__11 (registerOutputs_42__11), .inputs_42__10 (
            registerOutputs_42__10), .inputs_42__9 (registerOutputs_42__9), .inputs_42__8 (
            registerOutputs_42__8), .inputs_42__7 (registerOutputs_42__7), .inputs_42__6 (
            registerOutputs_42__6), .inputs_42__5 (registerOutputs_42__5), .inputs_42__4 (
            registerOutputs_42__4), .inputs_42__3 (registerOutputs_42__3), .inputs_42__2 (
            registerOutputs_42__2), .inputs_42__1 (registerOutputs_42__1), .inputs_42__0 (
            registerOutputs_42__0), .inputs_43__15 (registerOutputs_43__15), .inputs_43__14 (
            registerOutputs_43__14), .inputs_43__13 (registerOutputs_43__13), .inputs_43__12 (
            registerOutputs_43__12), .inputs_43__11 (registerOutputs_43__11), .inputs_43__10 (
            registerOutputs_43__10), .inputs_43__9 (registerOutputs_43__9), .inputs_43__8 (
            registerOutputs_43__8), .inputs_43__7 (registerOutputs_43__7), .inputs_43__6 (
            registerOutputs_43__6), .inputs_43__5 (registerOutputs_43__5), .inputs_43__4 (
            registerOutputs_43__4), .inputs_43__3 (registerOutputs_43__3), .inputs_43__2 (
            registerOutputs_43__2), .inputs_43__1 (registerOutputs_43__1), .inputs_43__0 (
            registerOutputs_43__0), .inputs_44__15 (registerOutputs_44__15), .inputs_44__14 (
            registerOutputs_44__14), .inputs_44__13 (registerOutputs_44__13), .inputs_44__12 (
            registerOutputs_44__12), .inputs_44__11 (registerOutputs_44__11), .inputs_44__10 (
            registerOutputs_44__10), .inputs_44__9 (registerOutputs_44__9), .inputs_44__8 (
            registerOutputs_44__8), .inputs_44__7 (registerOutputs_44__7), .inputs_44__6 (
            registerOutputs_44__6), .inputs_44__5 (registerOutputs_44__5), .inputs_44__4 (
            registerOutputs_44__4), .inputs_44__3 (registerOutputs_44__3), .inputs_44__2 (
            registerOutputs_44__2), .inputs_44__1 (registerOutputs_44__1), .inputs_44__0 (
            registerOutputs_44__0), .inputs_45__15 (registerOutputs_45__15), .inputs_45__14 (
            registerOutputs_45__14), .inputs_45__13 (registerOutputs_45__13), .inputs_45__12 (
            registerOutputs_45__12), .inputs_45__11 (registerOutputs_45__11), .inputs_45__10 (
            registerOutputs_45__10), .inputs_45__9 (registerOutputs_45__9), .inputs_45__8 (
            registerOutputs_45__8), .inputs_45__7 (registerOutputs_45__7), .inputs_45__6 (
            registerOutputs_45__6), .inputs_45__5 (registerOutputs_45__5), .inputs_45__4 (
            registerOutputs_45__4), .inputs_45__3 (registerOutputs_45__3), .inputs_45__2 (
            registerOutputs_45__2), .inputs_45__1 (registerOutputs_45__1), .inputs_45__0 (
            registerOutputs_45__0), .inputs_46__15 (registerOutputs_46__15), .inputs_46__14 (
            registerOutputs_46__14), .inputs_46__13 (registerOutputs_46__13), .inputs_46__12 (
            registerOutputs_46__12), .inputs_46__11 (registerOutputs_46__11), .inputs_46__10 (
            registerOutputs_46__10), .inputs_46__9 (registerOutputs_46__9), .inputs_46__8 (
            registerOutputs_46__8), .inputs_46__7 (registerOutputs_46__7), .inputs_46__6 (
            registerOutputs_46__6), .inputs_46__5 (registerOutputs_46__5), .inputs_46__4 (
            registerOutputs_46__4), .inputs_46__3 (registerOutputs_46__3), .inputs_46__2 (
            registerOutputs_46__2), .inputs_46__1 (registerOutputs_46__1), .inputs_46__0 (
            registerOutputs_46__0), .inputs_47__15 (registerOutputs_47__15), .inputs_47__14 (
            registerOutputs_47__14), .inputs_47__13 (registerOutputs_47__13), .inputs_47__12 (
            registerOutputs_47__12), .inputs_47__11 (registerOutputs_47__11), .inputs_47__10 (
            registerOutputs_47__10), .inputs_47__9 (registerOutputs_47__9), .inputs_47__8 (
            registerOutputs_47__8), .inputs_47__7 (registerOutputs_47__7), .inputs_47__6 (
            registerOutputs_47__6), .inputs_47__5 (registerOutputs_47__5), .inputs_47__4 (
            registerOutputs_47__4), .inputs_47__3 (registerOutputs_47__3), .inputs_47__2 (
            registerOutputs_47__2), .inputs_47__1 (registerOutputs_47__1), .inputs_47__0 (
            registerOutputs_47__0), .inputs_48__15 (registerOutputs_48__15), .inputs_48__14 (
            registerOutputs_48__14), .inputs_48__13 (registerOutputs_48__13), .inputs_48__12 (
            registerOutputs_48__12), .inputs_48__11 (registerOutputs_48__11), .inputs_48__10 (
            registerOutputs_48__10), .inputs_48__9 (registerOutputs_48__9), .inputs_48__8 (
            registerOutputs_48__8), .inputs_48__7 (registerOutputs_48__7), .inputs_48__6 (
            registerOutputs_48__6), .inputs_48__5 (registerOutputs_48__5), .inputs_48__4 (
            registerOutputs_48__4), .inputs_48__3 (registerOutputs_48__3), .inputs_48__2 (
            registerOutputs_48__2), .inputs_48__1 (registerOutputs_48__1), .inputs_48__0 (
            registerOutputs_48__0), .inputs_49__15 (registerOutputs_49__15), .inputs_49__14 (
            registerOutputs_49__14), .inputs_49__13 (registerOutputs_49__13), .inputs_49__12 (
            registerOutputs_49__12), .inputs_49__11 (registerOutputs_49__11), .inputs_49__10 (
            registerOutputs_49__10), .inputs_49__9 (registerOutputs_49__9), .inputs_49__8 (
            registerOutputs_49__8), .inputs_49__7 (registerOutputs_49__7), .inputs_49__6 (
            registerOutputs_49__6), .inputs_49__5 (registerOutputs_49__5), .inputs_49__4 (
            registerOutputs_49__4), .inputs_49__3 (registerOutputs_49__3), .inputs_49__2 (
            registerOutputs_49__2), .inputs_49__1 (registerOutputs_49__1), .inputs_49__0 (
            registerOutputs_49__0), .inputs_50__15 (registerOutputs_50__15), .inputs_50__14 (
            registerOutputs_50__14), .inputs_50__13 (registerOutputs_50__13), .inputs_50__12 (
            registerOutputs_50__12), .inputs_50__11 (registerOutputs_50__11), .inputs_50__10 (
            registerOutputs_50__10), .inputs_50__9 (registerOutputs_50__9), .inputs_50__8 (
            registerOutputs_50__8), .inputs_50__7 (registerOutputs_50__7), .inputs_50__6 (
            registerOutputs_50__6), .inputs_50__5 (registerOutputs_50__5), .inputs_50__4 (
            registerOutputs_50__4), .inputs_50__3 (registerOutputs_50__3), .inputs_50__2 (
            registerOutputs_50__2), .inputs_50__1 (registerOutputs_50__1), .inputs_50__0 (
            registerOutputs_50__0), .inputs_51__15 (registerOutputs_51__15), .inputs_51__14 (
            registerOutputs_51__14), .inputs_51__13 (registerOutputs_51__13), .inputs_51__12 (
            registerOutputs_51__12), .inputs_51__11 (registerOutputs_51__11), .inputs_51__10 (
            registerOutputs_51__10), .inputs_51__9 (registerOutputs_51__9), .inputs_51__8 (
            registerOutputs_51__8), .inputs_51__7 (registerOutputs_51__7), .inputs_51__6 (
            registerOutputs_51__6), .inputs_51__5 (registerOutputs_51__5), .inputs_51__4 (
            registerOutputs_51__4), .inputs_51__3 (registerOutputs_51__3), .inputs_51__2 (
            registerOutputs_51__2), .inputs_51__1 (registerOutputs_51__1), .inputs_51__0 (
            registerOutputs_51__0), .inputs_52__15 (registerOutputs_52__15), .inputs_52__14 (
            registerOutputs_52__14), .inputs_52__13 (registerOutputs_52__13), .inputs_52__12 (
            registerOutputs_52__12), .inputs_52__11 (registerOutputs_52__11), .inputs_52__10 (
            registerOutputs_52__10), .inputs_52__9 (registerOutputs_52__9), .inputs_52__8 (
            registerOutputs_52__8), .inputs_52__7 (registerOutputs_52__7), .inputs_52__6 (
            registerOutputs_52__6), .inputs_52__5 (registerOutputs_52__5), .inputs_52__4 (
            registerOutputs_52__4), .inputs_52__3 (registerOutputs_52__3), .inputs_52__2 (
            registerOutputs_52__2), .inputs_52__1 (registerOutputs_52__1), .inputs_52__0 (
            registerOutputs_52__0), .inputs_53__15 (registerOutputs_53__15), .inputs_53__14 (
            registerOutputs_53__14), .inputs_53__13 (registerOutputs_53__13), .inputs_53__12 (
            registerOutputs_53__12), .inputs_53__11 (registerOutputs_53__11), .inputs_53__10 (
            registerOutputs_53__10), .inputs_53__9 (registerOutputs_53__9), .inputs_53__8 (
            registerOutputs_53__8), .inputs_53__7 (registerOutputs_53__7), .inputs_53__6 (
            registerOutputs_53__6), .inputs_53__5 (registerOutputs_53__5), .inputs_53__4 (
            registerOutputs_53__4), .inputs_53__3 (registerOutputs_53__3), .inputs_53__2 (
            registerOutputs_53__2), .inputs_53__1 (registerOutputs_53__1), .inputs_53__0 (
            registerOutputs_53__0), .inputs_54__15 (registerOutputs_54__15), .inputs_54__14 (
            registerOutputs_54__14), .inputs_54__13 (registerOutputs_54__13), .inputs_54__12 (
            registerOutputs_54__12), .inputs_54__11 (registerOutputs_54__11), .inputs_54__10 (
            registerOutputs_54__10), .inputs_54__9 (registerOutputs_54__9), .inputs_54__8 (
            registerOutputs_54__8), .inputs_54__7 (registerOutputs_54__7), .inputs_54__6 (
            registerOutputs_54__6), .inputs_54__5 (registerOutputs_54__5), .inputs_54__4 (
            registerOutputs_54__4), .inputs_54__3 (registerOutputs_54__3), .inputs_54__2 (
            registerOutputs_54__2), .inputs_54__1 (registerOutputs_54__1), .inputs_54__0 (
            registerOutputs_54__0), .inputs_55__15 (registerOutputs_55__15), .inputs_55__14 (
            registerOutputs_55__14), .inputs_55__13 (registerOutputs_55__13), .inputs_55__12 (
            registerOutputs_55__12), .inputs_55__11 (registerOutputs_55__11), .inputs_55__10 (
            registerOutputs_55__10), .inputs_55__9 (registerOutputs_55__9), .inputs_55__8 (
            registerOutputs_55__8), .inputs_55__7 (registerOutputs_55__7), .inputs_55__6 (
            registerOutputs_55__6), .inputs_55__5 (registerOutputs_55__5), .inputs_55__4 (
            registerOutputs_55__4), .inputs_55__3 (registerOutputs_55__3), .inputs_55__2 (
            registerOutputs_55__2), .inputs_55__1 (registerOutputs_55__1), .inputs_55__0 (
            registerOutputs_55__0), .inputs_56__15 (registerOutputs_56__15), .inputs_56__14 (
            registerOutputs_56__14), .inputs_56__13 (registerOutputs_56__13), .inputs_56__12 (
            registerOutputs_56__12), .inputs_56__11 (registerOutputs_56__11), .inputs_56__10 (
            registerOutputs_56__10), .inputs_56__9 (registerOutputs_56__9), .inputs_56__8 (
            registerOutputs_56__8), .inputs_56__7 (registerOutputs_56__7), .inputs_56__6 (
            registerOutputs_56__6), .inputs_56__5 (registerOutputs_56__5), .inputs_56__4 (
            registerOutputs_56__4), .inputs_56__3 (registerOutputs_56__3), .inputs_56__2 (
            registerOutputs_56__2), .inputs_56__1 (registerOutputs_56__1), .inputs_56__0 (
            registerOutputs_56__0), .inputs_57__15 (registerOutputs_57__15), .inputs_57__14 (
            registerOutputs_57__14), .inputs_57__13 (registerOutputs_57__13), .inputs_57__12 (
            registerOutputs_57__12), .inputs_57__11 (registerOutputs_57__11), .inputs_57__10 (
            registerOutputs_57__10), .inputs_57__9 (registerOutputs_57__9), .inputs_57__8 (
            registerOutputs_57__8), .inputs_57__7 (registerOutputs_57__7), .inputs_57__6 (
            registerOutputs_57__6), .inputs_57__5 (registerOutputs_57__5), .inputs_57__4 (
            registerOutputs_57__4), .inputs_57__3 (registerOutputs_57__3), .inputs_57__2 (
            registerOutputs_57__2), .inputs_57__1 (registerOutputs_57__1), .inputs_57__0 (
            registerOutputs_57__0), .inputs_58__15 (registerOutputs_58__15), .inputs_58__14 (
            registerOutputs_58__14), .inputs_58__13 (registerOutputs_58__13), .inputs_58__12 (
            registerOutputs_58__12), .inputs_58__11 (registerOutputs_58__11), .inputs_58__10 (
            registerOutputs_58__10), .inputs_58__9 (registerOutputs_58__9), .inputs_58__8 (
            registerOutputs_58__8), .inputs_58__7 (registerOutputs_58__7), .inputs_58__6 (
            registerOutputs_58__6), .inputs_58__5 (registerOutputs_58__5), .inputs_58__4 (
            registerOutputs_58__4), .inputs_58__3 (registerOutputs_58__3), .inputs_58__2 (
            registerOutputs_58__2), .inputs_58__1 (registerOutputs_58__1), .inputs_58__0 (
            registerOutputs_58__0), .inputs_59__15 (registerOutputs_59__15), .inputs_59__14 (
            registerOutputs_59__14), .inputs_59__13 (registerOutputs_59__13), .inputs_59__12 (
            registerOutputs_59__12), .inputs_59__11 (registerOutputs_59__11), .inputs_59__10 (
            registerOutputs_59__10), .inputs_59__9 (registerOutputs_59__9), .inputs_59__8 (
            registerOutputs_59__8), .inputs_59__7 (registerOutputs_59__7), .inputs_59__6 (
            registerOutputs_59__6), .inputs_59__5 (registerOutputs_59__5), .inputs_59__4 (
            registerOutputs_59__4), .inputs_59__3 (registerOutputs_59__3), .inputs_59__2 (
            registerOutputs_59__2), .inputs_59__1 (registerOutputs_59__1), .inputs_59__0 (
            registerOutputs_59__0), .inputs_60__15 (registerOutputs_60__15), .inputs_60__14 (
            registerOutputs_60__14), .inputs_60__13 (registerOutputs_60__13), .inputs_60__12 (
            registerOutputs_60__12), .inputs_60__11 (registerOutputs_60__11), .inputs_60__10 (
            registerOutputs_60__10), .inputs_60__9 (registerOutputs_60__9), .inputs_60__8 (
            registerOutputs_60__8), .inputs_60__7 (registerOutputs_60__7), .inputs_60__6 (
            registerOutputs_60__6), .inputs_60__5 (registerOutputs_60__5), .inputs_60__4 (
            registerOutputs_60__4), .inputs_60__3 (registerOutputs_60__3), .inputs_60__2 (
            registerOutputs_60__2), .inputs_60__1 (registerOutputs_60__1), .inputs_60__0 (
            registerOutputs_60__0), .inputs_61__15 (registerOutputs_61__15), .inputs_61__14 (
            registerOutputs_61__14), .inputs_61__13 (registerOutputs_61__13), .inputs_61__12 (
            registerOutputs_61__12), .inputs_61__11 (registerOutputs_61__11), .inputs_61__10 (
            registerOutputs_61__10), .inputs_61__9 (registerOutputs_61__9), .inputs_61__8 (
            registerOutputs_61__8), .inputs_61__7 (registerOutputs_61__7), .inputs_61__6 (
            registerOutputs_61__6), .inputs_61__5 (registerOutputs_61__5), .inputs_61__4 (
            registerOutputs_61__4), .inputs_61__3 (registerOutputs_61__3), .inputs_61__2 (
            registerOutputs_61__2), .inputs_61__1 (registerOutputs_61__1), .inputs_61__0 (
            registerOutputs_61__0), .inputs_62__15 (registerOutputs_62__15), .inputs_62__14 (
            registerOutputs_62__14), .inputs_62__13 (registerOutputs_62__13), .inputs_62__12 (
            registerOutputs_62__12), .inputs_62__11 (registerOutputs_62__11), .inputs_62__10 (
            registerOutputs_62__10), .inputs_62__9 (registerOutputs_62__9), .inputs_62__8 (
            registerOutputs_62__8), .inputs_62__7 (registerOutputs_62__7), .inputs_62__6 (
            registerOutputs_62__6), .inputs_62__5 (registerOutputs_62__5), .inputs_62__4 (
            registerOutputs_62__4), .inputs_62__3 (registerOutputs_62__3), .inputs_62__2 (
            registerOutputs_62__2), .inputs_62__1 (registerOutputs_62__1), .inputs_62__0 (
            registerOutputs_62__0), .inputs_63__15 (registerOutputs_63__15), .inputs_63__14 (
            registerOutputs_63__14), .inputs_63__13 (registerOutputs_63__13), .inputs_63__12 (
            registerOutputs_63__12), .inputs_63__11 (registerOutputs_63__11), .inputs_63__10 (
            registerOutputs_63__10), .inputs_63__9 (registerOutputs_63__9), .inputs_63__8 (
            registerOutputs_63__8), .inputs_63__7 (registerOutputs_63__7), .inputs_63__6 (
            registerOutputs_63__6), .inputs_63__5 (registerOutputs_63__5), .inputs_63__4 (
            registerOutputs_63__4), .inputs_63__3 (registerOutputs_63__3), .inputs_63__2 (
            registerOutputs_63__2), .inputs_63__1 (registerOutputs_63__1), .inputs_63__0 (
            registerOutputs_63__0), .inputs_64__15 (registerOutputs_64__15), .inputs_64__14 (
            registerOutputs_64__14), .inputs_64__13 (registerOutputs_64__13), .inputs_64__12 (
            registerOutputs_64__12), .inputs_64__11 (registerOutputs_64__11), .inputs_64__10 (
            registerOutputs_64__10), .inputs_64__9 (registerOutputs_64__9), .inputs_64__8 (
            registerOutputs_64__8), .inputs_64__7 (registerOutputs_64__7), .inputs_64__6 (
            registerOutputs_64__6), .inputs_64__5 (registerOutputs_64__5), .inputs_64__4 (
            registerOutputs_64__4), .inputs_64__3 (registerOutputs_64__3), .inputs_64__2 (
            registerOutputs_64__2), .inputs_64__1 (registerOutputs_64__1), .inputs_64__0 (
            registerOutputs_64__0), .inputs_65__15 (registerOutputs_65__15), .inputs_65__14 (
            registerOutputs_65__14), .inputs_65__13 (registerOutputs_65__13), .inputs_65__12 (
            registerOutputs_65__12), .inputs_65__11 (registerOutputs_65__11), .inputs_65__10 (
            registerOutputs_65__10), .inputs_65__9 (registerOutputs_65__9), .inputs_65__8 (
            registerOutputs_65__8), .inputs_65__7 (registerOutputs_65__7), .inputs_65__6 (
            registerOutputs_65__6), .inputs_65__5 (registerOutputs_65__5), .inputs_65__4 (
            registerOutputs_65__4), .inputs_65__3 (registerOutputs_65__3), .inputs_65__2 (
            registerOutputs_65__2), .inputs_65__1 (registerOutputs_65__1), .inputs_65__0 (
            registerOutputs_65__0), .inputs_66__15 (registerOutputs_66__15), .inputs_66__14 (
            registerOutputs_66__14), .inputs_66__13 (registerOutputs_66__13), .inputs_66__12 (
            registerOutputs_66__12), .inputs_66__11 (registerOutputs_66__11), .inputs_66__10 (
            registerOutputs_66__10), .inputs_66__9 (registerOutputs_66__9), .inputs_66__8 (
            registerOutputs_66__8), .inputs_66__7 (registerOutputs_66__7), .inputs_66__6 (
            registerOutputs_66__6), .inputs_66__5 (registerOutputs_66__5), .inputs_66__4 (
            registerOutputs_66__4), .inputs_66__3 (registerOutputs_66__3), .inputs_66__2 (
            registerOutputs_66__2), .inputs_66__1 (registerOutputs_66__1), .inputs_66__0 (
            registerOutputs_66__0), .inputs_67__15 (registerOutputs_67__15), .inputs_67__14 (
            registerOutputs_67__14), .inputs_67__13 (registerOutputs_67__13), .inputs_67__12 (
            registerOutputs_67__12), .inputs_67__11 (registerOutputs_67__11), .inputs_67__10 (
            registerOutputs_67__10), .inputs_67__9 (registerOutputs_67__9), .inputs_67__8 (
            registerOutputs_67__8), .inputs_67__7 (registerOutputs_67__7), .inputs_67__6 (
            registerOutputs_67__6), .inputs_67__5 (registerOutputs_67__5), .inputs_67__4 (
            registerOutputs_67__4), .inputs_67__3 (registerOutputs_67__3), .inputs_67__2 (
            registerOutputs_67__2), .inputs_67__1 (registerOutputs_67__1), .inputs_67__0 (
            registerOutputs_67__0), .inputs_68__15 (registerOutputs_68__15), .inputs_68__14 (
            registerOutputs_68__14), .inputs_68__13 (registerOutputs_68__13), .inputs_68__12 (
            registerOutputs_68__12), .inputs_68__11 (registerOutputs_68__11), .inputs_68__10 (
            registerOutputs_68__10), .inputs_68__9 (registerOutputs_68__9), .inputs_68__8 (
            registerOutputs_68__8), .inputs_68__7 (registerOutputs_68__7), .inputs_68__6 (
            registerOutputs_68__6), .inputs_68__5 (registerOutputs_68__5), .inputs_68__4 (
            registerOutputs_68__4), .inputs_68__3 (registerOutputs_68__3), .inputs_68__2 (
            registerOutputs_68__2), .inputs_68__1 (registerOutputs_68__1), .inputs_68__0 (
            registerOutputs_68__0), .inputs_69__15 (registerOutputs_69__15), .inputs_69__14 (
            registerOutputs_69__14), .inputs_69__13 (registerOutputs_69__13), .inputs_69__12 (
            registerOutputs_69__12), .inputs_69__11 (registerOutputs_69__11), .inputs_69__10 (
            registerOutputs_69__10), .inputs_69__9 (registerOutputs_69__9), .inputs_69__8 (
            registerOutputs_69__8), .inputs_69__7 (registerOutputs_69__7), .inputs_69__6 (
            registerOutputs_69__6), .inputs_69__5 (registerOutputs_69__5), .inputs_69__4 (
            registerOutputs_69__4), .inputs_69__3 (registerOutputs_69__3), .inputs_69__2 (
            registerOutputs_69__2), .inputs_69__1 (registerOutputs_69__1), .inputs_69__0 (
            registerOutputs_69__0), .inputs_70__15 (registerOutputs_70__15), .inputs_70__14 (
            registerOutputs_70__14), .inputs_70__13 (registerOutputs_70__13), .inputs_70__12 (
            registerOutputs_70__12), .inputs_70__11 (registerOutputs_70__11), .inputs_70__10 (
            registerOutputs_70__10), .inputs_70__9 (registerOutputs_70__9), .inputs_70__8 (
            registerOutputs_70__8), .inputs_70__7 (registerOutputs_70__7), .inputs_70__6 (
            registerOutputs_70__6), .inputs_70__5 (registerOutputs_70__5), .inputs_70__4 (
            registerOutputs_70__4), .inputs_70__3 (registerOutputs_70__3), .inputs_70__2 (
            registerOutputs_70__2), .inputs_70__1 (registerOutputs_70__1), .inputs_70__0 (
            registerOutputs_70__0), .inputs_71__15 (registerOutputs_71__15), .inputs_71__14 (
            registerOutputs_71__14), .inputs_71__13 (registerOutputs_71__13), .inputs_71__12 (
            registerOutputs_71__12), .inputs_71__11 (registerOutputs_71__11), .inputs_71__10 (
            registerOutputs_71__10), .inputs_71__9 (registerOutputs_71__9), .inputs_71__8 (
            registerOutputs_71__8), .inputs_71__7 (registerOutputs_71__7), .inputs_71__6 (
            registerOutputs_71__6), .inputs_71__5 (registerOutputs_71__5), .inputs_71__4 (
            registerOutputs_71__4), .inputs_71__3 (registerOutputs_71__3), .inputs_71__2 (
            registerOutputs_71__2), .inputs_71__1 (registerOutputs_71__1), .inputs_71__0 (
            registerOutputs_71__0), .inputs_72__15 (registerOutputs_72__15), .inputs_72__14 (
            registerOutputs_72__14), .inputs_72__13 (registerOutputs_72__13), .inputs_72__12 (
            registerOutputs_72__12), .inputs_72__11 (registerOutputs_72__11), .inputs_72__10 (
            registerOutputs_72__10), .inputs_72__9 (registerOutputs_72__9), .inputs_72__8 (
            registerOutputs_72__8), .inputs_72__7 (registerOutputs_72__7), .inputs_72__6 (
            registerOutputs_72__6), .inputs_72__5 (registerOutputs_72__5), .inputs_72__4 (
            registerOutputs_72__4), .inputs_72__3 (registerOutputs_72__3), .inputs_72__2 (
            registerOutputs_72__2), .inputs_72__1 (registerOutputs_72__1), .inputs_72__0 (
            registerOutputs_72__0), .inputs_73__15 (registerOutputs_73__15), .inputs_73__14 (
            registerOutputs_73__14), .inputs_73__13 (registerOutputs_73__13), .inputs_73__12 (
            registerOutputs_73__12), .inputs_73__11 (registerOutputs_73__11), .inputs_73__10 (
            registerOutputs_73__10), .inputs_73__9 (registerOutputs_73__9), .inputs_73__8 (
            registerOutputs_73__8), .inputs_73__7 (registerOutputs_73__7), .inputs_73__6 (
            registerOutputs_73__6), .inputs_73__5 (registerOutputs_73__5), .inputs_73__4 (
            registerOutputs_73__4), .inputs_73__3 (registerOutputs_73__3), .inputs_73__2 (
            registerOutputs_73__2), .inputs_73__1 (registerOutputs_73__1), .inputs_73__0 (
            registerOutputs_73__0), .inputs_74__15 (registerOutputs_74__15), .inputs_74__14 (
            registerOutputs_74__14), .inputs_74__13 (registerOutputs_74__13), .inputs_74__12 (
            registerOutputs_74__12), .inputs_74__11 (registerOutputs_74__11), .inputs_74__10 (
            registerOutputs_74__10), .inputs_74__9 (registerOutputs_74__9), .inputs_74__8 (
            registerOutputs_74__8), .inputs_74__7 (registerOutputs_74__7), .inputs_74__6 (
            registerOutputs_74__6), .inputs_74__5 (registerOutputs_74__5), .inputs_74__4 (
            registerOutputs_74__4), .inputs_74__3 (registerOutputs_74__3), .inputs_74__2 (
            registerOutputs_74__2), .inputs_74__1 (registerOutputs_74__1), .inputs_74__0 (
            registerOutputs_74__0), .inputs_75__15 (registerOutputs_75__15), .inputs_75__14 (
            registerOutputs_75__14), .inputs_75__13 (registerOutputs_75__13), .inputs_75__12 (
            registerOutputs_75__12), .inputs_75__11 (registerOutputs_75__11), .inputs_75__10 (
            registerOutputs_75__10), .inputs_75__9 (registerOutputs_75__9), .inputs_75__8 (
            registerOutputs_75__8), .inputs_75__7 (registerOutputs_75__7), .inputs_75__6 (
            registerOutputs_75__6), .inputs_75__5 (registerOutputs_75__5), .inputs_75__4 (
            registerOutputs_75__4), .inputs_75__3 (registerOutputs_75__3), .inputs_75__2 (
            registerOutputs_75__2), .inputs_75__1 (registerOutputs_75__1), .inputs_75__0 (
            registerOutputs_75__0), .inputs_76__15 (registerOutputs_76__15), .inputs_76__14 (
            registerOutputs_76__14), .inputs_76__13 (registerOutputs_76__13), .inputs_76__12 (
            registerOutputs_76__12), .inputs_76__11 (registerOutputs_76__11), .inputs_76__10 (
            registerOutputs_76__10), .inputs_76__9 (registerOutputs_76__9), .inputs_76__8 (
            registerOutputs_76__8), .inputs_76__7 (registerOutputs_76__7), .inputs_76__6 (
            registerOutputs_76__6), .inputs_76__5 (registerOutputs_76__5), .inputs_76__4 (
            registerOutputs_76__4), .inputs_76__3 (registerOutputs_76__3), .inputs_76__2 (
            registerOutputs_76__2), .inputs_76__1 (registerOutputs_76__1), .inputs_76__0 (
            registerOutputs_76__0), .inputs_77__15 (registerOutputs_77__15), .inputs_77__14 (
            registerOutputs_77__14), .inputs_77__13 (registerOutputs_77__13), .inputs_77__12 (
            registerOutputs_77__12), .inputs_77__11 (registerOutputs_77__11), .inputs_77__10 (
            registerOutputs_77__10), .inputs_77__9 (registerOutputs_77__9), .inputs_77__8 (
            registerOutputs_77__8), .inputs_77__7 (registerOutputs_77__7), .inputs_77__6 (
            registerOutputs_77__6), .inputs_77__5 (registerOutputs_77__5), .inputs_77__4 (
            registerOutputs_77__4), .inputs_77__3 (registerOutputs_77__3), .inputs_77__2 (
            registerOutputs_77__2), .inputs_77__1 (registerOutputs_77__1), .inputs_77__0 (
            registerOutputs_77__0), .inputs_78__15 (registerOutputs_78__15), .inputs_78__14 (
            registerOutputs_78__14), .inputs_78__13 (registerOutputs_78__13), .inputs_78__12 (
            registerOutputs_78__12), .inputs_78__11 (registerOutputs_78__11), .inputs_78__10 (
            registerOutputs_78__10), .inputs_78__9 (registerOutputs_78__9), .inputs_78__8 (
            registerOutputs_78__8), .inputs_78__7 (registerOutputs_78__7), .inputs_78__6 (
            registerOutputs_78__6), .inputs_78__5 (registerOutputs_78__5), .inputs_78__4 (
            registerOutputs_78__4), .inputs_78__3 (registerOutputs_78__3), .inputs_78__2 (
            registerOutputs_78__2), .inputs_78__1 (registerOutputs_78__1), .inputs_78__0 (
            registerOutputs_78__0), .inputs_79__15 (registerOutputs_79__15), .inputs_79__14 (
            registerOutputs_79__14), .inputs_79__13 (registerOutputs_79__13), .inputs_79__12 (
            registerOutputs_79__12), .inputs_79__11 (registerOutputs_79__11), .inputs_79__10 (
            registerOutputs_79__10), .inputs_79__9 (registerOutputs_79__9), .inputs_79__8 (
            registerOutputs_79__8), .inputs_79__7 (registerOutputs_79__7), .inputs_79__6 (
            registerOutputs_79__6), .inputs_79__5 (registerOutputs_79__5), .inputs_79__4 (
            registerOutputs_79__4), .inputs_79__3 (registerOutputs_79__3), .inputs_79__2 (
            registerOutputs_79__2), .inputs_79__1 (registerOutputs_79__1), .inputs_79__0 (
            registerOutputs_79__0), .inputs_80__15 (registerOutputs_80__15), .inputs_80__14 (
            registerOutputs_80__14), .inputs_80__13 (registerOutputs_80__13), .inputs_80__12 (
            registerOutputs_80__12), .inputs_80__11 (registerOutputs_80__11), .inputs_80__10 (
            registerOutputs_80__10), .inputs_80__9 (registerOutputs_80__9), .inputs_80__8 (
            registerOutputs_80__8), .inputs_80__7 (registerOutputs_80__7), .inputs_80__6 (
            registerOutputs_80__6), .inputs_80__5 (registerOutputs_80__5), .inputs_80__4 (
            registerOutputs_80__4), .inputs_80__3 (registerOutputs_80__3), .inputs_80__2 (
            registerOutputs_80__2), .inputs_80__1 (registerOutputs_80__1), .inputs_80__0 (
            registerOutputs_80__0), .inputs_81__15 (registerOutputs_81__15), .inputs_81__14 (
            registerOutputs_81__14), .inputs_81__13 (registerOutputs_81__13), .inputs_81__12 (
            registerOutputs_81__12), .inputs_81__11 (registerOutputs_81__11), .inputs_81__10 (
            registerOutputs_81__10), .inputs_81__9 (registerOutputs_81__9), .inputs_81__8 (
            registerOutputs_81__8), .inputs_81__7 (registerOutputs_81__7), .inputs_81__6 (
            registerOutputs_81__6), .inputs_81__5 (registerOutputs_81__5), .inputs_81__4 (
            registerOutputs_81__4), .inputs_81__3 (registerOutputs_81__3), .inputs_81__2 (
            registerOutputs_81__2), .inputs_81__1 (registerOutputs_81__1), .inputs_81__0 (
            registerOutputs_81__0), .inputs_82__15 (registerOutputs_82__15), .inputs_82__14 (
            registerOutputs_82__14), .inputs_82__13 (registerOutputs_82__13), .inputs_82__12 (
            registerOutputs_82__12), .inputs_82__11 (registerOutputs_82__11), .inputs_82__10 (
            registerOutputs_82__10), .inputs_82__9 (registerOutputs_82__9), .inputs_82__8 (
            registerOutputs_82__8), .inputs_82__7 (registerOutputs_82__7), .inputs_82__6 (
            registerOutputs_82__6), .inputs_82__5 (registerOutputs_82__5), .inputs_82__4 (
            registerOutputs_82__4), .inputs_82__3 (registerOutputs_82__3), .inputs_82__2 (
            registerOutputs_82__2), .inputs_82__1 (registerOutputs_82__1), .inputs_82__0 (
            registerOutputs_82__0), .inputs_83__15 (registerOutputs_83__15), .inputs_83__14 (
            registerOutputs_83__14), .inputs_83__13 (registerOutputs_83__13), .inputs_83__12 (
            registerOutputs_83__12), .inputs_83__11 (registerOutputs_83__11), .inputs_83__10 (
            registerOutputs_83__10), .inputs_83__9 (registerOutputs_83__9), .inputs_83__8 (
            registerOutputs_83__8), .inputs_83__7 (registerOutputs_83__7), .inputs_83__6 (
            registerOutputs_83__6), .inputs_83__5 (registerOutputs_83__5), .inputs_83__4 (
            registerOutputs_83__4), .inputs_83__3 (registerOutputs_83__3), .inputs_83__2 (
            registerOutputs_83__2), .inputs_83__1 (registerOutputs_83__1), .inputs_83__0 (
            registerOutputs_83__0), .inputs_84__15 (registerOutputs_84__15), .inputs_84__14 (
            registerOutputs_84__14), .inputs_84__13 (registerOutputs_84__13), .inputs_84__12 (
            registerOutputs_84__12), .inputs_84__11 (registerOutputs_84__11), .inputs_84__10 (
            registerOutputs_84__10), .inputs_84__9 (registerOutputs_84__9), .inputs_84__8 (
            registerOutputs_84__8), .inputs_84__7 (registerOutputs_84__7), .inputs_84__6 (
            registerOutputs_84__6), .inputs_84__5 (registerOutputs_84__5), .inputs_84__4 (
            registerOutputs_84__4), .inputs_84__3 (registerOutputs_84__3), .inputs_84__2 (
            registerOutputs_84__2), .inputs_84__1 (registerOutputs_84__1), .inputs_84__0 (
            registerOutputs_84__0), .inputs_85__15 (registerOutputs_85__15), .inputs_85__14 (
            registerOutputs_85__14), .inputs_85__13 (registerOutputs_85__13), .inputs_85__12 (
            registerOutputs_85__12), .inputs_85__11 (registerOutputs_85__11), .inputs_85__10 (
            registerOutputs_85__10), .inputs_85__9 (registerOutputs_85__9), .inputs_85__8 (
            registerOutputs_85__8), .inputs_85__7 (registerOutputs_85__7), .inputs_85__6 (
            registerOutputs_85__6), .inputs_85__5 (registerOutputs_85__5), .inputs_85__4 (
            registerOutputs_85__4), .inputs_85__3 (registerOutputs_85__3), .inputs_85__2 (
            registerOutputs_85__2), .inputs_85__1 (registerOutputs_85__1), .inputs_85__0 (
            registerOutputs_85__0), .inputs_86__15 (registerOutputs_86__15), .inputs_86__14 (
            registerOutputs_86__14), .inputs_86__13 (registerOutputs_86__13), .inputs_86__12 (
            registerOutputs_86__12), .inputs_86__11 (registerOutputs_86__11), .inputs_86__10 (
            registerOutputs_86__10), .inputs_86__9 (registerOutputs_86__9), .inputs_86__8 (
            registerOutputs_86__8), .inputs_86__7 (registerOutputs_86__7), .inputs_86__6 (
            registerOutputs_86__6), .inputs_86__5 (registerOutputs_86__5), .inputs_86__4 (
            registerOutputs_86__4), .inputs_86__3 (registerOutputs_86__3), .inputs_86__2 (
            registerOutputs_86__2), .inputs_86__1 (registerOutputs_86__1), .inputs_86__0 (
            registerOutputs_86__0), .inputs_87__15 (registerOutputs_87__15), .inputs_87__14 (
            registerOutputs_87__14), .inputs_87__13 (registerOutputs_87__13), .inputs_87__12 (
            registerOutputs_87__12), .inputs_87__11 (registerOutputs_87__11), .inputs_87__10 (
            registerOutputs_87__10), .inputs_87__9 (registerOutputs_87__9), .inputs_87__8 (
            registerOutputs_87__8), .inputs_87__7 (registerOutputs_87__7), .inputs_87__6 (
            registerOutputs_87__6), .inputs_87__5 (registerOutputs_87__5), .inputs_87__4 (
            registerOutputs_87__4), .inputs_87__3 (registerOutputs_87__3), .inputs_87__2 (
            registerOutputs_87__2), .inputs_87__1 (registerOutputs_87__1), .inputs_87__0 (
            registerOutputs_87__0), .inputs_88__15 (registerOutputs_88__15), .inputs_88__14 (
            registerOutputs_88__14), .inputs_88__13 (registerOutputs_88__13), .inputs_88__12 (
            registerOutputs_88__12), .inputs_88__11 (registerOutputs_88__11), .inputs_88__10 (
            registerOutputs_88__10), .inputs_88__9 (registerOutputs_88__9), .inputs_88__8 (
            registerOutputs_88__8), .inputs_88__7 (registerOutputs_88__7), .inputs_88__6 (
            registerOutputs_88__6), .inputs_88__5 (registerOutputs_88__5), .inputs_88__4 (
            registerOutputs_88__4), .inputs_88__3 (registerOutputs_88__3), .inputs_88__2 (
            registerOutputs_88__2), .inputs_88__1 (registerOutputs_88__1), .inputs_88__0 (
            registerOutputs_88__0), .inputs_89__15 (registerOutputs_89__15), .inputs_89__14 (
            registerOutputs_89__14), .inputs_89__13 (registerOutputs_89__13), .inputs_89__12 (
            registerOutputs_89__12), .inputs_89__11 (registerOutputs_89__11), .inputs_89__10 (
            registerOutputs_89__10), .inputs_89__9 (registerOutputs_89__9), .inputs_89__8 (
            registerOutputs_89__8), .inputs_89__7 (registerOutputs_89__7), .inputs_89__6 (
            registerOutputs_89__6), .inputs_89__5 (registerOutputs_89__5), .inputs_89__4 (
            registerOutputs_89__4), .inputs_89__3 (registerOutputs_89__3), .inputs_89__2 (
            registerOutputs_89__2), .inputs_89__1 (registerOutputs_89__1), .inputs_89__0 (
            registerOutputs_89__0), .inputs_90__15 (registerOutputs_90__15), .inputs_90__14 (
            registerOutputs_90__14), .inputs_90__13 (registerOutputs_90__13), .inputs_90__12 (
            registerOutputs_90__12), .inputs_90__11 (registerOutputs_90__11), .inputs_90__10 (
            registerOutputs_90__10), .inputs_90__9 (registerOutputs_90__9), .inputs_90__8 (
            registerOutputs_90__8), .inputs_90__7 (registerOutputs_90__7), .inputs_90__6 (
            registerOutputs_90__6), .inputs_90__5 (registerOutputs_90__5), .inputs_90__4 (
            registerOutputs_90__4), .inputs_90__3 (registerOutputs_90__3), .inputs_90__2 (
            registerOutputs_90__2), .inputs_90__1 (registerOutputs_90__1), .inputs_90__0 (
            registerOutputs_90__0), .inputs_91__15 (registerOutputs_91__15), .inputs_91__14 (
            registerOutputs_91__14), .inputs_91__13 (registerOutputs_91__13), .inputs_91__12 (
            registerOutputs_91__12), .inputs_91__11 (registerOutputs_91__11), .inputs_91__10 (
            registerOutputs_91__10), .inputs_91__9 (registerOutputs_91__9), .inputs_91__8 (
            registerOutputs_91__8), .inputs_91__7 (registerOutputs_91__7), .inputs_91__6 (
            registerOutputs_91__6), .inputs_91__5 (registerOutputs_91__5), .inputs_91__4 (
            registerOutputs_91__4), .inputs_91__3 (registerOutputs_91__3), .inputs_91__2 (
            registerOutputs_91__2), .inputs_91__1 (registerOutputs_91__1), .inputs_91__0 (
            registerOutputs_91__0), .inputs_92__15 (registerOutputs_92__15), .inputs_92__14 (
            registerOutputs_92__14), .inputs_92__13 (registerOutputs_92__13), .inputs_92__12 (
            registerOutputs_92__12), .inputs_92__11 (registerOutputs_92__11), .inputs_92__10 (
            registerOutputs_92__10), .inputs_92__9 (registerOutputs_92__9), .inputs_92__8 (
            registerOutputs_92__8), .inputs_92__7 (registerOutputs_92__7), .inputs_92__6 (
            registerOutputs_92__6), .inputs_92__5 (registerOutputs_92__5), .inputs_92__4 (
            registerOutputs_92__4), .inputs_92__3 (registerOutputs_92__3), .inputs_92__2 (
            registerOutputs_92__2), .inputs_92__1 (registerOutputs_92__1), .inputs_92__0 (
            registerOutputs_92__0), .inputs_93__15 (registerOutputs_93__15), .inputs_93__14 (
            registerOutputs_93__14), .inputs_93__13 (registerOutputs_93__13), .inputs_93__12 (
            registerOutputs_93__12), .inputs_93__11 (registerOutputs_93__11), .inputs_93__10 (
            registerOutputs_93__10), .inputs_93__9 (registerOutputs_93__9), .inputs_93__8 (
            registerOutputs_93__8), .inputs_93__7 (registerOutputs_93__7), .inputs_93__6 (
            registerOutputs_93__6), .inputs_93__5 (registerOutputs_93__5), .inputs_93__4 (
            registerOutputs_93__4), .inputs_93__3 (registerOutputs_93__3), .inputs_93__2 (
            registerOutputs_93__2), .inputs_93__1 (registerOutputs_93__1), .inputs_93__0 (
            registerOutputs_93__0), .inputs_94__15 (registerOutputs_94__15), .inputs_94__14 (
            registerOutputs_94__14), .inputs_94__13 (registerOutputs_94__13), .inputs_94__12 (
            registerOutputs_94__12), .inputs_94__11 (registerOutputs_94__11), .inputs_94__10 (
            registerOutputs_94__10), .inputs_94__9 (registerOutputs_94__9), .inputs_94__8 (
            registerOutputs_94__8), .inputs_94__7 (registerOutputs_94__7), .inputs_94__6 (
            registerOutputs_94__6), .inputs_94__5 (registerOutputs_94__5), .inputs_94__4 (
            registerOutputs_94__4), .inputs_94__3 (registerOutputs_94__3), .inputs_94__2 (
            registerOutputs_94__2), .inputs_94__1 (registerOutputs_94__1), .inputs_94__0 (
            registerOutputs_94__0), .inputs_95__15 (registerOutputs_95__15), .inputs_95__14 (
            registerOutputs_95__14), .inputs_95__13 (registerOutputs_95__13), .inputs_95__12 (
            registerOutputs_95__12), .inputs_95__11 (registerOutputs_95__11), .inputs_95__10 (
            registerOutputs_95__10), .inputs_95__9 (registerOutputs_95__9), .inputs_95__8 (
            registerOutputs_95__8), .inputs_95__7 (registerOutputs_95__7), .inputs_95__6 (
            registerOutputs_95__6), .inputs_95__5 (registerOutputs_95__5), .inputs_95__4 (
            registerOutputs_95__4), .inputs_95__3 (registerOutputs_95__3), .inputs_95__2 (
            registerOutputs_95__2), .inputs_95__1 (registerOutputs_95__1), .inputs_95__0 (
            registerOutputs_95__0), .inputs_96__15 (registerOutputs_96__15), .inputs_96__14 (
            registerOutputs_96__14), .inputs_96__13 (registerOutputs_96__13), .inputs_96__12 (
            registerOutputs_96__12), .inputs_96__11 (registerOutputs_96__11), .inputs_96__10 (
            registerOutputs_96__10), .inputs_96__9 (registerOutputs_96__9), .inputs_96__8 (
            registerOutputs_96__8), .inputs_96__7 (registerOutputs_96__7), .inputs_96__6 (
            registerOutputs_96__6), .inputs_96__5 (registerOutputs_96__5), .inputs_96__4 (
            registerOutputs_96__4), .inputs_96__3 (registerOutputs_96__3), .inputs_96__2 (
            registerOutputs_96__2), .inputs_96__1 (registerOutputs_96__1), .inputs_96__0 (
            registerOutputs_96__0), .inputs_97__15 (registerOutputs_97__15), .inputs_97__14 (
            registerOutputs_97__14), .inputs_97__13 (registerOutputs_97__13), .inputs_97__12 (
            registerOutputs_97__12), .inputs_97__11 (registerOutputs_97__11), .inputs_97__10 (
            registerOutputs_97__10), .inputs_97__9 (registerOutputs_97__9), .inputs_97__8 (
            registerOutputs_97__8), .inputs_97__7 (registerOutputs_97__7), .inputs_97__6 (
            registerOutputs_97__6), .inputs_97__5 (registerOutputs_97__5), .inputs_97__4 (
            registerOutputs_97__4), .inputs_97__3 (registerOutputs_97__3), .inputs_97__2 (
            registerOutputs_97__2), .inputs_97__1 (registerOutputs_97__1), .inputs_97__0 (
            registerOutputs_97__0), .inputs_98__15 (registerOutputs_98__15), .inputs_98__14 (
            registerOutputs_98__14), .inputs_98__13 (registerOutputs_98__13), .inputs_98__12 (
            registerOutputs_98__12), .inputs_98__11 (registerOutputs_98__11), .inputs_98__10 (
            registerOutputs_98__10), .inputs_98__9 (registerOutputs_98__9), .inputs_98__8 (
            registerOutputs_98__8), .inputs_98__7 (registerOutputs_98__7), .inputs_98__6 (
            registerOutputs_98__6), .inputs_98__5 (registerOutputs_98__5), .inputs_98__4 (
            registerOutputs_98__4), .inputs_98__3 (registerOutputs_98__3), .inputs_98__2 (
            registerOutputs_98__2), .inputs_98__1 (registerOutputs_98__1), .inputs_98__0 (
            registerOutputs_98__0), .inputs_99__15 (registerOutputs_99__15), .inputs_99__14 (
            registerOutputs_99__14), .inputs_99__13 (registerOutputs_99__13), .inputs_99__12 (
            registerOutputs_99__12), .inputs_99__11 (registerOutputs_99__11), .inputs_99__10 (
            registerOutputs_99__10), .inputs_99__9 (registerOutputs_99__9), .inputs_99__8 (
            registerOutputs_99__8), .inputs_99__7 (registerOutputs_99__7), .inputs_99__6 (
            registerOutputs_99__6), .inputs_99__5 (registerOutputs_99__5), .inputs_99__4 (
            registerOutputs_99__4), .inputs_99__3 (registerOutputs_99__3), .inputs_99__2 (
            registerOutputs_99__2), .inputs_99__1 (registerOutputs_99__1), .inputs_99__0 (
            registerOutputs_99__0), .inputs_100__15 (registerOutputs_100__15), .inputs_100__14 (
            registerOutputs_100__14), .inputs_100__13 (registerOutputs_100__13)
            , .inputs_100__12 (registerOutputs_100__12), .inputs_100__11 (
            registerOutputs_100__11), .inputs_100__10 (registerOutputs_100__10)
            , .inputs_100__9 (registerOutputs_100__9), .inputs_100__8 (
            registerOutputs_100__8), .inputs_100__7 (registerOutputs_100__7), .inputs_100__6 (
            registerOutputs_100__6), .inputs_100__5 (registerOutputs_100__5), .inputs_100__4 (
            registerOutputs_100__4), .inputs_100__3 (registerOutputs_100__3), .inputs_100__2 (
            registerOutputs_100__2), .inputs_100__1 (registerOutputs_100__1), .inputs_100__0 (
            registerOutputs_100__0), .inputs_101__15 (registerOutputs_101__15), 
            .inputs_101__14 (registerOutputs_101__14), .inputs_101__13 (
            registerOutputs_101__13), .inputs_101__12 (registerOutputs_101__12)
            , .inputs_101__11 (registerOutputs_101__11), .inputs_101__10 (
            registerOutputs_101__10), .inputs_101__9 (registerOutputs_101__9), .inputs_101__8 (
            registerOutputs_101__8), .inputs_101__7 (registerOutputs_101__7), .inputs_101__6 (
            registerOutputs_101__6), .inputs_101__5 (registerOutputs_101__5), .inputs_101__4 (
            registerOutputs_101__4), .inputs_101__3 (registerOutputs_101__3), .inputs_101__2 (
            registerOutputs_101__2), .inputs_101__1 (registerOutputs_101__1), .inputs_101__0 (
            registerOutputs_101__0), .inputs_102__15 (registerOutputs_102__15), 
            .inputs_102__14 (registerOutputs_102__14), .inputs_102__13 (
            registerOutputs_102__13), .inputs_102__12 (registerOutputs_102__12)
            , .inputs_102__11 (registerOutputs_102__11), .inputs_102__10 (
            registerOutputs_102__10), .inputs_102__9 (registerOutputs_102__9), .inputs_102__8 (
            registerOutputs_102__8), .inputs_102__7 (registerOutputs_102__7), .inputs_102__6 (
            registerOutputs_102__6), .inputs_102__5 (registerOutputs_102__5), .inputs_102__4 (
            registerOutputs_102__4), .inputs_102__3 (registerOutputs_102__3), .inputs_102__2 (
            registerOutputs_102__2), .inputs_102__1 (registerOutputs_102__1), .inputs_102__0 (
            registerOutputs_102__0), .inputs_103__15 (registerOutputs_103__15), 
            .inputs_103__14 (registerOutputs_103__14), .inputs_103__13 (
            registerOutputs_103__13), .inputs_103__12 (registerOutputs_103__12)
            , .inputs_103__11 (registerOutputs_103__11), .inputs_103__10 (
            registerOutputs_103__10), .inputs_103__9 (registerOutputs_103__9), .inputs_103__8 (
            registerOutputs_103__8), .inputs_103__7 (registerOutputs_103__7), .inputs_103__6 (
            registerOutputs_103__6), .inputs_103__5 (registerOutputs_103__5), .inputs_103__4 (
            registerOutputs_103__4), .inputs_103__3 (registerOutputs_103__3), .inputs_103__2 (
            registerOutputs_103__2), .inputs_103__1 (registerOutputs_103__1), .inputs_103__0 (
            registerOutputs_103__0), .inputs_104__15 (registerOutputs_104__15), 
            .inputs_104__14 (registerOutputs_104__14), .inputs_104__13 (
            registerOutputs_104__13), .inputs_104__12 (registerOutputs_104__12)
            , .inputs_104__11 (registerOutputs_104__11), .inputs_104__10 (
            registerOutputs_104__10), .inputs_104__9 (registerOutputs_104__9), .inputs_104__8 (
            registerOutputs_104__8), .inputs_104__7 (registerOutputs_104__7), .inputs_104__6 (
            registerOutputs_104__6), .inputs_104__5 (registerOutputs_104__5), .inputs_104__4 (
            registerOutputs_104__4), .inputs_104__3 (registerOutputs_104__3), .inputs_104__2 (
            registerOutputs_104__2), .inputs_104__1 (registerOutputs_104__1), .inputs_104__0 (
            registerOutputs_104__0), .inputs_105__15 (registerOutputs_105__15), 
            .inputs_105__14 (registerOutputs_105__14), .inputs_105__13 (
            registerOutputs_105__13), .inputs_105__12 (registerOutputs_105__12)
            , .inputs_105__11 (registerOutputs_105__11), .inputs_105__10 (
            registerOutputs_105__10), .inputs_105__9 (registerOutputs_105__9), .inputs_105__8 (
            registerOutputs_105__8), .inputs_105__7 (registerOutputs_105__7), .inputs_105__6 (
            registerOutputs_105__6), .inputs_105__5 (registerOutputs_105__5), .inputs_105__4 (
            registerOutputs_105__4), .inputs_105__3 (registerOutputs_105__3), .inputs_105__2 (
            registerOutputs_105__2), .inputs_105__1 (registerOutputs_105__1), .inputs_105__0 (
            registerOutputs_105__0), .inputs_106__15 (registerOutputs_106__15), 
            .inputs_106__14 (registerOutputs_106__14), .inputs_106__13 (
            registerOutputs_106__13), .inputs_106__12 (registerOutputs_106__12)
            , .inputs_106__11 (registerOutputs_106__11), .inputs_106__10 (
            registerOutputs_106__10), .inputs_106__9 (registerOutputs_106__9), .inputs_106__8 (
            registerOutputs_106__8), .inputs_106__7 (registerOutputs_106__7), .inputs_106__6 (
            registerOutputs_106__6), .inputs_106__5 (registerOutputs_106__5), .inputs_106__4 (
            registerOutputs_106__4), .inputs_106__3 (registerOutputs_106__3), .inputs_106__2 (
            registerOutputs_106__2), .inputs_106__1 (registerOutputs_106__1), .inputs_106__0 (
            registerOutputs_106__0), .inputs_107__15 (registerOutputs_107__15), 
            .inputs_107__14 (registerOutputs_107__14), .inputs_107__13 (
            registerOutputs_107__13), .inputs_107__12 (registerOutputs_107__12)
            , .inputs_107__11 (registerOutputs_107__11), .inputs_107__10 (
            registerOutputs_107__10), .inputs_107__9 (registerOutputs_107__9), .inputs_107__8 (
            registerOutputs_107__8), .inputs_107__7 (registerOutputs_107__7), .inputs_107__6 (
            registerOutputs_107__6), .inputs_107__5 (registerOutputs_107__5), .inputs_107__4 (
            registerOutputs_107__4), .inputs_107__3 (registerOutputs_107__3), .inputs_107__2 (
            registerOutputs_107__2), .inputs_107__1 (registerOutputs_107__1), .inputs_107__0 (
            registerOutputs_107__0), .inputs_108__15 (registerOutputs_108__15), 
            .inputs_108__14 (registerOutputs_108__14), .inputs_108__13 (
            registerOutputs_108__13), .inputs_108__12 (registerOutputs_108__12)
            , .inputs_108__11 (registerOutputs_108__11), .inputs_108__10 (
            registerOutputs_108__10), .inputs_108__9 (registerOutputs_108__9), .inputs_108__8 (
            registerOutputs_108__8), .inputs_108__7 (registerOutputs_108__7), .inputs_108__6 (
            registerOutputs_108__6), .inputs_108__5 (registerOutputs_108__5), .inputs_108__4 (
            registerOutputs_108__4), .inputs_108__3 (registerOutputs_108__3), .inputs_108__2 (
            registerOutputs_108__2), .inputs_108__1 (registerOutputs_108__1), .inputs_108__0 (
            registerOutputs_108__0), .inputs_109__15 (registerOutputs_109__15), 
            .inputs_109__14 (registerOutputs_109__14), .inputs_109__13 (
            registerOutputs_109__13), .inputs_109__12 (registerOutputs_109__12)
            , .inputs_109__11 (registerOutputs_109__11), .inputs_109__10 (
            registerOutputs_109__10), .inputs_109__9 (registerOutputs_109__9), .inputs_109__8 (
            registerOutputs_109__8), .inputs_109__7 (registerOutputs_109__7), .inputs_109__6 (
            registerOutputs_109__6), .inputs_109__5 (registerOutputs_109__5), .inputs_109__4 (
            registerOutputs_109__4), .inputs_109__3 (registerOutputs_109__3), .inputs_109__2 (
            registerOutputs_109__2), .inputs_109__1 (registerOutputs_109__1), .inputs_109__0 (
            registerOutputs_109__0), .inputs_110__15 (registerOutputs_110__15), 
            .inputs_110__14 (registerOutputs_110__14), .inputs_110__13 (
            registerOutputs_110__13), .inputs_110__12 (registerOutputs_110__12)
            , .inputs_110__11 (registerOutputs_110__11), .inputs_110__10 (
            registerOutputs_110__10), .inputs_110__9 (registerOutputs_110__9), .inputs_110__8 (
            registerOutputs_110__8), .inputs_110__7 (registerOutputs_110__7), .inputs_110__6 (
            registerOutputs_110__6), .inputs_110__5 (registerOutputs_110__5), .inputs_110__4 (
            registerOutputs_110__4), .inputs_110__3 (registerOutputs_110__3), .inputs_110__2 (
            registerOutputs_110__2), .inputs_110__1 (registerOutputs_110__1), .inputs_110__0 (
            registerOutputs_110__0), .inputs_111__15 (registerOutputs_111__15), 
            .inputs_111__14 (registerOutputs_111__14), .inputs_111__13 (
            registerOutputs_111__13), .inputs_111__12 (registerOutputs_111__12)
            , .inputs_111__11 (registerOutputs_111__11), .inputs_111__10 (
            registerOutputs_111__10), .inputs_111__9 (registerOutputs_111__9), .inputs_111__8 (
            registerOutputs_111__8), .inputs_111__7 (registerOutputs_111__7), .inputs_111__6 (
            registerOutputs_111__6), .inputs_111__5 (registerOutputs_111__5), .inputs_111__4 (
            registerOutputs_111__4), .inputs_111__3 (registerOutputs_111__3), .inputs_111__2 (
            registerOutputs_111__2), .inputs_111__1 (registerOutputs_111__1), .inputs_111__0 (
            registerOutputs_111__0), .inputs_112__15 (registerOutputs_112__15), 
            .inputs_112__14 (registerOutputs_112__14), .inputs_112__13 (
            registerOutputs_112__13), .inputs_112__12 (registerOutputs_112__12)
            , .inputs_112__11 (registerOutputs_112__11), .inputs_112__10 (
            registerOutputs_112__10), .inputs_112__9 (registerOutputs_112__9), .inputs_112__8 (
            registerOutputs_112__8), .inputs_112__7 (registerOutputs_112__7), .inputs_112__6 (
            registerOutputs_112__6), .inputs_112__5 (registerOutputs_112__5), .inputs_112__4 (
            registerOutputs_112__4), .inputs_112__3 (registerOutputs_112__3), .inputs_112__2 (
            registerOutputs_112__2), .inputs_112__1 (registerOutputs_112__1), .inputs_112__0 (
            registerOutputs_112__0), .inputs_113__15 (registerOutputs_113__15), 
            .inputs_113__14 (registerOutputs_113__14), .inputs_113__13 (
            registerOutputs_113__13), .inputs_113__12 (registerOutputs_113__12)
            , .inputs_113__11 (registerOutputs_113__11), .inputs_113__10 (
            registerOutputs_113__10), .inputs_113__9 (registerOutputs_113__9), .inputs_113__8 (
            registerOutputs_113__8), .inputs_113__7 (registerOutputs_113__7), .inputs_113__6 (
            registerOutputs_113__6), .inputs_113__5 (registerOutputs_113__5), .inputs_113__4 (
            registerOutputs_113__4), .inputs_113__3 (registerOutputs_113__3), .inputs_113__2 (
            registerOutputs_113__2), .inputs_113__1 (registerOutputs_113__1), .inputs_113__0 (
            registerOutputs_113__0), .inputs_114__15 (registerOutputs_114__15), 
            .inputs_114__14 (registerOutputs_114__14), .inputs_114__13 (
            registerOutputs_114__13), .inputs_114__12 (registerOutputs_114__12)
            , .inputs_114__11 (registerOutputs_114__11), .inputs_114__10 (
            registerOutputs_114__10), .inputs_114__9 (registerOutputs_114__9), .inputs_114__8 (
            registerOutputs_114__8), .inputs_114__7 (registerOutputs_114__7), .inputs_114__6 (
            registerOutputs_114__6), .inputs_114__5 (registerOutputs_114__5), .inputs_114__4 (
            registerOutputs_114__4), .inputs_114__3 (registerOutputs_114__3), .inputs_114__2 (
            registerOutputs_114__2), .inputs_114__1 (registerOutputs_114__1), .inputs_114__0 (
            registerOutputs_114__0), .inputs_115__15 (registerOutputs_115__15), 
            .inputs_115__14 (registerOutputs_115__14), .inputs_115__13 (
            registerOutputs_115__13), .inputs_115__12 (registerOutputs_115__12)
            , .inputs_115__11 (registerOutputs_115__11), .inputs_115__10 (
            registerOutputs_115__10), .inputs_115__9 (registerOutputs_115__9), .inputs_115__8 (
            registerOutputs_115__8), .inputs_115__7 (registerOutputs_115__7), .inputs_115__6 (
            registerOutputs_115__6), .inputs_115__5 (registerOutputs_115__5), .inputs_115__4 (
            registerOutputs_115__4), .inputs_115__3 (registerOutputs_115__3), .inputs_115__2 (
            registerOutputs_115__2), .inputs_115__1 (registerOutputs_115__1), .inputs_115__0 (
            registerOutputs_115__0), .inputs_116__15 (registerOutputs_116__15), 
            .inputs_116__14 (registerOutputs_116__14), .inputs_116__13 (
            registerOutputs_116__13), .inputs_116__12 (registerOutputs_116__12)
            , .inputs_116__11 (registerOutputs_116__11), .inputs_116__10 (
            registerOutputs_116__10), .inputs_116__9 (registerOutputs_116__9), .inputs_116__8 (
            registerOutputs_116__8), .inputs_116__7 (registerOutputs_116__7), .inputs_116__6 (
            registerOutputs_116__6), .inputs_116__5 (registerOutputs_116__5), .inputs_116__4 (
            registerOutputs_116__4), .inputs_116__3 (registerOutputs_116__3), .inputs_116__2 (
            registerOutputs_116__2), .inputs_116__1 (registerOutputs_116__1), .inputs_116__0 (
            registerOutputs_116__0), .inputs_117__15 (registerOutputs_117__15), 
            .inputs_117__14 (registerOutputs_117__14), .inputs_117__13 (
            registerOutputs_117__13), .inputs_117__12 (registerOutputs_117__12)
            , .inputs_117__11 (registerOutputs_117__11), .inputs_117__10 (
            registerOutputs_117__10), .inputs_117__9 (registerOutputs_117__9), .inputs_117__8 (
            registerOutputs_117__8), .inputs_117__7 (registerOutputs_117__7), .inputs_117__6 (
            registerOutputs_117__6), .inputs_117__5 (registerOutputs_117__5), .inputs_117__4 (
            registerOutputs_117__4), .inputs_117__3 (registerOutputs_117__3), .inputs_117__2 (
            registerOutputs_117__2), .inputs_117__1 (registerOutputs_117__1), .inputs_117__0 (
            registerOutputs_117__0), .inputs_118__15 (registerOutputs_118__15), 
            .inputs_118__14 (registerOutputs_118__14), .inputs_118__13 (
            registerOutputs_118__13), .inputs_118__12 (registerOutputs_118__12)
            , .inputs_118__11 (registerOutputs_118__11), .inputs_118__10 (
            registerOutputs_118__10), .inputs_118__9 (registerOutputs_118__9), .inputs_118__8 (
            registerOutputs_118__8), .inputs_118__7 (registerOutputs_118__7), .inputs_118__6 (
            registerOutputs_118__6), .inputs_118__5 (registerOutputs_118__5), .inputs_118__4 (
            registerOutputs_118__4), .inputs_118__3 (registerOutputs_118__3), .inputs_118__2 (
            registerOutputs_118__2), .inputs_118__1 (registerOutputs_118__1), .inputs_118__0 (
            registerOutputs_118__0), .inputs_119__15 (registerOutputs_119__15), 
            .inputs_119__14 (registerOutputs_119__14), .inputs_119__13 (
            registerOutputs_119__13), .inputs_119__12 (registerOutputs_119__12)
            , .inputs_119__11 (registerOutputs_119__11), .inputs_119__10 (
            registerOutputs_119__10), .inputs_119__9 (registerOutputs_119__9), .inputs_119__8 (
            registerOutputs_119__8), .inputs_119__7 (registerOutputs_119__7), .inputs_119__6 (
            registerOutputs_119__6), .inputs_119__5 (registerOutputs_119__5), .inputs_119__4 (
            registerOutputs_119__4), .inputs_119__3 (registerOutputs_119__3), .inputs_119__2 (
            registerOutputs_119__2), .inputs_119__1 (registerOutputs_119__1), .inputs_119__0 (
            registerOutputs_119__0), .inputs_120__15 (registerOutputs_120__15), 
            .inputs_120__14 (registerOutputs_120__14), .inputs_120__13 (
            registerOutputs_120__13), .inputs_120__12 (registerOutputs_120__12)
            , .inputs_120__11 (registerOutputs_120__11), .inputs_120__10 (
            registerOutputs_120__10), .inputs_120__9 (registerOutputs_120__9), .inputs_120__8 (
            registerOutputs_120__8), .inputs_120__7 (registerOutputs_120__7), .inputs_120__6 (
            registerOutputs_120__6), .inputs_120__5 (registerOutputs_120__5), .inputs_120__4 (
            registerOutputs_120__4), .inputs_120__3 (registerOutputs_120__3), .inputs_120__2 (
            registerOutputs_120__2), .inputs_120__1 (registerOutputs_120__1), .inputs_120__0 (
            registerOutputs_120__0), .inputs_121__15 (registerOutputs_121__15), 
            .inputs_121__14 (registerOutputs_121__14), .inputs_121__13 (
            registerOutputs_121__13), .inputs_121__12 (registerOutputs_121__12)
            , .inputs_121__11 (registerOutputs_121__11), .inputs_121__10 (
            registerOutputs_121__10), .inputs_121__9 (registerOutputs_121__9), .inputs_121__8 (
            registerOutputs_121__8), .inputs_121__7 (registerOutputs_121__7), .inputs_121__6 (
            registerOutputs_121__6), .inputs_121__5 (registerOutputs_121__5), .inputs_121__4 (
            registerOutputs_121__4), .inputs_121__3 (registerOutputs_121__3), .inputs_121__2 (
            registerOutputs_121__2), .inputs_121__1 (registerOutputs_121__1), .inputs_121__0 (
            registerOutputs_121__0), .inputs_122__15 (registerOutputs_122__15), 
            .inputs_122__14 (registerOutputs_122__14), .inputs_122__13 (
            registerOutputs_122__13), .inputs_122__12 (registerOutputs_122__12)
            , .inputs_122__11 (registerOutputs_122__11), .inputs_122__10 (
            registerOutputs_122__10), .inputs_122__9 (registerOutputs_122__9), .inputs_122__8 (
            registerOutputs_122__8), .inputs_122__7 (registerOutputs_122__7), .inputs_122__6 (
            registerOutputs_122__6), .inputs_122__5 (registerOutputs_122__5), .inputs_122__4 (
            registerOutputs_122__4), .inputs_122__3 (registerOutputs_122__3), .inputs_122__2 (
            registerOutputs_122__2), .inputs_122__1 (registerOutputs_122__1), .inputs_122__0 (
            registerOutputs_122__0), .inputs_123__15 (registerOutputs_123__15), 
            .inputs_123__14 (registerOutputs_123__14), .inputs_123__13 (
            registerOutputs_123__13), .inputs_123__12 (registerOutputs_123__12)
            , .inputs_123__11 (registerOutputs_123__11), .inputs_123__10 (
            registerOutputs_123__10), .inputs_123__9 (registerOutputs_123__9), .inputs_123__8 (
            registerOutputs_123__8), .inputs_123__7 (registerOutputs_123__7), .inputs_123__6 (
            registerOutputs_123__6), .inputs_123__5 (registerOutputs_123__5), .inputs_123__4 (
            registerOutputs_123__4), .inputs_123__3 (registerOutputs_123__3), .inputs_123__2 (
            registerOutputs_123__2), .inputs_123__1 (registerOutputs_123__1), .inputs_123__0 (
            registerOutputs_123__0), .inputs_124__15 (registerOutputs_124__15), 
            .inputs_124__14 (registerOutputs_124__14), .inputs_124__13 (
            registerOutputs_124__13), .inputs_124__12 (registerOutputs_124__12)
            , .inputs_124__11 (registerOutputs_124__11), .inputs_124__10 (
            registerOutputs_124__10), .inputs_124__9 (registerOutputs_124__9), .inputs_124__8 (
            registerOutputs_124__8), .inputs_124__7 (registerOutputs_124__7), .inputs_124__6 (
            registerOutputs_124__6), .inputs_124__5 (registerOutputs_124__5), .inputs_124__4 (
            registerOutputs_124__4), .inputs_124__3 (registerOutputs_124__3), .inputs_124__2 (
            registerOutputs_124__2), .inputs_124__1 (registerOutputs_124__1), .inputs_124__0 (
            registerOutputs_124__0), .inputs_125__15 (registerOutputs_125__15), 
            .inputs_125__14 (registerOutputs_125__14), .inputs_125__13 (
            registerOutputs_125__13), .inputs_125__12 (registerOutputs_125__12)
            , .inputs_125__11 (registerOutputs_125__11), .inputs_125__10 (
            registerOutputs_125__10), .inputs_125__9 (registerOutputs_125__9), .inputs_125__8 (
            registerOutputs_125__8), .inputs_125__7 (registerOutputs_125__7), .inputs_125__6 (
            registerOutputs_125__6), .inputs_125__5 (registerOutputs_125__5), .inputs_125__4 (
            registerOutputs_125__4), .inputs_125__3 (registerOutputs_125__3), .inputs_125__2 (
            registerOutputs_125__2), .inputs_125__1 (registerOutputs_125__1), .inputs_125__0 (
            registerOutputs_125__0), .inputs_126__15 (registerOutputs_126__15), 
            .inputs_126__14 (registerOutputs_126__14), .inputs_126__13 (
            registerOutputs_126__13), .inputs_126__12 (registerOutputs_126__12)
            , .inputs_126__11 (registerOutputs_126__11), .inputs_126__10 (
            registerOutputs_126__10), .inputs_126__9 (registerOutputs_126__9), .inputs_126__8 (
            registerOutputs_126__8), .inputs_126__7 (registerOutputs_126__7), .inputs_126__6 (
            registerOutputs_126__6), .inputs_126__5 (registerOutputs_126__5), .inputs_126__4 (
            registerOutputs_126__4), .inputs_126__3 (registerOutputs_126__3), .inputs_126__2 (
            registerOutputs_126__2), .inputs_126__1 (registerOutputs_126__1), .inputs_126__0 (
            registerOutputs_126__0), .inputs_127__15 (registerOutputs_127__15), 
            .inputs_127__14 (registerOutputs_127__14), .inputs_127__13 (
            registerOutputs_127__13), .inputs_127__12 (registerOutputs_127__12)
            , .inputs_127__11 (registerOutputs_127__11), .inputs_127__10 (
            registerOutputs_127__10), .inputs_127__9 (registerOutputs_127__9), .inputs_127__8 (
            registerOutputs_127__8), .inputs_127__7 (registerOutputs_127__7), .inputs_127__6 (
            registerOutputs_127__6), .inputs_127__5 (registerOutputs_127__5), .inputs_127__4 (
            registerOutputs_127__4), .inputs_127__3 (registerOutputs_127__3), .inputs_127__2 (
            registerOutputs_127__2), .inputs_127__1 (registerOutputs_127__1), .inputs_127__0 (
            registerOutputs_127__0), .inputs_128__15 (registerOutputs_128__15), 
            .inputs_128__14 (registerOutputs_128__14), .inputs_128__13 (
            registerOutputs_128__13), .inputs_128__12 (registerOutputs_128__12)
            , .inputs_128__11 (registerOutputs_128__11), .inputs_128__10 (
            registerOutputs_128__10), .inputs_128__9 (registerOutputs_128__9), .inputs_128__8 (
            registerOutputs_128__8), .inputs_128__7 (registerOutputs_128__7), .inputs_128__6 (
            registerOutputs_128__6), .inputs_128__5 (registerOutputs_128__5), .inputs_128__4 (
            registerOutputs_128__4), .inputs_128__3 (registerOutputs_128__3), .inputs_128__2 (
            registerOutputs_128__2), .inputs_128__1 (registerOutputs_128__1), .inputs_128__0 (
            registerOutputs_128__0), .inputs_129__15 (registerOutputs_129__15), 
            .inputs_129__14 (registerOutputs_129__14), .inputs_129__13 (
            registerOutputs_129__13), .inputs_129__12 (registerOutputs_129__12)
            , .inputs_129__11 (registerOutputs_129__11), .inputs_129__10 (
            registerOutputs_129__10), .inputs_129__9 (registerOutputs_129__9), .inputs_129__8 (
            registerOutputs_129__8), .inputs_129__7 (registerOutputs_129__7), .inputs_129__6 (
            registerOutputs_129__6), .inputs_129__5 (registerOutputs_129__5), .inputs_129__4 (
            registerOutputs_129__4), .inputs_129__3 (registerOutputs_129__3), .inputs_129__2 (
            registerOutputs_129__2), .inputs_129__1 (registerOutputs_129__1), .inputs_129__0 (
            registerOutputs_129__0), .inputs_130__15 (registerOutputs_130__15), 
            .inputs_130__14 (registerOutputs_130__14), .inputs_130__13 (
            registerOutputs_130__13), .inputs_130__12 (registerOutputs_130__12)
            , .inputs_130__11 (registerOutputs_130__11), .inputs_130__10 (
            registerOutputs_130__10), .inputs_130__9 (registerOutputs_130__9), .inputs_130__8 (
            registerOutputs_130__8), .inputs_130__7 (registerOutputs_130__7), .inputs_130__6 (
            registerOutputs_130__6), .inputs_130__5 (registerOutputs_130__5), .inputs_130__4 (
            registerOutputs_130__4), .inputs_130__3 (registerOutputs_130__3), .inputs_130__2 (
            registerOutputs_130__2), .inputs_130__1 (registerOutputs_130__1), .inputs_130__0 (
            registerOutputs_130__0), .inputs_131__15 (registerOutputs_131__15), 
            .inputs_131__14 (registerOutputs_131__14), .inputs_131__13 (
            registerOutputs_131__13), .inputs_131__12 (registerOutputs_131__12)
            , .inputs_131__11 (registerOutputs_131__11), .inputs_131__10 (
            registerOutputs_131__10), .inputs_131__9 (registerOutputs_131__9), .inputs_131__8 (
            registerOutputs_131__8), .inputs_131__7 (registerOutputs_131__7), .inputs_131__6 (
            registerOutputs_131__6), .inputs_131__5 (registerOutputs_131__5), .inputs_131__4 (
            registerOutputs_131__4), .inputs_131__3 (registerOutputs_131__3), .inputs_131__2 (
            registerOutputs_131__2), .inputs_131__1 (registerOutputs_131__1), .inputs_131__0 (
            registerOutputs_131__0), .inputs_132__15 (registerOutputs_132__15), 
            .inputs_132__14 (registerOutputs_132__14), .inputs_132__13 (
            registerOutputs_132__13), .inputs_132__12 (registerOutputs_132__12)
            , .inputs_132__11 (registerOutputs_132__11), .inputs_132__10 (
            registerOutputs_132__10), .inputs_132__9 (registerOutputs_132__9), .inputs_132__8 (
            registerOutputs_132__8), .inputs_132__7 (registerOutputs_132__7), .inputs_132__6 (
            registerOutputs_132__6), .inputs_132__5 (registerOutputs_132__5), .inputs_132__4 (
            registerOutputs_132__4), .inputs_132__3 (registerOutputs_132__3), .inputs_132__2 (
            registerOutputs_132__2), .inputs_132__1 (registerOutputs_132__1), .inputs_132__0 (
            registerOutputs_132__0), .inputs_133__15 (registerOutputs_133__15), 
            .inputs_133__14 (registerOutputs_133__14), .inputs_133__13 (
            registerOutputs_133__13), .inputs_133__12 (registerOutputs_133__12)
            , .inputs_133__11 (registerOutputs_133__11), .inputs_133__10 (
            registerOutputs_133__10), .inputs_133__9 (registerOutputs_133__9), .inputs_133__8 (
            registerOutputs_133__8), .inputs_133__7 (registerOutputs_133__7), .inputs_133__6 (
            registerOutputs_133__6), .inputs_133__5 (registerOutputs_133__5), .inputs_133__4 (
            registerOutputs_133__4), .inputs_133__3 (registerOutputs_133__3), .inputs_133__2 (
            registerOutputs_133__2), .inputs_133__1 (registerOutputs_133__1), .inputs_133__0 (
            registerOutputs_133__0), .inputs_134__15 (registerOutputs_134__15), 
            .inputs_134__14 (registerOutputs_134__14), .inputs_134__13 (
            registerOutputs_134__13), .inputs_134__12 (registerOutputs_134__12)
            , .inputs_134__11 (registerOutputs_134__11), .inputs_134__10 (
            registerOutputs_134__10), .inputs_134__9 (registerOutputs_134__9), .inputs_134__8 (
            registerOutputs_134__8), .inputs_134__7 (registerOutputs_134__7), .inputs_134__6 (
            registerOutputs_134__6), .inputs_134__5 (registerOutputs_134__5), .inputs_134__4 (
            registerOutputs_134__4), .inputs_134__3 (registerOutputs_134__3), .inputs_134__2 (
            registerOutputs_134__2), .inputs_134__1 (registerOutputs_134__1), .inputs_134__0 (
            registerOutputs_134__0), .inputs_135__15 (registerOutputs_135__15), 
            .inputs_135__14 (registerOutputs_135__14), .inputs_135__13 (
            registerOutputs_135__13), .inputs_135__12 (registerOutputs_135__12)
            , .inputs_135__11 (registerOutputs_135__11), .inputs_135__10 (
            registerOutputs_135__10), .inputs_135__9 (registerOutputs_135__9), .inputs_135__8 (
            registerOutputs_135__8), .inputs_135__7 (registerOutputs_135__7), .inputs_135__6 (
            registerOutputs_135__6), .inputs_135__5 (registerOutputs_135__5), .inputs_135__4 (
            registerOutputs_135__4), .inputs_135__3 (registerOutputs_135__3), .inputs_135__2 (
            registerOutputs_135__2), .inputs_135__1 (registerOutputs_135__1), .inputs_135__0 (
            registerOutputs_135__0), .inputs_136__15 (registerOutputs_136__15), 
            .inputs_136__14 (registerOutputs_136__14), .inputs_136__13 (
            registerOutputs_136__13), .inputs_136__12 (registerOutputs_136__12)
            , .inputs_136__11 (registerOutputs_136__11), .inputs_136__10 (
            registerOutputs_136__10), .inputs_136__9 (registerOutputs_136__9), .inputs_136__8 (
            registerOutputs_136__8), .inputs_136__7 (registerOutputs_136__7), .inputs_136__6 (
            registerOutputs_136__6), .inputs_136__5 (registerOutputs_136__5), .inputs_136__4 (
            registerOutputs_136__4), .inputs_136__3 (registerOutputs_136__3), .inputs_136__2 (
            registerOutputs_136__2), .inputs_136__1 (registerOutputs_136__1), .inputs_136__0 (
            registerOutputs_136__0), .inputs_137__15 (registerOutputs_137__15), 
            .inputs_137__14 (registerOutputs_137__14), .inputs_137__13 (
            registerOutputs_137__13), .inputs_137__12 (registerOutputs_137__12)
            , .inputs_137__11 (registerOutputs_137__11), .inputs_137__10 (
            registerOutputs_137__10), .inputs_137__9 (registerOutputs_137__9), .inputs_137__8 (
            registerOutputs_137__8), .inputs_137__7 (registerOutputs_137__7), .inputs_137__6 (
            registerOutputs_137__6), .inputs_137__5 (registerOutputs_137__5), .inputs_137__4 (
            registerOutputs_137__4), .inputs_137__3 (registerOutputs_137__3), .inputs_137__2 (
            registerOutputs_137__2), .inputs_137__1 (registerOutputs_137__1), .inputs_137__0 (
            registerOutputs_137__0), .inputs_138__15 (registerOutputs_138__15), 
            .inputs_138__14 (registerOutputs_138__14), .inputs_138__13 (
            registerOutputs_138__13), .inputs_138__12 (registerOutputs_138__12)
            , .inputs_138__11 (registerOutputs_138__11), .inputs_138__10 (
            registerOutputs_138__10), .inputs_138__9 (registerOutputs_138__9), .inputs_138__8 (
            registerOutputs_138__8), .inputs_138__7 (registerOutputs_138__7), .inputs_138__6 (
            registerOutputs_138__6), .inputs_138__5 (registerOutputs_138__5), .inputs_138__4 (
            registerOutputs_138__4), .inputs_138__3 (registerOutputs_138__3), .inputs_138__2 (
            registerOutputs_138__2), .inputs_138__1 (registerOutputs_138__1), .inputs_138__0 (
            registerOutputs_138__0), .inputs_139__15 (registerOutputs_139__15), 
            .inputs_139__14 (registerOutputs_139__14), .inputs_139__13 (
            registerOutputs_139__13), .inputs_139__12 (registerOutputs_139__12)
            , .inputs_139__11 (registerOutputs_139__11), .inputs_139__10 (
            registerOutputs_139__10), .inputs_139__9 (registerOutputs_139__9), .inputs_139__8 (
            registerOutputs_139__8), .inputs_139__7 (registerOutputs_139__7), .inputs_139__6 (
            registerOutputs_139__6), .inputs_139__5 (registerOutputs_139__5), .inputs_139__4 (
            registerOutputs_139__4), .inputs_139__3 (registerOutputs_139__3), .inputs_139__2 (
            registerOutputs_139__2), .inputs_139__1 (registerOutputs_139__1), .inputs_139__0 (
            registerOutputs_139__0), .inputs_140__15 (registerOutputs_140__15), 
            .inputs_140__14 (registerOutputs_140__14), .inputs_140__13 (
            registerOutputs_140__13), .inputs_140__12 (registerOutputs_140__12)
            , .inputs_140__11 (registerOutputs_140__11), .inputs_140__10 (
            registerOutputs_140__10), .inputs_140__9 (registerOutputs_140__9), .inputs_140__8 (
            registerOutputs_140__8), .inputs_140__7 (registerOutputs_140__7), .inputs_140__6 (
            registerOutputs_140__6), .inputs_140__5 (registerOutputs_140__5), .inputs_140__4 (
            registerOutputs_140__4), .inputs_140__3 (registerOutputs_140__3), .inputs_140__2 (
            registerOutputs_140__2), .inputs_140__1 (registerOutputs_140__1), .inputs_140__0 (
            registerOutputs_140__0), .inputs_141__15 (registerOutputs_141__15), 
            .inputs_141__14 (registerOutputs_141__14), .inputs_141__13 (
            registerOutputs_141__13), .inputs_141__12 (registerOutputs_141__12)
            , .inputs_141__11 (registerOutputs_141__11), .inputs_141__10 (
            registerOutputs_141__10), .inputs_141__9 (registerOutputs_141__9), .inputs_141__8 (
            registerOutputs_141__8), .inputs_141__7 (registerOutputs_141__7), .inputs_141__6 (
            registerOutputs_141__6), .inputs_141__5 (registerOutputs_141__5), .inputs_141__4 (
            registerOutputs_141__4), .inputs_141__3 (registerOutputs_141__3), .inputs_141__2 (
            registerOutputs_141__2), .inputs_141__1 (registerOutputs_141__1), .inputs_141__0 (
            registerOutputs_141__0), .inputs_142__15 (registerOutputs_142__15), 
            .inputs_142__14 (registerOutputs_142__14), .inputs_142__13 (
            registerOutputs_142__13), .inputs_142__12 (registerOutputs_142__12)
            , .inputs_142__11 (registerOutputs_142__11), .inputs_142__10 (
            registerOutputs_142__10), .inputs_142__9 (registerOutputs_142__9), .inputs_142__8 (
            registerOutputs_142__8), .inputs_142__7 (registerOutputs_142__7), .inputs_142__6 (
            registerOutputs_142__6), .inputs_142__5 (registerOutputs_142__5), .inputs_142__4 (
            registerOutputs_142__4), .inputs_142__3 (registerOutputs_142__3), .inputs_142__2 (
            registerOutputs_142__2), .inputs_142__1 (registerOutputs_142__1), .inputs_142__0 (
            registerOutputs_142__0), .inputs_143__15 (registerOutputs_143__15), 
            .inputs_143__14 (registerOutputs_143__14), .inputs_143__13 (
            registerOutputs_143__13), .inputs_143__12 (registerOutputs_143__12)
            , .inputs_143__11 (registerOutputs_143__11), .inputs_143__10 (
            registerOutputs_143__10), .inputs_143__9 (registerOutputs_143__9), .inputs_143__8 (
            registerOutputs_143__8), .inputs_143__7 (registerOutputs_143__7), .inputs_143__6 (
            registerOutputs_143__6), .inputs_143__5 (registerOutputs_143__5), .inputs_143__4 (
            registerOutputs_143__4), .inputs_143__3 (registerOutputs_143__3), .inputs_143__2 (
            registerOutputs_143__2), .inputs_143__1 (registerOutputs_143__1), .inputs_143__0 (
            registerOutputs_143__0), .inputs_144__15 (registerOutputs_144__15), 
            .inputs_144__14 (registerOutputs_144__14), .inputs_144__13 (
            registerOutputs_144__13), .inputs_144__12 (registerOutputs_144__12)
            , .inputs_144__11 (registerOutputs_144__11), .inputs_144__10 (
            registerOutputs_144__10), .inputs_144__9 (registerOutputs_144__9), .inputs_144__8 (
            registerOutputs_144__8), .inputs_144__7 (registerOutputs_144__7), .inputs_144__6 (
            registerOutputs_144__6), .inputs_144__5 (registerOutputs_144__5), .inputs_144__4 (
            registerOutputs_144__4), .inputs_144__3 (registerOutputs_144__3), .inputs_144__2 (
            registerOutputs_144__2), .inputs_144__1 (registerOutputs_144__1), .inputs_144__0 (
            registerOutputs_144__0), .inputs_145__15 (registerOutputs_145__15), 
            .inputs_145__14 (registerOutputs_145__14), .inputs_145__13 (
            registerOutputs_145__13), .inputs_145__12 (registerOutputs_145__12)
            , .inputs_145__11 (registerOutputs_145__11), .inputs_145__10 (
            registerOutputs_145__10), .inputs_145__9 (registerOutputs_145__9), .inputs_145__8 (
            registerOutputs_145__8), .inputs_145__7 (registerOutputs_145__7), .inputs_145__6 (
            registerOutputs_145__6), .inputs_145__5 (registerOutputs_145__5), .inputs_145__4 (
            registerOutputs_145__4), .inputs_145__3 (registerOutputs_145__3), .inputs_145__2 (
            registerOutputs_145__2), .inputs_145__1 (registerOutputs_145__1), .inputs_145__0 (
            registerOutputs_145__0), .inputs_146__15 (registerOutputs_146__15), 
            .inputs_146__14 (registerOutputs_146__14), .inputs_146__13 (
            registerOutputs_146__13), .inputs_146__12 (registerOutputs_146__12)
            , .inputs_146__11 (registerOutputs_146__11), .inputs_146__10 (
            registerOutputs_146__10), .inputs_146__9 (registerOutputs_146__9), .inputs_146__8 (
            registerOutputs_146__8), .inputs_146__7 (registerOutputs_146__7), .inputs_146__6 (
            registerOutputs_146__6), .inputs_146__5 (registerOutputs_146__5), .inputs_146__4 (
            registerOutputs_146__4), .inputs_146__3 (registerOutputs_146__3), .inputs_146__2 (
            registerOutputs_146__2), .inputs_146__1 (registerOutputs_146__1), .inputs_146__0 (
            registerOutputs_146__0), .inputs_147__15 (registerOutputs_147__15), 
            .inputs_147__14 (registerOutputs_147__14), .inputs_147__13 (
            registerOutputs_147__13), .inputs_147__12 (registerOutputs_147__12)
            , .inputs_147__11 (registerOutputs_147__11), .inputs_147__10 (
            registerOutputs_147__10), .inputs_147__9 (registerOutputs_147__9), .inputs_147__8 (
            registerOutputs_147__8), .inputs_147__7 (registerOutputs_147__7), .inputs_147__6 (
            registerOutputs_147__6), .inputs_147__5 (registerOutputs_147__5), .inputs_147__4 (
            registerOutputs_147__4), .inputs_147__3 (registerOutputs_147__3), .inputs_147__2 (
            registerOutputs_147__2), .inputs_147__1 (registerOutputs_147__1), .inputs_147__0 (
            registerOutputs_147__0), .inputs_148__15 (registerOutputs_148__15), 
            .inputs_148__14 (registerOutputs_148__14), .inputs_148__13 (
            registerOutputs_148__13), .inputs_148__12 (registerOutputs_148__12)
            , .inputs_148__11 (registerOutputs_148__11), .inputs_148__10 (
            registerOutputs_148__10), .inputs_148__9 (registerOutputs_148__9), .inputs_148__8 (
            registerOutputs_148__8), .inputs_148__7 (registerOutputs_148__7), .inputs_148__6 (
            registerOutputs_148__6), .inputs_148__5 (registerOutputs_148__5), .inputs_148__4 (
            registerOutputs_148__4), .inputs_148__3 (registerOutputs_148__3), .inputs_148__2 (
            registerOutputs_148__2), .inputs_148__1 (registerOutputs_148__1), .inputs_148__0 (
            registerOutputs_148__0), .inputs_149__15 (registerOutputs_149__15), 
            .inputs_149__14 (registerOutputs_149__14), .inputs_149__13 (
            registerOutputs_149__13), .inputs_149__12 (registerOutputs_149__12)
            , .inputs_149__11 (registerOutputs_149__11), .inputs_149__10 (
            registerOutputs_149__10), .inputs_149__9 (registerOutputs_149__9), .inputs_149__8 (
            registerOutputs_149__8), .inputs_149__7 (registerOutputs_149__7), .inputs_149__6 (
            registerOutputs_149__6), .inputs_149__5 (registerOutputs_149__5), .inputs_149__4 (
            registerOutputs_149__4), .inputs_149__3 (registerOutputs_149__3), .inputs_149__2 (
            registerOutputs_149__2), .inputs_149__1 (registerOutputs_149__1), .inputs_149__0 (
            registerOutputs_149__0), .inputs_150__15 (registerOutputs_150__15), 
            .inputs_150__14 (registerOutputs_150__14), .inputs_150__13 (
            registerOutputs_150__13), .inputs_150__12 (registerOutputs_150__12)
            , .inputs_150__11 (registerOutputs_150__11), .inputs_150__10 (
            registerOutputs_150__10), .inputs_150__9 (registerOutputs_150__9), .inputs_150__8 (
            registerOutputs_150__8), .inputs_150__7 (registerOutputs_150__7), .inputs_150__6 (
            registerOutputs_150__6), .inputs_150__5 (registerOutputs_150__5), .inputs_150__4 (
            registerOutputs_150__4), .inputs_150__3 (registerOutputs_150__3), .inputs_150__2 (
            registerOutputs_150__2), .inputs_150__1 (registerOutputs_150__1), .inputs_150__0 (
            registerOutputs_150__0), .inputs_151__15 (registerOutputs_151__15), 
            .inputs_151__14 (registerOutputs_151__14), .inputs_151__13 (
            registerOutputs_151__13), .inputs_151__12 (registerOutputs_151__12)
            , .inputs_151__11 (registerOutputs_151__11), .inputs_151__10 (
            registerOutputs_151__10), .inputs_151__9 (registerOutputs_151__9), .inputs_151__8 (
            registerOutputs_151__8), .inputs_151__7 (registerOutputs_151__7), .inputs_151__6 (
            registerOutputs_151__6), .inputs_151__5 (registerOutputs_151__5), .inputs_151__4 (
            registerOutputs_151__4), .inputs_151__3 (registerOutputs_151__3), .inputs_151__2 (
            registerOutputs_151__2), .inputs_151__1 (registerOutputs_151__1), .inputs_151__0 (
            registerOutputs_151__0), .inputs_152__15 (registerOutputs_152__15), 
            .inputs_152__14 (registerOutputs_152__14), .inputs_152__13 (
            registerOutputs_152__13), .inputs_152__12 (registerOutputs_152__12)
            , .inputs_152__11 (registerOutputs_152__11), .inputs_152__10 (
            registerOutputs_152__10), .inputs_152__9 (registerOutputs_152__9), .inputs_152__8 (
            registerOutputs_152__8), .inputs_152__7 (registerOutputs_152__7), .inputs_152__6 (
            registerOutputs_152__6), .inputs_152__5 (registerOutputs_152__5), .inputs_152__4 (
            registerOutputs_152__4), .inputs_152__3 (registerOutputs_152__3), .inputs_152__2 (
            registerOutputs_152__2), .inputs_152__1 (registerOutputs_152__1), .inputs_152__0 (
            registerOutputs_152__0), .inputs_153__15 (registerOutputs_153__15), 
            .inputs_153__14 (registerOutputs_153__14), .inputs_153__13 (
            registerOutputs_153__13), .inputs_153__12 (registerOutputs_153__12)
            , .inputs_153__11 (registerOutputs_153__11), .inputs_153__10 (
            registerOutputs_153__10), .inputs_153__9 (registerOutputs_153__9), .inputs_153__8 (
            registerOutputs_153__8), .inputs_153__7 (registerOutputs_153__7), .inputs_153__6 (
            registerOutputs_153__6), .inputs_153__5 (registerOutputs_153__5), .inputs_153__4 (
            registerOutputs_153__4), .inputs_153__3 (registerOutputs_153__3), .inputs_153__2 (
            registerOutputs_153__2), .inputs_153__1 (registerOutputs_153__1), .inputs_153__0 (
            registerOutputs_153__0), .inputs_154__15 (registerOutputs_154__15), 
            .inputs_154__14 (registerOutputs_154__14), .inputs_154__13 (
            registerOutputs_154__13), .inputs_154__12 (registerOutputs_154__12)
            , .inputs_154__11 (registerOutputs_154__11), .inputs_154__10 (
            registerOutputs_154__10), .inputs_154__9 (registerOutputs_154__9), .inputs_154__8 (
            registerOutputs_154__8), .inputs_154__7 (registerOutputs_154__7), .inputs_154__6 (
            registerOutputs_154__6), .inputs_154__5 (registerOutputs_154__5), .inputs_154__4 (
            registerOutputs_154__4), .inputs_154__3 (registerOutputs_154__3), .inputs_154__2 (
            registerOutputs_154__2), .inputs_154__1 (registerOutputs_154__1), .inputs_154__0 (
            registerOutputs_154__0), .inputs_155__15 (registerOutputs_155__15), 
            .inputs_155__14 (registerOutputs_155__14), .inputs_155__13 (
            registerOutputs_155__13), .inputs_155__12 (registerOutputs_155__12)
            , .inputs_155__11 (registerOutputs_155__11), .inputs_155__10 (
            registerOutputs_155__10), .inputs_155__9 (registerOutputs_155__9), .inputs_155__8 (
            registerOutputs_155__8), .inputs_155__7 (registerOutputs_155__7), .inputs_155__6 (
            registerOutputs_155__6), .inputs_155__5 (registerOutputs_155__5), .inputs_155__4 (
            registerOutputs_155__4), .inputs_155__3 (registerOutputs_155__3), .inputs_155__2 (
            registerOutputs_155__2), .inputs_155__1 (registerOutputs_155__1), .inputs_155__0 (
            registerOutputs_155__0), .inputs_156__15 (registerOutputs_156__15), 
            .inputs_156__14 (registerOutputs_156__14), .inputs_156__13 (
            registerOutputs_156__13), .inputs_156__12 (registerOutputs_156__12)
            , .inputs_156__11 (registerOutputs_156__11), .inputs_156__10 (
            registerOutputs_156__10), .inputs_156__9 (registerOutputs_156__9), .inputs_156__8 (
            registerOutputs_156__8), .inputs_156__7 (registerOutputs_156__7), .inputs_156__6 (
            registerOutputs_156__6), .inputs_156__5 (registerOutputs_156__5), .inputs_156__4 (
            registerOutputs_156__4), .inputs_156__3 (registerOutputs_156__3), .inputs_156__2 (
            registerOutputs_156__2), .inputs_156__1 (registerOutputs_156__1), .inputs_156__0 (
            registerOutputs_156__0), .inputs_157__15 (registerOutputs_157__15), 
            .inputs_157__14 (registerOutputs_157__14), .inputs_157__13 (
            registerOutputs_157__13), .inputs_157__12 (registerOutputs_157__12)
            , .inputs_157__11 (registerOutputs_157__11), .inputs_157__10 (
            registerOutputs_157__10), .inputs_157__9 (registerOutputs_157__9), .inputs_157__8 (
            registerOutputs_157__8), .inputs_157__7 (registerOutputs_157__7), .inputs_157__6 (
            registerOutputs_157__6), .inputs_157__5 (registerOutputs_157__5), .inputs_157__4 (
            registerOutputs_157__4), .inputs_157__3 (registerOutputs_157__3), .inputs_157__2 (
            registerOutputs_157__2), .inputs_157__1 (registerOutputs_157__1), .inputs_157__0 (
            registerOutputs_157__0), .inputs_158__15 (registerOutputs_158__15), 
            .inputs_158__14 (registerOutputs_158__14), .inputs_158__13 (
            registerOutputs_158__13), .inputs_158__12 (registerOutputs_158__12)
            , .inputs_158__11 (registerOutputs_158__11), .inputs_158__10 (
            registerOutputs_158__10), .inputs_158__9 (registerOutputs_158__9), .inputs_158__8 (
            registerOutputs_158__8), .inputs_158__7 (registerOutputs_158__7), .inputs_158__6 (
            registerOutputs_158__6), .inputs_158__5 (registerOutputs_158__5), .inputs_158__4 (
            registerOutputs_158__4), .inputs_158__3 (registerOutputs_158__3), .inputs_158__2 (
            registerOutputs_158__2), .inputs_158__1 (registerOutputs_158__1), .inputs_158__0 (
            registerOutputs_158__0), .inputs_159__15 (registerOutputs_159__15), 
            .inputs_159__14 (registerOutputs_159__14), .inputs_159__13 (
            registerOutputs_159__13), .inputs_159__12 (registerOutputs_159__12)
            , .inputs_159__11 (registerOutputs_159__11), .inputs_159__10 (
            registerOutputs_159__10), .inputs_159__9 (registerOutputs_159__9), .inputs_159__8 (
            registerOutputs_159__8), .inputs_159__7 (registerOutputs_159__7), .inputs_159__6 (
            registerOutputs_159__6), .inputs_159__5 (registerOutputs_159__5), .inputs_159__4 (
            registerOutputs_159__4), .inputs_159__3 (registerOutputs_159__3), .inputs_159__2 (
            registerOutputs_159__2), .inputs_159__1 (registerOutputs_159__1), .inputs_159__0 (
            registerOutputs_159__0), .inputs_160__15 (registerOutputs_160__15), 
            .inputs_160__14 (registerOutputs_160__14), .inputs_160__13 (
            registerOutputs_160__13), .inputs_160__12 (registerOutputs_160__12)
            , .inputs_160__11 (registerOutputs_160__11), .inputs_160__10 (
            registerOutputs_160__10), .inputs_160__9 (registerOutputs_160__9), .inputs_160__8 (
            registerOutputs_160__8), .inputs_160__7 (registerOutputs_160__7), .inputs_160__6 (
            registerOutputs_160__6), .inputs_160__5 (registerOutputs_160__5), .inputs_160__4 (
            registerOutputs_160__4), .inputs_160__3 (registerOutputs_160__3), .inputs_160__2 (
            registerOutputs_160__2), .inputs_160__1 (registerOutputs_160__1), .inputs_160__0 (
            registerOutputs_160__0), .inputs_161__15 (registerOutputs_161__15), 
            .inputs_161__14 (registerOutputs_161__14), .inputs_161__13 (
            registerOutputs_161__13), .inputs_161__12 (registerOutputs_161__12)
            , .inputs_161__11 (registerOutputs_161__11), .inputs_161__10 (
            registerOutputs_161__10), .inputs_161__9 (registerOutputs_161__9), .inputs_161__8 (
            registerOutputs_161__8), .inputs_161__7 (registerOutputs_161__7), .inputs_161__6 (
            registerOutputs_161__6), .inputs_161__5 (registerOutputs_161__5), .inputs_161__4 (
            registerOutputs_161__4), .inputs_161__3 (registerOutputs_161__3), .inputs_161__2 (
            registerOutputs_161__2), .inputs_161__1 (registerOutputs_161__1), .inputs_161__0 (
            registerOutputs_161__0), .inputs_162__15 (registerOutputs_162__15), 
            .inputs_162__14 (registerOutputs_162__14), .inputs_162__13 (
            registerOutputs_162__13), .inputs_162__12 (registerOutputs_162__12)
            , .inputs_162__11 (registerOutputs_162__11), .inputs_162__10 (
            registerOutputs_162__10), .inputs_162__9 (registerOutputs_162__9), .inputs_162__8 (
            registerOutputs_162__8), .inputs_162__7 (registerOutputs_162__7), .inputs_162__6 (
            registerOutputs_162__6), .inputs_162__5 (registerOutputs_162__5), .inputs_162__4 (
            registerOutputs_162__4), .inputs_162__3 (registerOutputs_162__3), .inputs_162__2 (
            registerOutputs_162__2), .inputs_162__1 (registerOutputs_162__1), .inputs_162__0 (
            registerOutputs_162__0), .inputs_163__15 (registerOutputs_163__15), 
            .inputs_163__14 (registerOutputs_163__14), .inputs_163__13 (
            registerOutputs_163__13), .inputs_163__12 (registerOutputs_163__12)
            , .inputs_163__11 (registerOutputs_163__11), .inputs_163__10 (
            registerOutputs_163__10), .inputs_163__9 (registerOutputs_163__9), .inputs_163__8 (
            registerOutputs_163__8), .inputs_163__7 (registerOutputs_163__7), .inputs_163__6 (
            registerOutputs_163__6), .inputs_163__5 (registerOutputs_163__5), .inputs_163__4 (
            registerOutputs_163__4), .inputs_163__3 (registerOutputs_163__3), .inputs_163__2 (
            registerOutputs_163__2), .inputs_163__1 (registerOutputs_163__1), .inputs_163__0 (
            registerOutputs_163__0), .inputs_164__15 (registerOutputs_164__15), 
            .inputs_164__14 (registerOutputs_164__14), .inputs_164__13 (
            registerOutputs_164__13), .inputs_164__12 (registerOutputs_164__12)
            , .inputs_164__11 (registerOutputs_164__11), .inputs_164__10 (
            registerOutputs_164__10), .inputs_164__9 (registerOutputs_164__9), .inputs_164__8 (
            registerOutputs_164__8), .inputs_164__7 (registerOutputs_164__7), .inputs_164__6 (
            registerOutputs_164__6), .inputs_164__5 (registerOutputs_164__5), .inputs_164__4 (
            registerOutputs_164__4), .inputs_164__3 (registerOutputs_164__3), .inputs_164__2 (
            registerOutputs_164__2), .inputs_164__1 (registerOutputs_164__1), .inputs_164__0 (
            registerOutputs_164__0), .inputs_165__15 (registerOutputs_165__15), 
            .inputs_165__14 (registerOutputs_165__14), .inputs_165__13 (
            registerOutputs_165__13), .inputs_165__12 (registerOutputs_165__12)
            , .inputs_165__11 (registerOutputs_165__11), .inputs_165__10 (
            registerOutputs_165__10), .inputs_165__9 (registerOutputs_165__9), .inputs_165__8 (
            registerOutputs_165__8), .inputs_165__7 (registerOutputs_165__7), .inputs_165__6 (
            registerOutputs_165__6), .inputs_165__5 (registerOutputs_165__5), .inputs_165__4 (
            registerOutputs_165__4), .inputs_165__3 (registerOutputs_165__3), .inputs_165__2 (
            registerOutputs_165__2), .inputs_165__1 (registerOutputs_165__1), .inputs_165__0 (
            registerOutputs_165__0), .inputs_166__15 (registerOutputs_166__15), 
            .inputs_166__14 (registerOutputs_166__14), .inputs_166__13 (
            registerOutputs_166__13), .inputs_166__12 (registerOutputs_166__12)
            , .inputs_166__11 (registerOutputs_166__11), .inputs_166__10 (
            registerOutputs_166__10), .inputs_166__9 (registerOutputs_166__9), .inputs_166__8 (
            registerOutputs_166__8), .inputs_166__7 (registerOutputs_166__7), .inputs_166__6 (
            registerOutputs_166__6), .inputs_166__5 (registerOutputs_166__5), .inputs_166__4 (
            registerOutputs_166__4), .inputs_166__3 (registerOutputs_166__3), .inputs_166__2 (
            registerOutputs_166__2), .inputs_166__1 (registerOutputs_166__1), .inputs_166__0 (
            registerOutputs_166__0), .inputs_167__15 (registerOutputs_167__15), 
            .inputs_167__14 (registerOutputs_167__14), .inputs_167__13 (
            registerOutputs_167__13), .inputs_167__12 (registerOutputs_167__12)
            , .inputs_167__11 (registerOutputs_167__11), .inputs_167__10 (
            registerOutputs_167__10), .inputs_167__9 (registerOutputs_167__9), .inputs_167__8 (
            registerOutputs_167__8), .inputs_167__7 (registerOutputs_167__7), .inputs_167__6 (
            registerOutputs_167__6), .inputs_167__5 (registerOutputs_167__5), .inputs_167__4 (
            registerOutputs_167__4), .inputs_167__3 (registerOutputs_167__3), .inputs_167__2 (
            registerOutputs_167__2), .inputs_167__1 (registerOutputs_167__1), .inputs_167__0 (
            registerOutputs_167__0), .inputs_168__15 (registerOutputs_168__15), 
            .inputs_168__14 (registerOutputs_168__14), .inputs_168__13 (
            registerOutputs_168__13), .inputs_168__12 (registerOutputs_168__12)
            , .inputs_168__11 (registerOutputs_168__11), .inputs_168__10 (
            registerOutputs_168__10), .inputs_168__9 (registerOutputs_168__9), .inputs_168__8 (
            registerOutputs_168__8), .inputs_168__7 (registerOutputs_168__7), .inputs_168__6 (
            registerOutputs_168__6), .inputs_168__5 (registerOutputs_168__5), .inputs_168__4 (
            registerOutputs_168__4), .inputs_168__3 (registerOutputs_168__3), .inputs_168__2 (
            registerOutputs_168__2), .inputs_168__1 (registerOutputs_168__1), .inputs_168__0 (
            registerOutputs_168__0), .inputs_169__15 (registerOutputs_169__15), 
            .inputs_169__14 (registerOutputs_169__14), .inputs_169__13 (
            registerOutputs_169__13), .inputs_169__12 (registerOutputs_169__12)
            , .inputs_169__11 (registerOutputs_169__11), .inputs_169__10 (
            registerOutputs_169__10), .inputs_169__9 (registerOutputs_169__9), .inputs_169__8 (
            registerOutputs_169__8), .inputs_169__7 (registerOutputs_169__7), .inputs_169__6 (
            registerOutputs_169__6), .inputs_169__5 (registerOutputs_169__5), .inputs_169__4 (
            registerOutputs_169__4), .inputs_169__3 (registerOutputs_169__3), .inputs_169__2 (
            registerOutputs_169__2), .inputs_169__1 (registerOutputs_169__1), .inputs_169__0 (
            registerOutputs_169__0), .inputs_170__15 (registerOutputs_170__15), 
            .inputs_170__14 (registerOutputs_170__14), .inputs_170__13 (
            registerOutputs_170__13), .inputs_170__12 (registerOutputs_170__12)
            , .inputs_170__11 (registerOutputs_170__11), .inputs_170__10 (
            registerOutputs_170__10), .inputs_170__9 (registerOutputs_170__9), .inputs_170__8 (
            registerOutputs_170__8), .inputs_170__7 (registerOutputs_170__7), .inputs_170__6 (
            registerOutputs_170__6), .inputs_170__5 (registerOutputs_170__5), .inputs_170__4 (
            registerOutputs_170__4), .inputs_170__3 (registerOutputs_170__3), .inputs_170__2 (
            registerOutputs_170__2), .inputs_170__1 (registerOutputs_170__1), .inputs_170__0 (
            registerOutputs_170__0), .inputs_171__15 (registerOutputs_171__15), 
            .inputs_171__14 (registerOutputs_171__14), .inputs_171__13 (
            registerOutputs_171__13), .inputs_171__12 (registerOutputs_171__12)
            , .inputs_171__11 (registerOutputs_171__11), .inputs_171__10 (
            registerOutputs_171__10), .inputs_171__9 (registerOutputs_171__9), .inputs_171__8 (
            registerOutputs_171__8), .inputs_171__7 (registerOutputs_171__7), .inputs_171__6 (
            registerOutputs_171__6), .inputs_171__5 (registerOutputs_171__5), .inputs_171__4 (
            registerOutputs_171__4), .inputs_171__3 (registerOutputs_171__3), .inputs_171__2 (
            registerOutputs_171__2), .inputs_171__1 (registerOutputs_171__1), .inputs_171__0 (
            registerOutputs_171__0), .inputs_172__15 (registerOutputs_172__15), 
            .inputs_172__14 (registerOutputs_172__14), .inputs_172__13 (
            registerOutputs_172__13), .inputs_172__12 (registerOutputs_172__12)
            , .inputs_172__11 (registerOutputs_172__11), .inputs_172__10 (
            registerOutputs_172__10), .inputs_172__9 (registerOutputs_172__9), .inputs_172__8 (
            registerOutputs_172__8), .inputs_172__7 (registerOutputs_172__7), .inputs_172__6 (
            registerOutputs_172__6), .inputs_172__5 (registerOutputs_172__5), .inputs_172__4 (
            registerOutputs_172__4), .inputs_172__3 (registerOutputs_172__3), .inputs_172__2 (
            registerOutputs_172__2), .inputs_172__1 (registerOutputs_172__1), .inputs_172__0 (
            registerOutputs_172__0), .inputs_173__15 (registerOutputs_173__15), 
            .inputs_173__14 (registerOutputs_173__14), .inputs_173__13 (
            registerOutputs_173__13), .inputs_173__12 (registerOutputs_173__12)
            , .inputs_173__11 (registerOutputs_173__11), .inputs_173__10 (
            registerOutputs_173__10), .inputs_173__9 (registerOutputs_173__9), .inputs_173__8 (
            registerOutputs_173__8), .inputs_173__7 (registerOutputs_173__7), .inputs_173__6 (
            registerOutputs_173__6), .inputs_173__5 (registerOutputs_173__5), .inputs_173__4 (
            registerOutputs_173__4), .inputs_173__3 (registerOutputs_173__3), .inputs_173__2 (
            registerOutputs_173__2), .inputs_173__1 (registerOutputs_173__1), .inputs_173__0 (
            registerOutputs_173__0), .inputs_174__15 (registerOutputs_174__15), 
            .inputs_174__14 (registerOutputs_174__14), .inputs_174__13 (
            registerOutputs_174__13), .inputs_174__12 (registerOutputs_174__12)
            , .inputs_174__11 (registerOutputs_174__11), .inputs_174__10 (
            registerOutputs_174__10), .inputs_174__9 (registerOutputs_174__9), .inputs_174__8 (
            registerOutputs_174__8), .inputs_174__7 (registerOutputs_174__7), .inputs_174__6 (
            registerOutputs_174__6), .inputs_174__5 (registerOutputs_174__5), .inputs_174__4 (
            registerOutputs_174__4), .inputs_174__3 (registerOutputs_174__3), .inputs_174__2 (
            registerOutputs_174__2), .inputs_174__1 (registerOutputs_174__1), .inputs_174__0 (
            registerOutputs_174__0), .inputs_175__15 (registerOutputs_175__15), 
            .inputs_175__14 (registerOutputs_175__14), .inputs_175__13 (
            registerOutputs_175__13), .inputs_175__12 (registerOutputs_175__12)
            , .inputs_175__11 (registerOutputs_175__11), .inputs_175__10 (
            registerOutputs_175__10), .inputs_175__9 (registerOutputs_175__9), .inputs_175__8 (
            registerOutputs_175__8), .inputs_175__7 (registerOutputs_175__7), .inputs_175__6 (
            registerOutputs_175__6), .inputs_175__5 (registerOutputs_175__5), .inputs_175__4 (
            registerOutputs_175__4), .inputs_175__3 (registerOutputs_175__3), .inputs_175__2 (
            registerOutputs_175__2), .inputs_175__1 (registerOutputs_175__1), .inputs_175__0 (
            registerOutputs_175__0), .inputs_176__15 (registerOutputs_176__15), 
            .inputs_176__14 (registerOutputs_176__14), .inputs_176__13 (
            registerOutputs_176__13), .inputs_176__12 (registerOutputs_176__12)
            , .inputs_176__11 (registerOutputs_176__11), .inputs_176__10 (
            registerOutputs_176__10), .inputs_176__9 (registerOutputs_176__9), .inputs_176__8 (
            registerOutputs_176__8), .inputs_176__7 (registerOutputs_176__7), .inputs_176__6 (
            registerOutputs_176__6), .inputs_176__5 (registerOutputs_176__5), .inputs_176__4 (
            registerOutputs_176__4), .inputs_176__3 (registerOutputs_176__3), .inputs_176__2 (
            registerOutputs_176__2), .inputs_176__1 (registerOutputs_176__1), .inputs_176__0 (
            registerOutputs_176__0), .inputs_177__15 (registerOutputs_177__15), 
            .inputs_177__14 (registerOutputs_177__14), .inputs_177__13 (
            registerOutputs_177__13), .inputs_177__12 (registerOutputs_177__12)
            , .inputs_177__11 (registerOutputs_177__11), .inputs_177__10 (
            registerOutputs_177__10), .inputs_177__9 (registerOutputs_177__9), .inputs_177__8 (
            registerOutputs_177__8), .inputs_177__7 (registerOutputs_177__7), .inputs_177__6 (
            registerOutputs_177__6), .inputs_177__5 (registerOutputs_177__5), .inputs_177__4 (
            registerOutputs_177__4), .inputs_177__3 (registerOutputs_177__3), .inputs_177__2 (
            registerOutputs_177__2), .inputs_177__1 (registerOutputs_177__1), .inputs_177__0 (
            registerOutputs_177__0), .inputs_178__15 (registerOutputs_178__15), 
            .inputs_178__14 (registerOutputs_178__14), .inputs_178__13 (
            registerOutputs_178__13), .inputs_178__12 (registerOutputs_178__12)
            , .inputs_178__11 (registerOutputs_178__11), .inputs_178__10 (
            registerOutputs_178__10), .inputs_178__9 (registerOutputs_178__9), .inputs_178__8 (
            registerOutputs_178__8), .inputs_178__7 (registerOutputs_178__7), .inputs_178__6 (
            registerOutputs_178__6), .inputs_178__5 (registerOutputs_178__5), .inputs_178__4 (
            registerOutputs_178__4), .inputs_178__3 (registerOutputs_178__3), .inputs_178__2 (
            registerOutputs_178__2), .inputs_178__1 (registerOutputs_178__1), .inputs_178__0 (
            registerOutputs_178__0), .inputs_179__15 (registerOutputs_179__15), 
            .inputs_179__14 (registerOutputs_179__14), .inputs_179__13 (
            registerOutputs_179__13), .inputs_179__12 (registerOutputs_179__12)
            , .inputs_179__11 (registerOutputs_179__11), .inputs_179__10 (
            registerOutputs_179__10), .inputs_179__9 (registerOutputs_179__9), .inputs_179__8 (
            registerOutputs_179__8), .inputs_179__7 (registerOutputs_179__7), .inputs_179__6 (
            registerOutputs_179__6), .inputs_179__5 (registerOutputs_179__5), .inputs_179__4 (
            registerOutputs_179__4), .inputs_179__3 (registerOutputs_179__3), .inputs_179__2 (
            registerOutputs_179__2), .inputs_179__1 (registerOutputs_179__1), .inputs_179__0 (
            registerOutputs_179__0), .inputs_180__15 (registerOutputs_180__15), 
            .inputs_180__14 (registerOutputs_180__14), .inputs_180__13 (
            registerOutputs_180__13), .inputs_180__12 (registerOutputs_180__12)
            , .inputs_180__11 (registerOutputs_180__11), .inputs_180__10 (
            registerOutputs_180__10), .inputs_180__9 (registerOutputs_180__9), .inputs_180__8 (
            registerOutputs_180__8), .inputs_180__7 (registerOutputs_180__7), .inputs_180__6 (
            registerOutputs_180__6), .inputs_180__5 (registerOutputs_180__5), .inputs_180__4 (
            registerOutputs_180__4), .inputs_180__3 (registerOutputs_180__3), .inputs_180__2 (
            registerOutputs_180__2), .inputs_180__1 (registerOutputs_180__1), .inputs_180__0 (
            registerOutputs_180__0), .inputs_181__15 (registerOutputs_181__15), 
            .inputs_181__14 (registerOutputs_181__14), .inputs_181__13 (
            registerOutputs_181__13), .inputs_181__12 (registerOutputs_181__12)
            , .inputs_181__11 (registerOutputs_181__11), .inputs_181__10 (
            registerOutputs_181__10), .inputs_181__9 (registerOutputs_181__9), .inputs_181__8 (
            registerOutputs_181__8), .inputs_181__7 (registerOutputs_181__7), .inputs_181__6 (
            registerOutputs_181__6), .inputs_181__5 (registerOutputs_181__5), .inputs_181__4 (
            registerOutputs_181__4), .inputs_181__3 (registerOutputs_181__3), .inputs_181__2 (
            registerOutputs_181__2), .inputs_181__1 (registerOutputs_181__1), .inputs_181__0 (
            registerOutputs_181__0), .inputs_182__15 (registerOutputs_182__15), 
            .inputs_182__14 (registerOutputs_182__14), .inputs_182__13 (
            registerOutputs_182__13), .inputs_182__12 (registerOutputs_182__12)
            , .inputs_182__11 (registerOutputs_182__11), .inputs_182__10 (
            registerOutputs_182__10), .inputs_182__9 (registerOutputs_182__9), .inputs_182__8 (
            registerOutputs_182__8), .inputs_182__7 (registerOutputs_182__7), .inputs_182__6 (
            registerOutputs_182__6), .inputs_182__5 (registerOutputs_182__5), .inputs_182__4 (
            registerOutputs_182__4), .inputs_182__3 (registerOutputs_182__3), .inputs_182__2 (
            registerOutputs_182__2), .inputs_182__1 (registerOutputs_182__1), .inputs_182__0 (
            registerOutputs_182__0), .inputs_183__15 (registerOutputs_183__15), 
            .inputs_183__14 (registerOutputs_183__14), .inputs_183__13 (
            registerOutputs_183__13), .inputs_183__12 (registerOutputs_183__12)
            , .inputs_183__11 (registerOutputs_183__11), .inputs_183__10 (
            registerOutputs_183__10), .inputs_183__9 (registerOutputs_183__9), .inputs_183__8 (
            registerOutputs_183__8), .inputs_183__7 (registerOutputs_183__7), .inputs_183__6 (
            registerOutputs_183__6), .inputs_183__5 (registerOutputs_183__5), .inputs_183__4 (
            registerOutputs_183__4), .inputs_183__3 (registerOutputs_183__3), .inputs_183__2 (
            registerOutputs_183__2), .inputs_183__1 (registerOutputs_183__1), .inputs_183__0 (
            registerOutputs_183__0), .inputs_184__15 (registerOutputs_184__15), 
            .inputs_184__14 (registerOutputs_184__14), .inputs_184__13 (
            registerOutputs_184__13), .inputs_184__12 (registerOutputs_184__12)
            , .inputs_184__11 (registerOutputs_184__11), .inputs_184__10 (
            registerOutputs_184__10), .inputs_184__9 (registerOutputs_184__9), .inputs_184__8 (
            registerOutputs_184__8), .inputs_184__7 (registerOutputs_184__7), .inputs_184__6 (
            registerOutputs_184__6), .inputs_184__5 (registerOutputs_184__5), .inputs_184__4 (
            registerOutputs_184__4), .inputs_184__3 (registerOutputs_184__3), .inputs_184__2 (
            registerOutputs_184__2), .inputs_184__1 (registerOutputs_184__1), .inputs_184__0 (
            registerOutputs_184__0), .inputs_185__15 (registerOutputs_185__15), 
            .inputs_185__14 (registerOutputs_185__14), .inputs_185__13 (
            registerOutputs_185__13), .inputs_185__12 (registerOutputs_185__12)
            , .inputs_185__11 (registerOutputs_185__11), .inputs_185__10 (
            registerOutputs_185__10), .inputs_185__9 (registerOutputs_185__9), .inputs_185__8 (
            registerOutputs_185__8), .inputs_185__7 (registerOutputs_185__7), .inputs_185__6 (
            registerOutputs_185__6), .inputs_185__5 (registerOutputs_185__5), .inputs_185__4 (
            registerOutputs_185__4), .inputs_185__3 (registerOutputs_185__3), .inputs_185__2 (
            registerOutputs_185__2), .inputs_185__1 (registerOutputs_185__1), .inputs_185__0 (
            registerOutputs_185__0), .inputs_186__15 (registerOutputs_186__15), 
            .inputs_186__14 (registerOutputs_186__14), .inputs_186__13 (
            registerOutputs_186__13), .inputs_186__12 (registerOutputs_186__12)
            , .inputs_186__11 (registerOutputs_186__11), .inputs_186__10 (
            registerOutputs_186__10), .inputs_186__9 (registerOutputs_186__9), .inputs_186__8 (
            registerOutputs_186__8), .inputs_186__7 (registerOutputs_186__7), .inputs_186__6 (
            registerOutputs_186__6), .inputs_186__5 (registerOutputs_186__5), .inputs_186__4 (
            registerOutputs_186__4), .inputs_186__3 (registerOutputs_186__3), .inputs_186__2 (
            registerOutputs_186__2), .inputs_186__1 (registerOutputs_186__1), .inputs_186__0 (
            registerOutputs_186__0), .inputs_187__15 (registerOutputs_187__15), 
            .inputs_187__14 (registerOutputs_187__14), .inputs_187__13 (
            registerOutputs_187__13), .inputs_187__12 (registerOutputs_187__12)
            , .inputs_187__11 (registerOutputs_187__11), .inputs_187__10 (
            registerOutputs_187__10), .inputs_187__9 (registerOutputs_187__9), .inputs_187__8 (
            registerOutputs_187__8), .inputs_187__7 (registerOutputs_187__7), .inputs_187__6 (
            registerOutputs_187__6), .inputs_187__5 (registerOutputs_187__5), .inputs_187__4 (
            registerOutputs_187__4), .inputs_187__3 (registerOutputs_187__3), .inputs_187__2 (
            registerOutputs_187__2), .inputs_187__1 (registerOutputs_187__1), .inputs_187__0 (
            registerOutputs_187__0), .inputs_188__15 (registerOutputs_188__15), 
            .inputs_188__14 (registerOutputs_188__14), .inputs_188__13 (
            registerOutputs_188__13), .inputs_188__12 (registerOutputs_188__12)
            , .inputs_188__11 (registerOutputs_188__11), .inputs_188__10 (
            registerOutputs_188__10), .inputs_188__9 (registerOutputs_188__9), .inputs_188__8 (
            registerOutputs_188__8), .inputs_188__7 (registerOutputs_188__7), .inputs_188__6 (
            registerOutputs_188__6), .inputs_188__5 (registerOutputs_188__5), .inputs_188__4 (
            registerOutputs_188__4), .inputs_188__3 (registerOutputs_188__3), .inputs_188__2 (
            registerOutputs_188__2), .inputs_188__1 (registerOutputs_188__1), .inputs_188__0 (
            registerOutputs_188__0), .inputs_189__15 (registerOutputs_189__15), 
            .inputs_189__14 (registerOutputs_189__14), .inputs_189__13 (
            registerOutputs_189__13), .inputs_189__12 (registerOutputs_189__12)
            , .inputs_189__11 (registerOutputs_189__11), .inputs_189__10 (
            registerOutputs_189__10), .inputs_189__9 (registerOutputs_189__9), .inputs_189__8 (
            registerOutputs_189__8), .inputs_189__7 (registerOutputs_189__7), .inputs_189__6 (
            registerOutputs_189__6), .inputs_189__5 (registerOutputs_189__5), .inputs_189__4 (
            registerOutputs_189__4), .inputs_189__3 (registerOutputs_189__3), .inputs_189__2 (
            registerOutputs_189__2), .inputs_189__1 (registerOutputs_189__1), .inputs_189__0 (
            registerOutputs_189__0), .inputs_190__15 (registerOutputs_190__15), 
            .inputs_190__14 (registerOutputs_190__14), .inputs_190__13 (
            registerOutputs_190__13), .inputs_190__12 (registerOutputs_190__12)
            , .inputs_190__11 (registerOutputs_190__11), .inputs_190__10 (
            registerOutputs_190__10), .inputs_190__9 (registerOutputs_190__9), .inputs_190__8 (
            registerOutputs_190__8), .inputs_190__7 (registerOutputs_190__7), .inputs_190__6 (
            registerOutputs_190__6), .inputs_190__5 (registerOutputs_190__5), .inputs_190__4 (
            registerOutputs_190__4), .inputs_190__3 (registerOutputs_190__3), .inputs_190__2 (
            registerOutputs_190__2), .inputs_190__1 (registerOutputs_190__1), .inputs_190__0 (
            registerOutputs_190__0), .inputs_191__15 (registerOutputs_191__15), 
            .inputs_191__14 (registerOutputs_191__14), .inputs_191__13 (
            registerOutputs_191__13), .inputs_191__12 (registerOutputs_191__12)
            , .inputs_191__11 (registerOutputs_191__11), .inputs_191__10 (
            registerOutputs_191__10), .inputs_191__9 (registerOutputs_191__9), .inputs_191__8 (
            registerOutputs_191__8), .inputs_191__7 (registerOutputs_191__7), .inputs_191__6 (
            registerOutputs_191__6), .inputs_191__5 (registerOutputs_191__5), .inputs_191__4 (
            registerOutputs_191__4), .inputs_191__3 (registerOutputs_191__3), .inputs_191__2 (
            registerOutputs_191__2), .inputs_191__1 (registerOutputs_191__1), .inputs_191__0 (
            registerOutputs_191__0), .inputs_192__15 (registerOutputs_192__15), 
            .inputs_192__14 (registerOutputs_192__14), .inputs_192__13 (
            registerOutputs_192__13), .inputs_192__12 (registerOutputs_192__12)
            , .inputs_192__11 (registerOutputs_192__11), .inputs_192__10 (
            registerOutputs_192__10), .inputs_192__9 (registerOutputs_192__9), .inputs_192__8 (
            registerOutputs_192__8), .inputs_192__7 (registerOutputs_192__7), .inputs_192__6 (
            registerOutputs_192__6), .inputs_192__5 (registerOutputs_192__5), .inputs_192__4 (
            registerOutputs_192__4), .inputs_192__3 (registerOutputs_192__3), .inputs_192__2 (
            registerOutputs_192__2), .inputs_192__1 (registerOutputs_192__1), .inputs_192__0 (
            registerOutputs_192__0), .inputs_193__15 (registerOutputs_193__15), 
            .inputs_193__14 (registerOutputs_193__14), .inputs_193__13 (
            registerOutputs_193__13), .inputs_193__12 (registerOutputs_193__12)
            , .inputs_193__11 (registerOutputs_193__11), .inputs_193__10 (
            registerOutputs_193__10), .inputs_193__9 (registerOutputs_193__9), .inputs_193__8 (
            registerOutputs_193__8), .inputs_193__7 (registerOutputs_193__7), .inputs_193__6 (
            registerOutputs_193__6), .inputs_193__5 (registerOutputs_193__5), .inputs_193__4 (
            registerOutputs_193__4), .inputs_193__3 (registerOutputs_193__3), .inputs_193__2 (
            registerOutputs_193__2), .inputs_193__1 (registerOutputs_193__1), .inputs_193__0 (
            registerOutputs_193__0), .inputs_194__15 (registerOutputs_194__15), 
            .inputs_194__14 (registerOutputs_194__14), .inputs_194__13 (
            registerOutputs_194__13), .inputs_194__12 (registerOutputs_194__12)
            , .inputs_194__11 (registerOutputs_194__11), .inputs_194__10 (
            registerOutputs_194__10), .inputs_194__9 (registerOutputs_194__9), .inputs_194__8 (
            registerOutputs_194__8), .inputs_194__7 (registerOutputs_194__7), .inputs_194__6 (
            registerOutputs_194__6), .inputs_194__5 (registerOutputs_194__5), .inputs_194__4 (
            registerOutputs_194__4), .inputs_194__3 (registerOutputs_194__3), .inputs_194__2 (
            registerOutputs_194__2), .inputs_194__1 (registerOutputs_194__1), .inputs_194__0 (
            registerOutputs_194__0), .inputs_195__15 (registerOutputs_195__15), 
            .inputs_195__14 (registerOutputs_195__14), .inputs_195__13 (
            registerOutputs_195__13), .inputs_195__12 (registerOutputs_195__12)
            , .inputs_195__11 (registerOutputs_195__11), .inputs_195__10 (
            registerOutputs_195__10), .inputs_195__9 (registerOutputs_195__9), .inputs_195__8 (
            registerOutputs_195__8), .inputs_195__7 (registerOutputs_195__7), .inputs_195__6 (
            registerOutputs_195__6), .inputs_195__5 (registerOutputs_195__5), .inputs_195__4 (
            registerOutputs_195__4), .inputs_195__3 (registerOutputs_195__3), .inputs_195__2 (
            registerOutputs_195__2), .inputs_195__1 (registerOutputs_195__1), .inputs_195__0 (
            registerOutputs_195__0), .inputs_196__15 (registerOutputs_196__15), 
            .inputs_196__14 (registerOutputs_196__14), .inputs_196__13 (
            registerOutputs_196__13), .inputs_196__12 (registerOutputs_196__12)
            , .inputs_196__11 (registerOutputs_196__11), .inputs_196__10 (
            registerOutputs_196__10), .inputs_196__9 (registerOutputs_196__9), .inputs_196__8 (
            registerOutputs_196__8), .inputs_196__7 (registerOutputs_196__7), .inputs_196__6 (
            registerOutputs_196__6), .inputs_196__5 (registerOutputs_196__5), .inputs_196__4 (
            registerOutputs_196__4), .inputs_196__3 (registerOutputs_196__3), .inputs_196__2 (
            registerOutputs_196__2), .inputs_196__1 (registerOutputs_196__1), .inputs_196__0 (
            registerOutputs_196__0), .inputs_197__15 (registerOutputs_197__15), 
            .inputs_197__14 (registerOutputs_197__14), .inputs_197__13 (
            registerOutputs_197__13), .inputs_197__12 (registerOutputs_197__12)
            , .inputs_197__11 (registerOutputs_197__11), .inputs_197__10 (
            registerOutputs_197__10), .inputs_197__9 (registerOutputs_197__9), .inputs_197__8 (
            registerOutputs_197__8), .inputs_197__7 (registerOutputs_197__7), .inputs_197__6 (
            registerOutputs_197__6), .inputs_197__5 (registerOutputs_197__5), .inputs_197__4 (
            registerOutputs_197__4), .inputs_197__3 (registerOutputs_197__3), .inputs_197__2 (
            registerOutputs_197__2), .inputs_197__1 (registerOutputs_197__1), .inputs_197__0 (
            registerOutputs_197__0), .inputs_198__15 (registerOutputs_198__15), 
            .inputs_198__14 (registerOutputs_198__14), .inputs_198__13 (
            registerOutputs_198__13), .inputs_198__12 (registerOutputs_198__12)
            , .inputs_198__11 (registerOutputs_198__11), .inputs_198__10 (
            registerOutputs_198__10), .inputs_198__9 (registerOutputs_198__9), .inputs_198__8 (
            registerOutputs_198__8), .inputs_198__7 (registerOutputs_198__7), .inputs_198__6 (
            registerOutputs_198__6), .inputs_198__5 (registerOutputs_198__5), .inputs_198__4 (
            registerOutputs_198__4), .inputs_198__3 (registerOutputs_198__3), .inputs_198__2 (
            registerOutputs_198__2), .inputs_198__1 (registerOutputs_198__1), .inputs_198__0 (
            registerOutputs_198__0), .inputs_199__15 (registerOutputs_199__15), 
            .inputs_199__14 (registerOutputs_199__14), .inputs_199__13 (
            registerOutputs_199__13), .inputs_199__12 (registerOutputs_199__12)
            , .inputs_199__11 (registerOutputs_199__11), .inputs_199__10 (
            registerOutputs_199__10), .inputs_199__9 (registerOutputs_199__9), .inputs_199__8 (
            registerOutputs_199__8), .inputs_199__7 (registerOutputs_199__7), .inputs_199__6 (
            registerOutputs_199__6), .inputs_199__5 (registerOutputs_199__5), .inputs_199__4 (
            registerOutputs_199__4), .inputs_199__3 (registerOutputs_199__3), .inputs_199__2 (
            registerOutputs_199__2), .inputs_199__1 (registerOutputs_199__1), .inputs_199__0 (
            registerOutputs_199__0), .inputs_200__15 (registerOutputs_200__15), 
            .inputs_200__14 (registerOutputs_200__14), .inputs_200__13 (
            registerOutputs_200__13), .inputs_200__12 (registerOutputs_200__12)
            , .inputs_200__11 (registerOutputs_200__11), .inputs_200__10 (
            registerOutputs_200__10), .inputs_200__9 (registerOutputs_200__9), .inputs_200__8 (
            registerOutputs_200__8), .inputs_200__7 (registerOutputs_200__7), .inputs_200__6 (
            registerOutputs_200__6), .inputs_200__5 (registerOutputs_200__5), .inputs_200__4 (
            registerOutputs_200__4), .inputs_200__3 (registerOutputs_200__3), .inputs_200__2 (
            registerOutputs_200__2), .inputs_200__1 (registerOutputs_200__1), .inputs_200__0 (
            registerOutputs_200__0), .inputs_201__15 (registerOutputs_201__15), 
            .inputs_201__14 (registerOutputs_201__14), .inputs_201__13 (
            registerOutputs_201__13), .inputs_201__12 (registerOutputs_201__12)
            , .inputs_201__11 (registerOutputs_201__11), .inputs_201__10 (
            registerOutputs_201__10), .inputs_201__9 (registerOutputs_201__9), .inputs_201__8 (
            registerOutputs_201__8), .inputs_201__7 (registerOutputs_201__7), .inputs_201__6 (
            registerOutputs_201__6), .inputs_201__5 (registerOutputs_201__5), .inputs_201__4 (
            registerOutputs_201__4), .inputs_201__3 (registerOutputs_201__3), .inputs_201__2 (
            registerOutputs_201__2), .inputs_201__1 (registerOutputs_201__1), .inputs_201__0 (
            registerOutputs_201__0), .inputs_202__15 (registerOutputs_202__15), 
            .inputs_202__14 (registerOutputs_202__14), .inputs_202__13 (
            registerOutputs_202__13), .inputs_202__12 (registerOutputs_202__12)
            , .inputs_202__11 (registerOutputs_202__11), .inputs_202__10 (
            registerOutputs_202__10), .inputs_202__9 (registerOutputs_202__9), .inputs_202__8 (
            registerOutputs_202__8), .inputs_202__7 (registerOutputs_202__7), .inputs_202__6 (
            registerOutputs_202__6), .inputs_202__5 (registerOutputs_202__5), .inputs_202__4 (
            registerOutputs_202__4), .inputs_202__3 (registerOutputs_202__3), .inputs_202__2 (
            registerOutputs_202__2), .inputs_202__1 (registerOutputs_202__1), .inputs_202__0 (
            registerOutputs_202__0), .inputs_203__15 (registerOutputs_203__15), 
            .inputs_203__14 (registerOutputs_203__14), .inputs_203__13 (
            registerOutputs_203__13), .inputs_203__12 (registerOutputs_203__12)
            , .inputs_203__11 (registerOutputs_203__11), .inputs_203__10 (
            registerOutputs_203__10), .inputs_203__9 (registerOutputs_203__9), .inputs_203__8 (
            registerOutputs_203__8), .inputs_203__7 (registerOutputs_203__7), .inputs_203__6 (
            registerOutputs_203__6), .inputs_203__5 (registerOutputs_203__5), .inputs_203__4 (
            registerOutputs_203__4), .inputs_203__3 (registerOutputs_203__3), .inputs_203__2 (
            registerOutputs_203__2), .inputs_203__1 (registerOutputs_203__1), .inputs_203__0 (
            registerOutputs_203__0), .inputs_204__15 (registerOutputs_204__15), 
            .inputs_204__14 (registerOutputs_204__14), .inputs_204__13 (
            registerOutputs_204__13), .inputs_204__12 (registerOutputs_204__12)
            , .inputs_204__11 (registerOutputs_204__11), .inputs_204__10 (
            registerOutputs_204__10), .inputs_204__9 (registerOutputs_204__9), .inputs_204__8 (
            registerOutputs_204__8), .inputs_204__7 (registerOutputs_204__7), .inputs_204__6 (
            registerOutputs_204__6), .inputs_204__5 (registerOutputs_204__5), .inputs_204__4 (
            registerOutputs_204__4), .inputs_204__3 (registerOutputs_204__3), .inputs_204__2 (
            registerOutputs_204__2), .inputs_204__1 (registerOutputs_204__1), .inputs_204__0 (
            registerOutputs_204__0), .inputs_205__15 (registerOutputs_205__15), 
            .inputs_205__14 (registerOutputs_205__14), .inputs_205__13 (
            registerOutputs_205__13), .inputs_205__12 (registerOutputs_205__12)
            , .inputs_205__11 (registerOutputs_205__11), .inputs_205__10 (
            registerOutputs_205__10), .inputs_205__9 (registerOutputs_205__9), .inputs_205__8 (
            registerOutputs_205__8), .inputs_205__7 (registerOutputs_205__7), .inputs_205__6 (
            registerOutputs_205__6), .inputs_205__5 (registerOutputs_205__5), .inputs_205__4 (
            registerOutputs_205__4), .inputs_205__3 (registerOutputs_205__3), .inputs_205__2 (
            registerOutputs_205__2), .inputs_205__1 (registerOutputs_205__1), .inputs_205__0 (
            registerOutputs_205__0), .inputs_206__15 (registerOutputs_206__15), 
            .inputs_206__14 (registerOutputs_206__14), .inputs_206__13 (
            registerOutputs_206__13), .inputs_206__12 (registerOutputs_206__12)
            , .inputs_206__11 (registerOutputs_206__11), .inputs_206__10 (
            registerOutputs_206__10), .inputs_206__9 (registerOutputs_206__9), .inputs_206__8 (
            registerOutputs_206__8), .inputs_206__7 (registerOutputs_206__7), .inputs_206__6 (
            registerOutputs_206__6), .inputs_206__5 (registerOutputs_206__5), .inputs_206__4 (
            registerOutputs_206__4), .inputs_206__3 (registerOutputs_206__3), .inputs_206__2 (
            registerOutputs_206__2), .inputs_206__1 (registerOutputs_206__1), .inputs_206__0 (
            registerOutputs_206__0), .inputs_207__15 (registerOutputs_207__15), 
            .inputs_207__14 (registerOutputs_207__14), .inputs_207__13 (
            registerOutputs_207__13), .inputs_207__12 (registerOutputs_207__12)
            , .inputs_207__11 (registerOutputs_207__11), .inputs_207__10 (
            registerOutputs_207__10), .inputs_207__9 (registerOutputs_207__9), .inputs_207__8 (
            registerOutputs_207__8), .inputs_207__7 (registerOutputs_207__7), .inputs_207__6 (
            registerOutputs_207__6), .inputs_207__5 (registerOutputs_207__5), .inputs_207__4 (
            registerOutputs_207__4), .inputs_207__3 (registerOutputs_207__3), .inputs_207__2 (
            registerOutputs_207__2), .inputs_207__1 (registerOutputs_207__1), .inputs_207__0 (
            registerOutputs_207__0), .inputs_208__15 (registerOutputs_208__15), 
            .inputs_208__14 (registerOutputs_208__14), .inputs_208__13 (
            registerOutputs_208__13), .inputs_208__12 (registerOutputs_208__12)
            , .inputs_208__11 (registerOutputs_208__11), .inputs_208__10 (
            registerOutputs_208__10), .inputs_208__9 (registerOutputs_208__9), .inputs_208__8 (
            registerOutputs_208__8), .inputs_208__7 (registerOutputs_208__7), .inputs_208__6 (
            registerOutputs_208__6), .inputs_208__5 (registerOutputs_208__5), .inputs_208__4 (
            registerOutputs_208__4), .inputs_208__3 (registerOutputs_208__3), .inputs_208__2 (
            registerOutputs_208__2), .inputs_208__1 (registerOutputs_208__1), .inputs_208__0 (
            registerOutputs_208__0), .inputs_209__15 (registerOutputs_209__15), 
            .inputs_209__14 (registerOutputs_209__14), .inputs_209__13 (
            registerOutputs_209__13), .inputs_209__12 (registerOutputs_209__12)
            , .inputs_209__11 (registerOutputs_209__11), .inputs_209__10 (
            registerOutputs_209__10), .inputs_209__9 (registerOutputs_209__9), .inputs_209__8 (
            registerOutputs_209__8), .inputs_209__7 (registerOutputs_209__7), .inputs_209__6 (
            registerOutputs_209__6), .inputs_209__5 (registerOutputs_209__5), .inputs_209__4 (
            registerOutputs_209__4), .inputs_209__3 (registerOutputs_209__3), .inputs_209__2 (
            registerOutputs_209__2), .inputs_209__1 (registerOutputs_209__1), .inputs_209__0 (
            registerOutputs_209__0), .inputs_210__15 (registerOutputs_210__15), 
            .inputs_210__14 (registerOutputs_210__14), .inputs_210__13 (
            registerOutputs_210__13), .inputs_210__12 (registerOutputs_210__12)
            , .inputs_210__11 (registerOutputs_210__11), .inputs_210__10 (
            registerOutputs_210__10), .inputs_210__9 (registerOutputs_210__9), .inputs_210__8 (
            registerOutputs_210__8), .inputs_210__7 (registerOutputs_210__7), .inputs_210__6 (
            registerOutputs_210__6), .inputs_210__5 (registerOutputs_210__5), .inputs_210__4 (
            registerOutputs_210__4), .inputs_210__3 (registerOutputs_210__3), .inputs_210__2 (
            registerOutputs_210__2), .inputs_210__1 (registerOutputs_210__1), .inputs_210__0 (
            registerOutputs_210__0), .inputs_211__15 (registerOutputs_211__15), 
            .inputs_211__14 (registerOutputs_211__14), .inputs_211__13 (
            registerOutputs_211__13), .inputs_211__12 (registerOutputs_211__12)
            , .inputs_211__11 (registerOutputs_211__11), .inputs_211__10 (
            registerOutputs_211__10), .inputs_211__9 (registerOutputs_211__9), .inputs_211__8 (
            registerOutputs_211__8), .inputs_211__7 (registerOutputs_211__7), .inputs_211__6 (
            registerOutputs_211__6), .inputs_211__5 (registerOutputs_211__5), .inputs_211__4 (
            registerOutputs_211__4), .inputs_211__3 (registerOutputs_211__3), .inputs_211__2 (
            registerOutputs_211__2), .inputs_211__1 (registerOutputs_211__1), .inputs_211__0 (
            registerOutputs_211__0), .inputs_212__15 (registerOutputs_212__15), 
            .inputs_212__14 (registerOutputs_212__14), .inputs_212__13 (
            registerOutputs_212__13), .inputs_212__12 (registerOutputs_212__12)
            , .inputs_212__11 (registerOutputs_212__11), .inputs_212__10 (
            registerOutputs_212__10), .inputs_212__9 (registerOutputs_212__9), .inputs_212__8 (
            registerOutputs_212__8), .inputs_212__7 (registerOutputs_212__7), .inputs_212__6 (
            registerOutputs_212__6), .inputs_212__5 (registerOutputs_212__5), .inputs_212__4 (
            registerOutputs_212__4), .inputs_212__3 (registerOutputs_212__3), .inputs_212__2 (
            registerOutputs_212__2), .inputs_212__1 (registerOutputs_212__1), .inputs_212__0 (
            registerOutputs_212__0), .inputs_213__15 (registerOutputs_213__15), 
            .inputs_213__14 (registerOutputs_213__14), .inputs_213__13 (
            registerOutputs_213__13), .inputs_213__12 (registerOutputs_213__12)
            , .inputs_213__11 (registerOutputs_213__11), .inputs_213__10 (
            registerOutputs_213__10), .inputs_213__9 (registerOutputs_213__9), .inputs_213__8 (
            registerOutputs_213__8), .inputs_213__7 (registerOutputs_213__7), .inputs_213__6 (
            registerOutputs_213__6), .inputs_213__5 (registerOutputs_213__5), .inputs_213__4 (
            registerOutputs_213__4), .inputs_213__3 (registerOutputs_213__3), .inputs_213__2 (
            registerOutputs_213__2), .inputs_213__1 (registerOutputs_213__1), .inputs_213__0 (
            registerOutputs_213__0), .inputs_214__15 (registerOutputs_214__15), 
            .inputs_214__14 (registerOutputs_214__14), .inputs_214__13 (
            registerOutputs_214__13), .inputs_214__12 (registerOutputs_214__12)
            , .inputs_214__11 (registerOutputs_214__11), .inputs_214__10 (
            registerOutputs_214__10), .inputs_214__9 (registerOutputs_214__9), .inputs_214__8 (
            registerOutputs_214__8), .inputs_214__7 (registerOutputs_214__7), .inputs_214__6 (
            registerOutputs_214__6), .inputs_214__5 (registerOutputs_214__5), .inputs_214__4 (
            registerOutputs_214__4), .inputs_214__3 (registerOutputs_214__3), .inputs_214__2 (
            registerOutputs_214__2), .inputs_214__1 (registerOutputs_214__1), .inputs_214__0 (
            registerOutputs_214__0), .inputs_215__15 (registerOutputs_215__15), 
            .inputs_215__14 (registerOutputs_215__14), .inputs_215__13 (
            registerOutputs_215__13), .inputs_215__12 (registerOutputs_215__12)
            , .inputs_215__11 (registerOutputs_215__11), .inputs_215__10 (
            registerOutputs_215__10), .inputs_215__9 (registerOutputs_215__9), .inputs_215__8 (
            registerOutputs_215__8), .inputs_215__7 (registerOutputs_215__7), .inputs_215__6 (
            registerOutputs_215__6), .inputs_215__5 (registerOutputs_215__5), .inputs_215__4 (
            registerOutputs_215__4), .inputs_215__3 (registerOutputs_215__3), .inputs_215__2 (
            registerOutputs_215__2), .inputs_215__1 (registerOutputs_215__1), .inputs_215__0 (
            registerOutputs_215__0), .inputs_216__15 (registerOutputs_216__15), 
            .inputs_216__14 (registerOutputs_216__14), .inputs_216__13 (
            registerOutputs_216__13), .inputs_216__12 (registerOutputs_216__12)
            , .inputs_216__11 (registerOutputs_216__11), .inputs_216__10 (
            registerOutputs_216__10), .inputs_216__9 (registerOutputs_216__9), .inputs_216__8 (
            registerOutputs_216__8), .inputs_216__7 (registerOutputs_216__7), .inputs_216__6 (
            registerOutputs_216__6), .inputs_216__5 (registerOutputs_216__5), .inputs_216__4 (
            registerOutputs_216__4), .inputs_216__3 (registerOutputs_216__3), .inputs_216__2 (
            registerOutputs_216__2), .inputs_216__1 (registerOutputs_216__1), .inputs_216__0 (
            registerOutputs_216__0), .inputs_217__15 (registerOutputs_217__15), 
            .inputs_217__14 (registerOutputs_217__14), .inputs_217__13 (
            registerOutputs_217__13), .inputs_217__12 (registerOutputs_217__12)
            , .inputs_217__11 (registerOutputs_217__11), .inputs_217__10 (
            registerOutputs_217__10), .inputs_217__9 (registerOutputs_217__9), .inputs_217__8 (
            registerOutputs_217__8), .inputs_217__7 (registerOutputs_217__7), .inputs_217__6 (
            registerOutputs_217__6), .inputs_217__5 (registerOutputs_217__5), .inputs_217__4 (
            registerOutputs_217__4), .inputs_217__3 (registerOutputs_217__3), .inputs_217__2 (
            registerOutputs_217__2), .inputs_217__1 (registerOutputs_217__1), .inputs_217__0 (
            registerOutputs_217__0), .inputs_218__15 (registerOutputs_218__15), 
            .inputs_218__14 (registerOutputs_218__14), .inputs_218__13 (
            registerOutputs_218__13), .inputs_218__12 (registerOutputs_218__12)
            , .inputs_218__11 (registerOutputs_218__11), .inputs_218__10 (
            registerOutputs_218__10), .inputs_218__9 (registerOutputs_218__9), .inputs_218__8 (
            registerOutputs_218__8), .inputs_218__7 (registerOutputs_218__7), .inputs_218__6 (
            registerOutputs_218__6), .inputs_218__5 (registerOutputs_218__5), .inputs_218__4 (
            registerOutputs_218__4), .inputs_218__3 (registerOutputs_218__3), .inputs_218__2 (
            registerOutputs_218__2), .inputs_218__1 (registerOutputs_218__1), .inputs_218__0 (
            registerOutputs_218__0), .inputs_219__15 (registerOutputs_219__15), 
            .inputs_219__14 (registerOutputs_219__14), .inputs_219__13 (
            registerOutputs_219__13), .inputs_219__12 (registerOutputs_219__12)
            , .inputs_219__11 (registerOutputs_219__11), .inputs_219__10 (
            registerOutputs_219__10), .inputs_219__9 (registerOutputs_219__9), .inputs_219__8 (
            registerOutputs_219__8), .inputs_219__7 (registerOutputs_219__7), .inputs_219__6 (
            registerOutputs_219__6), .inputs_219__5 (registerOutputs_219__5), .inputs_219__4 (
            registerOutputs_219__4), .inputs_219__3 (registerOutputs_219__3), .inputs_219__2 (
            registerOutputs_219__2), .inputs_219__1 (registerOutputs_219__1), .inputs_219__0 (
            registerOutputs_219__0), .inputs_220__15 (registerOutputs_220__15), 
            .inputs_220__14 (registerOutputs_220__14), .inputs_220__13 (
            registerOutputs_220__13), .inputs_220__12 (registerOutputs_220__12)
            , .inputs_220__11 (registerOutputs_220__11), .inputs_220__10 (
            registerOutputs_220__10), .inputs_220__9 (registerOutputs_220__9), .inputs_220__8 (
            registerOutputs_220__8), .inputs_220__7 (registerOutputs_220__7), .inputs_220__6 (
            registerOutputs_220__6), .inputs_220__5 (registerOutputs_220__5), .inputs_220__4 (
            registerOutputs_220__4), .inputs_220__3 (registerOutputs_220__3), .inputs_220__2 (
            registerOutputs_220__2), .inputs_220__1 (registerOutputs_220__1), .inputs_220__0 (
            registerOutputs_220__0), .inputs_221__15 (registerOutputs_221__15), 
            .inputs_221__14 (registerOutputs_221__14), .inputs_221__13 (
            registerOutputs_221__13), .inputs_221__12 (registerOutputs_221__12)
            , .inputs_221__11 (registerOutputs_221__11), .inputs_221__10 (
            registerOutputs_221__10), .inputs_221__9 (registerOutputs_221__9), .inputs_221__8 (
            registerOutputs_221__8), .inputs_221__7 (registerOutputs_221__7), .inputs_221__6 (
            registerOutputs_221__6), .inputs_221__5 (registerOutputs_221__5), .inputs_221__4 (
            registerOutputs_221__4), .inputs_221__3 (registerOutputs_221__3), .inputs_221__2 (
            registerOutputs_221__2), .inputs_221__1 (registerOutputs_221__1), .inputs_221__0 (
            registerOutputs_221__0), .inputs_222__15 (registerOutputs_222__15), 
            .inputs_222__14 (registerOutputs_222__14), .inputs_222__13 (
            registerOutputs_222__13), .inputs_222__12 (registerOutputs_222__12)
            , .inputs_222__11 (registerOutputs_222__11), .inputs_222__10 (
            registerOutputs_222__10), .inputs_222__9 (registerOutputs_222__9), .inputs_222__8 (
            registerOutputs_222__8), .inputs_222__7 (registerOutputs_222__7), .inputs_222__6 (
            registerOutputs_222__6), .inputs_222__5 (registerOutputs_222__5), .inputs_222__4 (
            registerOutputs_222__4), .inputs_222__3 (registerOutputs_222__3), .inputs_222__2 (
            registerOutputs_222__2), .inputs_222__1 (registerOutputs_222__1), .inputs_222__0 (
            registerOutputs_222__0), .inputs_223__15 (registerOutputs_223__15), 
            .inputs_223__14 (registerOutputs_223__14), .inputs_223__13 (
            registerOutputs_223__13), .inputs_223__12 (registerOutputs_223__12)
            , .inputs_223__11 (registerOutputs_223__11), .inputs_223__10 (
            registerOutputs_223__10), .inputs_223__9 (registerOutputs_223__9), .inputs_223__8 (
            registerOutputs_223__8), .inputs_223__7 (registerOutputs_223__7), .inputs_223__6 (
            registerOutputs_223__6), .inputs_223__5 (registerOutputs_223__5), .inputs_223__4 (
            registerOutputs_223__4), .inputs_223__3 (registerOutputs_223__3), .inputs_223__2 (
            registerOutputs_223__2), .inputs_223__1 (registerOutputs_223__1), .inputs_223__0 (
            registerOutputs_223__0), .inputs_224__15 (registerOutputs_224__15), 
            .inputs_224__14 (registerOutputs_224__14), .inputs_224__13 (
            registerOutputs_224__13), .inputs_224__12 (registerOutputs_224__12)
            , .inputs_224__11 (registerOutputs_224__11), .inputs_224__10 (
            registerOutputs_224__10), .inputs_224__9 (registerOutputs_224__9), .inputs_224__8 (
            registerOutputs_224__8), .inputs_224__7 (registerOutputs_224__7), .inputs_224__6 (
            registerOutputs_224__6), .inputs_224__5 (registerOutputs_224__5), .inputs_224__4 (
            registerOutputs_224__4), .inputs_224__3 (registerOutputs_224__3), .inputs_224__2 (
            registerOutputs_224__2), .inputs_224__1 (registerOutputs_224__1), .inputs_224__0 (
            registerOutputs_224__0), .inputs_225__15 (registerOutputs_225__15), 
            .inputs_225__14 (registerOutputs_225__14), .inputs_225__13 (
            registerOutputs_225__13), .inputs_225__12 (registerOutputs_225__12)
            , .inputs_225__11 (registerOutputs_225__11), .inputs_225__10 (
            registerOutputs_225__10), .inputs_225__9 (registerOutputs_225__9), .inputs_225__8 (
            registerOutputs_225__8), .inputs_225__7 (registerOutputs_225__7), .inputs_225__6 (
            registerOutputs_225__6), .inputs_225__5 (registerOutputs_225__5), .inputs_225__4 (
            registerOutputs_225__4), .inputs_225__3 (registerOutputs_225__3), .inputs_225__2 (
            registerOutputs_225__2), .inputs_225__1 (registerOutputs_225__1), .inputs_225__0 (
            registerOutputs_225__0), .inputs_226__15 (registerOutputs_226__15), 
            .inputs_226__14 (registerOutputs_226__14), .inputs_226__13 (
            registerOutputs_226__13), .inputs_226__12 (registerOutputs_226__12)
            , .inputs_226__11 (registerOutputs_226__11), .inputs_226__10 (
            registerOutputs_226__10), .inputs_226__9 (registerOutputs_226__9), .inputs_226__8 (
            registerOutputs_226__8), .inputs_226__7 (registerOutputs_226__7), .inputs_226__6 (
            registerOutputs_226__6), .inputs_226__5 (registerOutputs_226__5), .inputs_226__4 (
            registerOutputs_226__4), .inputs_226__3 (registerOutputs_226__3), .inputs_226__2 (
            registerOutputs_226__2), .inputs_226__1 (registerOutputs_226__1), .inputs_226__0 (
            registerOutputs_226__0), .inputs_227__15 (registerOutputs_227__15), 
            .inputs_227__14 (registerOutputs_227__14), .inputs_227__13 (
            registerOutputs_227__13), .inputs_227__12 (registerOutputs_227__12)
            , .inputs_227__11 (registerOutputs_227__11), .inputs_227__10 (
            registerOutputs_227__10), .inputs_227__9 (registerOutputs_227__9), .inputs_227__8 (
            registerOutputs_227__8), .inputs_227__7 (registerOutputs_227__7), .inputs_227__6 (
            registerOutputs_227__6), .inputs_227__5 (registerOutputs_227__5), .inputs_227__4 (
            registerOutputs_227__4), .inputs_227__3 (registerOutputs_227__3), .inputs_227__2 (
            registerOutputs_227__2), .inputs_227__1 (registerOutputs_227__1), .inputs_227__0 (
            registerOutputs_227__0), .inputs_228__15 (registerOutputs_228__15), 
            .inputs_228__14 (registerOutputs_228__14), .inputs_228__13 (
            registerOutputs_228__13), .inputs_228__12 (registerOutputs_228__12)
            , .inputs_228__11 (registerOutputs_228__11), .inputs_228__10 (
            registerOutputs_228__10), .inputs_228__9 (registerOutputs_228__9), .inputs_228__8 (
            registerOutputs_228__8), .inputs_228__7 (registerOutputs_228__7), .inputs_228__6 (
            registerOutputs_228__6), .inputs_228__5 (registerOutputs_228__5), .inputs_228__4 (
            registerOutputs_228__4), .inputs_228__3 (registerOutputs_228__3), .inputs_228__2 (
            registerOutputs_228__2), .inputs_228__1 (registerOutputs_228__1), .inputs_228__0 (
            registerOutputs_228__0), .inputs_229__15 (registerOutputs_229__15), 
            .inputs_229__14 (registerOutputs_229__14), .inputs_229__13 (
            registerOutputs_229__13), .inputs_229__12 (registerOutputs_229__12)
            , .inputs_229__11 (registerOutputs_229__11), .inputs_229__10 (
            registerOutputs_229__10), .inputs_229__9 (registerOutputs_229__9), .inputs_229__8 (
            registerOutputs_229__8), .inputs_229__7 (registerOutputs_229__7), .inputs_229__6 (
            registerOutputs_229__6), .inputs_229__5 (registerOutputs_229__5), .inputs_229__4 (
            registerOutputs_229__4), .inputs_229__3 (registerOutputs_229__3), .inputs_229__2 (
            registerOutputs_229__2), .inputs_229__1 (registerOutputs_229__1), .inputs_229__0 (
            registerOutputs_229__0), .inputs_230__15 (registerOutputs_230__15), 
            .inputs_230__14 (registerOutputs_230__14), .inputs_230__13 (
            registerOutputs_230__13), .inputs_230__12 (registerOutputs_230__12)
            , .inputs_230__11 (registerOutputs_230__11), .inputs_230__10 (
            registerOutputs_230__10), .inputs_230__9 (registerOutputs_230__9), .inputs_230__8 (
            registerOutputs_230__8), .inputs_230__7 (registerOutputs_230__7), .inputs_230__6 (
            registerOutputs_230__6), .inputs_230__5 (registerOutputs_230__5), .inputs_230__4 (
            registerOutputs_230__4), .inputs_230__3 (registerOutputs_230__3), .inputs_230__2 (
            registerOutputs_230__2), .inputs_230__1 (registerOutputs_230__1), .inputs_230__0 (
            registerOutputs_230__0), .inputs_231__15 (registerOutputs_231__15), 
            .inputs_231__14 (registerOutputs_231__14), .inputs_231__13 (
            registerOutputs_231__13), .inputs_231__12 (registerOutputs_231__12)
            , .inputs_231__11 (registerOutputs_231__11), .inputs_231__10 (
            registerOutputs_231__10), .inputs_231__9 (registerOutputs_231__9), .inputs_231__8 (
            registerOutputs_231__8), .inputs_231__7 (registerOutputs_231__7), .inputs_231__6 (
            registerOutputs_231__6), .inputs_231__5 (registerOutputs_231__5), .inputs_231__4 (
            registerOutputs_231__4), .inputs_231__3 (registerOutputs_231__3), .inputs_231__2 (
            registerOutputs_231__2), .inputs_231__1 (registerOutputs_231__1), .inputs_231__0 (
            registerOutputs_231__0), .inputs_232__15 (registerOutputs_232__15), 
            .inputs_232__14 (registerOutputs_232__14), .inputs_232__13 (
            registerOutputs_232__13), .inputs_232__12 (registerOutputs_232__12)
            , .inputs_232__11 (registerOutputs_232__11), .inputs_232__10 (
            registerOutputs_232__10), .inputs_232__9 (registerOutputs_232__9), .inputs_232__8 (
            registerOutputs_232__8), .inputs_232__7 (registerOutputs_232__7), .inputs_232__6 (
            registerOutputs_232__6), .inputs_232__5 (registerOutputs_232__5), .inputs_232__4 (
            registerOutputs_232__4), .inputs_232__3 (registerOutputs_232__3), .inputs_232__2 (
            registerOutputs_232__2), .inputs_232__1 (registerOutputs_232__1), .inputs_232__0 (
            registerOutputs_232__0), .inputs_233__15 (registerOutputs_233__15), 
            .inputs_233__14 (registerOutputs_233__14), .inputs_233__13 (
            registerOutputs_233__13), .inputs_233__12 (registerOutputs_233__12)
            , .inputs_233__11 (registerOutputs_233__11), .inputs_233__10 (
            registerOutputs_233__10), .inputs_233__9 (registerOutputs_233__9), .inputs_233__8 (
            registerOutputs_233__8), .inputs_233__7 (registerOutputs_233__7), .inputs_233__6 (
            registerOutputs_233__6), .inputs_233__5 (registerOutputs_233__5), .inputs_233__4 (
            registerOutputs_233__4), .inputs_233__3 (registerOutputs_233__3), .inputs_233__2 (
            registerOutputs_233__2), .inputs_233__1 (registerOutputs_233__1), .inputs_233__0 (
            registerOutputs_233__0), .inputs_234__15 (registerOutputs_234__15), 
            .inputs_234__14 (registerOutputs_234__14), .inputs_234__13 (
            registerOutputs_234__13), .inputs_234__12 (registerOutputs_234__12)
            , .inputs_234__11 (registerOutputs_234__11), .inputs_234__10 (
            registerOutputs_234__10), .inputs_234__9 (registerOutputs_234__9), .inputs_234__8 (
            registerOutputs_234__8), .inputs_234__7 (registerOutputs_234__7), .inputs_234__6 (
            registerOutputs_234__6), .inputs_234__5 (registerOutputs_234__5), .inputs_234__4 (
            registerOutputs_234__4), .inputs_234__3 (registerOutputs_234__3), .inputs_234__2 (
            registerOutputs_234__2), .inputs_234__1 (registerOutputs_234__1), .inputs_234__0 (
            registerOutputs_234__0), .inputs_235__15 (registerOutputs_235__15), 
            .inputs_235__14 (registerOutputs_235__14), .inputs_235__13 (
            registerOutputs_235__13), .inputs_235__12 (registerOutputs_235__12)
            , .inputs_235__11 (registerOutputs_235__11), .inputs_235__10 (
            registerOutputs_235__10), .inputs_235__9 (registerOutputs_235__9), .inputs_235__8 (
            registerOutputs_235__8), .inputs_235__7 (registerOutputs_235__7), .inputs_235__6 (
            registerOutputs_235__6), .inputs_235__5 (registerOutputs_235__5), .inputs_235__4 (
            registerOutputs_235__4), .inputs_235__3 (registerOutputs_235__3), .inputs_235__2 (
            registerOutputs_235__2), .inputs_235__1 (registerOutputs_235__1), .inputs_235__0 (
            registerOutputs_235__0), .inputs_236__15 (registerOutputs_236__15), 
            .inputs_236__14 (registerOutputs_236__14), .inputs_236__13 (
            registerOutputs_236__13), .inputs_236__12 (registerOutputs_236__12)
            , .inputs_236__11 (registerOutputs_236__11), .inputs_236__10 (
            registerOutputs_236__10), .inputs_236__9 (registerOutputs_236__9), .inputs_236__8 (
            registerOutputs_236__8), .inputs_236__7 (registerOutputs_236__7), .inputs_236__6 (
            registerOutputs_236__6), .inputs_236__5 (registerOutputs_236__5), .inputs_236__4 (
            registerOutputs_236__4), .inputs_236__3 (registerOutputs_236__3), .inputs_236__2 (
            registerOutputs_236__2), .inputs_236__1 (registerOutputs_236__1), .inputs_236__0 (
            registerOutputs_236__0), .inputs_237__15 (registerOutputs_237__15), 
            .inputs_237__14 (registerOutputs_237__14), .inputs_237__13 (
            registerOutputs_237__13), .inputs_237__12 (registerOutputs_237__12)
            , .inputs_237__11 (registerOutputs_237__11), .inputs_237__10 (
            registerOutputs_237__10), .inputs_237__9 (registerOutputs_237__9), .inputs_237__8 (
            registerOutputs_237__8), .inputs_237__7 (registerOutputs_237__7), .inputs_237__6 (
            registerOutputs_237__6), .inputs_237__5 (registerOutputs_237__5), .inputs_237__4 (
            registerOutputs_237__4), .inputs_237__3 (registerOutputs_237__3), .inputs_237__2 (
            registerOutputs_237__2), .inputs_237__1 (registerOutputs_237__1), .inputs_237__0 (
            registerOutputs_237__0), .inputs_238__15 (registerOutputs_238__15), 
            .inputs_238__14 (registerOutputs_238__14), .inputs_238__13 (
            registerOutputs_238__13), .inputs_238__12 (registerOutputs_238__12)
            , .inputs_238__11 (registerOutputs_238__11), .inputs_238__10 (
            registerOutputs_238__10), .inputs_238__9 (registerOutputs_238__9), .inputs_238__8 (
            registerOutputs_238__8), .inputs_238__7 (registerOutputs_238__7), .inputs_238__6 (
            registerOutputs_238__6), .inputs_238__5 (registerOutputs_238__5), .inputs_238__4 (
            registerOutputs_238__4), .inputs_238__3 (registerOutputs_238__3), .inputs_238__2 (
            registerOutputs_238__2), .inputs_238__1 (registerOutputs_238__1), .inputs_238__0 (
            registerOutputs_238__0), .inputs_239__15 (registerOutputs_239__15), 
            .inputs_239__14 (registerOutputs_239__14), .inputs_239__13 (
            registerOutputs_239__13), .inputs_239__12 (registerOutputs_239__12)
            , .inputs_239__11 (registerOutputs_239__11), .inputs_239__10 (
            registerOutputs_239__10), .inputs_239__9 (registerOutputs_239__9), .inputs_239__8 (
            registerOutputs_239__8), .inputs_239__7 (registerOutputs_239__7), .inputs_239__6 (
            registerOutputs_239__6), .inputs_239__5 (registerOutputs_239__5), .inputs_239__4 (
            registerOutputs_239__4), .inputs_239__3 (registerOutputs_239__3), .inputs_239__2 (
            registerOutputs_239__2), .inputs_239__1 (registerOutputs_239__1), .inputs_239__0 (
            registerOutputs_239__0), .inputs_240__15 (registerOutputs_240__15), 
            .inputs_240__14 (registerOutputs_240__14), .inputs_240__13 (
            registerOutputs_240__13), .inputs_240__12 (registerOutputs_240__12)
            , .inputs_240__11 (registerOutputs_240__11), .inputs_240__10 (
            registerOutputs_240__10), .inputs_240__9 (registerOutputs_240__9), .inputs_240__8 (
            registerOutputs_240__8), .inputs_240__7 (registerOutputs_240__7), .inputs_240__6 (
            registerOutputs_240__6), .inputs_240__5 (registerOutputs_240__5), .inputs_240__4 (
            registerOutputs_240__4), .inputs_240__3 (registerOutputs_240__3), .inputs_240__2 (
            registerOutputs_240__2), .inputs_240__1 (registerOutputs_240__1), .inputs_240__0 (
            registerOutputs_240__0), .inputs_241__15 (registerOutputs_241__15), 
            .inputs_241__14 (registerOutputs_241__14), .inputs_241__13 (
            registerOutputs_241__13), .inputs_241__12 (registerOutputs_241__12)
            , .inputs_241__11 (registerOutputs_241__11), .inputs_241__10 (
            registerOutputs_241__10), .inputs_241__9 (registerOutputs_241__9), .inputs_241__8 (
            registerOutputs_241__8), .inputs_241__7 (registerOutputs_241__7), .inputs_241__6 (
            registerOutputs_241__6), .inputs_241__5 (registerOutputs_241__5), .inputs_241__4 (
            registerOutputs_241__4), .inputs_241__3 (registerOutputs_241__3), .inputs_241__2 (
            registerOutputs_241__2), .inputs_241__1 (registerOutputs_241__1), .inputs_241__0 (
            registerOutputs_241__0), .inputs_242__15 (registerOutputs_242__15), 
            .inputs_242__14 (registerOutputs_242__14), .inputs_242__13 (
            registerOutputs_242__13), .inputs_242__12 (registerOutputs_242__12)
            , .inputs_242__11 (registerOutputs_242__11), .inputs_242__10 (
            registerOutputs_242__10), .inputs_242__9 (registerOutputs_242__9), .inputs_242__8 (
            registerOutputs_242__8), .inputs_242__7 (registerOutputs_242__7), .inputs_242__6 (
            registerOutputs_242__6), .inputs_242__5 (registerOutputs_242__5), .inputs_242__4 (
            registerOutputs_242__4), .inputs_242__3 (registerOutputs_242__3), .inputs_242__2 (
            registerOutputs_242__2), .inputs_242__1 (registerOutputs_242__1), .inputs_242__0 (
            registerOutputs_242__0), .inputs_243__15 (registerOutputs_243__15), 
            .inputs_243__14 (registerOutputs_243__14), .inputs_243__13 (
            registerOutputs_243__13), .inputs_243__12 (registerOutputs_243__12)
            , .inputs_243__11 (registerOutputs_243__11), .inputs_243__10 (
            registerOutputs_243__10), .inputs_243__9 (registerOutputs_243__9), .inputs_243__8 (
            registerOutputs_243__8), .inputs_243__7 (registerOutputs_243__7), .inputs_243__6 (
            registerOutputs_243__6), .inputs_243__5 (registerOutputs_243__5), .inputs_243__4 (
            registerOutputs_243__4), .inputs_243__3 (registerOutputs_243__3), .inputs_243__2 (
            registerOutputs_243__2), .inputs_243__1 (registerOutputs_243__1), .inputs_243__0 (
            registerOutputs_243__0), .inputs_244__15 (registerOutputs_244__15), 
            .inputs_244__14 (registerOutputs_244__14), .inputs_244__13 (
            registerOutputs_244__13), .inputs_244__12 (registerOutputs_244__12)
            , .inputs_244__11 (registerOutputs_244__11), .inputs_244__10 (
            registerOutputs_244__10), .inputs_244__9 (registerOutputs_244__9), .inputs_244__8 (
            registerOutputs_244__8), .inputs_244__7 (registerOutputs_244__7), .inputs_244__6 (
            registerOutputs_244__6), .inputs_244__5 (registerOutputs_244__5), .inputs_244__4 (
            registerOutputs_244__4), .inputs_244__3 (registerOutputs_244__3), .inputs_244__2 (
            registerOutputs_244__2), .inputs_244__1 (registerOutputs_244__1), .inputs_244__0 (
            registerOutputs_244__0), .inputs_245__15 (registerOutputs_245__15), 
            .inputs_245__14 (registerOutputs_245__14), .inputs_245__13 (
            registerOutputs_245__13), .inputs_245__12 (registerOutputs_245__12)
            , .inputs_245__11 (registerOutputs_245__11), .inputs_245__10 (
            registerOutputs_245__10), .inputs_245__9 (registerOutputs_245__9), .inputs_245__8 (
            registerOutputs_245__8), .inputs_245__7 (registerOutputs_245__7), .inputs_245__6 (
            registerOutputs_245__6), .inputs_245__5 (registerOutputs_245__5), .inputs_245__4 (
            registerOutputs_245__4), .inputs_245__3 (registerOutputs_245__3), .inputs_245__2 (
            registerOutputs_245__2), .inputs_245__1 (registerOutputs_245__1), .inputs_245__0 (
            registerOutputs_245__0), .inputs_246__15 (registerOutputs_246__15), 
            .inputs_246__14 (registerOutputs_246__14), .inputs_246__13 (
            registerOutputs_246__13), .inputs_246__12 (registerOutputs_246__12)
            , .inputs_246__11 (registerOutputs_246__11), .inputs_246__10 (
            registerOutputs_246__10), .inputs_246__9 (registerOutputs_246__9), .inputs_246__8 (
            registerOutputs_246__8), .inputs_246__7 (registerOutputs_246__7), .inputs_246__6 (
            registerOutputs_246__6), .inputs_246__5 (registerOutputs_246__5), .inputs_246__4 (
            registerOutputs_246__4), .inputs_246__3 (registerOutputs_246__3), .inputs_246__2 (
            registerOutputs_246__2), .inputs_246__1 (registerOutputs_246__1), .inputs_246__0 (
            registerOutputs_246__0), .inputs_247__15 (registerOutputs_247__15), 
            .inputs_247__14 (registerOutputs_247__14), .inputs_247__13 (
            registerOutputs_247__13), .inputs_247__12 (registerOutputs_247__12)
            , .inputs_247__11 (registerOutputs_247__11), .inputs_247__10 (
            registerOutputs_247__10), .inputs_247__9 (registerOutputs_247__9), .inputs_247__8 (
            registerOutputs_247__8), .inputs_247__7 (registerOutputs_247__7), .inputs_247__6 (
            registerOutputs_247__6), .inputs_247__5 (registerOutputs_247__5), .inputs_247__4 (
            registerOutputs_247__4), .inputs_247__3 (registerOutputs_247__3), .inputs_247__2 (
            registerOutputs_247__2), .inputs_247__1 (registerOutputs_247__1), .inputs_247__0 (
            registerOutputs_247__0), .inputs_248__15 (registerOutputs_248__15), 
            .inputs_248__14 (registerOutputs_248__14), .inputs_248__13 (
            registerOutputs_248__13), .inputs_248__12 (registerOutputs_248__12)
            , .inputs_248__11 (registerOutputs_248__11), .inputs_248__10 (
            registerOutputs_248__10), .inputs_248__9 (registerOutputs_248__9), .inputs_248__8 (
            registerOutputs_248__8), .inputs_248__7 (registerOutputs_248__7), .inputs_248__6 (
            registerOutputs_248__6), .inputs_248__5 (registerOutputs_248__5), .inputs_248__4 (
            registerOutputs_248__4), .inputs_248__3 (registerOutputs_248__3), .inputs_248__2 (
            registerOutputs_248__2), .inputs_248__1 (registerOutputs_248__1), .inputs_248__0 (
            registerOutputs_248__0), .inputs_249__15 (registerOutputs_249__15), 
            .inputs_249__14 (registerOutputs_249__14), .inputs_249__13 (
            registerOutputs_249__13), .inputs_249__12 (registerOutputs_249__12)
            , .inputs_249__11 (registerOutputs_249__11), .inputs_249__10 (
            registerOutputs_249__10), .inputs_249__9 (registerOutputs_249__9), .inputs_249__8 (
            registerOutputs_249__8), .inputs_249__7 (registerOutputs_249__7), .inputs_249__6 (
            registerOutputs_249__6), .inputs_249__5 (registerOutputs_249__5), .inputs_249__4 (
            registerOutputs_249__4), .inputs_249__3 (registerOutputs_249__3), .inputs_249__2 (
            registerOutputs_249__2), .inputs_249__1 (registerOutputs_249__1), .inputs_249__0 (
            registerOutputs_249__0), .inputs_250__15 (registerOutputs_250__15), 
            .inputs_250__14 (registerOutputs_250__14), .inputs_250__13 (
            registerOutputs_250__13), .inputs_250__12 (registerOutputs_250__12)
            , .inputs_250__11 (registerOutputs_250__11), .inputs_250__10 (
            registerOutputs_250__10), .inputs_250__9 (registerOutputs_250__9), .inputs_250__8 (
            registerOutputs_250__8), .inputs_250__7 (registerOutputs_250__7), .inputs_250__6 (
            registerOutputs_250__6), .inputs_250__5 (registerOutputs_250__5), .inputs_250__4 (
            registerOutputs_250__4), .inputs_250__3 (registerOutputs_250__3), .inputs_250__2 (
            registerOutputs_250__2), .inputs_250__1 (registerOutputs_250__1), .inputs_250__0 (
            registerOutputs_250__0), .inputs_251__15 (registerOutputs_251__15), 
            .inputs_251__14 (registerOutputs_251__14), .inputs_251__13 (
            registerOutputs_251__13), .inputs_251__12 (registerOutputs_251__12)
            , .inputs_251__11 (registerOutputs_251__11), .inputs_251__10 (
            registerOutputs_251__10), .inputs_251__9 (registerOutputs_251__9), .inputs_251__8 (
            registerOutputs_251__8), .inputs_251__7 (registerOutputs_251__7), .inputs_251__6 (
            registerOutputs_251__6), .inputs_251__5 (registerOutputs_251__5), .inputs_251__4 (
            registerOutputs_251__4), .inputs_251__3 (registerOutputs_251__3), .inputs_251__2 (
            registerOutputs_251__2), .inputs_251__1 (registerOutputs_251__1), .inputs_251__0 (
            registerOutputs_251__0), .inputs_252__15 (registerOutputs_252__15), 
            .inputs_252__14 (registerOutputs_252__14), .inputs_252__13 (
            registerOutputs_252__13), .inputs_252__12 (registerOutputs_252__12)
            , .inputs_252__11 (registerOutputs_252__11), .inputs_252__10 (
            registerOutputs_252__10), .inputs_252__9 (registerOutputs_252__9), .inputs_252__8 (
            registerOutputs_252__8), .inputs_252__7 (registerOutputs_252__7), .inputs_252__6 (
            registerOutputs_252__6), .inputs_252__5 (registerOutputs_252__5), .inputs_252__4 (
            registerOutputs_252__4), .inputs_252__3 (registerOutputs_252__3), .inputs_252__2 (
            registerOutputs_252__2), .inputs_252__1 (registerOutputs_252__1), .inputs_252__0 (
            registerOutputs_252__0), .inputs_253__15 (registerOutputs_253__15), 
            .inputs_253__14 (registerOutputs_253__14), .inputs_253__13 (
            registerOutputs_253__13), .inputs_253__12 (registerOutputs_253__12)
            , .inputs_253__11 (registerOutputs_253__11), .inputs_253__10 (
            registerOutputs_253__10), .inputs_253__9 (registerOutputs_253__9), .inputs_253__8 (
            registerOutputs_253__8), .inputs_253__7 (registerOutputs_253__7), .inputs_253__6 (
            registerOutputs_253__6), .inputs_253__5 (registerOutputs_253__5), .inputs_253__4 (
            registerOutputs_253__4), .inputs_253__3 (registerOutputs_253__3), .inputs_253__2 (
            registerOutputs_253__2), .inputs_253__1 (registerOutputs_253__1), .inputs_253__0 (
            registerOutputs_253__0), .inputs_254__15 (registerOutputs_254__15), 
            .inputs_254__14 (registerOutputs_254__14), .inputs_254__13 (
            registerOutputs_254__13), .inputs_254__12 (registerOutputs_254__12)
            , .inputs_254__11 (registerOutputs_254__11), .inputs_254__10 (
            registerOutputs_254__10), .inputs_254__9 (registerOutputs_254__9), .inputs_254__8 (
            registerOutputs_254__8), .inputs_254__7 (registerOutputs_254__7), .inputs_254__6 (
            registerOutputs_254__6), .inputs_254__5 (registerOutputs_254__5), .inputs_254__4 (
            registerOutputs_254__4), .inputs_254__3 (registerOutputs_254__3), .inputs_254__2 (
            registerOutputs_254__2), .inputs_254__1 (registerOutputs_254__1), .inputs_254__0 (
            registerOutputs_254__0), .inputs_255__15 (registerOutputs_255__15), 
            .inputs_255__14 (registerOutputs_255__14), .inputs_255__13 (
            registerOutputs_255__13), .inputs_255__12 (registerOutputs_255__12)
            , .inputs_255__11 (registerOutputs_255__11), .inputs_255__10 (
            registerOutputs_255__10), .inputs_255__9 (registerOutputs_255__9), .inputs_255__8 (
            registerOutputs_255__8), .inputs_255__7 (registerOutputs_255__7), .inputs_255__6 (
            registerOutputs_255__6), .inputs_255__5 (registerOutputs_255__5), .inputs_255__4 (
            registerOutputs_255__4), .inputs_255__3 (registerOutputs_255__3), .inputs_255__2 (
            registerOutputs_255__2), .inputs_255__1 (registerOutputs_255__1), .inputs_255__0 (
            registerOutputs_255__0), .inputs_256__15 (registerOutputs_256__15), 
            .inputs_256__14 (registerOutputs_256__14), .inputs_256__13 (
            registerOutputs_256__13), .inputs_256__12 (registerOutputs_256__12)
            , .inputs_256__11 (registerOutputs_256__11), .inputs_256__10 (
            registerOutputs_256__10), .inputs_256__9 (registerOutputs_256__9), .inputs_256__8 (
            registerOutputs_256__8), .inputs_256__7 (registerOutputs_256__7), .inputs_256__6 (
            registerOutputs_256__6), .inputs_256__5 (registerOutputs_256__5), .inputs_256__4 (
            registerOutputs_256__4), .inputs_256__3 (registerOutputs_256__3), .inputs_256__2 (
            registerOutputs_256__2), .inputs_256__1 (registerOutputs_256__1), .inputs_256__0 (
            registerOutputs_256__0), .inputs_257__15 (registerOutputs_257__15), 
            .inputs_257__14 (registerOutputs_257__14), .inputs_257__13 (
            registerOutputs_257__13), .inputs_257__12 (registerOutputs_257__12)
            , .inputs_257__11 (registerOutputs_257__11), .inputs_257__10 (
            registerOutputs_257__10), .inputs_257__9 (registerOutputs_257__9), .inputs_257__8 (
            registerOutputs_257__8), .inputs_257__7 (registerOutputs_257__7), .inputs_257__6 (
            registerOutputs_257__6), .inputs_257__5 (registerOutputs_257__5), .inputs_257__4 (
            registerOutputs_257__4), .inputs_257__3 (registerOutputs_257__3), .inputs_257__2 (
            registerOutputs_257__2), .inputs_257__1 (registerOutputs_257__1), .inputs_257__0 (
            registerOutputs_257__0), .inputs_258__15 (registerOutputs_258__15), 
            .inputs_258__14 (registerOutputs_258__14), .inputs_258__13 (
            registerOutputs_258__13), .inputs_258__12 (registerOutputs_258__12)
            , .inputs_258__11 (registerOutputs_258__11), .inputs_258__10 (
            registerOutputs_258__10), .inputs_258__9 (registerOutputs_258__9), .inputs_258__8 (
            registerOutputs_258__8), .inputs_258__7 (registerOutputs_258__7), .inputs_258__6 (
            registerOutputs_258__6), .inputs_258__5 (registerOutputs_258__5), .inputs_258__4 (
            registerOutputs_258__4), .inputs_258__3 (registerOutputs_258__3), .inputs_258__2 (
            registerOutputs_258__2), .inputs_258__1 (registerOutputs_258__1), .inputs_258__0 (
            registerOutputs_258__0), .inputs_259__15 (registerOutputs_259__15), 
            .inputs_259__14 (registerOutputs_259__14), .inputs_259__13 (
            registerOutputs_259__13), .inputs_259__12 (registerOutputs_259__12)
            , .inputs_259__11 (registerOutputs_259__11), .inputs_259__10 (
            registerOutputs_259__10), .inputs_259__9 (registerOutputs_259__9), .inputs_259__8 (
            registerOutputs_259__8), .inputs_259__7 (registerOutputs_259__7), .inputs_259__6 (
            registerOutputs_259__6), .inputs_259__5 (registerOutputs_259__5), .inputs_259__4 (
            registerOutputs_259__4), .inputs_259__3 (registerOutputs_259__3), .inputs_259__2 (
            registerOutputs_259__2), .inputs_259__1 (registerOutputs_259__1), .inputs_259__0 (
            registerOutputs_259__0), .inputs_260__15 (registerOutputs_260__15), 
            .inputs_260__14 (registerOutputs_260__14), .inputs_260__13 (
            registerOutputs_260__13), .inputs_260__12 (registerOutputs_260__12)
            , .inputs_260__11 (registerOutputs_260__11), .inputs_260__10 (
            registerOutputs_260__10), .inputs_260__9 (registerOutputs_260__9), .inputs_260__8 (
            registerOutputs_260__8), .inputs_260__7 (registerOutputs_260__7), .inputs_260__6 (
            registerOutputs_260__6), .inputs_260__5 (registerOutputs_260__5), .inputs_260__4 (
            registerOutputs_260__4), .inputs_260__3 (registerOutputs_260__3), .inputs_260__2 (
            registerOutputs_260__2), .inputs_260__1 (registerOutputs_260__1), .inputs_260__0 (
            registerOutputs_260__0), .inputs_261__15 (registerOutputs_261__15), 
            .inputs_261__14 (registerOutputs_261__14), .inputs_261__13 (
            registerOutputs_261__13), .inputs_261__12 (registerOutputs_261__12)
            , .inputs_261__11 (registerOutputs_261__11), .inputs_261__10 (
            registerOutputs_261__10), .inputs_261__9 (registerOutputs_261__9), .inputs_261__8 (
            registerOutputs_261__8), .inputs_261__7 (registerOutputs_261__7), .inputs_261__6 (
            registerOutputs_261__6), .inputs_261__5 (registerOutputs_261__5), .inputs_261__4 (
            registerOutputs_261__4), .inputs_261__3 (registerOutputs_261__3), .inputs_261__2 (
            registerOutputs_261__2), .inputs_261__1 (registerOutputs_261__1), .inputs_261__0 (
            registerOutputs_261__0), .inputs_262__15 (registerOutputs_262__15), 
            .inputs_262__14 (registerOutputs_262__14), .inputs_262__13 (
            registerOutputs_262__13), .inputs_262__12 (registerOutputs_262__12)
            , .inputs_262__11 (registerOutputs_262__11), .inputs_262__10 (
            registerOutputs_262__10), .inputs_262__9 (registerOutputs_262__9), .inputs_262__8 (
            registerOutputs_262__8), .inputs_262__7 (registerOutputs_262__7), .inputs_262__6 (
            registerOutputs_262__6), .inputs_262__5 (registerOutputs_262__5), .inputs_262__4 (
            registerOutputs_262__4), .inputs_262__3 (registerOutputs_262__3), .inputs_262__2 (
            registerOutputs_262__2), .inputs_262__1 (registerOutputs_262__1), .inputs_262__0 (
            registerOutputs_262__0), .inputs_263__15 (registerOutputs_263__15), 
            .inputs_263__14 (registerOutputs_263__14), .inputs_263__13 (
            registerOutputs_263__13), .inputs_263__12 (registerOutputs_263__12)
            , .inputs_263__11 (registerOutputs_263__11), .inputs_263__10 (
            registerOutputs_263__10), .inputs_263__9 (registerOutputs_263__9), .inputs_263__8 (
            registerOutputs_263__8), .inputs_263__7 (registerOutputs_263__7), .inputs_263__6 (
            registerOutputs_263__6), .inputs_263__5 (registerOutputs_263__5), .inputs_263__4 (
            registerOutputs_263__4), .inputs_263__3 (registerOutputs_263__3), .inputs_263__2 (
            registerOutputs_263__2), .inputs_263__1 (registerOutputs_263__1), .inputs_263__0 (
            registerOutputs_263__0), .inputs_264__15 (registerOutputs_264__15), 
            .inputs_264__14 (registerOutputs_264__14), .inputs_264__13 (
            registerOutputs_264__13), .inputs_264__12 (registerOutputs_264__12)
            , .inputs_264__11 (registerOutputs_264__11), .inputs_264__10 (
            registerOutputs_264__10), .inputs_264__9 (registerOutputs_264__9), .inputs_264__8 (
            registerOutputs_264__8), .inputs_264__7 (registerOutputs_264__7), .inputs_264__6 (
            registerOutputs_264__6), .inputs_264__5 (registerOutputs_264__5), .inputs_264__4 (
            registerOutputs_264__4), .inputs_264__3 (registerOutputs_264__3), .inputs_264__2 (
            registerOutputs_264__2), .inputs_264__1 (registerOutputs_264__1), .inputs_264__0 (
            registerOutputs_264__0), .inputs_265__15 (registerOutputs_265__15), 
            .inputs_265__14 (registerOutputs_265__14), .inputs_265__13 (
            registerOutputs_265__13), .inputs_265__12 (registerOutputs_265__12)
            , .inputs_265__11 (registerOutputs_265__11), .inputs_265__10 (
            registerOutputs_265__10), .inputs_265__9 (registerOutputs_265__9), .inputs_265__8 (
            registerOutputs_265__8), .inputs_265__7 (registerOutputs_265__7), .inputs_265__6 (
            registerOutputs_265__6), .inputs_265__5 (registerOutputs_265__5), .inputs_265__4 (
            registerOutputs_265__4), .inputs_265__3 (registerOutputs_265__3), .inputs_265__2 (
            registerOutputs_265__2), .inputs_265__1 (registerOutputs_265__1), .inputs_265__0 (
            registerOutputs_265__0), .inputs_266__15 (registerOutputs_266__15), 
            .inputs_266__14 (registerOutputs_266__14), .inputs_266__13 (
            registerOutputs_266__13), .inputs_266__12 (registerOutputs_266__12)
            , .inputs_266__11 (registerOutputs_266__11), .inputs_266__10 (
            registerOutputs_266__10), .inputs_266__9 (registerOutputs_266__9), .inputs_266__8 (
            registerOutputs_266__8), .inputs_266__7 (registerOutputs_266__7), .inputs_266__6 (
            registerOutputs_266__6), .inputs_266__5 (registerOutputs_266__5), .inputs_266__4 (
            registerOutputs_266__4), .inputs_266__3 (registerOutputs_266__3), .inputs_266__2 (
            registerOutputs_266__2), .inputs_266__1 (registerOutputs_266__1), .inputs_266__0 (
            registerOutputs_266__0), .inputs_267__15 (registerOutputs_267__15), 
            .inputs_267__14 (registerOutputs_267__14), .inputs_267__13 (
            registerOutputs_267__13), .inputs_267__12 (registerOutputs_267__12)
            , .inputs_267__11 (registerOutputs_267__11), .inputs_267__10 (
            registerOutputs_267__10), .inputs_267__9 (registerOutputs_267__9), .inputs_267__8 (
            registerOutputs_267__8), .inputs_267__7 (registerOutputs_267__7), .inputs_267__6 (
            registerOutputs_267__6), .inputs_267__5 (registerOutputs_267__5), .inputs_267__4 (
            registerOutputs_267__4), .inputs_267__3 (registerOutputs_267__3), .inputs_267__2 (
            registerOutputs_267__2), .inputs_267__1 (registerOutputs_267__1), .inputs_267__0 (
            registerOutputs_267__0), .inputs_268__15 (registerOutputs_268__15), 
            .inputs_268__14 (registerOutputs_268__14), .inputs_268__13 (
            registerOutputs_268__13), .inputs_268__12 (registerOutputs_268__12)
            , .inputs_268__11 (registerOutputs_268__11), .inputs_268__10 (
            registerOutputs_268__10), .inputs_268__9 (registerOutputs_268__9), .inputs_268__8 (
            registerOutputs_268__8), .inputs_268__7 (registerOutputs_268__7), .inputs_268__6 (
            registerOutputs_268__6), .inputs_268__5 (registerOutputs_268__5), .inputs_268__4 (
            registerOutputs_268__4), .inputs_268__3 (registerOutputs_268__3), .inputs_268__2 (
            registerOutputs_268__2), .inputs_268__1 (registerOutputs_268__1), .inputs_268__0 (
            registerOutputs_268__0), .inputs_269__15 (registerOutputs_269__15), 
            .inputs_269__14 (registerOutputs_269__14), .inputs_269__13 (
            registerOutputs_269__13), .inputs_269__12 (registerOutputs_269__12)
            , .inputs_269__11 (registerOutputs_269__11), .inputs_269__10 (
            registerOutputs_269__10), .inputs_269__9 (registerOutputs_269__9), .inputs_269__8 (
            registerOutputs_269__8), .inputs_269__7 (registerOutputs_269__7), .inputs_269__6 (
            registerOutputs_269__6), .inputs_269__5 (registerOutputs_269__5), .inputs_269__4 (
            registerOutputs_269__4), .inputs_269__3 (registerOutputs_269__3), .inputs_269__2 (
            registerOutputs_269__2), .inputs_269__1 (registerOutputs_269__1), .inputs_269__0 (
            registerOutputs_269__0), .inputs_270__15 (registerOutputs_270__15), 
            .inputs_270__14 (registerOutputs_270__14), .inputs_270__13 (
            registerOutputs_270__13), .inputs_270__12 (registerOutputs_270__12)
            , .inputs_270__11 (registerOutputs_270__11), .inputs_270__10 (
            registerOutputs_270__10), .inputs_270__9 (registerOutputs_270__9), .inputs_270__8 (
            registerOutputs_270__8), .inputs_270__7 (registerOutputs_270__7), .inputs_270__6 (
            registerOutputs_270__6), .inputs_270__5 (registerOutputs_270__5), .inputs_270__4 (
            registerOutputs_270__4), .inputs_270__3 (registerOutputs_270__3), .inputs_270__2 (
            registerOutputs_270__2), .inputs_270__1 (registerOutputs_270__1), .inputs_270__0 (
            registerOutputs_270__0), .inputs_271__15 (registerOutputs_271__15), 
            .inputs_271__14 (registerOutputs_271__14), .inputs_271__13 (
            registerOutputs_271__13), .inputs_271__12 (registerOutputs_271__12)
            , .inputs_271__11 (registerOutputs_271__11), .inputs_271__10 (
            registerOutputs_271__10), .inputs_271__9 (registerOutputs_271__9), .inputs_271__8 (
            registerOutputs_271__8), .inputs_271__7 (registerOutputs_271__7), .inputs_271__6 (
            registerOutputs_271__6), .inputs_271__5 (registerOutputs_271__5), .inputs_271__4 (
            registerOutputs_271__4), .inputs_271__3 (registerOutputs_271__3), .inputs_271__2 (
            registerOutputs_271__2), .inputs_271__1 (registerOutputs_271__1), .inputs_271__0 (
            registerOutputs_271__0), .inputs_272__15 (registerOutputs_272__15), 
            .inputs_272__14 (registerOutputs_272__14), .inputs_272__13 (
            registerOutputs_272__13), .inputs_272__12 (registerOutputs_272__12)
            , .inputs_272__11 (registerOutputs_272__11), .inputs_272__10 (
            registerOutputs_272__10), .inputs_272__9 (registerOutputs_272__9), .inputs_272__8 (
            registerOutputs_272__8), .inputs_272__7 (registerOutputs_272__7), .inputs_272__6 (
            registerOutputs_272__6), .inputs_272__5 (registerOutputs_272__5), .inputs_272__4 (
            registerOutputs_272__4), .inputs_272__3 (registerOutputs_272__3), .inputs_272__2 (
            registerOutputs_272__2), .inputs_272__1 (registerOutputs_272__1), .inputs_272__0 (
            registerOutputs_272__0), .inputs_273__15 (registerOutputs_273__15), 
            .inputs_273__14 (registerOutputs_273__14), .inputs_273__13 (
            registerOutputs_273__13), .inputs_273__12 (registerOutputs_273__12)
            , .inputs_273__11 (registerOutputs_273__11), .inputs_273__10 (
            registerOutputs_273__10), .inputs_273__9 (registerOutputs_273__9), .inputs_273__8 (
            registerOutputs_273__8), .inputs_273__7 (registerOutputs_273__7), .inputs_273__6 (
            registerOutputs_273__6), .inputs_273__5 (registerOutputs_273__5), .inputs_273__4 (
            registerOutputs_273__4), .inputs_273__3 (registerOutputs_273__3), .inputs_273__2 (
            registerOutputs_273__2), .inputs_273__1 (registerOutputs_273__1), .inputs_273__0 (
            registerOutputs_273__0), .inputs_274__15 (registerOutputs_274__15), 
            .inputs_274__14 (registerOutputs_274__14), .inputs_274__13 (
            registerOutputs_274__13), .inputs_274__12 (registerOutputs_274__12)
            , .inputs_274__11 (registerOutputs_274__11), .inputs_274__10 (
            registerOutputs_274__10), .inputs_274__9 (registerOutputs_274__9), .inputs_274__8 (
            registerOutputs_274__8), .inputs_274__7 (registerOutputs_274__7), .inputs_274__6 (
            registerOutputs_274__6), .inputs_274__5 (registerOutputs_274__5), .inputs_274__4 (
            registerOutputs_274__4), .inputs_274__3 (registerOutputs_274__3), .inputs_274__2 (
            registerOutputs_274__2), .inputs_274__1 (registerOutputs_274__1), .inputs_274__0 (
            registerOutputs_274__0), .inputs_275__15 (registerOutputs_275__15), 
            .inputs_275__14 (registerOutputs_275__14), .inputs_275__13 (
            registerOutputs_275__13), .inputs_275__12 (registerOutputs_275__12)
            , .inputs_275__11 (registerOutputs_275__11), .inputs_275__10 (
            registerOutputs_275__10), .inputs_275__9 (registerOutputs_275__9), .inputs_275__8 (
            registerOutputs_275__8), .inputs_275__7 (registerOutputs_275__7), .inputs_275__6 (
            registerOutputs_275__6), .inputs_275__5 (registerOutputs_275__5), .inputs_275__4 (
            registerOutputs_275__4), .inputs_275__3 (registerOutputs_275__3), .inputs_275__2 (
            registerOutputs_275__2), .inputs_275__1 (registerOutputs_275__1), .inputs_275__0 (
            registerOutputs_275__0), .inputs_276__15 (registerOutputs_276__15), 
            .inputs_276__14 (registerOutputs_276__14), .inputs_276__13 (
            registerOutputs_276__13), .inputs_276__12 (registerOutputs_276__12)
            , .inputs_276__11 (registerOutputs_276__11), .inputs_276__10 (
            registerOutputs_276__10), .inputs_276__9 (registerOutputs_276__9), .inputs_276__8 (
            registerOutputs_276__8), .inputs_276__7 (registerOutputs_276__7), .inputs_276__6 (
            registerOutputs_276__6), .inputs_276__5 (registerOutputs_276__5), .inputs_276__4 (
            registerOutputs_276__4), .inputs_276__3 (registerOutputs_276__3), .inputs_276__2 (
            registerOutputs_276__2), .inputs_276__1 (registerOutputs_276__1), .inputs_276__0 (
            registerOutputs_276__0), .inputs_277__15 (registerOutputs_277__15), 
            .inputs_277__14 (registerOutputs_277__14), .inputs_277__13 (
            registerOutputs_277__13), .inputs_277__12 (registerOutputs_277__12)
            , .inputs_277__11 (registerOutputs_277__11), .inputs_277__10 (
            registerOutputs_277__10), .inputs_277__9 (registerOutputs_277__9), .inputs_277__8 (
            registerOutputs_277__8), .inputs_277__7 (registerOutputs_277__7), .inputs_277__6 (
            registerOutputs_277__6), .inputs_277__5 (registerOutputs_277__5), .inputs_277__4 (
            registerOutputs_277__4), .inputs_277__3 (registerOutputs_277__3), .inputs_277__2 (
            registerOutputs_277__2), .inputs_277__1 (registerOutputs_277__1), .inputs_277__0 (
            registerOutputs_277__0), .inputs_278__15 (registerOutputs_278__15), 
            .inputs_278__14 (registerOutputs_278__14), .inputs_278__13 (
            registerOutputs_278__13), .inputs_278__12 (registerOutputs_278__12)
            , .inputs_278__11 (registerOutputs_278__11), .inputs_278__10 (
            registerOutputs_278__10), .inputs_278__9 (registerOutputs_278__9), .inputs_278__8 (
            registerOutputs_278__8), .inputs_278__7 (registerOutputs_278__7), .inputs_278__6 (
            registerOutputs_278__6), .inputs_278__5 (registerOutputs_278__5), .inputs_278__4 (
            registerOutputs_278__4), .inputs_278__3 (registerOutputs_278__3), .inputs_278__2 (
            registerOutputs_278__2), .inputs_278__1 (registerOutputs_278__1), .inputs_278__0 (
            registerOutputs_278__0), .inputs_279__15 (registerOutputs_279__15), 
            .inputs_279__14 (registerOutputs_279__14), .inputs_279__13 (
            registerOutputs_279__13), .inputs_279__12 (registerOutputs_279__12)
            , .inputs_279__11 (registerOutputs_279__11), .inputs_279__10 (
            registerOutputs_279__10), .inputs_279__9 (registerOutputs_279__9), .inputs_279__8 (
            registerOutputs_279__8), .inputs_279__7 (registerOutputs_279__7), .inputs_279__6 (
            registerOutputs_279__6), .inputs_279__5 (registerOutputs_279__5), .inputs_279__4 (
            registerOutputs_279__4), .inputs_279__3 (registerOutputs_279__3), .inputs_279__2 (
            registerOutputs_279__2), .inputs_279__1 (registerOutputs_279__1), .inputs_279__0 (
            registerOutputs_279__0), .inputs_280__15 (registerOutputs_280__15), 
            .inputs_280__14 (registerOutputs_280__14), .inputs_280__13 (
            registerOutputs_280__13), .inputs_280__12 (registerOutputs_280__12)
            , .inputs_280__11 (registerOutputs_280__11), .inputs_280__10 (
            registerOutputs_280__10), .inputs_280__9 (registerOutputs_280__9), .inputs_280__8 (
            registerOutputs_280__8), .inputs_280__7 (registerOutputs_280__7), .inputs_280__6 (
            registerOutputs_280__6), .inputs_280__5 (registerOutputs_280__5), .inputs_280__4 (
            registerOutputs_280__4), .inputs_280__3 (registerOutputs_280__3), .inputs_280__2 (
            registerOutputs_280__2), .inputs_280__1 (registerOutputs_280__1), .inputs_280__0 (
            registerOutputs_280__0), .inputs_281__15 (registerOutputs_281__15), 
            .inputs_281__14 (registerOutputs_281__14), .inputs_281__13 (
            registerOutputs_281__13), .inputs_281__12 (registerOutputs_281__12)
            , .inputs_281__11 (registerOutputs_281__11), .inputs_281__10 (
            registerOutputs_281__10), .inputs_281__9 (registerOutputs_281__9), .inputs_281__8 (
            registerOutputs_281__8), .inputs_281__7 (registerOutputs_281__7), .inputs_281__6 (
            registerOutputs_281__6), .inputs_281__5 (registerOutputs_281__5), .inputs_281__4 (
            registerOutputs_281__4), .inputs_281__3 (registerOutputs_281__3), .inputs_281__2 (
            registerOutputs_281__2), .inputs_281__1 (registerOutputs_281__1), .inputs_281__0 (
            registerOutputs_281__0), .inputs_282__15 (registerOutputs_282__15), 
            .inputs_282__14 (registerOutputs_282__14), .inputs_282__13 (
            registerOutputs_282__13), .inputs_282__12 (registerOutputs_282__12)
            , .inputs_282__11 (registerOutputs_282__11), .inputs_282__10 (
            registerOutputs_282__10), .inputs_282__9 (registerOutputs_282__9), .inputs_282__8 (
            registerOutputs_282__8), .inputs_282__7 (registerOutputs_282__7), .inputs_282__6 (
            registerOutputs_282__6), .inputs_282__5 (registerOutputs_282__5), .inputs_282__4 (
            registerOutputs_282__4), .inputs_282__3 (registerOutputs_282__3), .inputs_282__2 (
            registerOutputs_282__2), .inputs_282__1 (registerOutputs_282__1), .inputs_282__0 (
            registerOutputs_282__0), .inputs_283__15 (registerOutputs_283__15), 
            .inputs_283__14 (registerOutputs_283__14), .inputs_283__13 (
            registerOutputs_283__13), .inputs_283__12 (registerOutputs_283__12)
            , .inputs_283__11 (registerOutputs_283__11), .inputs_283__10 (
            registerOutputs_283__10), .inputs_283__9 (registerOutputs_283__9), .inputs_283__8 (
            registerOutputs_283__8), .inputs_283__7 (registerOutputs_283__7), .inputs_283__6 (
            registerOutputs_283__6), .inputs_283__5 (registerOutputs_283__5), .inputs_283__4 (
            registerOutputs_283__4), .inputs_283__3 (registerOutputs_283__3), .inputs_283__2 (
            registerOutputs_283__2), .inputs_283__1 (registerOutputs_283__1), .inputs_283__0 (
            registerOutputs_283__0), .inputs_284__15 (registerOutputs_284__15), 
            .inputs_284__14 (registerOutputs_284__14), .inputs_284__13 (
            registerOutputs_284__13), .inputs_284__12 (registerOutputs_284__12)
            , .inputs_284__11 (registerOutputs_284__11), .inputs_284__10 (
            registerOutputs_284__10), .inputs_284__9 (registerOutputs_284__9), .inputs_284__8 (
            registerOutputs_284__8), .inputs_284__7 (registerOutputs_284__7), .inputs_284__6 (
            registerOutputs_284__6), .inputs_284__5 (registerOutputs_284__5), .inputs_284__4 (
            registerOutputs_284__4), .inputs_284__3 (registerOutputs_284__3), .inputs_284__2 (
            registerOutputs_284__2), .inputs_284__1 (registerOutputs_284__1), .inputs_284__0 (
            registerOutputs_284__0), .inputs_285__15 (registerOutputs_285__15), 
            .inputs_285__14 (registerOutputs_285__14), .inputs_285__13 (
            registerOutputs_285__13), .inputs_285__12 (registerOutputs_285__12)
            , .inputs_285__11 (registerOutputs_285__11), .inputs_285__10 (
            registerOutputs_285__10), .inputs_285__9 (registerOutputs_285__9), .inputs_285__8 (
            registerOutputs_285__8), .inputs_285__7 (registerOutputs_285__7), .inputs_285__6 (
            registerOutputs_285__6), .inputs_285__5 (registerOutputs_285__5), .inputs_285__4 (
            registerOutputs_285__4), .inputs_285__3 (registerOutputs_285__3), .inputs_285__2 (
            registerOutputs_285__2), .inputs_285__1 (registerOutputs_285__1), .inputs_285__0 (
            registerOutputs_285__0), .inputs_286__15 (registerOutputs_286__15), 
            .inputs_286__14 (registerOutputs_286__14), .inputs_286__13 (
            registerOutputs_286__13), .inputs_286__12 (registerOutputs_286__12)
            , .inputs_286__11 (registerOutputs_286__11), .inputs_286__10 (
            registerOutputs_286__10), .inputs_286__9 (registerOutputs_286__9), .inputs_286__8 (
            registerOutputs_286__8), .inputs_286__7 (registerOutputs_286__7), .inputs_286__6 (
            registerOutputs_286__6), .inputs_286__5 (registerOutputs_286__5), .inputs_286__4 (
            registerOutputs_286__4), .inputs_286__3 (registerOutputs_286__3), .inputs_286__2 (
            registerOutputs_286__2), .inputs_286__1 (registerOutputs_286__1), .inputs_286__0 (
            registerOutputs_286__0), .inputs_287__15 (registerOutputs_287__15), 
            .inputs_287__14 (registerOutputs_287__14), .inputs_287__13 (
            registerOutputs_287__13), .inputs_287__12 (registerOutputs_287__12)
            , .inputs_287__11 (registerOutputs_287__11), .inputs_287__10 (
            registerOutputs_287__10), .inputs_287__9 (registerOutputs_287__9), .inputs_287__8 (
            registerOutputs_287__8), .inputs_287__7 (registerOutputs_287__7), .inputs_287__6 (
            registerOutputs_287__6), .inputs_287__5 (registerOutputs_287__5), .inputs_287__4 (
            registerOutputs_287__4), .inputs_287__3 (registerOutputs_287__3), .inputs_287__2 (
            registerOutputs_287__2), .inputs_287__1 (registerOutputs_287__1), .inputs_287__0 (
            registerOutputs_287__0), .inputs_288__15 (registerOutputs_288__15), 
            .inputs_288__14 (registerOutputs_288__14), .inputs_288__13 (
            registerOutputs_288__13), .inputs_288__12 (registerOutputs_288__12)
            , .inputs_288__11 (registerOutputs_288__11), .inputs_288__10 (
            registerOutputs_288__10), .inputs_288__9 (registerOutputs_288__9), .inputs_288__8 (
            registerOutputs_288__8), .inputs_288__7 (registerOutputs_288__7), .inputs_288__6 (
            registerOutputs_288__6), .inputs_288__5 (registerOutputs_288__5), .inputs_288__4 (
            registerOutputs_288__4), .inputs_288__3 (registerOutputs_288__3), .inputs_288__2 (
            registerOutputs_288__2), .inputs_288__1 (registerOutputs_288__1), .inputs_288__0 (
            registerOutputs_288__0), .inputs_289__15 (registerOutputs_289__15), 
            .inputs_289__14 (registerOutputs_289__14), .inputs_289__13 (
            registerOutputs_289__13), .inputs_289__12 (registerOutputs_289__12)
            , .inputs_289__11 (registerOutputs_289__11), .inputs_289__10 (
            registerOutputs_289__10), .inputs_289__9 (registerOutputs_289__9), .inputs_289__8 (
            registerOutputs_289__8), .inputs_289__7 (registerOutputs_289__7), .inputs_289__6 (
            registerOutputs_289__6), .inputs_289__5 (registerOutputs_289__5), .inputs_289__4 (
            registerOutputs_289__4), .inputs_289__3 (registerOutputs_289__3), .inputs_289__2 (
            registerOutputs_289__2), .inputs_289__1 (registerOutputs_289__1), .inputs_289__0 (
            registerOutputs_289__0), .inputs_290__15 (registerOutputs_290__15), 
            .inputs_290__14 (registerOutputs_290__14), .inputs_290__13 (
            registerOutputs_290__13), .inputs_290__12 (registerOutputs_290__12)
            , .inputs_290__11 (registerOutputs_290__11), .inputs_290__10 (
            registerOutputs_290__10), .inputs_290__9 (registerOutputs_290__9), .inputs_290__8 (
            registerOutputs_290__8), .inputs_290__7 (registerOutputs_290__7), .inputs_290__6 (
            registerOutputs_290__6), .inputs_290__5 (registerOutputs_290__5), .inputs_290__4 (
            registerOutputs_290__4), .inputs_290__3 (registerOutputs_290__3), .inputs_290__2 (
            registerOutputs_290__2), .inputs_290__1 (registerOutputs_290__1), .inputs_290__0 (
            registerOutputs_290__0), .inputs_291__15 (registerOutputs_291__15), 
            .inputs_291__14 (registerOutputs_291__14), .inputs_291__13 (
            registerOutputs_291__13), .inputs_291__12 (registerOutputs_291__12)
            , .inputs_291__11 (registerOutputs_291__11), .inputs_291__10 (
            registerOutputs_291__10), .inputs_291__9 (registerOutputs_291__9), .inputs_291__8 (
            registerOutputs_291__8), .inputs_291__7 (registerOutputs_291__7), .inputs_291__6 (
            registerOutputs_291__6), .inputs_291__5 (registerOutputs_291__5), .inputs_291__4 (
            registerOutputs_291__4), .inputs_291__3 (registerOutputs_291__3), .inputs_291__2 (
            registerOutputs_291__2), .inputs_291__1 (registerOutputs_291__1), .inputs_291__0 (
            registerOutputs_291__0), .inputs_292__15 (registerOutputs_292__15), 
            .inputs_292__14 (registerOutputs_292__14), .inputs_292__13 (
            registerOutputs_292__13), .inputs_292__12 (registerOutputs_292__12)
            , .inputs_292__11 (registerOutputs_292__11), .inputs_292__10 (
            registerOutputs_292__10), .inputs_292__9 (registerOutputs_292__9), .inputs_292__8 (
            registerOutputs_292__8), .inputs_292__7 (registerOutputs_292__7), .inputs_292__6 (
            registerOutputs_292__6), .inputs_292__5 (registerOutputs_292__5), .inputs_292__4 (
            registerOutputs_292__4), .inputs_292__3 (registerOutputs_292__3), .inputs_292__2 (
            registerOutputs_292__2), .inputs_292__1 (registerOutputs_292__1), .inputs_292__0 (
            registerOutputs_292__0), .inputs_293__15 (registerOutputs_293__15), 
            .inputs_293__14 (registerOutputs_293__14), .inputs_293__13 (
            registerOutputs_293__13), .inputs_293__12 (registerOutputs_293__12)
            , .inputs_293__11 (registerOutputs_293__11), .inputs_293__10 (
            registerOutputs_293__10), .inputs_293__9 (registerOutputs_293__9), .inputs_293__8 (
            registerOutputs_293__8), .inputs_293__7 (registerOutputs_293__7), .inputs_293__6 (
            registerOutputs_293__6), .inputs_293__5 (registerOutputs_293__5), .inputs_293__4 (
            registerOutputs_293__4), .inputs_293__3 (registerOutputs_293__3), .inputs_293__2 (
            registerOutputs_293__2), .inputs_293__1 (registerOutputs_293__1), .inputs_293__0 (
            registerOutputs_293__0), .inputs_294__15 (registerOutputs_294__15), 
            .inputs_294__14 (registerOutputs_294__14), .inputs_294__13 (
            registerOutputs_294__13), .inputs_294__12 (registerOutputs_294__12)
            , .inputs_294__11 (registerOutputs_294__11), .inputs_294__10 (
            registerOutputs_294__10), .inputs_294__9 (registerOutputs_294__9), .inputs_294__8 (
            registerOutputs_294__8), .inputs_294__7 (registerOutputs_294__7), .inputs_294__6 (
            registerOutputs_294__6), .inputs_294__5 (registerOutputs_294__5), .inputs_294__4 (
            registerOutputs_294__4), .inputs_294__3 (registerOutputs_294__3), .inputs_294__2 (
            registerOutputs_294__2), .inputs_294__1 (registerOutputs_294__1), .inputs_294__0 (
            registerOutputs_294__0), .inputs_295__15 (registerOutputs_295__15), 
            .inputs_295__14 (registerOutputs_295__14), .inputs_295__13 (
            registerOutputs_295__13), .inputs_295__12 (registerOutputs_295__12)
            , .inputs_295__11 (registerOutputs_295__11), .inputs_295__10 (
            registerOutputs_295__10), .inputs_295__9 (registerOutputs_295__9), .inputs_295__8 (
            registerOutputs_295__8), .inputs_295__7 (registerOutputs_295__7), .inputs_295__6 (
            registerOutputs_295__6), .inputs_295__5 (registerOutputs_295__5), .inputs_295__4 (
            registerOutputs_295__4), .inputs_295__3 (registerOutputs_295__3), .inputs_295__2 (
            registerOutputs_295__2), .inputs_295__1 (registerOutputs_295__1), .inputs_295__0 (
            registerOutputs_295__0), .inputs_296__15 (registerOutputs_296__15), 
            .inputs_296__14 (registerOutputs_296__14), .inputs_296__13 (
            registerOutputs_296__13), .inputs_296__12 (registerOutputs_296__12)
            , .inputs_296__11 (registerOutputs_296__11), .inputs_296__10 (
            registerOutputs_296__10), .inputs_296__9 (registerOutputs_296__9), .inputs_296__8 (
            registerOutputs_296__8), .inputs_296__7 (registerOutputs_296__7), .inputs_296__6 (
            registerOutputs_296__6), .inputs_296__5 (registerOutputs_296__5), .inputs_296__4 (
            registerOutputs_296__4), .inputs_296__3 (registerOutputs_296__3), .inputs_296__2 (
            registerOutputs_296__2), .inputs_296__1 (registerOutputs_296__1), .inputs_296__0 (
            registerOutputs_296__0), .inputs_297__15 (registerOutputs_297__15), 
            .inputs_297__14 (registerOutputs_297__14), .inputs_297__13 (
            registerOutputs_297__13), .inputs_297__12 (registerOutputs_297__12)
            , .inputs_297__11 (registerOutputs_297__11), .inputs_297__10 (
            registerOutputs_297__10), .inputs_297__9 (registerOutputs_297__9), .inputs_297__8 (
            registerOutputs_297__8), .inputs_297__7 (registerOutputs_297__7), .inputs_297__6 (
            registerOutputs_297__6), .inputs_297__5 (registerOutputs_297__5), .inputs_297__4 (
            registerOutputs_297__4), .inputs_297__3 (registerOutputs_297__3), .inputs_297__2 (
            registerOutputs_297__2), .inputs_297__1 (registerOutputs_297__1), .inputs_297__0 (
            registerOutputs_297__0), .inputs_298__15 (registerOutputs_298__15), 
            .inputs_298__14 (registerOutputs_298__14), .inputs_298__13 (
            registerOutputs_298__13), .inputs_298__12 (registerOutputs_298__12)
            , .inputs_298__11 (registerOutputs_298__11), .inputs_298__10 (
            registerOutputs_298__10), .inputs_298__9 (registerOutputs_298__9), .inputs_298__8 (
            registerOutputs_298__8), .inputs_298__7 (registerOutputs_298__7), .inputs_298__6 (
            registerOutputs_298__6), .inputs_298__5 (registerOutputs_298__5), .inputs_298__4 (
            registerOutputs_298__4), .inputs_298__3 (registerOutputs_298__3), .inputs_298__2 (
            registerOutputs_298__2), .inputs_298__1 (registerOutputs_298__1), .inputs_298__0 (
            registerOutputs_298__0), .inputs_299__15 (registerOutputs_299__15), 
            .inputs_299__14 (registerOutputs_299__14), .inputs_299__13 (
            registerOutputs_299__13), .inputs_299__12 (registerOutputs_299__12)
            , .inputs_299__11 (registerOutputs_299__11), .inputs_299__10 (
            registerOutputs_299__10), .inputs_299__9 (registerOutputs_299__9), .inputs_299__8 (
            registerOutputs_299__8), .inputs_299__7 (registerOutputs_299__7), .inputs_299__6 (
            registerOutputs_299__6), .inputs_299__5 (registerOutputs_299__5), .inputs_299__4 (
            registerOutputs_299__4), .inputs_299__3 (registerOutputs_299__3), .inputs_299__2 (
            registerOutputs_299__2), .inputs_299__1 (registerOutputs_299__1), .inputs_299__0 (
            registerOutputs_299__0), .inputs_300__15 (registerOutputs_300__15), 
            .inputs_300__14 (registerOutputs_300__14), .inputs_300__13 (
            registerOutputs_300__13), .inputs_300__12 (registerOutputs_300__12)
            , .inputs_300__11 (registerOutputs_300__11), .inputs_300__10 (
            registerOutputs_300__10), .inputs_300__9 (registerOutputs_300__9), .inputs_300__8 (
            registerOutputs_300__8), .inputs_300__7 (registerOutputs_300__7), .inputs_300__6 (
            registerOutputs_300__6), .inputs_300__5 (registerOutputs_300__5), .inputs_300__4 (
            registerOutputs_300__4), .inputs_300__3 (registerOutputs_300__3), .inputs_300__2 (
            registerOutputs_300__2), .inputs_300__1 (registerOutputs_300__1), .inputs_300__0 (
            registerOutputs_300__0), .inputs_301__15 (registerOutputs_301__15), 
            .inputs_301__14 (registerOutputs_301__14), .inputs_301__13 (
            registerOutputs_301__13), .inputs_301__12 (registerOutputs_301__12)
            , .inputs_301__11 (registerOutputs_301__11), .inputs_301__10 (
            registerOutputs_301__10), .inputs_301__9 (registerOutputs_301__9), .inputs_301__8 (
            registerOutputs_301__8), .inputs_301__7 (registerOutputs_301__7), .inputs_301__6 (
            registerOutputs_301__6), .inputs_301__5 (registerOutputs_301__5), .inputs_301__4 (
            registerOutputs_301__4), .inputs_301__3 (registerOutputs_301__3), .inputs_301__2 (
            registerOutputs_301__2), .inputs_301__1 (registerOutputs_301__1), .inputs_301__0 (
            registerOutputs_301__0), .inputs_302__15 (registerOutputs_302__15), 
            .inputs_302__14 (registerOutputs_302__14), .inputs_302__13 (
            registerOutputs_302__13), .inputs_302__12 (registerOutputs_302__12)
            , .inputs_302__11 (registerOutputs_302__11), .inputs_302__10 (
            registerOutputs_302__10), .inputs_302__9 (registerOutputs_302__9), .inputs_302__8 (
            registerOutputs_302__8), .inputs_302__7 (registerOutputs_302__7), .inputs_302__6 (
            registerOutputs_302__6), .inputs_302__5 (registerOutputs_302__5), .inputs_302__4 (
            registerOutputs_302__4), .inputs_302__3 (registerOutputs_302__3), .inputs_302__2 (
            registerOutputs_302__2), .inputs_302__1 (registerOutputs_302__1), .inputs_302__0 (
            registerOutputs_302__0), .inputs_303__15 (registerOutputs_303__15), 
            .inputs_303__14 (registerOutputs_303__14), .inputs_303__13 (
            registerOutputs_303__13), .inputs_303__12 (registerOutputs_303__12)
            , .inputs_303__11 (registerOutputs_303__11), .inputs_303__10 (
            registerOutputs_303__10), .inputs_303__9 (registerOutputs_303__9), .inputs_303__8 (
            registerOutputs_303__8), .inputs_303__7 (registerOutputs_303__7), .inputs_303__6 (
            registerOutputs_303__6), .inputs_303__5 (registerOutputs_303__5), .inputs_303__4 (
            registerOutputs_303__4), .inputs_303__3 (registerOutputs_303__3), .inputs_303__2 (
            registerOutputs_303__2), .inputs_303__1 (registerOutputs_303__1), .inputs_303__0 (
            registerOutputs_303__0), .inputs_304__15 (registerOutputs_304__15), 
            .inputs_304__14 (registerOutputs_304__14), .inputs_304__13 (
            registerOutputs_304__13), .inputs_304__12 (registerOutputs_304__12)
            , .inputs_304__11 (registerOutputs_304__11), .inputs_304__10 (
            registerOutputs_304__10), .inputs_304__9 (registerOutputs_304__9), .inputs_304__8 (
            registerOutputs_304__8), .inputs_304__7 (registerOutputs_304__7), .inputs_304__6 (
            registerOutputs_304__6), .inputs_304__5 (registerOutputs_304__5), .inputs_304__4 (
            registerOutputs_304__4), .inputs_304__3 (registerOutputs_304__3), .inputs_304__2 (
            registerOutputs_304__2), .inputs_304__1 (registerOutputs_304__1), .inputs_304__0 (
            registerOutputs_304__0), .inputs_305__15 (registerOutputs_305__15), 
            .inputs_305__14 (registerOutputs_305__14), .inputs_305__13 (
            registerOutputs_305__13), .inputs_305__12 (registerOutputs_305__12)
            , .inputs_305__11 (registerOutputs_305__11), .inputs_305__10 (
            registerOutputs_305__10), .inputs_305__9 (registerOutputs_305__9), .inputs_305__8 (
            registerOutputs_305__8), .inputs_305__7 (registerOutputs_305__7), .inputs_305__6 (
            registerOutputs_305__6), .inputs_305__5 (registerOutputs_305__5), .inputs_305__4 (
            registerOutputs_305__4), .inputs_305__3 (registerOutputs_305__3), .inputs_305__2 (
            registerOutputs_305__2), .inputs_305__1 (registerOutputs_305__1), .inputs_305__0 (
            registerOutputs_305__0), .inputs_306__15 (registerOutputs_306__15), 
            .inputs_306__14 (registerOutputs_306__14), .inputs_306__13 (
            registerOutputs_306__13), .inputs_306__12 (registerOutputs_306__12)
            , .inputs_306__11 (registerOutputs_306__11), .inputs_306__10 (
            registerOutputs_306__10), .inputs_306__9 (registerOutputs_306__9), .inputs_306__8 (
            registerOutputs_306__8), .inputs_306__7 (registerOutputs_306__7), .inputs_306__6 (
            registerOutputs_306__6), .inputs_306__5 (registerOutputs_306__5), .inputs_306__4 (
            registerOutputs_306__4), .inputs_306__3 (registerOutputs_306__3), .inputs_306__2 (
            registerOutputs_306__2), .inputs_306__1 (registerOutputs_306__1), .inputs_306__0 (
            registerOutputs_306__0), .inputs_307__15 (registerOutputs_307__15), 
            .inputs_307__14 (registerOutputs_307__14), .inputs_307__13 (
            registerOutputs_307__13), .inputs_307__12 (registerOutputs_307__12)
            , .inputs_307__11 (registerOutputs_307__11), .inputs_307__10 (
            registerOutputs_307__10), .inputs_307__9 (registerOutputs_307__9), .inputs_307__8 (
            registerOutputs_307__8), .inputs_307__7 (registerOutputs_307__7), .inputs_307__6 (
            registerOutputs_307__6), .inputs_307__5 (registerOutputs_307__5), .inputs_307__4 (
            registerOutputs_307__4), .inputs_307__3 (registerOutputs_307__3), .inputs_307__2 (
            registerOutputs_307__2), .inputs_307__1 (registerOutputs_307__1), .inputs_307__0 (
            registerOutputs_307__0), .inputs_308__15 (registerOutputs_308__15), 
            .inputs_308__14 (registerOutputs_308__14), .inputs_308__13 (
            registerOutputs_308__13), .inputs_308__12 (registerOutputs_308__12)
            , .inputs_308__11 (registerOutputs_308__11), .inputs_308__10 (
            registerOutputs_308__10), .inputs_308__9 (registerOutputs_308__9), .inputs_308__8 (
            registerOutputs_308__8), .inputs_308__7 (registerOutputs_308__7), .inputs_308__6 (
            registerOutputs_308__6), .inputs_308__5 (registerOutputs_308__5), .inputs_308__4 (
            registerOutputs_308__4), .inputs_308__3 (registerOutputs_308__3), .inputs_308__2 (
            registerOutputs_308__2), .inputs_308__1 (registerOutputs_308__1), .inputs_308__0 (
            registerOutputs_308__0), .inputs_309__15 (registerOutputs_309__15), 
            .inputs_309__14 (registerOutputs_309__14), .inputs_309__13 (
            registerOutputs_309__13), .inputs_309__12 (registerOutputs_309__12)
            , .inputs_309__11 (registerOutputs_309__11), .inputs_309__10 (
            registerOutputs_309__10), .inputs_309__9 (registerOutputs_309__9), .inputs_309__8 (
            registerOutputs_309__8), .inputs_309__7 (registerOutputs_309__7), .inputs_309__6 (
            registerOutputs_309__6), .inputs_309__5 (registerOutputs_309__5), .inputs_309__4 (
            registerOutputs_309__4), .inputs_309__3 (registerOutputs_309__3), .inputs_309__2 (
            registerOutputs_309__2), .inputs_309__1 (registerOutputs_309__1), .inputs_309__0 (
            registerOutputs_309__0), .inputs_310__15 (registerOutputs_310__15), 
            .inputs_310__14 (registerOutputs_310__14), .inputs_310__13 (
            registerOutputs_310__13), .inputs_310__12 (registerOutputs_310__12)
            , .inputs_310__11 (registerOutputs_310__11), .inputs_310__10 (
            registerOutputs_310__10), .inputs_310__9 (registerOutputs_310__9), .inputs_310__8 (
            registerOutputs_310__8), .inputs_310__7 (registerOutputs_310__7), .inputs_310__6 (
            registerOutputs_310__6), .inputs_310__5 (registerOutputs_310__5), .inputs_310__4 (
            registerOutputs_310__4), .inputs_310__3 (registerOutputs_310__3), .inputs_310__2 (
            registerOutputs_310__2), .inputs_310__1 (registerOutputs_310__1), .inputs_310__0 (
            registerOutputs_310__0), .inputs_311__15 (registerOutputs_311__15), 
            .inputs_311__14 (registerOutputs_311__14), .inputs_311__13 (
            registerOutputs_311__13), .inputs_311__12 (registerOutputs_311__12)
            , .inputs_311__11 (registerOutputs_311__11), .inputs_311__10 (
            registerOutputs_311__10), .inputs_311__9 (registerOutputs_311__9), .inputs_311__8 (
            registerOutputs_311__8), .inputs_311__7 (registerOutputs_311__7), .inputs_311__6 (
            registerOutputs_311__6), .inputs_311__5 (registerOutputs_311__5), .inputs_311__4 (
            registerOutputs_311__4), .inputs_311__3 (registerOutputs_311__3), .inputs_311__2 (
            registerOutputs_311__2), .inputs_311__1 (registerOutputs_311__1), .inputs_311__0 (
            registerOutputs_311__0), .inputs_312__15 (registerOutputs_312__15), 
            .inputs_312__14 (registerOutputs_312__14), .inputs_312__13 (
            registerOutputs_312__13), .inputs_312__12 (registerOutputs_312__12)
            , .inputs_312__11 (registerOutputs_312__11), .inputs_312__10 (
            registerOutputs_312__10), .inputs_312__9 (registerOutputs_312__9), .inputs_312__8 (
            registerOutputs_312__8), .inputs_312__7 (registerOutputs_312__7), .inputs_312__6 (
            registerOutputs_312__6), .inputs_312__5 (registerOutputs_312__5), .inputs_312__4 (
            registerOutputs_312__4), .inputs_312__3 (registerOutputs_312__3), .inputs_312__2 (
            registerOutputs_312__2), .inputs_312__1 (registerOutputs_312__1), .inputs_312__0 (
            registerOutputs_312__0), .inputs_313__15 (registerOutputs_313__15), 
            .inputs_313__14 (registerOutputs_313__14), .inputs_313__13 (
            registerOutputs_313__13), .inputs_313__12 (registerOutputs_313__12)
            , .inputs_313__11 (registerOutputs_313__11), .inputs_313__10 (
            registerOutputs_313__10), .inputs_313__9 (registerOutputs_313__9), .inputs_313__8 (
            registerOutputs_313__8), .inputs_313__7 (registerOutputs_313__7), .inputs_313__6 (
            registerOutputs_313__6), .inputs_313__5 (registerOutputs_313__5), .inputs_313__4 (
            registerOutputs_313__4), .inputs_313__3 (registerOutputs_313__3), .inputs_313__2 (
            registerOutputs_313__2), .inputs_313__1 (registerOutputs_313__1), .inputs_313__0 (
            registerOutputs_313__0), .inputs_314__15 (registerOutputs_314__15), 
            .inputs_314__14 (registerOutputs_314__14), .inputs_314__13 (
            registerOutputs_314__13), .inputs_314__12 (registerOutputs_314__12)
            , .inputs_314__11 (registerOutputs_314__11), .inputs_314__10 (
            registerOutputs_314__10), .inputs_314__9 (registerOutputs_314__9), .inputs_314__8 (
            registerOutputs_314__8), .inputs_314__7 (registerOutputs_314__7), .inputs_314__6 (
            registerOutputs_314__6), .inputs_314__5 (registerOutputs_314__5), .inputs_314__4 (
            registerOutputs_314__4), .inputs_314__3 (registerOutputs_314__3), .inputs_314__2 (
            registerOutputs_314__2), .inputs_314__1 (registerOutputs_314__1), .inputs_314__0 (
            registerOutputs_314__0), .inputs_315__15 (registerOutputs_315__15), 
            .inputs_315__14 (registerOutputs_315__14), .inputs_315__13 (
            registerOutputs_315__13), .inputs_315__12 (registerOutputs_315__12)
            , .inputs_315__11 (registerOutputs_315__11), .inputs_315__10 (
            registerOutputs_315__10), .inputs_315__9 (registerOutputs_315__9), .inputs_315__8 (
            registerOutputs_315__8), .inputs_315__7 (registerOutputs_315__7), .inputs_315__6 (
            registerOutputs_315__6), .inputs_315__5 (registerOutputs_315__5), .inputs_315__4 (
            registerOutputs_315__4), .inputs_315__3 (registerOutputs_315__3), .inputs_315__2 (
            registerOutputs_315__2), .inputs_315__1 (registerOutputs_315__1), .inputs_315__0 (
            registerOutputs_315__0), .inputs_316__15 (registerOutputs_316__15), 
            .inputs_316__14 (registerOutputs_316__14), .inputs_316__13 (
            registerOutputs_316__13), .inputs_316__12 (registerOutputs_316__12)
            , .inputs_316__11 (registerOutputs_316__11), .inputs_316__10 (
            registerOutputs_316__10), .inputs_316__9 (registerOutputs_316__9), .inputs_316__8 (
            registerOutputs_316__8), .inputs_316__7 (registerOutputs_316__7), .inputs_316__6 (
            registerOutputs_316__6), .inputs_316__5 (registerOutputs_316__5), .inputs_316__4 (
            registerOutputs_316__4), .inputs_316__3 (registerOutputs_316__3), .inputs_316__2 (
            registerOutputs_316__2), .inputs_316__1 (registerOutputs_316__1), .inputs_316__0 (
            registerOutputs_316__0), .inputs_317__15 (registerOutputs_317__15), 
            .inputs_317__14 (registerOutputs_317__14), .inputs_317__13 (
            registerOutputs_317__13), .inputs_317__12 (registerOutputs_317__12)
            , .inputs_317__11 (registerOutputs_317__11), .inputs_317__10 (
            registerOutputs_317__10), .inputs_317__9 (registerOutputs_317__9), .inputs_317__8 (
            registerOutputs_317__8), .inputs_317__7 (registerOutputs_317__7), .inputs_317__6 (
            registerOutputs_317__6), .inputs_317__5 (registerOutputs_317__5), .inputs_317__4 (
            registerOutputs_317__4), .inputs_317__3 (registerOutputs_317__3), .inputs_317__2 (
            registerOutputs_317__2), .inputs_317__1 (registerOutputs_317__1), .inputs_317__0 (
            registerOutputs_317__0), .inputs_318__15 (registerOutputs_318__15), 
            .inputs_318__14 (registerOutputs_318__14), .inputs_318__13 (
            registerOutputs_318__13), .inputs_318__12 (registerOutputs_318__12)
            , .inputs_318__11 (registerOutputs_318__11), .inputs_318__10 (
            registerOutputs_318__10), .inputs_318__9 (registerOutputs_318__9), .inputs_318__8 (
            registerOutputs_318__8), .inputs_318__7 (registerOutputs_318__7), .inputs_318__6 (
            registerOutputs_318__6), .inputs_318__5 (registerOutputs_318__5), .inputs_318__4 (
            registerOutputs_318__4), .inputs_318__3 (registerOutputs_318__3), .inputs_318__2 (
            registerOutputs_318__2), .inputs_318__1 (registerOutputs_318__1), .inputs_318__0 (
            registerOutputs_318__0), .inputs_319__15 (registerOutputs_319__15), 
            .inputs_319__14 (registerOutputs_319__14), .inputs_319__13 (
            registerOutputs_319__13), .inputs_319__12 (registerOutputs_319__12)
            , .inputs_319__11 (registerOutputs_319__11), .inputs_319__10 (
            registerOutputs_319__10), .inputs_319__9 (registerOutputs_319__9), .inputs_319__8 (
            registerOutputs_319__8), .inputs_319__7 (registerOutputs_319__7), .inputs_319__6 (
            registerOutputs_319__6), .inputs_319__5 (registerOutputs_319__5), .inputs_319__4 (
            registerOutputs_319__4), .inputs_319__3 (registerOutputs_319__3), .inputs_319__2 (
            registerOutputs_319__2), .inputs_319__1 (registerOutputs_319__1), .inputs_319__0 (
            registerOutputs_319__0), .inputs_320__15 (registerOutputs_320__15), 
            .inputs_320__14 (registerOutputs_320__14), .inputs_320__13 (
            registerOutputs_320__13), .inputs_320__12 (registerOutputs_320__12)
            , .inputs_320__11 (registerOutputs_320__11), .inputs_320__10 (
            registerOutputs_320__10), .inputs_320__9 (registerOutputs_320__9), .inputs_320__8 (
            registerOutputs_320__8), .inputs_320__7 (registerOutputs_320__7), .inputs_320__6 (
            registerOutputs_320__6), .inputs_320__5 (registerOutputs_320__5), .inputs_320__4 (
            registerOutputs_320__4), .inputs_320__3 (registerOutputs_320__3), .inputs_320__2 (
            registerOutputs_320__2), .inputs_320__1 (registerOutputs_320__1), .inputs_320__0 (
            registerOutputs_320__0), .inputs_321__15 (registerOutputs_321__15), 
            .inputs_321__14 (registerOutputs_321__14), .inputs_321__13 (
            registerOutputs_321__13), .inputs_321__12 (registerOutputs_321__12)
            , .inputs_321__11 (registerOutputs_321__11), .inputs_321__10 (
            registerOutputs_321__10), .inputs_321__9 (registerOutputs_321__9), .inputs_321__8 (
            registerOutputs_321__8), .inputs_321__7 (registerOutputs_321__7), .inputs_321__6 (
            registerOutputs_321__6), .inputs_321__5 (registerOutputs_321__5), .inputs_321__4 (
            registerOutputs_321__4), .inputs_321__3 (registerOutputs_321__3), .inputs_321__2 (
            registerOutputs_321__2), .inputs_321__1 (registerOutputs_321__1), .inputs_321__0 (
            registerOutputs_321__0), .inputs_322__15 (registerOutputs_322__15), 
            .inputs_322__14 (registerOutputs_322__14), .inputs_322__13 (
            registerOutputs_322__13), .inputs_322__12 (registerOutputs_322__12)
            , .inputs_322__11 (registerOutputs_322__11), .inputs_322__10 (
            registerOutputs_322__10), .inputs_322__9 (registerOutputs_322__9), .inputs_322__8 (
            registerOutputs_322__8), .inputs_322__7 (registerOutputs_322__7), .inputs_322__6 (
            registerOutputs_322__6), .inputs_322__5 (registerOutputs_322__5), .inputs_322__4 (
            registerOutputs_322__4), .inputs_322__3 (registerOutputs_322__3), .inputs_322__2 (
            registerOutputs_322__2), .inputs_322__1 (registerOutputs_322__1), .inputs_322__0 (
            registerOutputs_322__0), .inputs_323__15 (registerOutputs_323__15), 
            .inputs_323__14 (registerOutputs_323__14), .inputs_323__13 (
            registerOutputs_323__13), .inputs_323__12 (registerOutputs_323__12)
            , .inputs_323__11 (registerOutputs_323__11), .inputs_323__10 (
            registerOutputs_323__10), .inputs_323__9 (registerOutputs_323__9), .inputs_323__8 (
            registerOutputs_323__8), .inputs_323__7 (registerOutputs_323__7), .inputs_323__6 (
            registerOutputs_323__6), .inputs_323__5 (registerOutputs_323__5), .inputs_323__4 (
            registerOutputs_323__4), .inputs_323__3 (registerOutputs_323__3), .inputs_323__2 (
            registerOutputs_323__2), .inputs_323__1 (registerOutputs_323__1), .inputs_323__0 (
            registerOutputs_323__0), .inputs_324__15 (registerOutputs_324__15), 
            .inputs_324__14 (registerOutputs_324__14), .inputs_324__13 (
            registerOutputs_324__13), .inputs_324__12 (registerOutputs_324__12)
            , .inputs_324__11 (registerOutputs_324__11), .inputs_324__10 (
            registerOutputs_324__10), .inputs_324__9 (registerOutputs_324__9), .inputs_324__8 (
            registerOutputs_324__8), .inputs_324__7 (registerOutputs_324__7), .inputs_324__6 (
            registerOutputs_324__6), .inputs_324__5 (registerOutputs_324__5), .inputs_324__4 (
            registerOutputs_324__4), .inputs_324__3 (registerOutputs_324__3), .inputs_324__2 (
            registerOutputs_324__2), .inputs_324__1 (registerOutputs_324__1), .inputs_324__0 (
            registerOutputs_324__0), .inputs_325__15 (registerOutputs_325__15), 
            .inputs_325__14 (registerOutputs_325__14), .inputs_325__13 (
            registerOutputs_325__13), .inputs_325__12 (registerOutputs_325__12)
            , .inputs_325__11 (registerOutputs_325__11), .inputs_325__10 (
            registerOutputs_325__10), .inputs_325__9 (registerOutputs_325__9), .inputs_325__8 (
            registerOutputs_325__8), .inputs_325__7 (registerOutputs_325__7), .inputs_325__6 (
            registerOutputs_325__6), .inputs_325__5 (registerOutputs_325__5), .inputs_325__4 (
            registerOutputs_325__4), .inputs_325__3 (registerOutputs_325__3), .inputs_325__2 (
            registerOutputs_325__2), .inputs_325__1 (registerOutputs_325__1), .inputs_325__0 (
            registerOutputs_325__0), .inputs_326__15 (registerOutputs_326__15), 
            .inputs_326__14 (registerOutputs_326__14), .inputs_326__13 (
            registerOutputs_326__13), .inputs_326__12 (registerOutputs_326__12)
            , .inputs_326__11 (registerOutputs_326__11), .inputs_326__10 (
            registerOutputs_326__10), .inputs_326__9 (registerOutputs_326__9), .inputs_326__8 (
            registerOutputs_326__8), .inputs_326__7 (registerOutputs_326__7), .inputs_326__6 (
            registerOutputs_326__6), .inputs_326__5 (registerOutputs_326__5), .inputs_326__4 (
            registerOutputs_326__4), .inputs_326__3 (registerOutputs_326__3), .inputs_326__2 (
            registerOutputs_326__2), .inputs_326__1 (registerOutputs_326__1), .inputs_326__0 (
            registerOutputs_326__0), .inputs_327__15 (registerOutputs_327__15), 
            .inputs_327__14 (registerOutputs_327__14), .inputs_327__13 (
            registerOutputs_327__13), .inputs_327__12 (registerOutputs_327__12)
            , .inputs_327__11 (registerOutputs_327__11), .inputs_327__10 (
            registerOutputs_327__10), .inputs_327__9 (registerOutputs_327__9), .inputs_327__8 (
            registerOutputs_327__8), .inputs_327__7 (registerOutputs_327__7), .inputs_327__6 (
            registerOutputs_327__6), .inputs_327__5 (registerOutputs_327__5), .inputs_327__4 (
            registerOutputs_327__4), .inputs_327__3 (registerOutputs_327__3), .inputs_327__2 (
            registerOutputs_327__2), .inputs_327__1 (registerOutputs_327__1), .inputs_327__0 (
            registerOutputs_327__0), .inputs_328__15 (registerOutputs_328__15), 
            .inputs_328__14 (registerOutputs_328__14), .inputs_328__13 (
            registerOutputs_328__13), .inputs_328__12 (registerOutputs_328__12)
            , .inputs_328__11 (registerOutputs_328__11), .inputs_328__10 (
            registerOutputs_328__10), .inputs_328__9 (registerOutputs_328__9), .inputs_328__8 (
            registerOutputs_328__8), .inputs_328__7 (registerOutputs_328__7), .inputs_328__6 (
            registerOutputs_328__6), .inputs_328__5 (registerOutputs_328__5), .inputs_328__4 (
            registerOutputs_328__4), .inputs_328__3 (registerOutputs_328__3), .inputs_328__2 (
            registerOutputs_328__2), .inputs_328__1 (registerOutputs_328__1), .inputs_328__0 (
            registerOutputs_328__0), .inputs_329__15 (registerOutputs_329__15), 
            .inputs_329__14 (registerOutputs_329__14), .inputs_329__13 (
            registerOutputs_329__13), .inputs_329__12 (registerOutputs_329__12)
            , .inputs_329__11 (registerOutputs_329__11), .inputs_329__10 (
            registerOutputs_329__10), .inputs_329__9 (registerOutputs_329__9), .inputs_329__8 (
            registerOutputs_329__8), .inputs_329__7 (registerOutputs_329__7), .inputs_329__6 (
            registerOutputs_329__6), .inputs_329__5 (registerOutputs_329__5), .inputs_329__4 (
            registerOutputs_329__4), .inputs_329__3 (registerOutputs_329__3), .inputs_329__2 (
            registerOutputs_329__2), .inputs_329__1 (registerOutputs_329__1), .inputs_329__0 (
            registerOutputs_329__0), .inputs_330__15 (registerOutputs_330__15), 
            .inputs_330__14 (registerOutputs_330__14), .inputs_330__13 (
            registerOutputs_330__13), .inputs_330__12 (registerOutputs_330__12)
            , .inputs_330__11 (registerOutputs_330__11), .inputs_330__10 (
            registerOutputs_330__10), .inputs_330__9 (registerOutputs_330__9), .inputs_330__8 (
            registerOutputs_330__8), .inputs_330__7 (registerOutputs_330__7), .inputs_330__6 (
            registerOutputs_330__6), .inputs_330__5 (registerOutputs_330__5), .inputs_330__4 (
            registerOutputs_330__4), .inputs_330__3 (registerOutputs_330__3), .inputs_330__2 (
            registerOutputs_330__2), .inputs_330__1 (registerOutputs_330__1), .inputs_330__0 (
            registerOutputs_330__0), .inputs_331__15 (registerOutputs_331__15), 
            .inputs_331__14 (registerOutputs_331__14), .inputs_331__13 (
            registerOutputs_331__13), .inputs_331__12 (registerOutputs_331__12)
            , .inputs_331__11 (registerOutputs_331__11), .inputs_331__10 (
            registerOutputs_331__10), .inputs_331__9 (registerOutputs_331__9), .inputs_331__8 (
            registerOutputs_331__8), .inputs_331__7 (registerOutputs_331__7), .inputs_331__6 (
            registerOutputs_331__6), .inputs_331__5 (registerOutputs_331__5), .inputs_331__4 (
            registerOutputs_331__4), .inputs_331__3 (registerOutputs_331__3), .inputs_331__2 (
            registerOutputs_331__2), .inputs_331__1 (registerOutputs_331__1), .inputs_331__0 (
            registerOutputs_331__0), .inputs_332__15 (registerOutputs_332__15), 
            .inputs_332__14 (registerOutputs_332__14), .inputs_332__13 (
            registerOutputs_332__13), .inputs_332__12 (registerOutputs_332__12)
            , .inputs_332__11 (registerOutputs_332__11), .inputs_332__10 (
            registerOutputs_332__10), .inputs_332__9 (registerOutputs_332__9), .inputs_332__8 (
            registerOutputs_332__8), .inputs_332__7 (registerOutputs_332__7), .inputs_332__6 (
            registerOutputs_332__6), .inputs_332__5 (registerOutputs_332__5), .inputs_332__4 (
            registerOutputs_332__4), .inputs_332__3 (registerOutputs_332__3), .inputs_332__2 (
            registerOutputs_332__2), .inputs_332__1 (registerOutputs_332__1), .inputs_332__0 (
            registerOutputs_332__0), .inputs_333__15 (registerOutputs_333__15), 
            .inputs_333__14 (registerOutputs_333__14), .inputs_333__13 (
            registerOutputs_333__13), .inputs_333__12 (registerOutputs_333__12)
            , .inputs_333__11 (registerOutputs_333__11), .inputs_333__10 (
            registerOutputs_333__10), .inputs_333__9 (registerOutputs_333__9), .inputs_333__8 (
            registerOutputs_333__8), .inputs_333__7 (registerOutputs_333__7), .inputs_333__6 (
            registerOutputs_333__6), .inputs_333__5 (registerOutputs_333__5), .inputs_333__4 (
            registerOutputs_333__4), .inputs_333__3 (registerOutputs_333__3), .inputs_333__2 (
            registerOutputs_333__2), .inputs_333__1 (registerOutputs_333__1), .inputs_333__0 (
            registerOutputs_333__0), .inputs_334__15 (registerOutputs_334__15), 
            .inputs_334__14 (registerOutputs_334__14), .inputs_334__13 (
            registerOutputs_334__13), .inputs_334__12 (registerOutputs_334__12)
            , .inputs_334__11 (registerOutputs_334__11), .inputs_334__10 (
            registerOutputs_334__10), .inputs_334__9 (registerOutputs_334__9), .inputs_334__8 (
            registerOutputs_334__8), .inputs_334__7 (registerOutputs_334__7), .inputs_334__6 (
            registerOutputs_334__6), .inputs_334__5 (registerOutputs_334__5), .inputs_334__4 (
            registerOutputs_334__4), .inputs_334__3 (registerOutputs_334__3), .inputs_334__2 (
            registerOutputs_334__2), .inputs_334__1 (registerOutputs_334__1), .inputs_334__0 (
            registerOutputs_334__0), .inputs_335__15 (registerOutputs_335__15), 
            .inputs_335__14 (registerOutputs_335__14), .inputs_335__13 (
            registerOutputs_335__13), .inputs_335__12 (registerOutputs_335__12)
            , .inputs_335__11 (registerOutputs_335__11), .inputs_335__10 (
            registerOutputs_335__10), .inputs_335__9 (registerOutputs_335__9), .inputs_335__8 (
            registerOutputs_335__8), .inputs_335__7 (registerOutputs_335__7), .inputs_335__6 (
            registerOutputs_335__6), .inputs_335__5 (registerOutputs_335__5), .inputs_335__4 (
            registerOutputs_335__4), .inputs_335__3 (registerOutputs_335__3), .inputs_335__2 (
            registerOutputs_335__2), .inputs_335__1 (registerOutputs_335__1), .inputs_335__0 (
            registerOutputs_335__0), .inputs_336__15 (registerOutputs_336__15), 
            .inputs_336__14 (registerOutputs_336__14), .inputs_336__13 (
            registerOutputs_336__13), .inputs_336__12 (registerOutputs_336__12)
            , .inputs_336__11 (registerOutputs_336__11), .inputs_336__10 (
            registerOutputs_336__10), .inputs_336__9 (registerOutputs_336__9), .inputs_336__8 (
            registerOutputs_336__8), .inputs_336__7 (registerOutputs_336__7), .inputs_336__6 (
            registerOutputs_336__6), .inputs_336__5 (registerOutputs_336__5), .inputs_336__4 (
            registerOutputs_336__4), .inputs_336__3 (registerOutputs_336__3), .inputs_336__2 (
            registerOutputs_336__2), .inputs_336__1 (registerOutputs_336__1), .inputs_336__0 (
            registerOutputs_336__0), .inputs_337__15 (registerOutputs_337__15), 
            .inputs_337__14 (registerOutputs_337__14), .inputs_337__13 (
            registerOutputs_337__13), .inputs_337__12 (registerOutputs_337__12)
            , .inputs_337__11 (registerOutputs_337__11), .inputs_337__10 (
            registerOutputs_337__10), .inputs_337__9 (registerOutputs_337__9), .inputs_337__8 (
            registerOutputs_337__8), .inputs_337__7 (registerOutputs_337__7), .inputs_337__6 (
            registerOutputs_337__6), .inputs_337__5 (registerOutputs_337__5), .inputs_337__4 (
            registerOutputs_337__4), .inputs_337__3 (registerOutputs_337__3), .inputs_337__2 (
            registerOutputs_337__2), .inputs_337__1 (registerOutputs_337__1), .inputs_337__0 (
            registerOutputs_337__0), .inputs_338__15 (registerOutputs_338__15), 
            .inputs_338__14 (registerOutputs_338__14), .inputs_338__13 (
            registerOutputs_338__13), .inputs_338__12 (registerOutputs_338__12)
            , .inputs_338__11 (registerOutputs_338__11), .inputs_338__10 (
            registerOutputs_338__10), .inputs_338__9 (registerOutputs_338__9), .inputs_338__8 (
            registerOutputs_338__8), .inputs_338__7 (registerOutputs_338__7), .inputs_338__6 (
            registerOutputs_338__6), .inputs_338__5 (registerOutputs_338__5), .inputs_338__4 (
            registerOutputs_338__4), .inputs_338__3 (registerOutputs_338__3), .inputs_338__2 (
            registerOutputs_338__2), .inputs_338__1 (registerOutputs_338__1), .inputs_338__0 (
            registerOutputs_338__0), .inputs_339__15 (registerOutputs_339__15), 
            .inputs_339__14 (registerOutputs_339__14), .inputs_339__13 (
            registerOutputs_339__13), .inputs_339__12 (registerOutputs_339__12)
            , .inputs_339__11 (registerOutputs_339__11), .inputs_339__10 (
            registerOutputs_339__10), .inputs_339__9 (registerOutputs_339__9), .inputs_339__8 (
            registerOutputs_339__8), .inputs_339__7 (registerOutputs_339__7), .inputs_339__6 (
            registerOutputs_339__6), .inputs_339__5 (registerOutputs_339__5), .inputs_339__4 (
            registerOutputs_339__4), .inputs_339__3 (registerOutputs_339__3), .inputs_339__2 (
            registerOutputs_339__2), .inputs_339__1 (registerOutputs_339__1), .inputs_339__0 (
            registerOutputs_339__0), .inputs_340__15 (registerOutputs_340__15), 
            .inputs_340__14 (registerOutputs_340__14), .inputs_340__13 (
            registerOutputs_340__13), .inputs_340__12 (registerOutputs_340__12)
            , .inputs_340__11 (registerOutputs_340__11), .inputs_340__10 (
            registerOutputs_340__10), .inputs_340__9 (registerOutputs_340__9), .inputs_340__8 (
            registerOutputs_340__8), .inputs_340__7 (registerOutputs_340__7), .inputs_340__6 (
            registerOutputs_340__6), .inputs_340__5 (registerOutputs_340__5), .inputs_340__4 (
            registerOutputs_340__4), .inputs_340__3 (registerOutputs_340__3), .inputs_340__2 (
            registerOutputs_340__2), .inputs_340__1 (registerOutputs_340__1), .inputs_340__0 (
            registerOutputs_340__0), .inputs_341__15 (registerOutputs_341__15), 
            .inputs_341__14 (registerOutputs_341__14), .inputs_341__13 (
            registerOutputs_341__13), .inputs_341__12 (registerOutputs_341__12)
            , .inputs_341__11 (registerOutputs_341__11), .inputs_341__10 (
            registerOutputs_341__10), .inputs_341__9 (registerOutputs_341__9), .inputs_341__8 (
            registerOutputs_341__8), .inputs_341__7 (registerOutputs_341__7), .inputs_341__6 (
            registerOutputs_341__6), .inputs_341__5 (registerOutputs_341__5), .inputs_341__4 (
            registerOutputs_341__4), .inputs_341__3 (registerOutputs_341__3), .inputs_341__2 (
            registerOutputs_341__2), .inputs_341__1 (registerOutputs_341__1), .inputs_341__0 (
            registerOutputs_341__0), .inputs_342__15 (registerOutputs_342__15), 
            .inputs_342__14 (registerOutputs_342__14), .inputs_342__13 (
            registerOutputs_342__13), .inputs_342__12 (registerOutputs_342__12)
            , .inputs_342__11 (registerOutputs_342__11), .inputs_342__10 (
            registerOutputs_342__10), .inputs_342__9 (registerOutputs_342__9), .inputs_342__8 (
            registerOutputs_342__8), .inputs_342__7 (registerOutputs_342__7), .inputs_342__6 (
            registerOutputs_342__6), .inputs_342__5 (registerOutputs_342__5), .inputs_342__4 (
            registerOutputs_342__4), .inputs_342__3 (registerOutputs_342__3), .inputs_342__2 (
            registerOutputs_342__2), .inputs_342__1 (registerOutputs_342__1), .inputs_342__0 (
            registerOutputs_342__0), .inputs_343__15 (registerOutputs_343__15), 
            .inputs_343__14 (registerOutputs_343__14), .inputs_343__13 (
            registerOutputs_343__13), .inputs_343__12 (registerOutputs_343__12)
            , .inputs_343__11 (registerOutputs_343__11), .inputs_343__10 (
            registerOutputs_343__10), .inputs_343__9 (registerOutputs_343__9), .inputs_343__8 (
            registerOutputs_343__8), .inputs_343__7 (registerOutputs_343__7), .inputs_343__6 (
            registerOutputs_343__6), .inputs_343__5 (registerOutputs_343__5), .inputs_343__4 (
            registerOutputs_343__4), .inputs_343__3 (registerOutputs_343__3), .inputs_343__2 (
            registerOutputs_343__2), .inputs_343__1 (registerOutputs_343__1), .inputs_343__0 (
            registerOutputs_343__0), .inputs_344__15 (registerOutputs_344__15), 
            .inputs_344__14 (registerOutputs_344__14), .inputs_344__13 (
            registerOutputs_344__13), .inputs_344__12 (registerOutputs_344__12)
            , .inputs_344__11 (registerOutputs_344__11), .inputs_344__10 (
            registerOutputs_344__10), .inputs_344__9 (registerOutputs_344__9), .inputs_344__8 (
            registerOutputs_344__8), .inputs_344__7 (registerOutputs_344__7), .inputs_344__6 (
            registerOutputs_344__6), .inputs_344__5 (registerOutputs_344__5), .inputs_344__4 (
            registerOutputs_344__4), .inputs_344__3 (registerOutputs_344__3), .inputs_344__2 (
            registerOutputs_344__2), .inputs_344__1 (registerOutputs_344__1), .inputs_344__0 (
            registerOutputs_344__0), .inputs_345__15 (registerOutputs_345__15), 
            .inputs_345__14 (registerOutputs_345__14), .inputs_345__13 (
            registerOutputs_345__13), .inputs_345__12 (registerOutputs_345__12)
            , .inputs_345__11 (registerOutputs_345__11), .inputs_345__10 (
            registerOutputs_345__10), .inputs_345__9 (registerOutputs_345__9), .inputs_345__8 (
            registerOutputs_345__8), .inputs_345__7 (registerOutputs_345__7), .inputs_345__6 (
            registerOutputs_345__6), .inputs_345__5 (registerOutputs_345__5), .inputs_345__4 (
            registerOutputs_345__4), .inputs_345__3 (registerOutputs_345__3), .inputs_345__2 (
            registerOutputs_345__2), .inputs_345__1 (registerOutputs_345__1), .inputs_345__0 (
            registerOutputs_345__0), .inputs_346__15 (registerOutputs_346__15), 
            .inputs_346__14 (registerOutputs_346__14), .inputs_346__13 (
            registerOutputs_346__13), .inputs_346__12 (registerOutputs_346__12)
            , .inputs_346__11 (registerOutputs_346__11), .inputs_346__10 (
            registerOutputs_346__10), .inputs_346__9 (registerOutputs_346__9), .inputs_346__8 (
            registerOutputs_346__8), .inputs_346__7 (registerOutputs_346__7), .inputs_346__6 (
            registerOutputs_346__6), .inputs_346__5 (registerOutputs_346__5), .inputs_346__4 (
            registerOutputs_346__4), .inputs_346__3 (registerOutputs_346__3), .inputs_346__2 (
            registerOutputs_346__2), .inputs_346__1 (registerOutputs_346__1), .inputs_346__0 (
            registerOutputs_346__0), .inputs_347__15 (registerOutputs_347__15), 
            .inputs_347__14 (registerOutputs_347__14), .inputs_347__13 (
            registerOutputs_347__13), .inputs_347__12 (registerOutputs_347__12)
            , .inputs_347__11 (registerOutputs_347__11), .inputs_347__10 (
            registerOutputs_347__10), .inputs_347__9 (registerOutputs_347__9), .inputs_347__8 (
            registerOutputs_347__8), .inputs_347__7 (registerOutputs_347__7), .inputs_347__6 (
            registerOutputs_347__6), .inputs_347__5 (registerOutputs_347__5), .inputs_347__4 (
            registerOutputs_347__4), .inputs_347__3 (registerOutputs_347__3), .inputs_347__2 (
            registerOutputs_347__2), .inputs_347__1 (registerOutputs_347__1), .inputs_347__0 (
            registerOutputs_347__0), .inputs_348__15 (registerOutputs_348__15), 
            .inputs_348__14 (registerOutputs_348__14), .inputs_348__13 (
            registerOutputs_348__13), .inputs_348__12 (registerOutputs_348__12)
            , .inputs_348__11 (registerOutputs_348__11), .inputs_348__10 (
            registerOutputs_348__10), .inputs_348__9 (registerOutputs_348__9), .inputs_348__8 (
            registerOutputs_348__8), .inputs_348__7 (registerOutputs_348__7), .inputs_348__6 (
            registerOutputs_348__6), .inputs_348__5 (registerOutputs_348__5), .inputs_348__4 (
            registerOutputs_348__4), .inputs_348__3 (registerOutputs_348__3), .inputs_348__2 (
            registerOutputs_348__2), .inputs_348__1 (registerOutputs_348__1), .inputs_348__0 (
            registerOutputs_348__0), .inputs_349__15 (registerOutputs_349__15), 
            .inputs_349__14 (registerOutputs_349__14), .inputs_349__13 (
            registerOutputs_349__13), .inputs_349__12 (registerOutputs_349__12)
            , .inputs_349__11 (registerOutputs_349__11), .inputs_349__10 (
            registerOutputs_349__10), .inputs_349__9 (registerOutputs_349__9), .inputs_349__8 (
            registerOutputs_349__8), .inputs_349__7 (registerOutputs_349__7), .inputs_349__6 (
            registerOutputs_349__6), .inputs_349__5 (registerOutputs_349__5), .inputs_349__4 (
            registerOutputs_349__4), .inputs_349__3 (registerOutputs_349__3), .inputs_349__2 (
            registerOutputs_349__2), .inputs_349__1 (registerOutputs_349__1), .inputs_349__0 (
            registerOutputs_349__0), .inputs_350__15 (registerOutputs_350__15), 
            .inputs_350__14 (registerOutputs_350__14), .inputs_350__13 (
            registerOutputs_350__13), .inputs_350__12 (registerOutputs_350__12)
            , .inputs_350__11 (registerOutputs_350__11), .inputs_350__10 (
            registerOutputs_350__10), .inputs_350__9 (registerOutputs_350__9), .inputs_350__8 (
            registerOutputs_350__8), .inputs_350__7 (registerOutputs_350__7), .inputs_350__6 (
            registerOutputs_350__6), .inputs_350__5 (registerOutputs_350__5), .inputs_350__4 (
            registerOutputs_350__4), .inputs_350__3 (registerOutputs_350__3), .inputs_350__2 (
            registerOutputs_350__2), .inputs_350__1 (registerOutputs_350__1), .inputs_350__0 (
            registerOutputs_350__0), .inputs_351__15 (registerOutputs_351__15), 
            .inputs_351__14 (registerOutputs_351__14), .inputs_351__13 (
            registerOutputs_351__13), .inputs_351__12 (registerOutputs_351__12)
            , .inputs_351__11 (registerOutputs_351__11), .inputs_351__10 (
            registerOutputs_351__10), .inputs_351__9 (registerOutputs_351__9), .inputs_351__8 (
            registerOutputs_351__8), .inputs_351__7 (registerOutputs_351__7), .inputs_351__6 (
            registerOutputs_351__6), .inputs_351__5 (registerOutputs_351__5), .inputs_351__4 (
            registerOutputs_351__4), .inputs_351__3 (registerOutputs_351__3), .inputs_351__2 (
            registerOutputs_351__2), .inputs_351__1 (registerOutputs_351__1), .inputs_351__0 (
            registerOutputs_351__0), .inputs_352__15 (registerOutputs_352__15), 
            .inputs_352__14 (registerOutputs_352__14), .inputs_352__13 (
            registerOutputs_352__13), .inputs_352__12 (registerOutputs_352__12)
            , .inputs_352__11 (registerOutputs_352__11), .inputs_352__10 (
            registerOutputs_352__10), .inputs_352__9 (registerOutputs_352__9), .inputs_352__8 (
            registerOutputs_352__8), .inputs_352__7 (registerOutputs_352__7), .inputs_352__6 (
            registerOutputs_352__6), .inputs_352__5 (registerOutputs_352__5), .inputs_352__4 (
            registerOutputs_352__4), .inputs_352__3 (registerOutputs_352__3), .inputs_352__2 (
            registerOutputs_352__2), .inputs_352__1 (registerOutputs_352__1), .inputs_352__0 (
            registerOutputs_352__0), .inputs_353__15 (registerOutputs_353__15), 
            .inputs_353__14 (registerOutputs_353__14), .inputs_353__13 (
            registerOutputs_353__13), .inputs_353__12 (registerOutputs_353__12)
            , .inputs_353__11 (registerOutputs_353__11), .inputs_353__10 (
            registerOutputs_353__10), .inputs_353__9 (registerOutputs_353__9), .inputs_353__8 (
            registerOutputs_353__8), .inputs_353__7 (registerOutputs_353__7), .inputs_353__6 (
            registerOutputs_353__6), .inputs_353__5 (registerOutputs_353__5), .inputs_353__4 (
            registerOutputs_353__4), .inputs_353__3 (registerOutputs_353__3), .inputs_353__2 (
            registerOutputs_353__2), .inputs_353__1 (registerOutputs_353__1), .inputs_353__0 (
            registerOutputs_353__0), .inputs_354__15 (registerOutputs_354__15), 
            .inputs_354__14 (registerOutputs_354__14), .inputs_354__13 (
            registerOutputs_354__13), .inputs_354__12 (registerOutputs_354__12)
            , .inputs_354__11 (registerOutputs_354__11), .inputs_354__10 (
            registerOutputs_354__10), .inputs_354__9 (registerOutputs_354__9), .inputs_354__8 (
            registerOutputs_354__8), .inputs_354__7 (registerOutputs_354__7), .inputs_354__6 (
            registerOutputs_354__6), .inputs_354__5 (registerOutputs_354__5), .inputs_354__4 (
            registerOutputs_354__4), .inputs_354__3 (registerOutputs_354__3), .inputs_354__2 (
            registerOutputs_354__2), .inputs_354__1 (registerOutputs_354__1), .inputs_354__0 (
            registerOutputs_354__0), .inputs_355__15 (registerOutputs_355__15), 
            .inputs_355__14 (registerOutputs_355__14), .inputs_355__13 (
            registerOutputs_355__13), .inputs_355__12 (registerOutputs_355__12)
            , .inputs_355__11 (registerOutputs_355__11), .inputs_355__10 (
            registerOutputs_355__10), .inputs_355__9 (registerOutputs_355__9), .inputs_355__8 (
            registerOutputs_355__8), .inputs_355__7 (registerOutputs_355__7), .inputs_355__6 (
            registerOutputs_355__6), .inputs_355__5 (registerOutputs_355__5), .inputs_355__4 (
            registerOutputs_355__4), .inputs_355__3 (registerOutputs_355__3), .inputs_355__2 (
            registerOutputs_355__2), .inputs_355__1 (registerOutputs_355__1), .inputs_355__0 (
            registerOutputs_355__0), .inputs_356__15 (registerOutputs_356__15), 
            .inputs_356__14 (registerOutputs_356__14), .inputs_356__13 (
            registerOutputs_356__13), .inputs_356__12 (registerOutputs_356__12)
            , .inputs_356__11 (registerOutputs_356__11), .inputs_356__10 (
            registerOutputs_356__10), .inputs_356__9 (registerOutputs_356__9), .inputs_356__8 (
            registerOutputs_356__8), .inputs_356__7 (registerOutputs_356__7), .inputs_356__6 (
            registerOutputs_356__6), .inputs_356__5 (registerOutputs_356__5), .inputs_356__4 (
            registerOutputs_356__4), .inputs_356__3 (registerOutputs_356__3), .inputs_356__2 (
            registerOutputs_356__2), .inputs_356__1 (registerOutputs_356__1), .inputs_356__0 (
            registerOutputs_356__0), .inputs_357__15 (registerOutputs_357__15), 
            .inputs_357__14 (registerOutputs_357__14), .inputs_357__13 (
            registerOutputs_357__13), .inputs_357__12 (registerOutputs_357__12)
            , .inputs_357__11 (registerOutputs_357__11), .inputs_357__10 (
            registerOutputs_357__10), .inputs_357__9 (registerOutputs_357__9), .inputs_357__8 (
            registerOutputs_357__8), .inputs_357__7 (registerOutputs_357__7), .inputs_357__6 (
            registerOutputs_357__6), .inputs_357__5 (registerOutputs_357__5), .inputs_357__4 (
            registerOutputs_357__4), .inputs_357__3 (registerOutputs_357__3), .inputs_357__2 (
            registerOutputs_357__2), .inputs_357__1 (registerOutputs_357__1), .inputs_357__0 (
            registerOutputs_357__0), .inputs_358__15 (registerOutputs_358__15), 
            .inputs_358__14 (registerOutputs_358__14), .inputs_358__13 (
            registerOutputs_358__13), .inputs_358__12 (registerOutputs_358__12)
            , .inputs_358__11 (registerOutputs_358__11), .inputs_358__10 (
            registerOutputs_358__10), .inputs_358__9 (registerOutputs_358__9), .inputs_358__8 (
            registerOutputs_358__8), .inputs_358__7 (registerOutputs_358__7), .inputs_358__6 (
            registerOutputs_358__6), .inputs_358__5 (registerOutputs_358__5), .inputs_358__4 (
            registerOutputs_358__4), .inputs_358__3 (registerOutputs_358__3), .inputs_358__2 (
            registerOutputs_358__2), .inputs_358__1 (registerOutputs_358__1), .inputs_358__0 (
            registerOutputs_358__0), .inputs_359__15 (registerOutputs_359__15), 
            .inputs_359__14 (registerOutputs_359__14), .inputs_359__13 (
            registerOutputs_359__13), .inputs_359__12 (registerOutputs_359__12)
            , .inputs_359__11 (registerOutputs_359__11), .inputs_359__10 (
            registerOutputs_359__10), .inputs_359__9 (registerOutputs_359__9), .inputs_359__8 (
            registerOutputs_359__8), .inputs_359__7 (registerOutputs_359__7), .inputs_359__6 (
            registerOutputs_359__6), .inputs_359__5 (registerOutputs_359__5), .inputs_359__4 (
            registerOutputs_359__4), .inputs_359__3 (registerOutputs_359__3), .inputs_359__2 (
            registerOutputs_359__2), .inputs_359__1 (registerOutputs_359__1), .inputs_359__0 (
            registerOutputs_359__0), .inputs_360__15 (registerOutputs_360__15), 
            .inputs_360__14 (registerOutputs_360__14), .inputs_360__13 (
            registerOutputs_360__13), .inputs_360__12 (registerOutputs_360__12)
            , .inputs_360__11 (registerOutputs_360__11), .inputs_360__10 (
            registerOutputs_360__10), .inputs_360__9 (registerOutputs_360__9), .inputs_360__8 (
            registerOutputs_360__8), .inputs_360__7 (registerOutputs_360__7), .inputs_360__6 (
            registerOutputs_360__6), .inputs_360__5 (registerOutputs_360__5), .inputs_360__4 (
            registerOutputs_360__4), .inputs_360__3 (registerOutputs_360__3), .inputs_360__2 (
            registerOutputs_360__2), .inputs_360__1 (registerOutputs_360__1), .inputs_360__0 (
            registerOutputs_360__0), .inputs_361__15 (registerOutputs_361__15), 
            .inputs_361__14 (registerOutputs_361__14), .inputs_361__13 (
            registerOutputs_361__13), .inputs_361__12 (registerOutputs_361__12)
            , .inputs_361__11 (registerOutputs_361__11), .inputs_361__10 (
            registerOutputs_361__10), .inputs_361__9 (registerOutputs_361__9), .inputs_361__8 (
            registerOutputs_361__8), .inputs_361__7 (registerOutputs_361__7), .inputs_361__6 (
            registerOutputs_361__6), .inputs_361__5 (registerOutputs_361__5), .inputs_361__4 (
            registerOutputs_361__4), .inputs_361__3 (registerOutputs_361__3), .inputs_361__2 (
            registerOutputs_361__2), .inputs_361__1 (registerOutputs_361__1), .inputs_361__0 (
            registerOutputs_361__0), .inputs_362__15 (registerOutputs_362__15), 
            .inputs_362__14 (registerOutputs_362__14), .inputs_362__13 (
            registerOutputs_362__13), .inputs_362__12 (registerOutputs_362__12)
            , .inputs_362__11 (registerOutputs_362__11), .inputs_362__10 (
            registerOutputs_362__10), .inputs_362__9 (registerOutputs_362__9), .inputs_362__8 (
            registerOutputs_362__8), .inputs_362__7 (registerOutputs_362__7), .inputs_362__6 (
            registerOutputs_362__6), .inputs_362__5 (registerOutputs_362__5), .inputs_362__4 (
            registerOutputs_362__4), .inputs_362__3 (registerOutputs_362__3), .inputs_362__2 (
            registerOutputs_362__2), .inputs_362__1 (registerOutputs_362__1), .inputs_362__0 (
            registerOutputs_362__0), .inputs_363__15 (registerOutputs_363__15), 
            .inputs_363__14 (registerOutputs_363__14), .inputs_363__13 (
            registerOutputs_363__13), .inputs_363__12 (registerOutputs_363__12)
            , .inputs_363__11 (registerOutputs_363__11), .inputs_363__10 (
            registerOutputs_363__10), .inputs_363__9 (registerOutputs_363__9), .inputs_363__8 (
            registerOutputs_363__8), .inputs_363__7 (registerOutputs_363__7), .inputs_363__6 (
            registerOutputs_363__6), .inputs_363__5 (registerOutputs_363__5), .inputs_363__4 (
            registerOutputs_363__4), .inputs_363__3 (registerOutputs_363__3), .inputs_363__2 (
            registerOutputs_363__2), .inputs_363__1 (registerOutputs_363__1), .inputs_363__0 (
            registerOutputs_363__0), .inputs_364__15 (registerOutputs_364__15), 
            .inputs_364__14 (registerOutputs_364__14), .inputs_364__13 (
            registerOutputs_364__13), .inputs_364__12 (registerOutputs_364__12)
            , .inputs_364__11 (registerOutputs_364__11), .inputs_364__10 (
            registerOutputs_364__10), .inputs_364__9 (registerOutputs_364__9), .inputs_364__8 (
            registerOutputs_364__8), .inputs_364__7 (registerOutputs_364__7), .inputs_364__6 (
            registerOutputs_364__6), .inputs_364__5 (registerOutputs_364__5), .inputs_364__4 (
            registerOutputs_364__4), .inputs_364__3 (registerOutputs_364__3), .inputs_364__2 (
            registerOutputs_364__2), .inputs_364__1 (registerOutputs_364__1), .inputs_364__0 (
            registerOutputs_364__0), .inputs_365__15 (registerOutputs_365__15), 
            .inputs_365__14 (registerOutputs_365__14), .inputs_365__13 (
            registerOutputs_365__13), .inputs_365__12 (registerOutputs_365__12)
            , .inputs_365__11 (registerOutputs_365__11), .inputs_365__10 (
            registerOutputs_365__10), .inputs_365__9 (registerOutputs_365__9), .inputs_365__8 (
            registerOutputs_365__8), .inputs_365__7 (registerOutputs_365__7), .inputs_365__6 (
            registerOutputs_365__6), .inputs_365__5 (registerOutputs_365__5), .inputs_365__4 (
            registerOutputs_365__4), .inputs_365__3 (registerOutputs_365__3), .inputs_365__2 (
            registerOutputs_365__2), .inputs_365__1 (registerOutputs_365__1), .inputs_365__0 (
            registerOutputs_365__0), .inputs_366__15 (registerOutputs_366__15), 
            .inputs_366__14 (registerOutputs_366__14), .inputs_366__13 (
            registerOutputs_366__13), .inputs_366__12 (registerOutputs_366__12)
            , .inputs_366__11 (registerOutputs_366__11), .inputs_366__10 (
            registerOutputs_366__10), .inputs_366__9 (registerOutputs_366__9), .inputs_366__8 (
            registerOutputs_366__8), .inputs_366__7 (registerOutputs_366__7), .inputs_366__6 (
            registerOutputs_366__6), .inputs_366__5 (registerOutputs_366__5), .inputs_366__4 (
            registerOutputs_366__4), .inputs_366__3 (registerOutputs_366__3), .inputs_366__2 (
            registerOutputs_366__2), .inputs_366__1 (registerOutputs_366__1), .inputs_366__0 (
            registerOutputs_366__0), .inputs_367__15 (registerOutputs_367__15), 
            .inputs_367__14 (registerOutputs_367__14), .inputs_367__13 (
            registerOutputs_367__13), .inputs_367__12 (registerOutputs_367__12)
            , .inputs_367__11 (registerOutputs_367__11), .inputs_367__10 (
            registerOutputs_367__10), .inputs_367__9 (registerOutputs_367__9), .inputs_367__8 (
            registerOutputs_367__8), .inputs_367__7 (registerOutputs_367__7), .inputs_367__6 (
            registerOutputs_367__6), .inputs_367__5 (registerOutputs_367__5), .inputs_367__4 (
            registerOutputs_367__4), .inputs_367__3 (registerOutputs_367__3), .inputs_367__2 (
            registerOutputs_367__2), .inputs_367__1 (registerOutputs_367__1), .inputs_367__0 (
            registerOutputs_367__0), .inputs_368__15 (registerOutputs_368__15), 
            .inputs_368__14 (registerOutputs_368__14), .inputs_368__13 (
            registerOutputs_368__13), .inputs_368__12 (registerOutputs_368__12)
            , .inputs_368__11 (registerOutputs_368__11), .inputs_368__10 (
            registerOutputs_368__10), .inputs_368__9 (registerOutputs_368__9), .inputs_368__8 (
            registerOutputs_368__8), .inputs_368__7 (registerOutputs_368__7), .inputs_368__6 (
            registerOutputs_368__6), .inputs_368__5 (registerOutputs_368__5), .inputs_368__4 (
            registerOutputs_368__4), .inputs_368__3 (registerOutputs_368__3), .inputs_368__2 (
            registerOutputs_368__2), .inputs_368__1 (registerOutputs_368__1), .inputs_368__0 (
            registerOutputs_368__0), .inputs_369__15 (registerOutputs_369__15), 
            .inputs_369__14 (registerOutputs_369__14), .inputs_369__13 (
            registerOutputs_369__13), .inputs_369__12 (registerOutputs_369__12)
            , .inputs_369__11 (registerOutputs_369__11), .inputs_369__10 (
            registerOutputs_369__10), .inputs_369__9 (registerOutputs_369__9), .inputs_369__8 (
            registerOutputs_369__8), .inputs_369__7 (registerOutputs_369__7), .inputs_369__6 (
            registerOutputs_369__6), .inputs_369__5 (registerOutputs_369__5), .inputs_369__4 (
            registerOutputs_369__4), .inputs_369__3 (registerOutputs_369__3), .inputs_369__2 (
            registerOutputs_369__2), .inputs_369__1 (registerOutputs_369__1), .inputs_369__0 (
            registerOutputs_369__0), .inputs_370__15 (registerOutputs_370__15), 
            .inputs_370__14 (registerOutputs_370__14), .inputs_370__13 (
            registerOutputs_370__13), .inputs_370__12 (registerOutputs_370__12)
            , .inputs_370__11 (registerOutputs_370__11), .inputs_370__10 (
            registerOutputs_370__10), .inputs_370__9 (registerOutputs_370__9), .inputs_370__8 (
            registerOutputs_370__8), .inputs_370__7 (registerOutputs_370__7), .inputs_370__6 (
            registerOutputs_370__6), .inputs_370__5 (registerOutputs_370__5), .inputs_370__4 (
            registerOutputs_370__4), .inputs_370__3 (registerOutputs_370__3), .inputs_370__2 (
            registerOutputs_370__2), .inputs_370__1 (registerOutputs_370__1), .inputs_370__0 (
            registerOutputs_370__0), .inputs_371__15 (registerOutputs_371__15), 
            .inputs_371__14 (registerOutputs_371__14), .inputs_371__13 (
            registerOutputs_371__13), .inputs_371__12 (registerOutputs_371__12)
            , .inputs_371__11 (registerOutputs_371__11), .inputs_371__10 (
            registerOutputs_371__10), .inputs_371__9 (registerOutputs_371__9), .inputs_371__8 (
            registerOutputs_371__8), .inputs_371__7 (registerOutputs_371__7), .inputs_371__6 (
            registerOutputs_371__6), .inputs_371__5 (registerOutputs_371__5), .inputs_371__4 (
            registerOutputs_371__4), .inputs_371__3 (registerOutputs_371__3), .inputs_371__2 (
            registerOutputs_371__2), .inputs_371__1 (registerOutputs_371__1), .inputs_371__0 (
            registerOutputs_371__0), .inputs_372__15 (registerOutputs_372__15), 
            .inputs_372__14 (registerOutputs_372__14), .inputs_372__13 (
            registerOutputs_372__13), .inputs_372__12 (registerOutputs_372__12)
            , .inputs_372__11 (registerOutputs_372__11), .inputs_372__10 (
            registerOutputs_372__10), .inputs_372__9 (registerOutputs_372__9), .inputs_372__8 (
            registerOutputs_372__8), .inputs_372__7 (registerOutputs_372__7), .inputs_372__6 (
            registerOutputs_372__6), .inputs_372__5 (registerOutputs_372__5), .inputs_372__4 (
            registerOutputs_372__4), .inputs_372__3 (registerOutputs_372__3), .inputs_372__2 (
            registerOutputs_372__2), .inputs_372__1 (registerOutputs_372__1), .inputs_372__0 (
            registerOutputs_372__0), .inputs_373__15 (registerOutputs_373__15), 
            .inputs_373__14 (registerOutputs_373__14), .inputs_373__13 (
            registerOutputs_373__13), .inputs_373__12 (registerOutputs_373__12)
            , .inputs_373__11 (registerOutputs_373__11), .inputs_373__10 (
            registerOutputs_373__10), .inputs_373__9 (registerOutputs_373__9), .inputs_373__8 (
            registerOutputs_373__8), .inputs_373__7 (registerOutputs_373__7), .inputs_373__6 (
            registerOutputs_373__6), .inputs_373__5 (registerOutputs_373__5), .inputs_373__4 (
            registerOutputs_373__4), .inputs_373__3 (registerOutputs_373__3), .inputs_373__2 (
            registerOutputs_373__2), .inputs_373__1 (registerOutputs_373__1), .inputs_373__0 (
            registerOutputs_373__0), .inputs_374__15 (registerOutputs_374__15), 
            .inputs_374__14 (registerOutputs_374__14), .inputs_374__13 (
            registerOutputs_374__13), .inputs_374__12 (registerOutputs_374__12)
            , .inputs_374__11 (registerOutputs_374__11), .inputs_374__10 (
            registerOutputs_374__10), .inputs_374__9 (registerOutputs_374__9), .inputs_374__8 (
            registerOutputs_374__8), .inputs_374__7 (registerOutputs_374__7), .inputs_374__6 (
            registerOutputs_374__6), .inputs_374__5 (registerOutputs_374__5), .inputs_374__4 (
            registerOutputs_374__4), .inputs_374__3 (registerOutputs_374__3), .inputs_374__2 (
            registerOutputs_374__2), .inputs_374__1 (registerOutputs_374__1), .inputs_374__0 (
            registerOutputs_374__0), .inputs_375__15 (registerOutputs_375__15), 
            .inputs_375__14 (registerOutputs_375__14), .inputs_375__13 (
            registerOutputs_375__13), .inputs_375__12 (registerOutputs_375__12)
            , .inputs_375__11 (registerOutputs_375__11), .inputs_375__10 (
            registerOutputs_375__10), .inputs_375__9 (registerOutputs_375__9), .inputs_375__8 (
            registerOutputs_375__8), .inputs_375__7 (registerOutputs_375__7), .inputs_375__6 (
            registerOutputs_375__6), .inputs_375__5 (registerOutputs_375__5), .inputs_375__4 (
            registerOutputs_375__4), .inputs_375__3 (registerOutputs_375__3), .inputs_375__2 (
            registerOutputs_375__2), .inputs_375__1 (registerOutputs_375__1), .inputs_375__0 (
            registerOutputs_375__0), .inputs_376__15 (registerOutputs_376__15), 
            .inputs_376__14 (registerOutputs_376__14), .inputs_376__13 (
            registerOutputs_376__13), .inputs_376__12 (registerOutputs_376__12)
            , .inputs_376__11 (registerOutputs_376__11), .inputs_376__10 (
            registerOutputs_376__10), .inputs_376__9 (registerOutputs_376__9), .inputs_376__8 (
            registerOutputs_376__8), .inputs_376__7 (registerOutputs_376__7), .inputs_376__6 (
            registerOutputs_376__6), .inputs_376__5 (registerOutputs_376__5), .inputs_376__4 (
            registerOutputs_376__4), .inputs_376__3 (registerOutputs_376__3), .inputs_376__2 (
            registerOutputs_376__2), .inputs_376__1 (registerOutputs_376__1), .inputs_376__0 (
            registerOutputs_376__0), .inputs_377__15 (registerOutputs_377__15), 
            .inputs_377__14 (registerOutputs_377__14), .inputs_377__13 (
            registerOutputs_377__13), .inputs_377__12 (registerOutputs_377__12)
            , .inputs_377__11 (registerOutputs_377__11), .inputs_377__10 (
            registerOutputs_377__10), .inputs_377__9 (registerOutputs_377__9), .inputs_377__8 (
            registerOutputs_377__8), .inputs_377__7 (registerOutputs_377__7), .inputs_377__6 (
            registerOutputs_377__6), .inputs_377__5 (registerOutputs_377__5), .inputs_377__4 (
            registerOutputs_377__4), .inputs_377__3 (registerOutputs_377__3), .inputs_377__2 (
            registerOutputs_377__2), .inputs_377__1 (registerOutputs_377__1), .inputs_377__0 (
            registerOutputs_377__0), .inputs_378__15 (registerOutputs_378__15), 
            .inputs_378__14 (registerOutputs_378__14), .inputs_378__13 (
            registerOutputs_378__13), .inputs_378__12 (registerOutputs_378__12)
            , .inputs_378__11 (registerOutputs_378__11), .inputs_378__10 (
            registerOutputs_378__10), .inputs_378__9 (registerOutputs_378__9), .inputs_378__8 (
            registerOutputs_378__8), .inputs_378__7 (registerOutputs_378__7), .inputs_378__6 (
            registerOutputs_378__6), .inputs_378__5 (registerOutputs_378__5), .inputs_378__4 (
            registerOutputs_378__4), .inputs_378__3 (registerOutputs_378__3), .inputs_378__2 (
            registerOutputs_378__2), .inputs_378__1 (registerOutputs_378__1), .inputs_378__0 (
            registerOutputs_378__0), .inputs_379__15 (registerOutputs_379__15), 
            .inputs_379__14 (registerOutputs_379__14), .inputs_379__13 (
            registerOutputs_379__13), .inputs_379__12 (registerOutputs_379__12)
            , .inputs_379__11 (registerOutputs_379__11), .inputs_379__10 (
            registerOutputs_379__10), .inputs_379__9 (registerOutputs_379__9), .inputs_379__8 (
            registerOutputs_379__8), .inputs_379__7 (registerOutputs_379__7), .inputs_379__6 (
            registerOutputs_379__6), .inputs_379__5 (registerOutputs_379__5), .inputs_379__4 (
            registerOutputs_379__4), .inputs_379__3 (registerOutputs_379__3), .inputs_379__2 (
            registerOutputs_379__2), .inputs_379__1 (registerOutputs_379__1), .inputs_379__0 (
            registerOutputs_379__0), .inputs_380__15 (registerOutputs_380__15), 
            .inputs_380__14 (registerOutputs_380__14), .inputs_380__13 (
            registerOutputs_380__13), .inputs_380__12 (registerOutputs_380__12)
            , .inputs_380__11 (registerOutputs_380__11), .inputs_380__10 (
            registerOutputs_380__10), .inputs_380__9 (registerOutputs_380__9), .inputs_380__8 (
            registerOutputs_380__8), .inputs_380__7 (registerOutputs_380__7), .inputs_380__6 (
            registerOutputs_380__6), .inputs_380__5 (registerOutputs_380__5), .inputs_380__4 (
            registerOutputs_380__4), .inputs_380__3 (registerOutputs_380__3), .inputs_380__2 (
            registerOutputs_380__2), .inputs_380__1 (registerOutputs_380__1), .inputs_380__0 (
            registerOutputs_380__0), .inputs_381__15 (registerOutputs_381__15), 
            .inputs_381__14 (registerOutputs_381__14), .inputs_381__13 (
            registerOutputs_381__13), .inputs_381__12 (registerOutputs_381__12)
            , .inputs_381__11 (registerOutputs_381__11), .inputs_381__10 (
            registerOutputs_381__10), .inputs_381__9 (registerOutputs_381__9), .inputs_381__8 (
            registerOutputs_381__8), .inputs_381__7 (registerOutputs_381__7), .inputs_381__6 (
            registerOutputs_381__6), .inputs_381__5 (registerOutputs_381__5), .inputs_381__4 (
            registerOutputs_381__4), .inputs_381__3 (registerOutputs_381__3), .inputs_381__2 (
            registerOutputs_381__2), .inputs_381__1 (registerOutputs_381__1), .inputs_381__0 (
            registerOutputs_381__0), .inputs_382__15 (registerOutputs_382__15), 
            .inputs_382__14 (registerOutputs_382__14), .inputs_382__13 (
            registerOutputs_382__13), .inputs_382__12 (registerOutputs_382__12)
            , .inputs_382__11 (registerOutputs_382__11), .inputs_382__10 (
            registerOutputs_382__10), .inputs_382__9 (registerOutputs_382__9), .inputs_382__8 (
            registerOutputs_382__8), .inputs_382__7 (registerOutputs_382__7), .inputs_382__6 (
            registerOutputs_382__6), .inputs_382__5 (registerOutputs_382__5), .inputs_382__4 (
            registerOutputs_382__4), .inputs_382__3 (registerOutputs_382__3), .inputs_382__2 (
            registerOutputs_382__2), .inputs_382__1 (registerOutputs_382__1), .inputs_382__0 (
            registerOutputs_382__0), .inputs_383__15 (registerOutputs_383__15), 
            .inputs_383__14 (registerOutputs_383__14), .inputs_383__13 (
            registerOutputs_383__13), .inputs_383__12 (registerOutputs_383__12)
            , .inputs_383__11 (registerOutputs_383__11), .inputs_383__10 (
            registerOutputs_383__10), .inputs_383__9 (registerOutputs_383__9), .inputs_383__8 (
            registerOutputs_383__8), .inputs_383__7 (registerOutputs_383__7), .inputs_383__6 (
            registerOutputs_383__6), .inputs_383__5 (registerOutputs_383__5), .inputs_383__4 (
            registerOutputs_383__4), .inputs_383__3 (registerOutputs_383__3), .inputs_383__2 (
            registerOutputs_383__2), .inputs_383__1 (registerOutputs_383__1), .inputs_383__0 (
            registerOutputs_383__0), .inputs_384__15 (registerOutputs_384__15), 
            .inputs_384__14 (registerOutputs_384__14), .inputs_384__13 (
            registerOutputs_384__13), .inputs_384__12 (registerOutputs_384__12)
            , .inputs_384__11 (registerOutputs_384__11), .inputs_384__10 (
            registerOutputs_384__10), .inputs_384__9 (registerOutputs_384__9), .inputs_384__8 (
            registerOutputs_384__8), .inputs_384__7 (registerOutputs_384__7), .inputs_384__6 (
            registerOutputs_384__6), .inputs_384__5 (registerOutputs_384__5), .inputs_384__4 (
            registerOutputs_384__4), .inputs_384__3 (registerOutputs_384__3), .inputs_384__2 (
            registerOutputs_384__2), .inputs_384__1 (registerOutputs_384__1), .inputs_384__0 (
            registerOutputs_384__0), .inputs_385__15 (registerOutputs_385__15), 
            .inputs_385__14 (registerOutputs_385__14), .inputs_385__13 (
            registerOutputs_385__13), .inputs_385__12 (registerOutputs_385__12)
            , .inputs_385__11 (registerOutputs_385__11), .inputs_385__10 (
            registerOutputs_385__10), .inputs_385__9 (registerOutputs_385__9), .inputs_385__8 (
            registerOutputs_385__8), .inputs_385__7 (registerOutputs_385__7), .inputs_385__6 (
            registerOutputs_385__6), .inputs_385__5 (registerOutputs_385__5), .inputs_385__4 (
            registerOutputs_385__4), .inputs_385__3 (registerOutputs_385__3), .inputs_385__2 (
            registerOutputs_385__2), .inputs_385__1 (registerOutputs_385__1), .inputs_385__0 (
            registerOutputs_385__0), .inputs_386__15 (registerOutputs_386__15), 
            .inputs_386__14 (registerOutputs_386__14), .inputs_386__13 (
            registerOutputs_386__13), .inputs_386__12 (registerOutputs_386__12)
            , .inputs_386__11 (registerOutputs_386__11), .inputs_386__10 (
            registerOutputs_386__10), .inputs_386__9 (registerOutputs_386__9), .inputs_386__8 (
            registerOutputs_386__8), .inputs_386__7 (registerOutputs_386__7), .inputs_386__6 (
            registerOutputs_386__6), .inputs_386__5 (registerOutputs_386__5), .inputs_386__4 (
            registerOutputs_386__4), .inputs_386__3 (registerOutputs_386__3), .inputs_386__2 (
            registerOutputs_386__2), .inputs_386__1 (registerOutputs_386__1), .inputs_386__0 (
            registerOutputs_386__0), .inputs_387__15 (registerOutputs_387__15), 
            .inputs_387__14 (registerOutputs_387__14), .inputs_387__13 (
            registerOutputs_387__13), .inputs_387__12 (registerOutputs_387__12)
            , .inputs_387__11 (registerOutputs_387__11), .inputs_387__10 (
            registerOutputs_387__10), .inputs_387__9 (registerOutputs_387__9), .inputs_387__8 (
            registerOutputs_387__8), .inputs_387__7 (registerOutputs_387__7), .inputs_387__6 (
            registerOutputs_387__6), .inputs_387__5 (registerOutputs_387__5), .inputs_387__4 (
            registerOutputs_387__4), .inputs_387__3 (registerOutputs_387__3), .inputs_387__2 (
            registerOutputs_387__2), .inputs_387__1 (registerOutputs_387__1), .inputs_387__0 (
            registerOutputs_387__0), .inputs_388__15 (registerOutputs_388__15), 
            .inputs_388__14 (registerOutputs_388__14), .inputs_388__13 (
            registerOutputs_388__13), .inputs_388__12 (registerOutputs_388__12)
            , .inputs_388__11 (registerOutputs_388__11), .inputs_388__10 (
            registerOutputs_388__10), .inputs_388__9 (registerOutputs_388__9), .inputs_388__8 (
            registerOutputs_388__8), .inputs_388__7 (registerOutputs_388__7), .inputs_388__6 (
            registerOutputs_388__6), .inputs_388__5 (registerOutputs_388__5), .inputs_388__4 (
            registerOutputs_388__4), .inputs_388__3 (registerOutputs_388__3), .inputs_388__2 (
            registerOutputs_388__2), .inputs_388__1 (registerOutputs_388__1), .inputs_388__0 (
            registerOutputs_388__0), .inputs_389__15 (registerOutputs_389__15), 
            .inputs_389__14 (registerOutputs_389__14), .inputs_389__13 (
            registerOutputs_389__13), .inputs_389__12 (registerOutputs_389__12)
            , .inputs_389__11 (registerOutputs_389__11), .inputs_389__10 (
            registerOutputs_389__10), .inputs_389__9 (registerOutputs_389__9), .inputs_389__8 (
            registerOutputs_389__8), .inputs_389__7 (registerOutputs_389__7), .inputs_389__6 (
            registerOutputs_389__6), .inputs_389__5 (registerOutputs_389__5), .inputs_389__4 (
            registerOutputs_389__4), .inputs_389__3 (registerOutputs_389__3), .inputs_389__2 (
            registerOutputs_389__2), .inputs_389__1 (registerOutputs_389__1), .inputs_389__0 (
            registerOutputs_389__0), .inputs_390__15 (registerOutputs_390__15), 
            .inputs_390__14 (registerOutputs_390__14), .inputs_390__13 (
            registerOutputs_390__13), .inputs_390__12 (registerOutputs_390__12)
            , .inputs_390__11 (registerOutputs_390__11), .inputs_390__10 (
            registerOutputs_390__10), .inputs_390__9 (registerOutputs_390__9), .inputs_390__8 (
            registerOutputs_390__8), .inputs_390__7 (registerOutputs_390__7), .inputs_390__6 (
            registerOutputs_390__6), .inputs_390__5 (registerOutputs_390__5), .inputs_390__4 (
            registerOutputs_390__4), .inputs_390__3 (registerOutputs_390__3), .inputs_390__2 (
            registerOutputs_390__2), .inputs_390__1 (registerOutputs_390__1), .inputs_390__0 (
            registerOutputs_390__0), .inputs_391__15 (registerOutputs_391__15), 
            .inputs_391__14 (registerOutputs_391__14), .inputs_391__13 (
            registerOutputs_391__13), .inputs_391__12 (registerOutputs_391__12)
            , .inputs_391__11 (registerOutputs_391__11), .inputs_391__10 (
            registerOutputs_391__10), .inputs_391__9 (registerOutputs_391__9), .inputs_391__8 (
            registerOutputs_391__8), .inputs_391__7 (registerOutputs_391__7), .inputs_391__6 (
            registerOutputs_391__6), .inputs_391__5 (registerOutputs_391__5), .inputs_391__4 (
            registerOutputs_391__4), .inputs_391__3 (registerOutputs_391__3), .inputs_391__2 (
            registerOutputs_391__2), .inputs_391__1 (registerOutputs_391__1), .inputs_391__0 (
            registerOutputs_391__0), .inputs_392__15 (registerOutputs_392__15), 
            .inputs_392__14 (registerOutputs_392__14), .inputs_392__13 (
            registerOutputs_392__13), .inputs_392__12 (registerOutputs_392__12)
            , .inputs_392__11 (registerOutputs_392__11), .inputs_392__10 (
            registerOutputs_392__10), .inputs_392__9 (registerOutputs_392__9), .inputs_392__8 (
            registerOutputs_392__8), .inputs_392__7 (registerOutputs_392__7), .inputs_392__6 (
            registerOutputs_392__6), .inputs_392__5 (registerOutputs_392__5), .inputs_392__4 (
            registerOutputs_392__4), .inputs_392__3 (registerOutputs_392__3), .inputs_392__2 (
            registerOutputs_392__2), .inputs_392__1 (registerOutputs_392__1), .inputs_392__0 (
            registerOutputs_392__0), .inputs_393__15 (registerOutputs_393__15), 
            .inputs_393__14 (registerOutputs_393__14), .inputs_393__13 (
            registerOutputs_393__13), .inputs_393__12 (registerOutputs_393__12)
            , .inputs_393__11 (registerOutputs_393__11), .inputs_393__10 (
            registerOutputs_393__10), .inputs_393__9 (registerOutputs_393__9), .inputs_393__8 (
            registerOutputs_393__8), .inputs_393__7 (registerOutputs_393__7), .inputs_393__6 (
            registerOutputs_393__6), .inputs_393__5 (registerOutputs_393__5), .inputs_393__4 (
            registerOutputs_393__4), .inputs_393__3 (registerOutputs_393__3), .inputs_393__2 (
            registerOutputs_393__2), .inputs_393__1 (registerOutputs_393__1), .inputs_393__0 (
            registerOutputs_393__0), .inputs_394__15 (registerOutputs_394__15), 
            .inputs_394__14 (registerOutputs_394__14), .inputs_394__13 (
            registerOutputs_394__13), .inputs_394__12 (registerOutputs_394__12)
            , .inputs_394__11 (registerOutputs_394__11), .inputs_394__10 (
            registerOutputs_394__10), .inputs_394__9 (registerOutputs_394__9), .inputs_394__8 (
            registerOutputs_394__8), .inputs_394__7 (registerOutputs_394__7), .inputs_394__6 (
            registerOutputs_394__6), .inputs_394__5 (registerOutputs_394__5), .inputs_394__4 (
            registerOutputs_394__4), .inputs_394__3 (registerOutputs_394__3), .inputs_394__2 (
            registerOutputs_394__2), .inputs_394__1 (registerOutputs_394__1), .inputs_394__0 (
            registerOutputs_394__0), .inputs_395__15 (registerOutputs_395__15), 
            .inputs_395__14 (registerOutputs_395__14), .inputs_395__13 (
            registerOutputs_395__13), .inputs_395__12 (registerOutputs_395__12)
            , .inputs_395__11 (registerOutputs_395__11), .inputs_395__10 (
            registerOutputs_395__10), .inputs_395__9 (registerOutputs_395__9), .inputs_395__8 (
            registerOutputs_395__8), .inputs_395__7 (registerOutputs_395__7), .inputs_395__6 (
            registerOutputs_395__6), .inputs_395__5 (registerOutputs_395__5), .inputs_395__4 (
            registerOutputs_395__4), .inputs_395__3 (registerOutputs_395__3), .inputs_395__2 (
            registerOutputs_395__2), .inputs_395__1 (registerOutputs_395__1), .inputs_395__0 (
            registerOutputs_395__0), .inputs_396__15 (registerOutputs_396__15), 
            .inputs_396__14 (registerOutputs_396__14), .inputs_396__13 (
            registerOutputs_396__13), .inputs_396__12 (registerOutputs_396__12)
            , .inputs_396__11 (registerOutputs_396__11), .inputs_396__10 (
            registerOutputs_396__10), .inputs_396__9 (registerOutputs_396__9), .inputs_396__8 (
            registerOutputs_396__8), .inputs_396__7 (registerOutputs_396__7), .inputs_396__6 (
            registerOutputs_396__6), .inputs_396__5 (registerOutputs_396__5), .inputs_396__4 (
            registerOutputs_396__4), .inputs_396__3 (registerOutputs_396__3), .inputs_396__2 (
            registerOutputs_396__2), .inputs_396__1 (registerOutputs_396__1), .inputs_396__0 (
            registerOutputs_396__0), .inputs_397__15 (registerOutputs_397__15), 
            .inputs_397__14 (registerOutputs_397__14), .inputs_397__13 (
            registerOutputs_397__13), .inputs_397__12 (registerOutputs_397__12)
            , .inputs_397__11 (registerOutputs_397__11), .inputs_397__10 (
            registerOutputs_397__10), .inputs_397__9 (registerOutputs_397__9), .inputs_397__8 (
            registerOutputs_397__8), .inputs_397__7 (registerOutputs_397__7), .inputs_397__6 (
            registerOutputs_397__6), .inputs_397__5 (registerOutputs_397__5), .inputs_397__4 (
            registerOutputs_397__4), .inputs_397__3 (registerOutputs_397__3), .inputs_397__2 (
            registerOutputs_397__2), .inputs_397__1 (registerOutputs_397__1), .inputs_397__0 (
            registerOutputs_397__0), .inputs_398__15 (registerOutputs_398__15), 
            .inputs_398__14 (registerOutputs_398__14), .inputs_398__13 (
            registerOutputs_398__13), .inputs_398__12 (registerOutputs_398__12)
            , .inputs_398__11 (registerOutputs_398__11), .inputs_398__10 (
            registerOutputs_398__10), .inputs_398__9 (registerOutputs_398__9), .inputs_398__8 (
            registerOutputs_398__8), .inputs_398__7 (registerOutputs_398__7), .inputs_398__6 (
            registerOutputs_398__6), .inputs_398__5 (registerOutputs_398__5), .inputs_398__4 (
            registerOutputs_398__4), .inputs_398__3 (registerOutputs_398__3), .inputs_398__2 (
            registerOutputs_398__2), .inputs_398__1 (registerOutputs_398__1), .inputs_398__0 (
            registerOutputs_398__0), .inputs_399__15 (registerOutputs_399__15), 
            .inputs_399__14 (registerOutputs_399__14), .inputs_399__13 (
            registerOutputs_399__13), .inputs_399__12 (registerOutputs_399__12)
            , .inputs_399__11 (registerOutputs_399__11), .inputs_399__10 (
            registerOutputs_399__10), .inputs_399__9 (registerOutputs_399__9), .inputs_399__8 (
            registerOutputs_399__8), .inputs_399__7 (registerOutputs_399__7), .inputs_399__6 (
            registerOutputs_399__6), .inputs_399__5 (registerOutputs_399__5), .inputs_399__4 (
            registerOutputs_399__4), .inputs_399__3 (registerOutputs_399__3), .inputs_399__2 (
            registerOutputs_399__2), .inputs_399__1 (registerOutputs_399__1), .inputs_399__0 (
            registerOutputs_399__0), .inputs_400__15 (registerOutputs_400__15), 
            .inputs_400__14 (registerOutputs_400__14), .inputs_400__13 (
            registerOutputs_400__13), .inputs_400__12 (registerOutputs_400__12)
            , .inputs_400__11 (registerOutputs_400__11), .inputs_400__10 (
            registerOutputs_400__10), .inputs_400__9 (registerOutputs_400__9), .inputs_400__8 (
            registerOutputs_400__8), .inputs_400__7 (registerOutputs_400__7), .inputs_400__6 (
            registerOutputs_400__6), .inputs_400__5 (registerOutputs_400__5), .inputs_400__4 (
            registerOutputs_400__4), .inputs_400__3 (registerOutputs_400__3), .inputs_400__2 (
            registerOutputs_400__2), .inputs_400__1 (registerOutputs_400__1), .inputs_400__0 (
            registerOutputs_400__0), .inputs_401__15 (registerOutputs_401__15), 
            .inputs_401__14 (registerOutputs_401__14), .inputs_401__13 (
            registerOutputs_401__13), .inputs_401__12 (registerOutputs_401__12)
            , .inputs_401__11 (registerOutputs_401__11), .inputs_401__10 (
            registerOutputs_401__10), .inputs_401__9 (registerOutputs_401__9), .inputs_401__8 (
            registerOutputs_401__8), .inputs_401__7 (registerOutputs_401__7), .inputs_401__6 (
            registerOutputs_401__6), .inputs_401__5 (registerOutputs_401__5), .inputs_401__4 (
            registerOutputs_401__4), .inputs_401__3 (registerOutputs_401__3), .inputs_401__2 (
            registerOutputs_401__2), .inputs_401__1 (registerOutputs_401__1), .inputs_401__0 (
            registerOutputs_401__0), .inputs_402__15 (registerOutputs_402__15), 
            .inputs_402__14 (registerOutputs_402__14), .inputs_402__13 (
            registerOutputs_402__13), .inputs_402__12 (registerOutputs_402__12)
            , .inputs_402__11 (registerOutputs_402__11), .inputs_402__10 (
            registerOutputs_402__10), .inputs_402__9 (registerOutputs_402__9), .inputs_402__8 (
            registerOutputs_402__8), .inputs_402__7 (registerOutputs_402__7), .inputs_402__6 (
            registerOutputs_402__6), .inputs_402__5 (registerOutputs_402__5), .inputs_402__4 (
            registerOutputs_402__4), .inputs_402__3 (registerOutputs_402__3), .inputs_402__2 (
            registerOutputs_402__2), .inputs_402__1 (registerOutputs_402__1), .inputs_402__0 (
            registerOutputs_402__0), .inputs_403__15 (registerOutputs_403__15), 
            .inputs_403__14 (registerOutputs_403__14), .inputs_403__13 (
            registerOutputs_403__13), .inputs_403__12 (registerOutputs_403__12)
            , .inputs_403__11 (registerOutputs_403__11), .inputs_403__10 (
            registerOutputs_403__10), .inputs_403__9 (registerOutputs_403__9), .inputs_403__8 (
            registerOutputs_403__8), .inputs_403__7 (registerOutputs_403__7), .inputs_403__6 (
            registerOutputs_403__6), .inputs_403__5 (registerOutputs_403__5), .inputs_403__4 (
            registerOutputs_403__4), .inputs_403__3 (registerOutputs_403__3), .inputs_403__2 (
            registerOutputs_403__2), .inputs_403__1 (registerOutputs_403__1), .inputs_403__0 (
            registerOutputs_403__0), .inputs_404__15 (registerOutputs_404__15), 
            .inputs_404__14 (registerOutputs_404__14), .inputs_404__13 (
            registerOutputs_404__13), .inputs_404__12 (registerOutputs_404__12)
            , .inputs_404__11 (registerOutputs_404__11), .inputs_404__10 (
            registerOutputs_404__10), .inputs_404__9 (registerOutputs_404__9), .inputs_404__8 (
            registerOutputs_404__8), .inputs_404__7 (registerOutputs_404__7), .inputs_404__6 (
            registerOutputs_404__6), .inputs_404__5 (registerOutputs_404__5), .inputs_404__4 (
            registerOutputs_404__4), .inputs_404__3 (registerOutputs_404__3), .inputs_404__2 (
            registerOutputs_404__2), .inputs_404__1 (registerOutputs_404__1), .inputs_404__0 (
            registerOutputs_404__0), .inputs_405__15 (registerOutputs_405__15), 
            .inputs_405__14 (registerOutputs_405__14), .inputs_405__13 (
            registerOutputs_405__13), .inputs_405__12 (registerOutputs_405__12)
            , .inputs_405__11 (registerOutputs_405__11), .inputs_405__10 (
            registerOutputs_405__10), .inputs_405__9 (registerOutputs_405__9), .inputs_405__8 (
            registerOutputs_405__8), .inputs_405__7 (registerOutputs_405__7), .inputs_405__6 (
            registerOutputs_405__6), .inputs_405__5 (registerOutputs_405__5), .inputs_405__4 (
            registerOutputs_405__4), .inputs_405__3 (registerOutputs_405__3), .inputs_405__2 (
            registerOutputs_405__2), .inputs_405__1 (registerOutputs_405__1), .inputs_405__0 (
            registerOutputs_405__0), .inputs_406__15 (registerOutputs_406__15), 
            .inputs_406__14 (registerOutputs_406__14), .inputs_406__13 (
            registerOutputs_406__13), .inputs_406__12 (registerOutputs_406__12)
            , .inputs_406__11 (registerOutputs_406__11), .inputs_406__10 (
            registerOutputs_406__10), .inputs_406__9 (registerOutputs_406__9), .inputs_406__8 (
            registerOutputs_406__8), .inputs_406__7 (registerOutputs_406__7), .inputs_406__6 (
            registerOutputs_406__6), .inputs_406__5 (registerOutputs_406__5), .inputs_406__4 (
            registerOutputs_406__4), .inputs_406__3 (registerOutputs_406__3), .inputs_406__2 (
            registerOutputs_406__2), .inputs_406__1 (registerOutputs_406__1), .inputs_406__0 (
            registerOutputs_406__0), .inputs_407__15 (registerOutputs_407__15), 
            .inputs_407__14 (registerOutputs_407__14), .inputs_407__13 (
            registerOutputs_407__13), .inputs_407__12 (registerOutputs_407__12)
            , .inputs_407__11 (registerOutputs_407__11), .inputs_407__10 (
            registerOutputs_407__10), .inputs_407__9 (registerOutputs_407__9), .inputs_407__8 (
            registerOutputs_407__8), .inputs_407__7 (registerOutputs_407__7), .inputs_407__6 (
            registerOutputs_407__6), .inputs_407__5 (registerOutputs_407__5), .inputs_407__4 (
            registerOutputs_407__4), .inputs_407__3 (registerOutputs_407__3), .inputs_407__2 (
            registerOutputs_407__2), .inputs_407__1 (registerOutputs_407__1), .inputs_407__0 (
            registerOutputs_407__0), .inputs_408__15 (registerOutputs_408__15), 
            .inputs_408__14 (registerOutputs_408__14), .inputs_408__13 (
            registerOutputs_408__13), .inputs_408__12 (registerOutputs_408__12)
            , .inputs_408__11 (registerOutputs_408__11), .inputs_408__10 (
            registerOutputs_408__10), .inputs_408__9 (registerOutputs_408__9), .inputs_408__8 (
            registerOutputs_408__8), .inputs_408__7 (registerOutputs_408__7), .inputs_408__6 (
            registerOutputs_408__6), .inputs_408__5 (registerOutputs_408__5), .inputs_408__4 (
            registerOutputs_408__4), .inputs_408__3 (registerOutputs_408__3), .inputs_408__2 (
            registerOutputs_408__2), .inputs_408__1 (registerOutputs_408__1), .inputs_408__0 (
            registerOutputs_408__0), .inputs_409__15 (registerOutputs_409__15), 
            .inputs_409__14 (registerOutputs_409__14), .inputs_409__13 (
            registerOutputs_409__13), .inputs_409__12 (registerOutputs_409__12)
            , .inputs_409__11 (registerOutputs_409__11), .inputs_409__10 (
            registerOutputs_409__10), .inputs_409__9 (registerOutputs_409__9), .inputs_409__8 (
            registerOutputs_409__8), .inputs_409__7 (registerOutputs_409__7), .inputs_409__6 (
            registerOutputs_409__6), .inputs_409__5 (registerOutputs_409__5), .inputs_409__4 (
            registerOutputs_409__4), .inputs_409__3 (registerOutputs_409__3), .inputs_409__2 (
            registerOutputs_409__2), .inputs_409__1 (registerOutputs_409__1), .inputs_409__0 (
            registerOutputs_409__0), .inputs_410__15 (registerOutputs_410__15), 
            .inputs_410__14 (registerOutputs_410__14), .inputs_410__13 (
            registerOutputs_410__13), .inputs_410__12 (registerOutputs_410__12)
            , .inputs_410__11 (registerOutputs_410__11), .inputs_410__10 (
            registerOutputs_410__10), .inputs_410__9 (registerOutputs_410__9), .inputs_410__8 (
            registerOutputs_410__8), .inputs_410__7 (registerOutputs_410__7), .inputs_410__6 (
            registerOutputs_410__6), .inputs_410__5 (registerOutputs_410__5), .inputs_410__4 (
            registerOutputs_410__4), .inputs_410__3 (registerOutputs_410__3), .inputs_410__2 (
            registerOutputs_410__2), .inputs_410__1 (registerOutputs_410__1), .inputs_410__0 (
            registerOutputs_410__0), .inputs_411__15 (registerOutputs_411__15), 
            .inputs_411__14 (registerOutputs_411__14), .inputs_411__13 (
            registerOutputs_411__13), .inputs_411__12 (registerOutputs_411__12)
            , .inputs_411__11 (registerOutputs_411__11), .inputs_411__10 (
            registerOutputs_411__10), .inputs_411__9 (registerOutputs_411__9), .inputs_411__8 (
            registerOutputs_411__8), .inputs_411__7 (registerOutputs_411__7), .inputs_411__6 (
            registerOutputs_411__6), .inputs_411__5 (registerOutputs_411__5), .inputs_411__4 (
            registerOutputs_411__4), .inputs_411__3 (registerOutputs_411__3), .inputs_411__2 (
            registerOutputs_411__2), .inputs_411__1 (registerOutputs_411__1), .inputs_411__0 (
            registerOutputs_411__0), .inputs_412__15 (registerOutputs_412__15), 
            .inputs_412__14 (registerOutputs_412__14), .inputs_412__13 (
            registerOutputs_412__13), .inputs_412__12 (registerOutputs_412__12)
            , .inputs_412__11 (registerOutputs_412__11), .inputs_412__10 (
            registerOutputs_412__10), .inputs_412__9 (registerOutputs_412__9), .inputs_412__8 (
            registerOutputs_412__8), .inputs_412__7 (registerOutputs_412__7), .inputs_412__6 (
            registerOutputs_412__6), .inputs_412__5 (registerOutputs_412__5), .inputs_412__4 (
            registerOutputs_412__4), .inputs_412__3 (registerOutputs_412__3), .inputs_412__2 (
            registerOutputs_412__2), .inputs_412__1 (registerOutputs_412__1), .inputs_412__0 (
            registerOutputs_412__0), .inputs_413__15 (registerOutputs_413__15), 
            .inputs_413__14 (registerOutputs_413__14), .inputs_413__13 (
            registerOutputs_413__13), .inputs_413__12 (registerOutputs_413__12)
            , .inputs_413__11 (registerOutputs_413__11), .inputs_413__10 (
            registerOutputs_413__10), .inputs_413__9 (registerOutputs_413__9), .inputs_413__8 (
            registerOutputs_413__8), .inputs_413__7 (registerOutputs_413__7), .inputs_413__6 (
            registerOutputs_413__6), .inputs_413__5 (registerOutputs_413__5), .inputs_413__4 (
            registerOutputs_413__4), .inputs_413__3 (registerOutputs_413__3), .inputs_413__2 (
            registerOutputs_413__2), .inputs_413__1 (registerOutputs_413__1), .inputs_413__0 (
            registerOutputs_413__0), .inputs_414__15 (registerOutputs_414__15), 
            .inputs_414__14 (registerOutputs_414__14), .inputs_414__13 (
            registerOutputs_414__13), .inputs_414__12 (registerOutputs_414__12)
            , .inputs_414__11 (registerOutputs_414__11), .inputs_414__10 (
            registerOutputs_414__10), .inputs_414__9 (registerOutputs_414__9), .inputs_414__8 (
            registerOutputs_414__8), .inputs_414__7 (registerOutputs_414__7), .inputs_414__6 (
            registerOutputs_414__6), .inputs_414__5 (registerOutputs_414__5), .inputs_414__4 (
            registerOutputs_414__4), .inputs_414__3 (registerOutputs_414__3), .inputs_414__2 (
            registerOutputs_414__2), .inputs_414__1 (registerOutputs_414__1), .inputs_414__0 (
            registerOutputs_414__0), .inputs_415__15 (registerOutputs_415__15), 
            .inputs_415__14 (registerOutputs_415__14), .inputs_415__13 (
            registerOutputs_415__13), .inputs_415__12 (registerOutputs_415__12)
            , .inputs_415__11 (registerOutputs_415__11), .inputs_415__10 (
            registerOutputs_415__10), .inputs_415__9 (registerOutputs_415__9), .inputs_415__8 (
            registerOutputs_415__8), .inputs_415__7 (registerOutputs_415__7), .inputs_415__6 (
            registerOutputs_415__6), .inputs_415__5 (registerOutputs_415__5), .inputs_415__4 (
            registerOutputs_415__4), .inputs_415__3 (registerOutputs_415__3), .inputs_415__2 (
            registerOutputs_415__2), .inputs_415__1 (registerOutputs_415__1), .inputs_415__0 (
            registerOutputs_415__0), .inputs_416__15 (registerOutputs_416__15), 
            .inputs_416__14 (registerOutputs_416__14), .inputs_416__13 (
            registerOutputs_416__13), .inputs_416__12 (registerOutputs_416__12)
            , .inputs_416__11 (registerOutputs_416__11), .inputs_416__10 (
            registerOutputs_416__10), .inputs_416__9 (registerOutputs_416__9), .inputs_416__8 (
            registerOutputs_416__8), .inputs_416__7 (registerOutputs_416__7), .inputs_416__6 (
            registerOutputs_416__6), .inputs_416__5 (registerOutputs_416__5), .inputs_416__4 (
            registerOutputs_416__4), .inputs_416__3 (registerOutputs_416__3), .inputs_416__2 (
            registerOutputs_416__2), .inputs_416__1 (registerOutputs_416__1), .inputs_416__0 (
            registerOutputs_416__0), .inputs_417__15 (registerOutputs_417__15), 
            .inputs_417__14 (registerOutputs_417__14), .inputs_417__13 (
            registerOutputs_417__13), .inputs_417__12 (registerOutputs_417__12)
            , .inputs_417__11 (registerOutputs_417__11), .inputs_417__10 (
            registerOutputs_417__10), .inputs_417__9 (registerOutputs_417__9), .inputs_417__8 (
            registerOutputs_417__8), .inputs_417__7 (registerOutputs_417__7), .inputs_417__6 (
            registerOutputs_417__6), .inputs_417__5 (registerOutputs_417__5), .inputs_417__4 (
            registerOutputs_417__4), .inputs_417__3 (registerOutputs_417__3), .inputs_417__2 (
            registerOutputs_417__2), .inputs_417__1 (registerOutputs_417__1), .inputs_417__0 (
            registerOutputs_417__0), .inputs_418__15 (registerOutputs_418__15), 
            .inputs_418__14 (registerOutputs_418__14), .inputs_418__13 (
            registerOutputs_418__13), .inputs_418__12 (registerOutputs_418__12)
            , .inputs_418__11 (registerOutputs_418__11), .inputs_418__10 (
            registerOutputs_418__10), .inputs_418__9 (registerOutputs_418__9), .inputs_418__8 (
            registerOutputs_418__8), .inputs_418__7 (registerOutputs_418__7), .inputs_418__6 (
            registerOutputs_418__6), .inputs_418__5 (registerOutputs_418__5), .inputs_418__4 (
            registerOutputs_418__4), .inputs_418__3 (registerOutputs_418__3), .inputs_418__2 (
            registerOutputs_418__2), .inputs_418__1 (registerOutputs_418__1), .inputs_418__0 (
            registerOutputs_418__0), .inputs_419__15 (registerOutputs_419__15), 
            .inputs_419__14 (registerOutputs_419__14), .inputs_419__13 (
            registerOutputs_419__13), .inputs_419__12 (registerOutputs_419__12)
            , .inputs_419__11 (registerOutputs_419__11), .inputs_419__10 (
            registerOutputs_419__10), .inputs_419__9 (registerOutputs_419__9), .inputs_419__8 (
            registerOutputs_419__8), .inputs_419__7 (registerOutputs_419__7), .inputs_419__6 (
            registerOutputs_419__6), .inputs_419__5 (registerOutputs_419__5), .inputs_419__4 (
            registerOutputs_419__4), .inputs_419__3 (registerOutputs_419__3), .inputs_419__2 (
            registerOutputs_419__2), .inputs_419__1 (registerOutputs_419__1), .inputs_419__0 (
            registerOutputs_419__0), .inputs_420__15 (registerOutputs_420__15), 
            .inputs_420__14 (registerOutputs_420__14), .inputs_420__13 (
            registerOutputs_420__13), .inputs_420__12 (registerOutputs_420__12)
            , .inputs_420__11 (registerOutputs_420__11), .inputs_420__10 (
            registerOutputs_420__10), .inputs_420__9 (registerOutputs_420__9), .inputs_420__8 (
            registerOutputs_420__8), .inputs_420__7 (registerOutputs_420__7), .inputs_420__6 (
            registerOutputs_420__6), .inputs_420__5 (registerOutputs_420__5), .inputs_420__4 (
            registerOutputs_420__4), .inputs_420__3 (registerOutputs_420__3), .inputs_420__2 (
            registerOutputs_420__2), .inputs_420__1 (registerOutputs_420__1), .inputs_420__0 (
            registerOutputs_420__0), .inputs_421__15 (registerOutputs_421__15), 
            .inputs_421__14 (registerOutputs_421__14), .inputs_421__13 (
            registerOutputs_421__13), .inputs_421__12 (registerOutputs_421__12)
            , .inputs_421__11 (registerOutputs_421__11), .inputs_421__10 (
            registerOutputs_421__10), .inputs_421__9 (registerOutputs_421__9), .inputs_421__8 (
            registerOutputs_421__8), .inputs_421__7 (registerOutputs_421__7), .inputs_421__6 (
            registerOutputs_421__6), .inputs_421__5 (registerOutputs_421__5), .inputs_421__4 (
            registerOutputs_421__4), .inputs_421__3 (registerOutputs_421__3), .inputs_421__2 (
            registerOutputs_421__2), .inputs_421__1 (registerOutputs_421__1), .inputs_421__0 (
            registerOutputs_421__0), .inputs_422__15 (registerOutputs_422__15), 
            .inputs_422__14 (registerOutputs_422__14), .inputs_422__13 (
            registerOutputs_422__13), .inputs_422__12 (registerOutputs_422__12)
            , .inputs_422__11 (registerOutputs_422__11), .inputs_422__10 (
            registerOutputs_422__10), .inputs_422__9 (registerOutputs_422__9), .inputs_422__8 (
            registerOutputs_422__8), .inputs_422__7 (registerOutputs_422__7), .inputs_422__6 (
            registerOutputs_422__6), .inputs_422__5 (registerOutputs_422__5), .inputs_422__4 (
            registerOutputs_422__4), .inputs_422__3 (registerOutputs_422__3), .inputs_422__2 (
            registerOutputs_422__2), .inputs_422__1 (registerOutputs_422__1), .inputs_422__0 (
            registerOutputs_422__0), .inputs_423__15 (registerOutputs_423__15), 
            .inputs_423__14 (registerOutputs_423__14), .inputs_423__13 (
            registerOutputs_423__13), .inputs_423__12 (registerOutputs_423__12)
            , .inputs_423__11 (registerOutputs_423__11), .inputs_423__10 (
            registerOutputs_423__10), .inputs_423__9 (registerOutputs_423__9), .inputs_423__8 (
            registerOutputs_423__8), .inputs_423__7 (registerOutputs_423__7), .inputs_423__6 (
            registerOutputs_423__6), .inputs_423__5 (registerOutputs_423__5), .inputs_423__4 (
            registerOutputs_423__4), .inputs_423__3 (registerOutputs_423__3), .inputs_423__2 (
            registerOutputs_423__2), .inputs_423__1 (registerOutputs_423__1), .inputs_423__0 (
            registerOutputs_423__0), .inputs_424__15 (registerOutputs_424__15), 
            .inputs_424__14 (registerOutputs_424__14), .inputs_424__13 (
            registerOutputs_424__13), .inputs_424__12 (registerOutputs_424__12)
            , .inputs_424__11 (registerOutputs_424__11), .inputs_424__10 (
            registerOutputs_424__10), .inputs_424__9 (registerOutputs_424__9), .inputs_424__8 (
            registerOutputs_424__8), .inputs_424__7 (registerOutputs_424__7), .inputs_424__6 (
            registerOutputs_424__6), .inputs_424__5 (registerOutputs_424__5), .inputs_424__4 (
            registerOutputs_424__4), .inputs_424__3 (registerOutputs_424__3), .inputs_424__2 (
            registerOutputs_424__2), .inputs_424__1 (registerOutputs_424__1), .inputs_424__0 (
            registerOutputs_424__0), .inputs_425__15 (registerOutputs_425__15), 
            .inputs_425__14 (registerOutputs_425__14), .inputs_425__13 (
            registerOutputs_425__13), .inputs_425__12 (registerOutputs_425__12)
            , .inputs_425__11 (registerOutputs_425__11), .inputs_425__10 (
            registerOutputs_425__10), .inputs_425__9 (registerOutputs_425__9), .inputs_425__8 (
            registerOutputs_425__8), .inputs_425__7 (registerOutputs_425__7), .inputs_425__6 (
            registerOutputs_425__6), .inputs_425__5 (registerOutputs_425__5), .inputs_425__4 (
            registerOutputs_425__4), .inputs_425__3 (registerOutputs_425__3), .inputs_425__2 (
            registerOutputs_425__2), .inputs_425__1 (registerOutputs_425__1), .inputs_425__0 (
            registerOutputs_425__0), .inputs_426__15 (registerOutputs_426__15), 
            .inputs_426__14 (registerOutputs_426__14), .inputs_426__13 (
            registerOutputs_426__13), .inputs_426__12 (registerOutputs_426__12)
            , .inputs_426__11 (registerOutputs_426__11), .inputs_426__10 (
            registerOutputs_426__10), .inputs_426__9 (registerOutputs_426__9), .inputs_426__8 (
            registerOutputs_426__8), .inputs_426__7 (registerOutputs_426__7), .inputs_426__6 (
            registerOutputs_426__6), .inputs_426__5 (registerOutputs_426__5), .inputs_426__4 (
            registerOutputs_426__4), .inputs_426__3 (registerOutputs_426__3), .inputs_426__2 (
            registerOutputs_426__2), .inputs_426__1 (registerOutputs_426__1), .inputs_426__0 (
            registerOutputs_426__0), .inputs_427__15 (registerOutputs_427__15), 
            .inputs_427__14 (registerOutputs_427__14), .inputs_427__13 (
            registerOutputs_427__13), .inputs_427__12 (registerOutputs_427__12)
            , .inputs_427__11 (registerOutputs_427__11), .inputs_427__10 (
            registerOutputs_427__10), .inputs_427__9 (registerOutputs_427__9), .inputs_427__8 (
            registerOutputs_427__8), .inputs_427__7 (registerOutputs_427__7), .inputs_427__6 (
            registerOutputs_427__6), .inputs_427__5 (registerOutputs_427__5), .inputs_427__4 (
            registerOutputs_427__4), .inputs_427__3 (registerOutputs_427__3), .inputs_427__2 (
            registerOutputs_427__2), .inputs_427__1 (registerOutputs_427__1), .inputs_427__0 (
            registerOutputs_427__0), .inputs_428__15 (registerOutputs_428__15), 
            .inputs_428__14 (registerOutputs_428__14), .inputs_428__13 (
            registerOutputs_428__13), .inputs_428__12 (registerOutputs_428__12)
            , .inputs_428__11 (registerOutputs_428__11), .inputs_428__10 (
            registerOutputs_428__10), .inputs_428__9 (registerOutputs_428__9), .inputs_428__8 (
            registerOutputs_428__8), .inputs_428__7 (registerOutputs_428__7), .inputs_428__6 (
            registerOutputs_428__6), .inputs_428__5 (registerOutputs_428__5), .inputs_428__4 (
            registerOutputs_428__4), .inputs_428__3 (registerOutputs_428__3), .inputs_428__2 (
            registerOutputs_428__2), .inputs_428__1 (registerOutputs_428__1), .inputs_428__0 (
            registerOutputs_428__0), .inputs_429__15 (registerOutputs_429__15), 
            .inputs_429__14 (registerOutputs_429__14), .inputs_429__13 (
            registerOutputs_429__13), .inputs_429__12 (registerOutputs_429__12)
            , .inputs_429__11 (registerOutputs_429__11), .inputs_429__10 (
            registerOutputs_429__10), .inputs_429__9 (registerOutputs_429__9), .inputs_429__8 (
            registerOutputs_429__8), .inputs_429__7 (registerOutputs_429__7), .inputs_429__6 (
            registerOutputs_429__6), .inputs_429__5 (registerOutputs_429__5), .inputs_429__4 (
            registerOutputs_429__4), .inputs_429__3 (registerOutputs_429__3), .inputs_429__2 (
            registerOutputs_429__2), .inputs_429__1 (registerOutputs_429__1), .inputs_429__0 (
            registerOutputs_429__0), .inputs_430__15 (registerOutputs_430__15), 
            .inputs_430__14 (registerOutputs_430__14), .inputs_430__13 (
            registerOutputs_430__13), .inputs_430__12 (registerOutputs_430__12)
            , .inputs_430__11 (registerOutputs_430__11), .inputs_430__10 (
            registerOutputs_430__10), .inputs_430__9 (registerOutputs_430__9), .inputs_430__8 (
            registerOutputs_430__8), .inputs_430__7 (registerOutputs_430__7), .inputs_430__6 (
            registerOutputs_430__6), .inputs_430__5 (registerOutputs_430__5), .inputs_430__4 (
            registerOutputs_430__4), .inputs_430__3 (registerOutputs_430__3), .inputs_430__2 (
            registerOutputs_430__2), .inputs_430__1 (registerOutputs_430__1), .inputs_430__0 (
            registerOutputs_430__0), .inputs_431__15 (registerOutputs_431__15), 
            .inputs_431__14 (registerOutputs_431__14), .inputs_431__13 (
            registerOutputs_431__13), .inputs_431__12 (registerOutputs_431__12)
            , .inputs_431__11 (registerOutputs_431__11), .inputs_431__10 (
            registerOutputs_431__10), .inputs_431__9 (registerOutputs_431__9), .inputs_431__8 (
            registerOutputs_431__8), .inputs_431__7 (registerOutputs_431__7), .inputs_431__6 (
            registerOutputs_431__6), .inputs_431__5 (registerOutputs_431__5), .inputs_431__4 (
            registerOutputs_431__4), .inputs_431__3 (registerOutputs_431__3), .inputs_431__2 (
            registerOutputs_431__2), .inputs_431__1 (registerOutputs_431__1), .inputs_431__0 (
            registerOutputs_431__0), .inputs_432__15 (registerOutputs_432__15), 
            .inputs_432__14 (registerOutputs_432__14), .inputs_432__13 (
            registerOutputs_432__13), .inputs_432__12 (registerOutputs_432__12)
            , .inputs_432__11 (registerOutputs_432__11), .inputs_432__10 (
            registerOutputs_432__10), .inputs_432__9 (registerOutputs_432__9), .inputs_432__8 (
            registerOutputs_432__8), .inputs_432__7 (registerOutputs_432__7), .inputs_432__6 (
            registerOutputs_432__6), .inputs_432__5 (registerOutputs_432__5), .inputs_432__4 (
            registerOutputs_432__4), .inputs_432__3 (registerOutputs_432__3), .inputs_432__2 (
            registerOutputs_432__2), .inputs_432__1 (registerOutputs_432__1), .inputs_432__0 (
            registerOutputs_432__0), .inputs_433__15 (registerOutputs_433__15), 
            .inputs_433__14 (registerOutputs_433__14), .inputs_433__13 (
            registerOutputs_433__13), .inputs_433__12 (registerOutputs_433__12)
            , .inputs_433__11 (registerOutputs_433__11), .inputs_433__10 (
            registerOutputs_433__10), .inputs_433__9 (registerOutputs_433__9), .inputs_433__8 (
            registerOutputs_433__8), .inputs_433__7 (registerOutputs_433__7), .inputs_433__6 (
            registerOutputs_433__6), .inputs_433__5 (registerOutputs_433__5), .inputs_433__4 (
            registerOutputs_433__4), .inputs_433__3 (registerOutputs_433__3), .inputs_433__2 (
            registerOutputs_433__2), .inputs_433__1 (registerOutputs_433__1), .inputs_433__0 (
            registerOutputs_433__0), .inputs_434__15 (registerOutputs_434__15), 
            .inputs_434__14 (registerOutputs_434__14), .inputs_434__13 (
            registerOutputs_434__13), .inputs_434__12 (registerOutputs_434__12)
            , .inputs_434__11 (registerOutputs_434__11), .inputs_434__10 (
            registerOutputs_434__10), .inputs_434__9 (registerOutputs_434__9), .inputs_434__8 (
            registerOutputs_434__8), .inputs_434__7 (registerOutputs_434__7), .inputs_434__6 (
            registerOutputs_434__6), .inputs_434__5 (registerOutputs_434__5), .inputs_434__4 (
            registerOutputs_434__4), .inputs_434__3 (registerOutputs_434__3), .inputs_434__2 (
            registerOutputs_434__2), .inputs_434__1 (registerOutputs_434__1), .inputs_434__0 (
            registerOutputs_434__0), .inputs_435__15 (registerOutputs_435__15), 
            .inputs_435__14 (registerOutputs_435__14), .inputs_435__13 (
            registerOutputs_435__13), .inputs_435__12 (registerOutputs_435__12)
            , .inputs_435__11 (registerOutputs_435__11), .inputs_435__10 (
            registerOutputs_435__10), .inputs_435__9 (registerOutputs_435__9), .inputs_435__8 (
            registerOutputs_435__8), .inputs_435__7 (registerOutputs_435__7), .inputs_435__6 (
            registerOutputs_435__6), .inputs_435__5 (registerOutputs_435__5), .inputs_435__4 (
            registerOutputs_435__4), .inputs_435__3 (registerOutputs_435__3), .inputs_435__2 (
            registerOutputs_435__2), .inputs_435__1 (registerOutputs_435__1), .inputs_435__0 (
            registerOutputs_435__0), .inputs_436__15 (registerOutputs_436__15), 
            .inputs_436__14 (registerOutputs_436__14), .inputs_436__13 (
            registerOutputs_436__13), .inputs_436__12 (registerOutputs_436__12)
            , .inputs_436__11 (registerOutputs_436__11), .inputs_436__10 (
            registerOutputs_436__10), .inputs_436__9 (registerOutputs_436__9), .inputs_436__8 (
            registerOutputs_436__8), .inputs_436__7 (registerOutputs_436__7), .inputs_436__6 (
            registerOutputs_436__6), .inputs_436__5 (registerOutputs_436__5), .inputs_436__4 (
            registerOutputs_436__4), .inputs_436__3 (registerOutputs_436__3), .inputs_436__2 (
            registerOutputs_436__2), .inputs_436__1 (registerOutputs_436__1), .inputs_436__0 (
            registerOutputs_436__0), .inputs_437__15 (registerOutputs_437__15), 
            .inputs_437__14 (registerOutputs_437__14), .inputs_437__13 (
            registerOutputs_437__13), .inputs_437__12 (registerOutputs_437__12)
            , .inputs_437__11 (registerOutputs_437__11), .inputs_437__10 (
            registerOutputs_437__10), .inputs_437__9 (registerOutputs_437__9), .inputs_437__8 (
            registerOutputs_437__8), .inputs_437__7 (registerOutputs_437__7), .inputs_437__6 (
            registerOutputs_437__6), .inputs_437__5 (registerOutputs_437__5), .inputs_437__4 (
            registerOutputs_437__4), .inputs_437__3 (registerOutputs_437__3), .inputs_437__2 (
            registerOutputs_437__2), .inputs_437__1 (registerOutputs_437__1), .inputs_437__0 (
            registerOutputs_437__0), .inputs_438__15 (registerOutputs_438__15), 
            .inputs_438__14 (registerOutputs_438__14), .inputs_438__13 (
            registerOutputs_438__13), .inputs_438__12 (registerOutputs_438__12)
            , .inputs_438__11 (registerOutputs_438__11), .inputs_438__10 (
            registerOutputs_438__10), .inputs_438__9 (registerOutputs_438__9), .inputs_438__8 (
            registerOutputs_438__8), .inputs_438__7 (registerOutputs_438__7), .inputs_438__6 (
            registerOutputs_438__6), .inputs_438__5 (registerOutputs_438__5), .inputs_438__4 (
            registerOutputs_438__4), .inputs_438__3 (registerOutputs_438__3), .inputs_438__2 (
            registerOutputs_438__2), .inputs_438__1 (registerOutputs_438__1), .inputs_438__0 (
            registerOutputs_438__0), .inputs_439__15 (registerOutputs_439__15), 
            .inputs_439__14 (registerOutputs_439__14), .inputs_439__13 (
            registerOutputs_439__13), .inputs_439__12 (registerOutputs_439__12)
            , .inputs_439__11 (registerOutputs_439__11), .inputs_439__10 (
            registerOutputs_439__10), .inputs_439__9 (registerOutputs_439__9), .inputs_439__8 (
            registerOutputs_439__8), .inputs_439__7 (registerOutputs_439__7), .inputs_439__6 (
            registerOutputs_439__6), .inputs_439__5 (registerOutputs_439__5), .inputs_439__4 (
            registerOutputs_439__4), .inputs_439__3 (registerOutputs_439__3), .inputs_439__2 (
            registerOutputs_439__2), .inputs_439__1 (registerOutputs_439__1), .inputs_439__0 (
            registerOutputs_439__0), .inputs_440__15 (registerOutputs_440__15), 
            .inputs_440__14 (registerOutputs_440__14), .inputs_440__13 (
            registerOutputs_440__13), .inputs_440__12 (registerOutputs_440__12)
            , .inputs_440__11 (registerOutputs_440__11), .inputs_440__10 (
            registerOutputs_440__10), .inputs_440__9 (registerOutputs_440__9), .inputs_440__8 (
            registerOutputs_440__8), .inputs_440__7 (registerOutputs_440__7), .inputs_440__6 (
            registerOutputs_440__6), .inputs_440__5 (registerOutputs_440__5), .inputs_440__4 (
            registerOutputs_440__4), .inputs_440__3 (registerOutputs_440__3), .inputs_440__2 (
            registerOutputs_440__2), .inputs_440__1 (registerOutputs_440__1), .inputs_440__0 (
            registerOutputs_440__0), .inputs_441__15 (registerOutputs_441__15), 
            .inputs_441__14 (registerOutputs_441__14), .inputs_441__13 (
            registerOutputs_441__13), .inputs_441__12 (registerOutputs_441__12)
            , .inputs_441__11 (registerOutputs_441__11), .inputs_441__10 (
            registerOutputs_441__10), .inputs_441__9 (registerOutputs_441__9), .inputs_441__8 (
            registerOutputs_441__8), .inputs_441__7 (registerOutputs_441__7), .inputs_441__6 (
            registerOutputs_441__6), .inputs_441__5 (registerOutputs_441__5), .inputs_441__4 (
            registerOutputs_441__4), .inputs_441__3 (registerOutputs_441__3), .inputs_441__2 (
            registerOutputs_441__2), .inputs_441__1 (registerOutputs_441__1), .inputs_441__0 (
            registerOutputs_441__0), .inputs_442__15 (registerOutputs_442__15), 
            .inputs_442__14 (registerOutputs_442__14), .inputs_442__13 (
            registerOutputs_442__13), .inputs_442__12 (registerOutputs_442__12)
            , .inputs_442__11 (registerOutputs_442__11), .inputs_442__10 (
            registerOutputs_442__10), .inputs_442__9 (registerOutputs_442__9), .inputs_442__8 (
            registerOutputs_442__8), .inputs_442__7 (registerOutputs_442__7), .inputs_442__6 (
            registerOutputs_442__6), .inputs_442__5 (registerOutputs_442__5), .inputs_442__4 (
            registerOutputs_442__4), .inputs_442__3 (registerOutputs_442__3), .inputs_442__2 (
            registerOutputs_442__2), .inputs_442__1 (registerOutputs_442__1), .inputs_442__0 (
            registerOutputs_442__0), .inputs_443__15 (registerOutputs_443__15), 
            .inputs_443__14 (registerOutputs_443__14), .inputs_443__13 (
            registerOutputs_443__13), .inputs_443__12 (registerOutputs_443__12)
            , .inputs_443__11 (registerOutputs_443__11), .inputs_443__10 (
            registerOutputs_443__10), .inputs_443__9 (registerOutputs_443__9), .inputs_443__8 (
            registerOutputs_443__8), .inputs_443__7 (registerOutputs_443__7), .inputs_443__6 (
            registerOutputs_443__6), .inputs_443__5 (registerOutputs_443__5), .inputs_443__4 (
            registerOutputs_443__4), .inputs_443__3 (registerOutputs_443__3), .inputs_443__2 (
            registerOutputs_443__2), .inputs_443__1 (registerOutputs_443__1), .inputs_443__0 (
            registerOutputs_443__0), .inputs_444__15 (registerOutputs_444__15), 
            .inputs_444__14 (registerOutputs_444__14), .inputs_444__13 (
            registerOutputs_444__13), .inputs_444__12 (registerOutputs_444__12)
            , .inputs_444__11 (registerOutputs_444__11), .inputs_444__10 (
            registerOutputs_444__10), .inputs_444__9 (registerOutputs_444__9), .inputs_444__8 (
            registerOutputs_444__8), .inputs_444__7 (registerOutputs_444__7), .inputs_444__6 (
            registerOutputs_444__6), .inputs_444__5 (registerOutputs_444__5), .inputs_444__4 (
            registerOutputs_444__4), .inputs_444__3 (registerOutputs_444__3), .inputs_444__2 (
            registerOutputs_444__2), .inputs_444__1 (registerOutputs_444__1), .inputs_444__0 (
            registerOutputs_444__0), .inputs_445__15 (registerOutputs_445__15), 
            .inputs_445__14 (registerOutputs_445__14), .inputs_445__13 (
            registerOutputs_445__13), .inputs_445__12 (registerOutputs_445__12)
            , .inputs_445__11 (registerOutputs_445__11), .inputs_445__10 (
            registerOutputs_445__10), .inputs_445__9 (registerOutputs_445__9), .inputs_445__8 (
            registerOutputs_445__8), .inputs_445__7 (registerOutputs_445__7), .inputs_445__6 (
            registerOutputs_445__6), .inputs_445__5 (registerOutputs_445__5), .inputs_445__4 (
            registerOutputs_445__4), .inputs_445__3 (registerOutputs_445__3), .inputs_445__2 (
            registerOutputs_445__2), .inputs_445__1 (registerOutputs_445__1), .inputs_445__0 (
            registerOutputs_445__0), .inputs_446__15 (registerOutputs_446__15), 
            .inputs_446__14 (registerOutputs_446__14), .inputs_446__13 (
            registerOutputs_446__13), .inputs_446__12 (registerOutputs_446__12)
            , .inputs_446__11 (registerOutputs_446__11), .inputs_446__10 (
            registerOutputs_446__10), .inputs_446__9 (registerOutputs_446__9), .inputs_446__8 (
            registerOutputs_446__8), .inputs_446__7 (registerOutputs_446__7), .inputs_446__6 (
            registerOutputs_446__6), .inputs_446__5 (registerOutputs_446__5), .inputs_446__4 (
            registerOutputs_446__4), .inputs_446__3 (registerOutputs_446__3), .inputs_446__2 (
            registerOutputs_446__2), .inputs_446__1 (registerOutputs_446__1), .inputs_446__0 (
            registerOutputs_446__0), .inputs_447__15 (registerOutputs_447__15), 
            .inputs_447__14 (registerOutputs_447__14), .inputs_447__13 (
            registerOutputs_447__13), .inputs_447__12 (registerOutputs_447__12)
            , .inputs_447__11 (registerOutputs_447__11), .inputs_447__10 (
            registerOutputs_447__10), .inputs_447__9 (registerOutputs_447__9), .inputs_447__8 (
            registerOutputs_447__8), .inputs_447__7 (registerOutputs_447__7), .inputs_447__6 (
            registerOutputs_447__6), .inputs_447__5 (registerOutputs_447__5), .inputs_447__4 (
            registerOutputs_447__4), .inputs_447__3 (registerOutputs_447__3), .inputs_447__2 (
            registerOutputs_447__2), .inputs_447__1 (registerOutputs_447__1), .inputs_447__0 (
            registerOutputs_447__0), .inputs_448__15 (registerOutputs_448__15), 
            .inputs_448__14 (registerOutputs_448__14), .inputs_448__13 (
            registerOutputs_448__13), .inputs_448__12 (registerOutputs_448__12)
            , .inputs_448__11 (registerOutputs_448__11), .inputs_448__10 (
            registerOutputs_448__10), .inputs_448__9 (registerOutputs_448__9), .inputs_448__8 (
            registerOutputs_448__8), .inputs_448__7 (registerOutputs_448__7), .inputs_448__6 (
            registerOutputs_448__6), .inputs_448__5 (registerOutputs_448__5), .inputs_448__4 (
            registerOutputs_448__4), .inputs_448__3 (registerOutputs_448__3), .inputs_448__2 (
            registerOutputs_448__2), .inputs_448__1 (registerOutputs_448__1), .inputs_448__0 (
            registerOutputs_448__0), .inputs_449__15 (registerOutputs_449__15), 
            .inputs_449__14 (registerOutputs_449__14), .inputs_449__13 (
            registerOutputs_449__13), .inputs_449__12 (registerOutputs_449__12)
            , .inputs_449__11 (registerOutputs_449__11), .inputs_449__10 (
            registerOutputs_449__10), .inputs_449__9 (registerOutputs_449__9), .inputs_449__8 (
            registerOutputs_449__8), .inputs_449__7 (registerOutputs_449__7), .inputs_449__6 (
            registerOutputs_449__6), .inputs_449__5 (registerOutputs_449__5), .inputs_449__4 (
            registerOutputs_449__4), .inputs_449__3 (registerOutputs_449__3), .inputs_449__2 (
            registerOutputs_449__2), .inputs_449__1 (registerOutputs_449__1), .inputs_449__0 (
            registerOutputs_449__0), .inputs_450__15 (registerOutputs_450__15), 
            .inputs_450__14 (registerOutputs_450__14), .inputs_450__13 (
            registerOutputs_450__13), .inputs_450__12 (registerOutputs_450__12)
            , .inputs_450__11 (registerOutputs_450__11), .inputs_450__10 (
            registerOutputs_450__10), .inputs_450__9 (registerOutputs_450__9), .inputs_450__8 (
            registerOutputs_450__8), .inputs_450__7 (registerOutputs_450__7), .inputs_450__6 (
            registerOutputs_450__6), .inputs_450__5 (registerOutputs_450__5), .inputs_450__4 (
            registerOutputs_450__4), .inputs_450__3 (registerOutputs_450__3), .inputs_450__2 (
            registerOutputs_450__2), .inputs_450__1 (registerOutputs_450__1), .inputs_450__0 (
            registerOutputs_450__0), .inputs_451__15 (registerOutputs_451__15), 
            .inputs_451__14 (registerOutputs_451__14), .inputs_451__13 (
            registerOutputs_451__13), .inputs_451__12 (registerOutputs_451__12)
            , .inputs_451__11 (registerOutputs_451__11), .inputs_451__10 (
            registerOutputs_451__10), .inputs_451__9 (registerOutputs_451__9), .inputs_451__8 (
            registerOutputs_451__8), .inputs_451__7 (registerOutputs_451__7), .inputs_451__6 (
            registerOutputs_451__6), .inputs_451__5 (registerOutputs_451__5), .inputs_451__4 (
            registerOutputs_451__4), .inputs_451__3 (registerOutputs_451__3), .inputs_451__2 (
            registerOutputs_451__2), .inputs_451__1 (registerOutputs_451__1), .inputs_451__0 (
            registerOutputs_451__0), .inputs_452__15 (registerOutputs_452__15), 
            .inputs_452__14 (registerOutputs_452__14), .inputs_452__13 (
            registerOutputs_452__13), .inputs_452__12 (registerOutputs_452__12)
            , .inputs_452__11 (registerOutputs_452__11), .inputs_452__10 (
            registerOutputs_452__10), .inputs_452__9 (registerOutputs_452__9), .inputs_452__8 (
            registerOutputs_452__8), .inputs_452__7 (registerOutputs_452__7), .inputs_452__6 (
            registerOutputs_452__6), .inputs_452__5 (registerOutputs_452__5), .inputs_452__4 (
            registerOutputs_452__4), .inputs_452__3 (registerOutputs_452__3), .inputs_452__2 (
            registerOutputs_452__2), .inputs_452__1 (registerOutputs_452__1), .inputs_452__0 (
            registerOutputs_452__0), .inputs_453__15 (registerOutputs_453__15), 
            .inputs_453__14 (registerOutputs_453__14), .inputs_453__13 (
            registerOutputs_453__13), .inputs_453__12 (registerOutputs_453__12)
            , .inputs_453__11 (registerOutputs_453__11), .inputs_453__10 (
            registerOutputs_453__10), .inputs_453__9 (registerOutputs_453__9), .inputs_453__8 (
            registerOutputs_453__8), .inputs_453__7 (registerOutputs_453__7), .inputs_453__6 (
            registerOutputs_453__6), .inputs_453__5 (registerOutputs_453__5), .inputs_453__4 (
            registerOutputs_453__4), .inputs_453__3 (registerOutputs_453__3), .inputs_453__2 (
            registerOutputs_453__2), .inputs_453__1 (registerOutputs_453__1), .inputs_453__0 (
            registerOutputs_453__0), .inputs_454__15 (registerOutputs_454__15), 
            .inputs_454__14 (registerOutputs_454__14), .inputs_454__13 (
            registerOutputs_454__13), .inputs_454__12 (registerOutputs_454__12)
            , .inputs_454__11 (registerOutputs_454__11), .inputs_454__10 (
            registerOutputs_454__10), .inputs_454__9 (registerOutputs_454__9), .inputs_454__8 (
            registerOutputs_454__8), .inputs_454__7 (registerOutputs_454__7), .inputs_454__6 (
            registerOutputs_454__6), .inputs_454__5 (registerOutputs_454__5), .inputs_454__4 (
            registerOutputs_454__4), .inputs_454__3 (registerOutputs_454__3), .inputs_454__2 (
            registerOutputs_454__2), .inputs_454__1 (registerOutputs_454__1), .inputs_454__0 (
            registerOutputs_454__0), .inputs_455__15 (registerOutputs_455__15), 
            .inputs_455__14 (registerOutputs_455__14), .inputs_455__13 (
            registerOutputs_455__13), .inputs_455__12 (registerOutputs_455__12)
            , .inputs_455__11 (registerOutputs_455__11), .inputs_455__10 (
            registerOutputs_455__10), .inputs_455__9 (registerOutputs_455__9), .inputs_455__8 (
            registerOutputs_455__8), .inputs_455__7 (registerOutputs_455__7), .inputs_455__6 (
            registerOutputs_455__6), .inputs_455__5 (registerOutputs_455__5), .inputs_455__4 (
            registerOutputs_455__4), .inputs_455__3 (registerOutputs_455__3), .inputs_455__2 (
            registerOutputs_455__2), .inputs_455__1 (registerOutputs_455__1), .inputs_455__0 (
            registerOutputs_455__0), .inputs_456__15 (registerOutputs_456__15), 
            .inputs_456__14 (registerOutputs_456__14), .inputs_456__13 (
            registerOutputs_456__13), .inputs_456__12 (registerOutputs_456__12)
            , .inputs_456__11 (registerOutputs_456__11), .inputs_456__10 (
            registerOutputs_456__10), .inputs_456__9 (registerOutputs_456__9), .inputs_456__8 (
            registerOutputs_456__8), .inputs_456__7 (registerOutputs_456__7), .inputs_456__6 (
            registerOutputs_456__6), .inputs_456__5 (registerOutputs_456__5), .inputs_456__4 (
            registerOutputs_456__4), .inputs_456__3 (registerOutputs_456__3), .inputs_456__2 (
            registerOutputs_456__2), .inputs_456__1 (registerOutputs_456__1), .inputs_456__0 (
            registerOutputs_456__0), .inputs_457__15 (registerOutputs_457__15), 
            .inputs_457__14 (registerOutputs_457__14), .inputs_457__13 (
            registerOutputs_457__13), .inputs_457__12 (registerOutputs_457__12)
            , .inputs_457__11 (registerOutputs_457__11), .inputs_457__10 (
            registerOutputs_457__10), .inputs_457__9 (registerOutputs_457__9), .inputs_457__8 (
            registerOutputs_457__8), .inputs_457__7 (registerOutputs_457__7), .inputs_457__6 (
            registerOutputs_457__6), .inputs_457__5 (registerOutputs_457__5), .inputs_457__4 (
            registerOutputs_457__4), .inputs_457__3 (registerOutputs_457__3), .inputs_457__2 (
            registerOutputs_457__2), .inputs_457__1 (registerOutputs_457__1), .inputs_457__0 (
            registerOutputs_457__0), .inputs_458__15 (registerOutputs_458__15), 
            .inputs_458__14 (registerOutputs_458__14), .inputs_458__13 (
            registerOutputs_458__13), .inputs_458__12 (registerOutputs_458__12)
            , .inputs_458__11 (registerOutputs_458__11), .inputs_458__10 (
            registerOutputs_458__10), .inputs_458__9 (registerOutputs_458__9), .inputs_458__8 (
            registerOutputs_458__8), .inputs_458__7 (registerOutputs_458__7), .inputs_458__6 (
            registerOutputs_458__6), .inputs_458__5 (registerOutputs_458__5), .inputs_458__4 (
            registerOutputs_458__4), .inputs_458__3 (registerOutputs_458__3), .inputs_458__2 (
            registerOutputs_458__2), .inputs_458__1 (registerOutputs_458__1), .inputs_458__0 (
            registerOutputs_458__0), .inputs_459__15 (registerOutputs_459__15), 
            .inputs_459__14 (registerOutputs_459__14), .inputs_459__13 (
            registerOutputs_459__13), .inputs_459__12 (registerOutputs_459__12)
            , .inputs_459__11 (registerOutputs_459__11), .inputs_459__10 (
            registerOutputs_459__10), .inputs_459__9 (registerOutputs_459__9), .inputs_459__8 (
            registerOutputs_459__8), .inputs_459__7 (registerOutputs_459__7), .inputs_459__6 (
            registerOutputs_459__6), .inputs_459__5 (registerOutputs_459__5), .inputs_459__4 (
            registerOutputs_459__4), .inputs_459__3 (registerOutputs_459__3), .inputs_459__2 (
            registerOutputs_459__2), .inputs_459__1 (registerOutputs_459__1), .inputs_459__0 (
            registerOutputs_459__0), .inputs_460__15 (registerOutputs_460__15), 
            .inputs_460__14 (registerOutputs_460__14), .inputs_460__13 (
            registerOutputs_460__13), .inputs_460__12 (registerOutputs_460__12)
            , .inputs_460__11 (registerOutputs_460__11), .inputs_460__10 (
            registerOutputs_460__10), .inputs_460__9 (registerOutputs_460__9), .inputs_460__8 (
            registerOutputs_460__8), .inputs_460__7 (registerOutputs_460__7), .inputs_460__6 (
            registerOutputs_460__6), .inputs_460__5 (registerOutputs_460__5), .inputs_460__4 (
            registerOutputs_460__4), .inputs_460__3 (registerOutputs_460__3), .inputs_460__2 (
            registerOutputs_460__2), .inputs_460__1 (registerOutputs_460__1), .inputs_460__0 (
            registerOutputs_460__0), .inputs_461__15 (registerOutputs_461__15), 
            .inputs_461__14 (registerOutputs_461__14), .inputs_461__13 (
            registerOutputs_461__13), .inputs_461__12 (registerOutputs_461__12)
            , .inputs_461__11 (registerOutputs_461__11), .inputs_461__10 (
            registerOutputs_461__10), .inputs_461__9 (registerOutputs_461__9), .inputs_461__8 (
            registerOutputs_461__8), .inputs_461__7 (registerOutputs_461__7), .inputs_461__6 (
            registerOutputs_461__6), .inputs_461__5 (registerOutputs_461__5), .inputs_461__4 (
            registerOutputs_461__4), .inputs_461__3 (registerOutputs_461__3), .inputs_461__2 (
            registerOutputs_461__2), .inputs_461__1 (registerOutputs_461__1), .inputs_461__0 (
            registerOutputs_461__0), .inputs_462__15 (registerOutputs_462__15), 
            .inputs_462__14 (registerOutputs_462__14), .inputs_462__13 (
            registerOutputs_462__13), .inputs_462__12 (registerOutputs_462__12)
            , .inputs_462__11 (registerOutputs_462__11), .inputs_462__10 (
            registerOutputs_462__10), .inputs_462__9 (registerOutputs_462__9), .inputs_462__8 (
            registerOutputs_462__8), .inputs_462__7 (registerOutputs_462__7), .inputs_462__6 (
            registerOutputs_462__6), .inputs_462__5 (registerOutputs_462__5), .inputs_462__4 (
            registerOutputs_462__4), .inputs_462__3 (registerOutputs_462__3), .inputs_462__2 (
            registerOutputs_462__2), .inputs_462__1 (registerOutputs_462__1), .inputs_462__0 (
            registerOutputs_462__0), .inputs_463__15 (registerOutputs_463__15), 
            .inputs_463__14 (registerOutputs_463__14), .inputs_463__13 (
            registerOutputs_463__13), .inputs_463__12 (registerOutputs_463__12)
            , .inputs_463__11 (registerOutputs_463__11), .inputs_463__10 (
            registerOutputs_463__10), .inputs_463__9 (registerOutputs_463__9), .inputs_463__8 (
            registerOutputs_463__8), .inputs_463__7 (registerOutputs_463__7), .inputs_463__6 (
            registerOutputs_463__6), .inputs_463__5 (registerOutputs_463__5), .inputs_463__4 (
            registerOutputs_463__4), .inputs_463__3 (registerOutputs_463__3), .inputs_463__2 (
            registerOutputs_463__2), .inputs_463__1 (registerOutputs_463__1), .inputs_463__0 (
            registerOutputs_463__0), .inputs_464__15 (registerOutputs_464__15), 
            .inputs_464__14 (registerOutputs_464__14), .inputs_464__13 (
            registerOutputs_464__13), .inputs_464__12 (registerOutputs_464__12)
            , .inputs_464__11 (registerOutputs_464__11), .inputs_464__10 (
            registerOutputs_464__10), .inputs_464__9 (registerOutputs_464__9), .inputs_464__8 (
            registerOutputs_464__8), .inputs_464__7 (registerOutputs_464__7), .inputs_464__6 (
            registerOutputs_464__6), .inputs_464__5 (registerOutputs_464__5), .inputs_464__4 (
            registerOutputs_464__4), .inputs_464__3 (registerOutputs_464__3), .inputs_464__2 (
            registerOutputs_464__2), .inputs_464__1 (registerOutputs_464__1), .inputs_464__0 (
            registerOutputs_464__0), .inputs_465__15 (registerOutputs_465__15), 
            .inputs_465__14 (registerOutputs_465__14), .inputs_465__13 (
            registerOutputs_465__13), .inputs_465__12 (registerOutputs_465__12)
            , .inputs_465__11 (registerOutputs_465__11), .inputs_465__10 (
            registerOutputs_465__10), .inputs_465__9 (registerOutputs_465__9), .inputs_465__8 (
            registerOutputs_465__8), .inputs_465__7 (registerOutputs_465__7), .inputs_465__6 (
            registerOutputs_465__6), .inputs_465__5 (registerOutputs_465__5), .inputs_465__4 (
            registerOutputs_465__4), .inputs_465__3 (registerOutputs_465__3), .inputs_465__2 (
            registerOutputs_465__2), .inputs_465__1 (registerOutputs_465__1), .inputs_465__0 (
            registerOutputs_465__0), .inputs_466__15 (registerOutputs_466__15), 
            .inputs_466__14 (registerOutputs_466__14), .inputs_466__13 (
            registerOutputs_466__13), .inputs_466__12 (registerOutputs_466__12)
            , .inputs_466__11 (registerOutputs_466__11), .inputs_466__10 (
            registerOutputs_466__10), .inputs_466__9 (registerOutputs_466__9), .inputs_466__8 (
            registerOutputs_466__8), .inputs_466__7 (registerOutputs_466__7), .inputs_466__6 (
            registerOutputs_466__6), .inputs_466__5 (registerOutputs_466__5), .inputs_466__4 (
            registerOutputs_466__4), .inputs_466__3 (registerOutputs_466__3), .inputs_466__2 (
            registerOutputs_466__2), .inputs_466__1 (registerOutputs_466__1), .inputs_466__0 (
            registerOutputs_466__0), .inputs_467__15 (registerOutputs_467__15), 
            .inputs_467__14 (registerOutputs_467__14), .inputs_467__13 (
            registerOutputs_467__13), .inputs_467__12 (registerOutputs_467__12)
            , .inputs_467__11 (registerOutputs_467__11), .inputs_467__10 (
            registerOutputs_467__10), .inputs_467__9 (registerOutputs_467__9), .inputs_467__8 (
            registerOutputs_467__8), .inputs_467__7 (registerOutputs_467__7), .inputs_467__6 (
            registerOutputs_467__6), .inputs_467__5 (registerOutputs_467__5), .inputs_467__4 (
            registerOutputs_467__4), .inputs_467__3 (registerOutputs_467__3), .inputs_467__2 (
            registerOutputs_467__2), .inputs_467__1 (registerOutputs_467__1), .inputs_467__0 (
            registerOutputs_467__0), .inputs_468__15 (registerOutputs_468__15), 
            .inputs_468__14 (registerOutputs_468__14), .inputs_468__13 (
            registerOutputs_468__13), .inputs_468__12 (registerOutputs_468__12)
            , .inputs_468__11 (registerOutputs_468__11), .inputs_468__10 (
            registerOutputs_468__10), .inputs_468__9 (registerOutputs_468__9), .inputs_468__8 (
            registerOutputs_468__8), .inputs_468__7 (registerOutputs_468__7), .inputs_468__6 (
            registerOutputs_468__6), .inputs_468__5 (registerOutputs_468__5), .inputs_468__4 (
            registerOutputs_468__4), .inputs_468__3 (registerOutputs_468__3), .inputs_468__2 (
            registerOutputs_468__2), .inputs_468__1 (registerOutputs_468__1), .inputs_468__0 (
            registerOutputs_468__0), .inputs_469__15 (registerOutputs_469__15), 
            .inputs_469__14 (registerOutputs_469__14), .inputs_469__13 (
            registerOutputs_469__13), .inputs_469__12 (registerOutputs_469__12)
            , .inputs_469__11 (registerOutputs_469__11), .inputs_469__10 (
            registerOutputs_469__10), .inputs_469__9 (registerOutputs_469__9), .inputs_469__8 (
            registerOutputs_469__8), .inputs_469__7 (registerOutputs_469__7), .inputs_469__6 (
            registerOutputs_469__6), .inputs_469__5 (registerOutputs_469__5), .inputs_469__4 (
            registerOutputs_469__4), .inputs_469__3 (registerOutputs_469__3), .inputs_469__2 (
            registerOutputs_469__2), .inputs_469__1 (registerOutputs_469__1), .inputs_469__0 (
            registerOutputs_469__0), .inputs_470__15 (registerOutputs_470__15), 
            .inputs_470__14 (registerOutputs_470__14), .inputs_470__13 (
            registerOutputs_470__13), .inputs_470__12 (registerOutputs_470__12)
            , .inputs_470__11 (registerOutputs_470__11), .inputs_470__10 (
            registerOutputs_470__10), .inputs_470__9 (registerOutputs_470__9), .inputs_470__8 (
            registerOutputs_470__8), .inputs_470__7 (registerOutputs_470__7), .inputs_470__6 (
            registerOutputs_470__6), .inputs_470__5 (registerOutputs_470__5), .inputs_470__4 (
            registerOutputs_470__4), .inputs_470__3 (registerOutputs_470__3), .inputs_470__2 (
            registerOutputs_470__2), .inputs_470__1 (registerOutputs_470__1), .inputs_470__0 (
            registerOutputs_470__0), .inputs_471__15 (registerOutputs_471__15), 
            .inputs_471__14 (registerOutputs_471__14), .inputs_471__13 (
            registerOutputs_471__13), .inputs_471__12 (registerOutputs_471__12)
            , .inputs_471__11 (registerOutputs_471__11), .inputs_471__10 (
            registerOutputs_471__10), .inputs_471__9 (registerOutputs_471__9), .inputs_471__8 (
            registerOutputs_471__8), .inputs_471__7 (registerOutputs_471__7), .inputs_471__6 (
            registerOutputs_471__6), .inputs_471__5 (registerOutputs_471__5), .inputs_471__4 (
            registerOutputs_471__4), .inputs_471__3 (registerOutputs_471__3), .inputs_471__2 (
            registerOutputs_471__2), .inputs_471__1 (registerOutputs_471__1), .inputs_471__0 (
            registerOutputs_471__0), .inputs_472__15 (registerOutputs_472__15), 
            .inputs_472__14 (registerOutputs_472__14), .inputs_472__13 (
            registerOutputs_472__13), .inputs_472__12 (registerOutputs_472__12)
            , .inputs_472__11 (registerOutputs_472__11), .inputs_472__10 (
            registerOutputs_472__10), .inputs_472__9 (registerOutputs_472__9), .inputs_472__8 (
            registerOutputs_472__8), .inputs_472__7 (registerOutputs_472__7), .inputs_472__6 (
            registerOutputs_472__6), .inputs_472__5 (registerOutputs_472__5), .inputs_472__4 (
            registerOutputs_472__4), .inputs_472__3 (registerOutputs_472__3), .inputs_472__2 (
            registerOutputs_472__2), .inputs_472__1 (registerOutputs_472__1), .inputs_472__0 (
            registerOutputs_472__0), .inputs_473__15 (registerOutputs_473__15), 
            .inputs_473__14 (registerOutputs_473__14), .inputs_473__13 (
            registerOutputs_473__13), .inputs_473__12 (registerOutputs_473__12)
            , .inputs_473__11 (registerOutputs_473__11), .inputs_473__10 (
            registerOutputs_473__10), .inputs_473__9 (registerOutputs_473__9), .inputs_473__8 (
            registerOutputs_473__8), .inputs_473__7 (registerOutputs_473__7), .inputs_473__6 (
            registerOutputs_473__6), .inputs_473__5 (registerOutputs_473__5), .inputs_473__4 (
            registerOutputs_473__4), .inputs_473__3 (registerOutputs_473__3), .inputs_473__2 (
            registerOutputs_473__2), .inputs_473__1 (registerOutputs_473__1), .inputs_473__0 (
            registerOutputs_473__0), .inputs_474__15 (registerOutputs_474__15), 
            .inputs_474__14 (registerOutputs_474__14), .inputs_474__13 (
            registerOutputs_474__13), .inputs_474__12 (registerOutputs_474__12)
            , .inputs_474__11 (registerOutputs_474__11), .inputs_474__10 (
            registerOutputs_474__10), .inputs_474__9 (registerOutputs_474__9), .inputs_474__8 (
            registerOutputs_474__8), .inputs_474__7 (registerOutputs_474__7), .inputs_474__6 (
            registerOutputs_474__6), .inputs_474__5 (registerOutputs_474__5), .inputs_474__4 (
            registerOutputs_474__4), .inputs_474__3 (registerOutputs_474__3), .inputs_474__2 (
            registerOutputs_474__2), .inputs_474__1 (registerOutputs_474__1), .inputs_474__0 (
            registerOutputs_474__0), .inputs_475__15 (registerOutputs_475__15), 
            .inputs_475__14 (registerOutputs_475__14), .inputs_475__13 (
            registerOutputs_475__13), .inputs_475__12 (registerOutputs_475__12)
            , .inputs_475__11 (registerOutputs_475__11), .inputs_475__10 (
            registerOutputs_475__10), .inputs_475__9 (registerOutputs_475__9), .inputs_475__8 (
            registerOutputs_475__8), .inputs_475__7 (registerOutputs_475__7), .inputs_475__6 (
            registerOutputs_475__6), .inputs_475__5 (registerOutputs_475__5), .inputs_475__4 (
            registerOutputs_475__4), .inputs_475__3 (registerOutputs_475__3), .inputs_475__2 (
            registerOutputs_475__2), .inputs_475__1 (registerOutputs_475__1), .inputs_475__0 (
            registerOutputs_475__0), .inputs_476__15 (registerOutputs_476__15), 
            .inputs_476__14 (registerOutputs_476__14), .inputs_476__13 (
            registerOutputs_476__13), .inputs_476__12 (registerOutputs_476__12)
            , .inputs_476__11 (registerOutputs_476__11), .inputs_476__10 (
            registerOutputs_476__10), .inputs_476__9 (registerOutputs_476__9), .inputs_476__8 (
            registerOutputs_476__8), .inputs_476__7 (registerOutputs_476__7), .inputs_476__6 (
            registerOutputs_476__6), .inputs_476__5 (registerOutputs_476__5), .inputs_476__4 (
            registerOutputs_476__4), .inputs_476__3 (registerOutputs_476__3), .inputs_476__2 (
            registerOutputs_476__2), .inputs_476__1 (registerOutputs_476__1), .inputs_476__0 (
            registerOutputs_476__0), .inputs_477__15 (registerOutputs_477__15), 
            .inputs_477__14 (registerOutputs_477__14), .inputs_477__13 (
            registerOutputs_477__13), .inputs_477__12 (registerOutputs_477__12)
            , .inputs_477__11 (registerOutputs_477__11), .inputs_477__10 (
            registerOutputs_477__10), .inputs_477__9 (registerOutputs_477__9), .inputs_477__8 (
            registerOutputs_477__8), .inputs_477__7 (registerOutputs_477__7), .inputs_477__6 (
            registerOutputs_477__6), .inputs_477__5 (registerOutputs_477__5), .inputs_477__4 (
            registerOutputs_477__4), .inputs_477__3 (registerOutputs_477__3), .inputs_477__2 (
            registerOutputs_477__2), .inputs_477__1 (registerOutputs_477__1), .inputs_477__0 (
            registerOutputs_477__0), .inputs_478__15 (registerOutputs_478__15), 
            .inputs_478__14 (registerOutputs_478__14), .inputs_478__13 (
            registerOutputs_478__13), .inputs_478__12 (registerOutputs_478__12)
            , .inputs_478__11 (registerOutputs_478__11), .inputs_478__10 (
            registerOutputs_478__10), .inputs_478__9 (registerOutputs_478__9), .inputs_478__8 (
            registerOutputs_478__8), .inputs_478__7 (registerOutputs_478__7), .inputs_478__6 (
            registerOutputs_478__6), .inputs_478__5 (registerOutputs_478__5), .inputs_478__4 (
            registerOutputs_478__4), .inputs_478__3 (registerOutputs_478__3), .inputs_478__2 (
            registerOutputs_478__2), .inputs_478__1 (registerOutputs_478__1), .inputs_478__0 (
            registerOutputs_478__0), .inputs_479__15 (registerOutputs_479__15), 
            .inputs_479__14 (registerOutputs_479__14), .inputs_479__13 (
            registerOutputs_479__13), .inputs_479__12 (registerOutputs_479__12)
            , .inputs_479__11 (registerOutputs_479__11), .inputs_479__10 (
            registerOutputs_479__10), .inputs_479__9 (registerOutputs_479__9), .inputs_479__8 (
            registerOutputs_479__8), .inputs_479__7 (registerOutputs_479__7), .inputs_479__6 (
            registerOutputs_479__6), .inputs_479__5 (registerOutputs_479__5), .inputs_479__4 (
            registerOutputs_479__4), .inputs_479__3 (registerOutputs_479__3), .inputs_479__2 (
            registerOutputs_479__2), .inputs_479__1 (registerOutputs_479__1), .inputs_479__0 (
            registerOutputs_479__0), .inputs_480__15 (registerOutputs_480__15), 
            .inputs_480__14 (registerOutputs_480__14), .inputs_480__13 (
            registerOutputs_480__13), .inputs_480__12 (registerOutputs_480__12)
            , .inputs_480__11 (registerOutputs_480__11), .inputs_480__10 (
            registerOutputs_480__10), .inputs_480__9 (registerOutputs_480__9), .inputs_480__8 (
            registerOutputs_480__8), .inputs_480__7 (registerOutputs_480__7), .inputs_480__6 (
            registerOutputs_480__6), .inputs_480__5 (registerOutputs_480__5), .inputs_480__4 (
            registerOutputs_480__4), .inputs_480__3 (registerOutputs_480__3), .inputs_480__2 (
            registerOutputs_480__2), .inputs_480__1 (registerOutputs_480__1), .inputs_480__0 (
            registerOutputs_480__0), .inputs_481__15 (registerOutputs_481__15), 
            .inputs_481__14 (registerOutputs_481__14), .inputs_481__13 (
            registerOutputs_481__13), .inputs_481__12 (registerOutputs_481__12)
            , .inputs_481__11 (registerOutputs_481__11), .inputs_481__10 (
            registerOutputs_481__10), .inputs_481__9 (registerOutputs_481__9), .inputs_481__8 (
            registerOutputs_481__8), .inputs_481__7 (registerOutputs_481__7), .inputs_481__6 (
            registerOutputs_481__6), .inputs_481__5 (registerOutputs_481__5), .inputs_481__4 (
            registerOutputs_481__4), .inputs_481__3 (registerOutputs_481__3), .inputs_481__2 (
            registerOutputs_481__2), .inputs_481__1 (registerOutputs_481__1), .inputs_481__0 (
            registerOutputs_481__0), .inputs_482__15 (registerOutputs_482__15), 
            .inputs_482__14 (registerOutputs_482__14), .inputs_482__13 (
            registerOutputs_482__13), .inputs_482__12 (registerOutputs_482__12)
            , .inputs_482__11 (registerOutputs_482__11), .inputs_482__10 (
            registerOutputs_482__10), .inputs_482__9 (registerOutputs_482__9), .inputs_482__8 (
            registerOutputs_482__8), .inputs_482__7 (registerOutputs_482__7), .inputs_482__6 (
            registerOutputs_482__6), .inputs_482__5 (registerOutputs_482__5), .inputs_482__4 (
            registerOutputs_482__4), .inputs_482__3 (registerOutputs_482__3), .inputs_482__2 (
            registerOutputs_482__2), .inputs_482__1 (registerOutputs_482__1), .inputs_482__0 (
            registerOutputs_482__0), .inputs_483__15 (registerOutputs_483__15), 
            .inputs_483__14 (registerOutputs_483__14), .inputs_483__13 (
            registerOutputs_483__13), .inputs_483__12 (registerOutputs_483__12)
            , .inputs_483__11 (registerOutputs_483__11), .inputs_483__10 (
            registerOutputs_483__10), .inputs_483__9 (registerOutputs_483__9), .inputs_483__8 (
            registerOutputs_483__8), .inputs_483__7 (registerOutputs_483__7), .inputs_483__6 (
            registerOutputs_483__6), .inputs_483__5 (registerOutputs_483__5), .inputs_483__4 (
            registerOutputs_483__4), .inputs_483__3 (registerOutputs_483__3), .inputs_483__2 (
            registerOutputs_483__2), .inputs_483__1 (registerOutputs_483__1), .inputs_483__0 (
            registerOutputs_483__0), .inputs_484__15 (registerOutputs_484__15), 
            .inputs_484__14 (registerOutputs_484__15), .inputs_484__13 (
            registerOutputs_484__15), .inputs_484__12 (registerOutputs_484__15)
            , .inputs_484__11 (registerOutputs_484__15), .inputs_484__10 (
            registerOutputs_484__15), .inputs_484__9 (registerOutputs_484__15), 
            .inputs_484__8 (registerOutputs_484__15), .inputs_484__7 (
            registerOutputs_484__15), .inputs_484__6 (registerOutputs_484__15), 
            .inputs_484__5 (registerOutputs_484__15), .inputs_484__4 (
            registerOutputs_484__15), .inputs_484__3 (registerOutputs_484__15), 
            .inputs_484__2 (registerOutputs_484__15), .inputs_484__1 (
            registerOutputs_484__15), .inputs_484__0 (registerOutputs_484__15), 
            .inputs_485__15 (registerOutputs_484__15), .inputs_485__14 (
            registerOutputs_484__15), .inputs_485__13 (registerOutputs_484__15)
            , .inputs_485__12 (registerOutputs_484__15), .inputs_485__11 (
            registerOutputs_484__15), .inputs_485__10 (registerOutputs_484__15)
            , .inputs_485__9 (registerOutputs_484__15), .inputs_485__8 (
            registerOutputs_484__15), .inputs_485__7 (registerOutputs_484__15), 
            .inputs_485__6 (registerOutputs_484__15), .inputs_485__5 (
            registerOutputs_484__15), .inputs_485__4 (registerOutputs_484__15), 
            .inputs_485__3 (registerOutputs_484__15), .inputs_485__2 (
            registerOutputs_484__15), .inputs_485__1 (registerOutputs_484__15), 
            .inputs_485__0 (registerOutputs_484__15), .inputs_486__15 (
            registerOutputs_484__15), .inputs_486__14 (registerOutputs_484__15)
            , .inputs_486__13 (registerOutputs_484__15), .inputs_486__12 (
            registerOutputs_484__15), .inputs_486__11 (registerOutputs_484__15)
            , .inputs_486__10 (registerOutputs_484__15), .inputs_486__9 (
            registerOutputs_484__15), .inputs_486__8 (registerOutputs_484__15), 
            .inputs_486__7 (registerOutputs_484__15), .inputs_486__6 (
            registerOutputs_484__15), .inputs_486__5 (registerOutputs_484__15), 
            .inputs_486__4 (registerOutputs_484__15), .inputs_486__3 (
            registerOutputs_484__15), .inputs_486__2 (registerOutputs_484__15), 
            .inputs_486__1 (registerOutputs_484__15), .inputs_486__0 (
            registerOutputs_484__15), .inputs_487__15 (registerOutputs_484__15)
            , .inputs_487__14 (registerOutputs_484__15), .inputs_487__13 (
            registerOutputs_484__15), .inputs_487__12 (registerOutputs_484__15)
            , .inputs_487__11 (registerOutputs_484__15), .inputs_487__10 (
            registerOutputs_484__15), .inputs_487__9 (registerOutputs_484__15), 
            .inputs_487__8 (registerOutputs_484__15), .inputs_487__7 (
            registerOutputs_484__15), .inputs_487__6 (registerOutputs_484__15), 
            .inputs_487__5 (registerOutputs_484__15), .inputs_487__4 (
            registerOutputs_484__15), .inputs_487__3 (registerOutputs_484__15), 
            .inputs_487__2 (registerOutputs_484__15), .inputs_487__1 (
            registerOutputs_484__15), .inputs_487__0 (registerOutputs_484__15), 
            .inputs_488__15 (registerOutputs_484__15), .inputs_488__14 (
            registerOutputs_484__15), .inputs_488__13 (registerOutputs_484__15)
            , .inputs_488__12 (registerOutputs_484__15), .inputs_488__11 (
            registerOutputs_484__15), .inputs_488__10 (registerOutputs_484__15)
            , .inputs_488__9 (registerOutputs_484__15), .inputs_488__8 (
            registerOutputs_484__15), .inputs_488__7 (registerOutputs_484__15), 
            .inputs_488__6 (registerOutputs_484__15), .inputs_488__5 (
            registerOutputs_484__15), .inputs_488__4 (registerOutputs_484__15), 
            .inputs_488__3 (registerOutputs_484__15), .inputs_488__2 (
            registerOutputs_484__15), .inputs_488__1 (registerOutputs_484__15), 
            .inputs_488__0 (registerOutputs_484__15), .inputs_489__15 (
            registerOutputs_484__15), .inputs_489__14 (registerOutputs_484__15)
            , .inputs_489__13 (registerOutputs_484__15), .inputs_489__12 (
            registerOutputs_484__15), .inputs_489__11 (registerOutputs_484__15)
            , .inputs_489__10 (registerOutputs_484__15), .inputs_489__9 (
            registerOutputs_484__15), .inputs_489__8 (registerOutputs_484__15), 
            .inputs_489__7 (registerOutputs_484__15), .inputs_489__6 (
            registerOutputs_484__15), .inputs_489__5 (registerOutputs_484__15), 
            .inputs_489__4 (registerOutputs_484__15), .inputs_489__3 (
            registerOutputs_484__15), .inputs_489__2 (registerOutputs_484__15), 
            .inputs_489__1 (registerOutputs_484__15), .inputs_489__0 (
            registerOutputs_484__15), .inputs_490__15 (registerOutputs_484__15)
            , .inputs_490__14 (registerOutputs_484__15), .inputs_490__13 (
            registerOutputs_484__15), .inputs_490__12 (registerOutputs_484__15)
            , .inputs_490__11 (registerOutputs_484__15), .inputs_490__10 (
            registerOutputs_484__15), .inputs_490__9 (registerOutputs_484__15), 
            .inputs_490__8 (registerOutputs_484__15), .inputs_490__7 (
            registerOutputs_484__15), .inputs_490__6 (registerOutputs_484__15), 
            .inputs_490__5 (registerOutputs_484__15), .inputs_490__4 (
            registerOutputs_484__15), .inputs_490__3 (registerOutputs_484__15), 
            .inputs_490__2 (registerOutputs_484__15), .inputs_490__1 (
            registerOutputs_484__15), .inputs_490__0 (registerOutputs_484__15), 
            .inputs_491__15 (registerOutputs_484__15), .inputs_491__14 (
            registerOutputs_484__15), .inputs_491__13 (registerOutputs_484__15)
            , .inputs_491__12 (registerOutputs_484__15), .inputs_491__11 (
            registerOutputs_484__15), .inputs_491__10 (registerOutputs_484__15)
            , .inputs_491__9 (registerOutputs_484__15), .inputs_491__8 (
            registerOutputs_484__15), .inputs_491__7 (registerOutputs_484__15), 
            .inputs_491__6 (registerOutputs_484__15), .inputs_491__5 (
            registerOutputs_484__15), .inputs_491__4 (registerOutputs_484__15), 
            .inputs_491__3 (registerOutputs_484__15), .inputs_491__2 (
            registerOutputs_484__15), .inputs_491__1 (registerOutputs_484__15), 
            .inputs_491__0 (registerOutputs_484__15), .inputs_492__15 (
            registerOutputs_484__15), .inputs_492__14 (registerOutputs_484__15)
            , .inputs_492__13 (registerOutputs_484__15), .inputs_492__12 (
            registerOutputs_484__15), .inputs_492__11 (registerOutputs_484__15)
            , .inputs_492__10 (registerOutputs_484__15), .inputs_492__9 (
            registerOutputs_484__15), .inputs_492__8 (registerOutputs_484__15), 
            .inputs_492__7 (registerOutputs_484__15), .inputs_492__6 (
            registerOutputs_484__15), .inputs_492__5 (registerOutputs_484__15), 
            .inputs_492__4 (registerOutputs_484__15), .inputs_492__3 (
            registerOutputs_484__15), .inputs_492__2 (registerOutputs_484__15), 
            .inputs_492__1 (registerOutputs_484__15), .inputs_492__0 (
            registerOutputs_484__15), .inputs_493__15 (registerOutputs_484__15)
            , .inputs_493__14 (registerOutputs_484__15), .inputs_493__13 (
            registerOutputs_484__15), .inputs_493__12 (registerOutputs_484__15)
            , .inputs_493__11 (registerOutputs_484__15), .inputs_493__10 (
            registerOutputs_484__15), .inputs_493__9 (registerOutputs_484__15), 
            .inputs_493__8 (registerOutputs_484__15), .inputs_493__7 (
            registerOutputs_484__15), .inputs_493__6 (registerOutputs_484__15), 
            .inputs_493__5 (registerOutputs_484__15), .inputs_493__4 (
            registerOutputs_484__15), .inputs_493__3 (registerOutputs_484__15), 
            .inputs_493__2 (registerOutputs_484__15), .inputs_493__1 (
            registerOutputs_484__15), .inputs_493__0 (registerOutputs_484__15), 
            .inputs_494__15 (registerOutputs_484__15), .inputs_494__14 (
            registerOutputs_484__15), .inputs_494__13 (registerOutputs_484__15)
            , .inputs_494__12 (registerOutputs_484__15), .inputs_494__11 (
            registerOutputs_484__15), .inputs_494__10 (registerOutputs_484__15)
            , .inputs_494__9 (registerOutputs_484__15), .inputs_494__8 (
            registerOutputs_484__15), .inputs_494__7 (registerOutputs_484__15), 
            .inputs_494__6 (registerOutputs_484__15), .inputs_494__5 (
            registerOutputs_484__15), .inputs_494__4 (registerOutputs_484__15), 
            .inputs_494__3 (registerOutputs_484__15), .inputs_494__2 (
            registerOutputs_484__15), .inputs_494__1 (registerOutputs_484__15), 
            .inputs_494__0 (registerOutputs_484__15), .inputs_495__15 (
            registerOutputs_484__15), .inputs_495__14 (registerOutputs_484__15)
            , .inputs_495__13 (registerOutputs_484__15), .inputs_495__12 (
            registerOutputs_484__15), .inputs_495__11 (registerOutputs_484__15)
            , .inputs_495__10 (registerOutputs_484__15), .inputs_495__9 (
            registerOutputs_484__15), .inputs_495__8 (registerOutputs_484__15), 
            .inputs_495__7 (registerOutputs_484__15), .inputs_495__6 (
            registerOutputs_484__15), .inputs_495__5 (registerOutputs_484__15), 
            .inputs_495__4 (registerOutputs_484__15), .inputs_495__3 (
            registerOutputs_484__15), .inputs_495__2 (registerOutputs_484__15), 
            .inputs_495__1 (registerOutputs_484__15), .inputs_495__0 (
            registerOutputs_484__15), .inputs_496__15 (registerOutputs_484__15)
            , .inputs_496__14 (registerOutputs_484__15), .inputs_496__13 (
            registerOutputs_484__15), .inputs_496__12 (registerOutputs_484__15)
            , .inputs_496__11 (registerOutputs_484__15), .inputs_496__10 (
            registerOutputs_484__15), .inputs_496__9 (registerOutputs_484__15), 
            .inputs_496__8 (registerOutputs_484__15), .inputs_496__7 (
            registerOutputs_484__15), .inputs_496__6 (registerOutputs_484__15), 
            .inputs_496__5 (registerOutputs_484__15), .inputs_496__4 (
            registerOutputs_484__15), .inputs_496__3 (registerOutputs_484__15), 
            .inputs_496__2 (registerOutputs_484__15), .inputs_496__1 (
            registerOutputs_484__15), .inputs_496__0 (registerOutputs_484__15), 
            .inputs_497__15 (registerOutputs_484__15), .inputs_497__14 (
            registerOutputs_484__15), .inputs_497__13 (registerOutputs_484__15)
            , .inputs_497__12 (registerOutputs_484__15), .inputs_497__11 (
            registerOutputs_484__15), .inputs_497__10 (registerOutputs_484__15)
            , .inputs_497__9 (registerOutputs_484__15), .inputs_497__8 (
            registerOutputs_484__15), .inputs_497__7 (registerOutputs_484__15), 
            .inputs_497__6 (registerOutputs_484__15), .inputs_497__5 (
            registerOutputs_484__15), .inputs_497__4 (registerOutputs_484__15), 
            .inputs_497__3 (registerOutputs_484__15), .inputs_497__2 (
            registerOutputs_484__15), .inputs_497__1 (registerOutputs_484__15), 
            .inputs_497__0 (registerOutputs_484__15), .inputs_498__15 (
            registerOutputs_484__15), .inputs_498__14 (registerOutputs_484__15)
            , .inputs_498__13 (registerOutputs_484__15), .inputs_498__12 (
            registerOutputs_484__15), .inputs_498__11 (registerOutputs_484__15)
            , .inputs_498__10 (registerOutputs_484__15), .inputs_498__9 (
            registerOutputs_484__15), .inputs_498__8 (registerOutputs_484__15), 
            .inputs_498__7 (registerOutputs_484__15), .inputs_498__6 (
            registerOutputs_484__15), .inputs_498__5 (registerOutputs_484__15), 
            .inputs_498__4 (registerOutputs_484__15), .inputs_498__3 (
            registerOutputs_484__15), .inputs_498__2 (registerOutputs_484__15), 
            .inputs_498__1 (registerOutputs_484__15), .inputs_498__0 (
            registerOutputs_484__15), .inputs_499__15 (registerOutputs_484__15)
            , .inputs_499__14 (registerOutputs_484__15), .inputs_499__13 (
            registerOutputs_484__15), .inputs_499__12 (registerOutputs_484__15)
            , .inputs_499__11 (registerOutputs_484__15), .inputs_499__10 (
            registerOutputs_484__15), .inputs_499__9 (registerOutputs_484__15), 
            .inputs_499__8 (registerOutputs_484__15), .inputs_499__7 (
            registerOutputs_484__15), .inputs_499__6 (registerOutputs_484__15), 
            .inputs_499__5 (registerOutputs_484__15), .inputs_499__4 (
            registerOutputs_484__15), .inputs_499__3 (registerOutputs_484__15), 
            .inputs_499__2 (registerOutputs_484__15), .inputs_499__1 (
            registerOutputs_484__15), .inputs_499__0 (registerOutputs_484__15), 
            .inputs_500__15 (registerOutputs_484__15), .inputs_500__14 (
            registerOutputs_484__15), .inputs_500__13 (registerOutputs_484__15)
            , .inputs_500__12 (registerOutputs_484__15), .inputs_500__11 (
            registerOutputs_484__15), .inputs_500__10 (registerOutputs_484__15)
            , .inputs_500__9 (registerOutputs_484__15), .inputs_500__8 (
            registerOutputs_484__15), .inputs_500__7 (registerOutputs_484__15), 
            .inputs_500__6 (registerOutputs_484__15), .inputs_500__5 (
            registerOutputs_484__15), .inputs_500__4 (registerOutputs_484__15), 
            .inputs_500__3 (registerOutputs_484__15), .inputs_500__2 (
            registerOutputs_484__15), .inputs_500__1 (registerOutputs_484__15), 
            .inputs_500__0 (registerOutputs_484__15), .inputs_501__15 (
            registerOutputs_484__15), .inputs_501__14 (registerOutputs_484__15)
            , .inputs_501__13 (registerOutputs_484__15), .inputs_501__12 (
            registerOutputs_484__15), .inputs_501__11 (registerOutputs_484__15)
            , .inputs_501__10 (registerOutputs_484__15), .inputs_501__9 (
            registerOutputs_484__15), .inputs_501__8 (registerOutputs_484__15), 
            .inputs_501__7 (registerOutputs_484__15), .inputs_501__6 (
            registerOutputs_484__15), .inputs_501__5 (registerOutputs_484__15), 
            .inputs_501__4 (registerOutputs_484__15), .inputs_501__3 (
            registerOutputs_484__15), .inputs_501__2 (registerOutputs_484__15), 
            .inputs_501__1 (registerOutputs_484__15), .inputs_501__0 (
            registerOutputs_484__15), .inputs_502__15 (registerOutputs_484__15)
            , .inputs_502__14 (registerOutputs_484__15), .inputs_502__13 (
            registerOutputs_484__15), .inputs_502__12 (registerOutputs_484__15)
            , .inputs_502__11 (registerOutputs_484__15), .inputs_502__10 (
            registerOutputs_484__15), .inputs_502__9 (registerOutputs_484__15), 
            .inputs_502__8 (registerOutputs_484__15), .inputs_502__7 (
            registerOutputs_484__15), .inputs_502__6 (registerOutputs_484__15), 
            .inputs_502__5 (registerOutputs_484__15), .inputs_502__4 (
            registerOutputs_484__15), .inputs_502__3 (registerOutputs_484__15), 
            .inputs_502__2 (registerOutputs_484__15), .inputs_502__1 (
            registerOutputs_484__15), .inputs_502__0 (registerOutputs_484__15), 
            .inputs_503__15 (registerOutputs_484__15), .inputs_503__14 (
            registerOutputs_484__15), .inputs_503__13 (registerOutputs_484__15)
            , .inputs_503__12 (registerOutputs_484__15), .inputs_503__11 (
            registerOutputs_484__15), .inputs_503__10 (registerOutputs_484__15)
            , .inputs_503__9 (registerOutputs_484__15), .inputs_503__8 (
            registerOutputs_484__15), .inputs_503__7 (registerOutputs_484__15), 
            .inputs_503__6 (registerOutputs_484__15), .inputs_503__5 (
            registerOutputs_484__15), .inputs_503__4 (registerOutputs_484__15), 
            .inputs_503__3 (registerOutputs_484__15), .inputs_503__2 (
            registerOutputs_484__15), .inputs_503__1 (registerOutputs_484__15), 
            .inputs_503__0 (registerOutputs_484__15), .inputs_504__15 (
            registerOutputs_484__15), .inputs_504__14 (registerOutputs_484__15)
            , .inputs_504__13 (registerOutputs_484__15), .inputs_504__12 (
            registerOutputs_484__15), .inputs_504__11 (registerOutputs_484__15)
            , .inputs_504__10 (registerOutputs_484__15), .inputs_504__9 (
            registerOutputs_484__15), .inputs_504__8 (registerOutputs_484__15), 
            .inputs_504__7 (registerOutputs_484__15), .inputs_504__6 (
            registerOutputs_484__15), .inputs_504__5 (registerOutputs_484__15), 
            .inputs_504__4 (registerOutputs_484__15), .inputs_504__3 (
            registerOutputs_484__15), .inputs_504__2 (registerOutputs_484__15), 
            .inputs_504__1 (registerOutputs_484__15), .inputs_504__0 (
            registerOutputs_484__15), .inputs_505__15 (registerOutputs_484__15)
            , .inputs_505__14 (registerOutputs_484__15), .inputs_505__13 (
            registerOutputs_484__15), .inputs_505__12 (registerOutputs_484__15)
            , .inputs_505__11 (registerOutputs_484__15), .inputs_505__10 (
            registerOutputs_484__15), .inputs_505__9 (registerOutputs_484__15), 
            .inputs_505__8 (registerOutputs_484__15), .inputs_505__7 (
            registerOutputs_484__15), .inputs_505__6 (registerOutputs_484__15), 
            .inputs_505__5 (registerOutputs_484__15), .inputs_505__4 (
            registerOutputs_484__15), .inputs_505__3 (registerOutputs_484__15), 
            .inputs_505__2 (registerOutputs_484__15), .inputs_505__1 (
            registerOutputs_484__15), .inputs_505__0 (registerOutputs_484__15), 
            .inputs_506__15 (registerOutputs_484__15), .inputs_506__14 (
            registerOutputs_484__15), .inputs_506__13 (registerOutputs_484__15)
            , .inputs_506__12 (registerOutputs_484__15), .inputs_506__11 (
            registerOutputs_484__15), .inputs_506__10 (registerOutputs_484__15)
            , .inputs_506__9 (registerOutputs_484__15), .inputs_506__8 (
            registerOutputs_484__15), .inputs_506__7 (registerOutputs_484__15), 
            .inputs_506__6 (registerOutputs_484__15), .inputs_506__5 (
            registerOutputs_484__15), .inputs_506__4 (registerOutputs_484__15), 
            .inputs_506__3 (registerOutputs_484__15), .inputs_506__2 (
            registerOutputs_484__15), .inputs_506__1 (registerOutputs_484__15), 
            .inputs_506__0 (registerOutputs_484__15), .inputs_507__15 (
            registerOutputs_484__15), .inputs_507__14 (registerOutputs_484__15)
            , .inputs_507__13 (registerOutputs_484__15), .inputs_507__12 (
            registerOutputs_484__15), .inputs_507__11 (registerOutputs_484__15)
            , .inputs_507__10 (registerOutputs_484__15), .inputs_507__9 (
            registerOutputs_484__15), .inputs_507__8 (registerOutputs_484__15), 
            .inputs_507__7 (registerOutputs_484__15), .inputs_507__6 (
            registerOutputs_484__15), .inputs_507__5 (registerOutputs_484__15), 
            .inputs_507__4 (registerOutputs_484__15), .inputs_507__3 (
            registerOutputs_484__15), .inputs_507__2 (registerOutputs_484__15), 
            .inputs_507__1 (registerOutputs_484__15), .inputs_507__0 (
            registerOutputs_484__15), .inputs_508__15 (registerOutputs_484__15)
            , .inputs_508__14 (registerOutputs_484__15), .inputs_508__13 (
            registerOutputs_484__15), .inputs_508__12 (registerOutputs_484__15)
            , .inputs_508__11 (registerOutputs_484__15), .inputs_508__10 (
            registerOutputs_484__15), .inputs_508__9 (registerOutputs_484__15), 
            .inputs_508__8 (registerOutputs_484__15), .inputs_508__7 (
            registerOutputs_484__15), .inputs_508__6 (registerOutputs_484__15), 
            .inputs_508__5 (registerOutputs_484__15), .inputs_508__4 (
            registerOutputs_484__15), .inputs_508__3 (registerOutputs_484__15), 
            .inputs_508__2 (registerOutputs_484__15), .inputs_508__1 (
            registerOutputs_484__15), .inputs_508__0 (registerOutputs_484__15), 
            .inputs_509__15 (registerOutputs_484__15), .inputs_509__14 (
            registerOutputs_484__15), .inputs_509__13 (registerOutputs_484__15)
            , .inputs_509__12 (registerOutputs_484__15), .inputs_509__11 (
            registerOutputs_484__15), .inputs_509__10 (registerOutputs_484__15)
            , .inputs_509__9 (registerOutputs_484__15), .inputs_509__8 (
            registerOutputs_484__15), .inputs_509__7 (registerOutputs_484__15), 
            .inputs_509__6 (registerOutputs_484__15), .inputs_509__5 (
            registerOutputs_484__15), .inputs_509__4 (registerOutputs_484__15), 
            .inputs_509__3 (registerOutputs_484__15), .inputs_509__2 (
            registerOutputs_484__15), .inputs_509__1 (registerOutputs_484__15), 
            .inputs_509__0 (registerOutputs_484__15), .inputs_510__15 (
            registerOutputs_484__15), .inputs_510__14 (registerOutputs_484__15)
            , .inputs_510__13 (registerOutputs_484__15), .inputs_510__12 (
            registerOutputs_484__15), .inputs_510__11 (registerOutputs_484__15)
            , .inputs_510__10 (registerOutputs_484__15), .inputs_510__9 (
            registerOutputs_484__15), .inputs_510__8 (registerOutputs_484__15), 
            .inputs_510__7 (registerOutputs_484__15), .inputs_510__6 (
            registerOutputs_484__15), .inputs_510__5 (registerOutputs_484__15), 
            .inputs_510__4 (registerOutputs_484__15), .inputs_510__3 (
            registerOutputs_484__15), .inputs_510__2 (registerOutputs_484__15), 
            .inputs_510__1 (registerOutputs_484__15), .inputs_510__0 (
            registerOutputs_484__15), .inputs_511__15 (registerOutputs_484__15)
            , .inputs_511__14 (registerOutputs_484__15), .inputs_511__13 (
            registerOutputs_484__15), .inputs_511__12 (registerOutputs_484__15)
            , .inputs_511__11 (registerOutputs_484__15), .inputs_511__10 (
            registerOutputs_484__15), .inputs_511__9 (registerOutputs_484__15), 
            .inputs_511__8 (registerOutputs_484__15), .inputs_511__7 (
            registerOutputs_484__15), .inputs_511__6 (registerOutputs_484__15), 
            .inputs_511__5 (registerOutputs_484__15), .inputs_511__4 (
            registerOutputs_484__15), .inputs_511__3 (registerOutputs_484__15), 
            .inputs_511__2 (registerOutputs_484__15), .inputs_511__1 (
            registerOutputs_484__15), .inputs_511__0 (registerOutputs_484__15), 
            .selectionLines ({nx33625,registerSelector_7,nx38155,
            registerSelector_5,registerSelector_4,nx38157,nx33629,
            registerSelector_1,nx33633}), .\output  ({
            selectedRegisterMuxOutput[15],selectedRegisterMuxOutput[14],
            selectedRegisterMuxOutput[13],selectedRegisterMuxOutput[12],
            selectedRegisterMuxOutput[11],selectedRegisterMuxOutput[10],
            selectedRegisterMuxOutput[9],selectedRegisterMuxOutput[8],
            selectedRegisterMuxOutput[7],selectedRegisterMuxOutput[6],
            selectedRegisterMuxOutput[5],selectedRegisterMuxOutput[4],
            selectedRegisterMuxOutput[3],selectedRegisterMuxOutput[2],
            selectedRegisterMuxOutput[1],selectedRegisterMuxOutput[0]})) ;
    Mux2_16 reluMUX (.A ({outToRam_15,outToRam_14,outToRam_13,outToRam_12,
            outToRam_11,outToRam_10,outToRam_9,outToRam_8,outToRam_7,outToRam_6,
            outToRam_5,outToRam_4,outToRam_3,outToRam_2,outToRam_1,outToRam_0})
            , .B ({registerOutputs_484__15,registerOutputs_484__15,
            registerOutputs_484__15,registerOutputs_484__15,
            registerOutputs_484__15,registerOutputs_484__15,
            registerOutputs_484__15,registerOutputs_484__15,
            registerOutputs_484__15,registerOutputs_484__15,
            registerOutputs_484__15,registerOutputs_484__15,
            registerOutputs_484__15,registerOutputs_484__15,
            registerOutputs_484__15,registerOutputs_484__15}), .S (isRelu), .C (
            {reluMuxOutuput_15,reluMuxOutuput_14,reluMuxOutuput_13,
            reluMuxOutuput_12,reluMuxOutuput_11,reluMuxOutuput_10,
            reluMuxOutuput_9,reluMuxOutuput_8,reluMuxOutuput_7,reluMuxOutuput_6,
            reluMuxOutuput_5,reluMuxOutuput_4,reluMuxOutuput_3,reluMuxOutuput_2,
            reluMuxOutuput_1,reluMuxOutuput_0})) ;
    Tristate_16 tristateBuffer (.\input  ({reluMuxOutuput_15,reluMuxOutuput_14,
                reluMuxOutuput_13,reluMuxOutuput_12,reluMuxOutuput_11,
                reluMuxOutuput_10,reluMuxOutuput_9,reluMuxOutuput_8,
                reluMuxOutuput_7,reluMuxOutuput_6,reluMuxOutuput_5,
                reluMuxOutuput_4,reluMuxOutuput_3,reluMuxOutuput_2,
                reluMuxOutuput_1,reluMuxOutuput_0}), .en (tristateEnable), .\output  (
                {writeBus[15],writeBus[14],writeBus[13],writeBus[12],
                writeBus[11],writeBus[10],writeBus[9],writeBus[8],writeBus[7],
                writeBus[6],writeBus[5],writeBus[4],writeBus[3],writeBus[2],
                writeBus[1],writeBus[0]})) ;
    Counter_9 counterSelector (.en (counterEnable), .reset (resetCounter), .clk (
              notClk), .count ({registerSelector_8,registerSelector_7,
              registerSelector_6,registerSelector_5,registerSelector_4,
              registerSelector_3,registerSelector_2,registerSelector_1,
              registerSelector_0})) ;
    Reg_16 outputRegMap (.D ({nx36023,nx36165,nx36307,nx36449,nx36591,nx36733,
           nx36875,nx37017,nx37159,nx37301,nx37443,nx37585,nx37727,nx37869,
           nx38011,nx38153}), .en (enableDecoder), .clk (clk), .rst (
           resetRegisters), .Q ({outToRam_15,outToRam_14,outToRam_13,outToRam_12
           ,outToRam_11,outToRam_10,outToRam_9,outToRam_8,outToRam_7,outToRam_6,
           outToRam_5,outToRam_4,outToRam_3,outToRam_2,outToRam_1,outToRam_0})
           ) ;
    fake_gnd ix32635 (.Y (registerOutputs_484__15)) ;
    nor02ii ix975 (.Y (isRelu), .A0 (isPool), .A1 (outToRam_15)) ;
    or02 ix1 (.Y (resetCounter), .A0 (finishSlice), .A1 (resetRegisters)) ;
    inv01 ix33135 (.Y (notClk), .A (clk)) ;
    or02 ix5 (.Y (enableRegister_0), .A0 (nx35743), .A1 (decoderOutput_0)) ;
    or02 ix7 (.Y (enableRegister_1), .A0 (nx35743), .A1 (decoderOutput_1)) ;
    or02 ix9 (.Y (enableRegister_2), .A0 (nx35743), .A1 (decoderOutput_2)) ;
    or02 ix11 (.Y (enableRegister_3), .A0 (nx35743), .A1 (decoderOutput_3)) ;
    or02 ix13 (.Y (enableRegister_4), .A0 (nx35743), .A1 (decoderOutput_4)) ;
    or02 ix15 (.Y (enableRegister_5), .A0 (nx35743), .A1 (decoderOutput_5)) ;
    or02 ix17 (.Y (enableRegister_6), .A0 (nx35745), .A1 (decoderOutput_6)) ;
    or02 ix19 (.Y (enableRegister_7), .A0 (nx35745), .A1 (decoderOutput_7)) ;
    or02 ix21 (.Y (enableRegister_8), .A0 (nx35745), .A1 (decoderOutput_8)) ;
    or02 ix23 (.Y (enableRegister_9), .A0 (nx35745), .A1 (decoderOutput_9)) ;
    or02 ix25 (.Y (enableRegister_10), .A0 (nx35745), .A1 (decoderOutput_10)) ;
    or02 ix27 (.Y (enableRegister_11), .A0 (nx35745), .A1 (decoderOutput_11)) ;
    or02 ix29 (.Y (enableRegister_12), .A0 (nx35745), .A1 (decoderOutput_12)) ;
    or02 ix31 (.Y (enableRegister_13), .A0 (nx35747), .A1 (decoderOutput_13)) ;
    or02 ix33 (.Y (enableRegister_14), .A0 (nx35747), .A1 (decoderOutput_14)) ;
    or02 ix35 (.Y (enableRegister_15), .A0 (nx35747), .A1 (decoderOutput_15)) ;
    or02 ix37 (.Y (enableRegister_16), .A0 (nx35747), .A1 (decoderOutput_16)) ;
    or02 ix39 (.Y (enableRegister_17), .A0 (nx35747), .A1 (decoderOutput_17)) ;
    or02 ix41 (.Y (enableRegister_18), .A0 (nx35747), .A1 (decoderOutput_18)) ;
    or02 ix43 (.Y (enableRegister_19), .A0 (nx35747), .A1 (decoderOutput_19)) ;
    or02 ix45 (.Y (enableRegister_20), .A0 (nx35749), .A1 (decoderOutput_20)) ;
    or02 ix47 (.Y (enableRegister_21), .A0 (nx35749), .A1 (decoderOutput_21)) ;
    or02 ix49 (.Y (enableRegister_22), .A0 (nx35749), .A1 (decoderOutput_22)) ;
    or02 ix51 (.Y (enableRegister_23), .A0 (nx35749), .A1 (decoderOutput_23)) ;
    or02 ix53 (.Y (enableRegister_24), .A0 (nx35749), .A1 (decoderOutput_24)) ;
    or02 ix55 (.Y (enableRegister_25), .A0 (nx35749), .A1 (decoderOutput_25)) ;
    or02 ix57 (.Y (enableRegister_26), .A0 (nx35749), .A1 (decoderOutput_26)) ;
    or02 ix59 (.Y (enableRegister_27), .A0 (nx35751), .A1 (decoderOutput_27)) ;
    or02 ix61 (.Y (enableRegister_28), .A0 (nx35751), .A1 (decoderOutput_28)) ;
    or02 ix63 (.Y (enableRegister_29), .A0 (nx35751), .A1 (decoderOutput_29)) ;
    or02 ix65 (.Y (enableRegister_30), .A0 (nx35751), .A1 (decoderOutput_30)) ;
    or02 ix67 (.Y (enableRegister_31), .A0 (nx35751), .A1 (decoderOutput_31)) ;
    or02 ix69 (.Y (enableRegister_32), .A0 (nx35751), .A1 (decoderOutput_32)) ;
    or02 ix71 (.Y (enableRegister_33), .A0 (nx35751), .A1 (decoderOutput_33)) ;
    or02 ix73 (.Y (enableRegister_34), .A0 (nx35753), .A1 (decoderOutput_34)) ;
    or02 ix75 (.Y (enableRegister_35), .A0 (nx35753), .A1 (decoderOutput_35)) ;
    or02 ix77 (.Y (enableRegister_36), .A0 (nx35753), .A1 (decoderOutput_36)) ;
    or02 ix79 (.Y (enableRegister_37), .A0 (nx35753), .A1 (decoderOutput_37)) ;
    or02 ix81 (.Y (enableRegister_38), .A0 (nx35753), .A1 (decoderOutput_38)) ;
    or02 ix83 (.Y (enableRegister_39), .A0 (nx35753), .A1 (decoderOutput_39)) ;
    or02 ix85 (.Y (enableRegister_40), .A0 (nx35753), .A1 (decoderOutput_40)) ;
    or02 ix87 (.Y (enableRegister_41), .A0 (nx35755), .A1 (decoderOutput_41)) ;
    or02 ix89 (.Y (enableRegister_42), .A0 (nx35755), .A1 (decoderOutput_42)) ;
    or02 ix91 (.Y (enableRegister_43), .A0 (nx35755), .A1 (decoderOutput_43)) ;
    or02 ix93 (.Y (enableRegister_44), .A0 (nx35755), .A1 (decoderOutput_44)) ;
    or02 ix95 (.Y (enableRegister_45), .A0 (nx35755), .A1 (decoderOutput_45)) ;
    or02 ix97 (.Y (enableRegister_46), .A0 (nx35755), .A1 (decoderOutput_46)) ;
    or02 ix99 (.Y (enableRegister_47), .A0 (nx35755), .A1 (decoderOutput_47)) ;
    or02 ix101 (.Y (enableRegister_48), .A0 (nx35757), .A1 (decoderOutput_48)) ;
    or02 ix103 (.Y (enableRegister_49), .A0 (nx35757), .A1 (decoderOutput_49)) ;
    or02 ix105 (.Y (enableRegister_50), .A0 (nx35757), .A1 (decoderOutput_50)) ;
    or02 ix107 (.Y (enableRegister_51), .A0 (nx35757), .A1 (decoderOutput_51)) ;
    or02 ix109 (.Y (enableRegister_52), .A0 (nx35757), .A1 (decoderOutput_52)) ;
    or02 ix111 (.Y (enableRegister_53), .A0 (nx35757), .A1 (decoderOutput_53)) ;
    or02 ix113 (.Y (enableRegister_54), .A0 (nx35757), .A1 (decoderOutput_54)) ;
    or02 ix115 (.Y (enableRegister_55), .A0 (nx35759), .A1 (decoderOutput_55)) ;
    or02 ix117 (.Y (enableRegister_56), .A0 (nx35759), .A1 (decoderOutput_56)) ;
    or02 ix119 (.Y (enableRegister_57), .A0 (nx35759), .A1 (decoderOutput_57)) ;
    or02 ix121 (.Y (enableRegister_58), .A0 (nx35759), .A1 (decoderOutput_58)) ;
    or02 ix123 (.Y (enableRegister_59), .A0 (nx35759), .A1 (decoderOutput_59)) ;
    or02 ix125 (.Y (enableRegister_60), .A0 (nx35759), .A1 (decoderOutput_60)) ;
    or02 ix127 (.Y (enableRegister_61), .A0 (nx35759), .A1 (decoderOutput_61)) ;
    or02 ix129 (.Y (enableRegister_62), .A0 (nx35761), .A1 (decoderOutput_62)) ;
    or02 ix131 (.Y (enableRegister_63), .A0 (nx35761), .A1 (decoderOutput_63)) ;
    or02 ix133 (.Y (enableRegister_64), .A0 (nx35761), .A1 (decoderOutput_64)) ;
    or02 ix135 (.Y (enableRegister_65), .A0 (nx35761), .A1 (decoderOutput_65)) ;
    or02 ix137 (.Y (enableRegister_66), .A0 (nx35761), .A1 (decoderOutput_66)) ;
    or02 ix139 (.Y (enableRegister_67), .A0 (nx35761), .A1 (decoderOutput_67)) ;
    or02 ix141 (.Y (enableRegister_68), .A0 (nx35761), .A1 (decoderOutput_68)) ;
    or02 ix143 (.Y (enableRegister_69), .A0 (nx35763), .A1 (decoderOutput_69)) ;
    or02 ix145 (.Y (enableRegister_70), .A0 (nx35763), .A1 (decoderOutput_70)) ;
    or02 ix147 (.Y (enableRegister_71), .A0 (nx35763), .A1 (decoderOutput_71)) ;
    or02 ix149 (.Y (enableRegister_72), .A0 (nx35763), .A1 (decoderOutput_72)) ;
    or02 ix151 (.Y (enableRegister_73), .A0 (nx35763), .A1 (decoderOutput_73)) ;
    or02 ix153 (.Y (enableRegister_74), .A0 (nx35763), .A1 (decoderOutput_74)) ;
    or02 ix155 (.Y (enableRegister_75), .A0 (nx35763), .A1 (decoderOutput_75)) ;
    or02 ix157 (.Y (enableRegister_76), .A0 (nx35765), .A1 (decoderOutput_76)) ;
    or02 ix159 (.Y (enableRegister_77), .A0 (nx35765), .A1 (decoderOutput_77)) ;
    or02 ix161 (.Y (enableRegister_78), .A0 (nx35765), .A1 (decoderOutput_78)) ;
    or02 ix163 (.Y (enableRegister_79), .A0 (nx35765), .A1 (decoderOutput_79)) ;
    or02 ix165 (.Y (enableRegister_80), .A0 (nx35765), .A1 (decoderOutput_80)) ;
    or02 ix167 (.Y (enableRegister_81), .A0 (nx35765), .A1 (decoderOutput_81)) ;
    or02 ix169 (.Y (enableRegister_82), .A0 (nx35765), .A1 (decoderOutput_82)) ;
    or02 ix171 (.Y (enableRegister_83), .A0 (nx35767), .A1 (decoderOutput_83)) ;
    or02 ix173 (.Y (enableRegister_84), .A0 (nx35767), .A1 (decoderOutput_84)) ;
    or02 ix175 (.Y (enableRegister_85), .A0 (nx35767), .A1 (decoderOutput_85)) ;
    or02 ix177 (.Y (enableRegister_86), .A0 (nx35767), .A1 (decoderOutput_86)) ;
    or02 ix179 (.Y (enableRegister_87), .A0 (nx35767), .A1 (decoderOutput_87)) ;
    or02 ix181 (.Y (enableRegister_88), .A0 (nx35767), .A1 (decoderOutput_88)) ;
    or02 ix183 (.Y (enableRegister_89), .A0 (nx35767), .A1 (decoderOutput_89)) ;
    or02 ix185 (.Y (enableRegister_90), .A0 (nx35769), .A1 (decoderOutput_90)) ;
    or02 ix187 (.Y (enableRegister_91), .A0 (nx35769), .A1 (decoderOutput_91)) ;
    or02 ix189 (.Y (enableRegister_92), .A0 (nx35769), .A1 (decoderOutput_92)) ;
    or02 ix191 (.Y (enableRegister_93), .A0 (nx35769), .A1 (decoderOutput_93)) ;
    or02 ix193 (.Y (enableRegister_94), .A0 (nx35769), .A1 (decoderOutput_94)) ;
    or02 ix195 (.Y (enableRegister_95), .A0 (nx35769), .A1 (decoderOutput_95)) ;
    or02 ix197 (.Y (enableRegister_96), .A0 (nx35769), .A1 (decoderOutput_96)) ;
    or02 ix199 (.Y (enableRegister_97), .A0 (nx35771), .A1 (decoderOutput_97)) ;
    or02 ix201 (.Y (enableRegister_98), .A0 (nx35771), .A1 (decoderOutput_98)) ;
    or02 ix203 (.Y (enableRegister_99), .A0 (nx35771), .A1 (decoderOutput_99)) ;
    or02 ix205 (.Y (enableRegister_100), .A0 (nx35771), .A1 (decoderOutput_100)
         ) ;
    or02 ix207 (.Y (enableRegister_101), .A0 (nx35771), .A1 (decoderOutput_101)
         ) ;
    or02 ix209 (.Y (enableRegister_102), .A0 (nx35771), .A1 (decoderOutput_102)
         ) ;
    or02 ix211 (.Y (enableRegister_103), .A0 (nx35771), .A1 (decoderOutput_103)
         ) ;
    or02 ix213 (.Y (enableRegister_104), .A0 (nx35773), .A1 (decoderOutput_104)
         ) ;
    or02 ix215 (.Y (enableRegister_105), .A0 (nx35773), .A1 (decoderOutput_105)
         ) ;
    or02 ix217 (.Y (enableRegister_106), .A0 (nx35773), .A1 (decoderOutput_106)
         ) ;
    or02 ix219 (.Y (enableRegister_107), .A0 (nx35773), .A1 (decoderOutput_107)
         ) ;
    or02 ix221 (.Y (enableRegister_108), .A0 (nx35773), .A1 (decoderOutput_108)
         ) ;
    or02 ix223 (.Y (enableRegister_109), .A0 (nx35773), .A1 (decoderOutput_109)
         ) ;
    or02 ix225 (.Y (enableRegister_110), .A0 (nx35773), .A1 (decoderOutput_110)
         ) ;
    or02 ix227 (.Y (enableRegister_111), .A0 (nx35775), .A1 (decoderOutput_111)
         ) ;
    or02 ix229 (.Y (enableRegister_112), .A0 (nx35775), .A1 (decoderOutput_112)
         ) ;
    or02 ix231 (.Y (enableRegister_113), .A0 (nx35775), .A1 (decoderOutput_113)
         ) ;
    or02 ix233 (.Y (enableRegister_114), .A0 (nx35775), .A1 (decoderOutput_114)
         ) ;
    or02 ix235 (.Y (enableRegister_115), .A0 (nx35775), .A1 (decoderOutput_115)
         ) ;
    or02 ix237 (.Y (enableRegister_116), .A0 (nx35775), .A1 (decoderOutput_116)
         ) ;
    or02 ix239 (.Y (enableRegister_117), .A0 (nx35775), .A1 (decoderOutput_117)
         ) ;
    or02 ix241 (.Y (enableRegister_118), .A0 (nx35777), .A1 (decoderOutput_118)
         ) ;
    or02 ix243 (.Y (enableRegister_119), .A0 (nx35777), .A1 (decoderOutput_119)
         ) ;
    or02 ix245 (.Y (enableRegister_120), .A0 (nx35777), .A1 (decoderOutput_120)
         ) ;
    or02 ix247 (.Y (enableRegister_121), .A0 (nx35777), .A1 (decoderOutput_121)
         ) ;
    or02 ix249 (.Y (enableRegister_122), .A0 (nx35777), .A1 (decoderOutput_122)
         ) ;
    or02 ix251 (.Y (enableRegister_123), .A0 (nx35777), .A1 (decoderOutput_123)
         ) ;
    or02 ix253 (.Y (enableRegister_124), .A0 (nx35777), .A1 (decoderOutput_124)
         ) ;
    or02 ix255 (.Y (enableRegister_125), .A0 (nx35779), .A1 (decoderOutput_125)
         ) ;
    or02 ix257 (.Y (enableRegister_126), .A0 (nx35779), .A1 (decoderOutput_126)
         ) ;
    or02 ix259 (.Y (enableRegister_127), .A0 (nx35779), .A1 (decoderOutput_127)
         ) ;
    or02 ix261 (.Y (enableRegister_128), .A0 (nx35779), .A1 (decoderOutput_128)
         ) ;
    or02 ix263 (.Y (enableRegister_129), .A0 (nx35779), .A1 (decoderOutput_129)
         ) ;
    or02 ix265 (.Y (enableRegister_130), .A0 (nx35779), .A1 (decoderOutput_130)
         ) ;
    or02 ix267 (.Y (enableRegister_131), .A0 (nx35779), .A1 (decoderOutput_131)
         ) ;
    or02 ix269 (.Y (enableRegister_132), .A0 (nx35781), .A1 (decoderOutput_132)
         ) ;
    or02 ix271 (.Y (enableRegister_133), .A0 (nx35781), .A1 (decoderOutput_133)
         ) ;
    or02 ix273 (.Y (enableRegister_134), .A0 (nx35781), .A1 (decoderOutput_134)
         ) ;
    or02 ix275 (.Y (enableRegister_135), .A0 (nx35781), .A1 (decoderOutput_135)
         ) ;
    or02 ix277 (.Y (enableRegister_136), .A0 (nx35781), .A1 (decoderOutput_136)
         ) ;
    or02 ix279 (.Y (enableRegister_137), .A0 (nx35781), .A1 (decoderOutput_137)
         ) ;
    or02 ix281 (.Y (enableRegister_138), .A0 (nx35781), .A1 (decoderOutput_138)
         ) ;
    or02 ix283 (.Y (enableRegister_139), .A0 (nx35783), .A1 (decoderOutput_139)
         ) ;
    or02 ix285 (.Y (enableRegister_140), .A0 (nx35783), .A1 (decoderOutput_140)
         ) ;
    or02 ix287 (.Y (enableRegister_141), .A0 (nx35783), .A1 (decoderOutput_141)
         ) ;
    or02 ix289 (.Y (enableRegister_142), .A0 (nx35783), .A1 (decoderOutput_142)
         ) ;
    or02 ix291 (.Y (enableRegister_143), .A0 (nx35783), .A1 (decoderOutput_143)
         ) ;
    or02 ix293 (.Y (enableRegister_144), .A0 (nx35783), .A1 (decoderOutput_144)
         ) ;
    or02 ix295 (.Y (enableRegister_145), .A0 (nx35783), .A1 (decoderOutput_145)
         ) ;
    or02 ix297 (.Y (enableRegister_146), .A0 (nx35785), .A1 (decoderOutput_146)
         ) ;
    or02 ix299 (.Y (enableRegister_147), .A0 (nx35785), .A1 (decoderOutput_147)
         ) ;
    or02 ix301 (.Y (enableRegister_148), .A0 (nx35785), .A1 (decoderOutput_148)
         ) ;
    or02 ix303 (.Y (enableRegister_149), .A0 (nx35785), .A1 (decoderOutput_149)
         ) ;
    or02 ix305 (.Y (enableRegister_150), .A0 (nx35785), .A1 (decoderOutput_150)
         ) ;
    or02 ix307 (.Y (enableRegister_151), .A0 (nx35785), .A1 (decoderOutput_151)
         ) ;
    or02 ix309 (.Y (enableRegister_152), .A0 (nx35785), .A1 (decoderOutput_152)
         ) ;
    or02 ix311 (.Y (enableRegister_153), .A0 (nx35787), .A1 (decoderOutput_153)
         ) ;
    or02 ix313 (.Y (enableRegister_154), .A0 (nx35787), .A1 (decoderOutput_154)
         ) ;
    or02 ix315 (.Y (enableRegister_155), .A0 (nx35787), .A1 (decoderOutput_155)
         ) ;
    or02 ix317 (.Y (enableRegister_156), .A0 (nx35787), .A1 (decoderOutput_156)
         ) ;
    or02 ix319 (.Y (enableRegister_157), .A0 (nx35787), .A1 (decoderOutput_157)
         ) ;
    or02 ix321 (.Y (enableRegister_158), .A0 (nx35787), .A1 (decoderOutput_158)
         ) ;
    or02 ix323 (.Y (enableRegister_159), .A0 (nx35787), .A1 (decoderOutput_159)
         ) ;
    or02 ix325 (.Y (enableRegister_160), .A0 (nx35789), .A1 (decoderOutput_160)
         ) ;
    or02 ix327 (.Y (enableRegister_161), .A0 (nx35789), .A1 (decoderOutput_161)
         ) ;
    or02 ix329 (.Y (enableRegister_162), .A0 (nx35789), .A1 (decoderOutput_162)
         ) ;
    or02 ix331 (.Y (enableRegister_163), .A0 (nx35789), .A1 (decoderOutput_163)
         ) ;
    or02 ix333 (.Y (enableRegister_164), .A0 (nx35789), .A1 (decoderOutput_164)
         ) ;
    or02 ix335 (.Y (enableRegister_165), .A0 (nx35789), .A1 (decoderOutput_165)
         ) ;
    or02 ix337 (.Y (enableRegister_166), .A0 (nx35789), .A1 (decoderOutput_166)
         ) ;
    or02 ix339 (.Y (enableRegister_167), .A0 (nx35791), .A1 (decoderOutput_167)
         ) ;
    or02 ix341 (.Y (enableRegister_168), .A0 (nx35791), .A1 (decoderOutput_168)
         ) ;
    or02 ix343 (.Y (enableRegister_169), .A0 (nx35791), .A1 (decoderOutput_169)
         ) ;
    or02 ix345 (.Y (enableRegister_170), .A0 (nx35791), .A1 (decoderOutput_170)
         ) ;
    or02 ix347 (.Y (enableRegister_171), .A0 (nx35791), .A1 (decoderOutput_171)
         ) ;
    or02 ix349 (.Y (enableRegister_172), .A0 (nx35791), .A1 (decoderOutput_172)
         ) ;
    or02 ix351 (.Y (enableRegister_173), .A0 (nx35791), .A1 (decoderOutput_173)
         ) ;
    or02 ix353 (.Y (enableRegister_174), .A0 (nx35793), .A1 (decoderOutput_174)
         ) ;
    or02 ix355 (.Y (enableRegister_175), .A0 (nx35793), .A1 (decoderOutput_175)
         ) ;
    or02 ix357 (.Y (enableRegister_176), .A0 (nx35793), .A1 (decoderOutput_176)
         ) ;
    or02 ix359 (.Y (enableRegister_177), .A0 (nx35793), .A1 (decoderOutput_177)
         ) ;
    or02 ix361 (.Y (enableRegister_178), .A0 (nx35793), .A1 (decoderOutput_178)
         ) ;
    or02 ix363 (.Y (enableRegister_179), .A0 (nx35793), .A1 (decoderOutput_179)
         ) ;
    or02 ix365 (.Y (enableRegister_180), .A0 (nx35793), .A1 (decoderOutput_180)
         ) ;
    or02 ix367 (.Y (enableRegister_181), .A0 (nx35795), .A1 (decoderOutput_181)
         ) ;
    or02 ix369 (.Y (enableRegister_182), .A0 (nx35795), .A1 (decoderOutput_182)
         ) ;
    or02 ix371 (.Y (enableRegister_183), .A0 (nx35795), .A1 (decoderOutput_183)
         ) ;
    or02 ix373 (.Y (enableRegister_184), .A0 (nx35795), .A1 (decoderOutput_184)
         ) ;
    or02 ix375 (.Y (enableRegister_185), .A0 (nx35795), .A1 (decoderOutput_185)
         ) ;
    or02 ix377 (.Y (enableRegister_186), .A0 (nx35795), .A1 (decoderOutput_186)
         ) ;
    or02 ix379 (.Y (enableRegister_187), .A0 (nx35795), .A1 (decoderOutput_187)
         ) ;
    or02 ix381 (.Y (enableRegister_188), .A0 (nx35797), .A1 (decoderOutput_188)
         ) ;
    or02 ix383 (.Y (enableRegister_189), .A0 (nx35797), .A1 (decoderOutput_189)
         ) ;
    or02 ix385 (.Y (enableRegister_190), .A0 (nx35797), .A1 (decoderOutput_190)
         ) ;
    or02 ix387 (.Y (enableRegister_191), .A0 (nx35797), .A1 (decoderOutput_191)
         ) ;
    or02 ix389 (.Y (enableRegister_192), .A0 (nx35797), .A1 (decoderOutput_192)
         ) ;
    or02 ix391 (.Y (enableRegister_193), .A0 (nx35797), .A1 (decoderOutput_193)
         ) ;
    or02 ix393 (.Y (enableRegister_194), .A0 (nx35797), .A1 (decoderOutput_194)
         ) ;
    or02 ix395 (.Y (enableRegister_195), .A0 (nx35799), .A1 (decoderOutput_195)
         ) ;
    or02 ix397 (.Y (enableRegister_196), .A0 (nx35799), .A1 (decoderOutput_196)
         ) ;
    or02 ix399 (.Y (enableRegister_197), .A0 (nx35799), .A1 (decoderOutput_197)
         ) ;
    or02 ix401 (.Y (enableRegister_198), .A0 (nx35799), .A1 (decoderOutput_198)
         ) ;
    or02 ix403 (.Y (enableRegister_199), .A0 (nx35799), .A1 (decoderOutput_199)
         ) ;
    or02 ix405 (.Y (enableRegister_200), .A0 (nx35799), .A1 (decoderOutput_200)
         ) ;
    or02 ix407 (.Y (enableRegister_201), .A0 (nx35799), .A1 (decoderOutput_201)
         ) ;
    or02 ix409 (.Y (enableRegister_202), .A0 (nx35801), .A1 (decoderOutput_202)
         ) ;
    or02 ix411 (.Y (enableRegister_203), .A0 (nx35801), .A1 (decoderOutput_203)
         ) ;
    or02 ix413 (.Y (enableRegister_204), .A0 (nx35801), .A1 (decoderOutput_204)
         ) ;
    or02 ix415 (.Y (enableRegister_205), .A0 (nx35801), .A1 (decoderOutput_205)
         ) ;
    or02 ix417 (.Y (enableRegister_206), .A0 (nx35801), .A1 (decoderOutput_206)
         ) ;
    or02 ix419 (.Y (enableRegister_207), .A0 (nx35801), .A1 (decoderOutput_207)
         ) ;
    or02 ix421 (.Y (enableRegister_208), .A0 (nx35801), .A1 (decoderOutput_208)
         ) ;
    or02 ix423 (.Y (enableRegister_209), .A0 (nx35803), .A1 (decoderOutput_209)
         ) ;
    or02 ix425 (.Y (enableRegister_210), .A0 (nx35803), .A1 (decoderOutput_210)
         ) ;
    or02 ix427 (.Y (enableRegister_211), .A0 (nx35803), .A1 (decoderOutput_211)
         ) ;
    or02 ix429 (.Y (enableRegister_212), .A0 (nx35803), .A1 (decoderOutput_212)
         ) ;
    or02 ix431 (.Y (enableRegister_213), .A0 (nx35803), .A1 (decoderOutput_213)
         ) ;
    or02 ix433 (.Y (enableRegister_214), .A0 (nx35803), .A1 (decoderOutput_214)
         ) ;
    or02 ix435 (.Y (enableRegister_215), .A0 (nx35803), .A1 (decoderOutput_215)
         ) ;
    or02 ix437 (.Y (enableRegister_216), .A0 (nx35805), .A1 (decoderOutput_216)
         ) ;
    or02 ix439 (.Y (enableRegister_217), .A0 (nx35805), .A1 (decoderOutput_217)
         ) ;
    or02 ix441 (.Y (enableRegister_218), .A0 (nx35805), .A1 (decoderOutput_218)
         ) ;
    or02 ix443 (.Y (enableRegister_219), .A0 (nx35805), .A1 (decoderOutput_219)
         ) ;
    or02 ix445 (.Y (enableRegister_220), .A0 (nx35805), .A1 (decoderOutput_220)
         ) ;
    or02 ix447 (.Y (enableRegister_221), .A0 (nx35805), .A1 (decoderOutput_221)
         ) ;
    or02 ix449 (.Y (enableRegister_222), .A0 (nx35805), .A1 (decoderOutput_222)
         ) ;
    or02 ix451 (.Y (enableRegister_223), .A0 (nx35807), .A1 (decoderOutput_223)
         ) ;
    or02 ix453 (.Y (enableRegister_224), .A0 (nx35807), .A1 (decoderOutput_224)
         ) ;
    or02 ix455 (.Y (enableRegister_225), .A0 (nx35807), .A1 (decoderOutput_225)
         ) ;
    or02 ix457 (.Y (enableRegister_226), .A0 (nx35807), .A1 (decoderOutput_226)
         ) ;
    or02 ix459 (.Y (enableRegister_227), .A0 (nx35807), .A1 (decoderOutput_227)
         ) ;
    or02 ix461 (.Y (enableRegister_228), .A0 (nx35807), .A1 (decoderOutput_228)
         ) ;
    or02 ix463 (.Y (enableRegister_229), .A0 (nx35807), .A1 (decoderOutput_229)
         ) ;
    or02 ix465 (.Y (enableRegister_230), .A0 (nx35809), .A1 (decoderOutput_230)
         ) ;
    or02 ix467 (.Y (enableRegister_231), .A0 (nx35809), .A1 (decoderOutput_231)
         ) ;
    or02 ix469 (.Y (enableRegister_232), .A0 (nx35809), .A1 (decoderOutput_232)
         ) ;
    or02 ix471 (.Y (enableRegister_233), .A0 (nx35809), .A1 (decoderOutput_233)
         ) ;
    or02 ix473 (.Y (enableRegister_234), .A0 (nx35809), .A1 (decoderOutput_234)
         ) ;
    or02 ix475 (.Y (enableRegister_235), .A0 (nx35809), .A1 (decoderOutput_235)
         ) ;
    or02 ix477 (.Y (enableRegister_236), .A0 (nx35809), .A1 (decoderOutput_236)
         ) ;
    or02 ix479 (.Y (enableRegister_237), .A0 (nx35811), .A1 (decoderOutput_237)
         ) ;
    or02 ix481 (.Y (enableRegister_238), .A0 (nx35811), .A1 (decoderOutput_238)
         ) ;
    or02 ix483 (.Y (enableRegister_239), .A0 (nx35811), .A1 (decoderOutput_239)
         ) ;
    or02 ix485 (.Y (enableRegister_240), .A0 (nx35811), .A1 (decoderOutput_240)
         ) ;
    or02 ix487 (.Y (enableRegister_241), .A0 (nx35811), .A1 (decoderOutput_241)
         ) ;
    or02 ix489 (.Y (enableRegister_242), .A0 (nx35811), .A1 (decoderOutput_242)
         ) ;
    or02 ix491 (.Y (enableRegister_243), .A0 (nx35811), .A1 (decoderOutput_243)
         ) ;
    or02 ix493 (.Y (enableRegister_244), .A0 (nx35813), .A1 (decoderOutput_244)
         ) ;
    or02 ix495 (.Y (enableRegister_245), .A0 (nx35813), .A1 (decoderOutput_245)
         ) ;
    or02 ix497 (.Y (enableRegister_246), .A0 (nx35813), .A1 (decoderOutput_246)
         ) ;
    or02 ix499 (.Y (enableRegister_247), .A0 (nx35813), .A1 (decoderOutput_247)
         ) ;
    or02 ix501 (.Y (enableRegister_248), .A0 (nx35813), .A1 (decoderOutput_248)
         ) ;
    or02 ix503 (.Y (enableRegister_249), .A0 (nx35813), .A1 (decoderOutput_249)
         ) ;
    or02 ix505 (.Y (enableRegister_250), .A0 (nx35813), .A1 (decoderOutput_250)
         ) ;
    or02 ix507 (.Y (enableRegister_251), .A0 (nx35815), .A1 (decoderOutput_251)
         ) ;
    or02 ix509 (.Y (enableRegister_252), .A0 (nx35815), .A1 (decoderOutput_252)
         ) ;
    or02 ix511 (.Y (enableRegister_253), .A0 (nx35815), .A1 (decoderOutput_253)
         ) ;
    or02 ix513 (.Y (enableRegister_254), .A0 (nx35815), .A1 (decoderOutput_254)
         ) ;
    or02 ix515 (.Y (enableRegister_255), .A0 (nx35815), .A1 (decoderOutput_255)
         ) ;
    or02 ix517 (.Y (enableRegister_256), .A0 (nx35815), .A1 (decoderOutput_256)
         ) ;
    or02 ix519 (.Y (enableRegister_257), .A0 (nx35815), .A1 (decoderOutput_257)
         ) ;
    or02 ix521 (.Y (enableRegister_258), .A0 (nx35817), .A1 (decoderOutput_258)
         ) ;
    or02 ix523 (.Y (enableRegister_259), .A0 (nx35817), .A1 (decoderOutput_259)
         ) ;
    or02 ix525 (.Y (enableRegister_260), .A0 (nx35817), .A1 (decoderOutput_260)
         ) ;
    or02 ix527 (.Y (enableRegister_261), .A0 (nx35817), .A1 (decoderOutput_261)
         ) ;
    or02 ix529 (.Y (enableRegister_262), .A0 (nx35817), .A1 (decoderOutput_262)
         ) ;
    or02 ix531 (.Y (enableRegister_263), .A0 (nx35817), .A1 (decoderOutput_263)
         ) ;
    or02 ix533 (.Y (enableRegister_264), .A0 (nx35817), .A1 (decoderOutput_264)
         ) ;
    or02 ix535 (.Y (enableRegister_265), .A0 (nx35819), .A1 (decoderOutput_265)
         ) ;
    or02 ix537 (.Y (enableRegister_266), .A0 (nx35819), .A1 (decoderOutput_266)
         ) ;
    or02 ix539 (.Y (enableRegister_267), .A0 (nx35819), .A1 (decoderOutput_267)
         ) ;
    or02 ix541 (.Y (enableRegister_268), .A0 (nx35819), .A1 (decoderOutput_268)
         ) ;
    or02 ix543 (.Y (enableRegister_269), .A0 (nx35819), .A1 (decoderOutput_269)
         ) ;
    or02 ix545 (.Y (enableRegister_270), .A0 (nx35819), .A1 (decoderOutput_270)
         ) ;
    or02 ix547 (.Y (enableRegister_271), .A0 (nx35819), .A1 (decoderOutput_271)
         ) ;
    or02 ix549 (.Y (enableRegister_272), .A0 (nx35821), .A1 (decoderOutput_272)
         ) ;
    or02 ix551 (.Y (enableRegister_273), .A0 (nx35821), .A1 (decoderOutput_273)
         ) ;
    or02 ix553 (.Y (enableRegister_274), .A0 (nx35821), .A1 (decoderOutput_274)
         ) ;
    or02 ix555 (.Y (enableRegister_275), .A0 (nx35821), .A1 (decoderOutput_275)
         ) ;
    or02 ix557 (.Y (enableRegister_276), .A0 (nx35821), .A1 (decoderOutput_276)
         ) ;
    or02 ix559 (.Y (enableRegister_277), .A0 (nx35821), .A1 (decoderOutput_277)
         ) ;
    or02 ix561 (.Y (enableRegister_278), .A0 (nx35821), .A1 (decoderOutput_278)
         ) ;
    or02 ix563 (.Y (enableRegister_279), .A0 (nx35823), .A1 (decoderOutput_279)
         ) ;
    or02 ix565 (.Y (enableRegister_280), .A0 (nx35823), .A1 (decoderOutput_280)
         ) ;
    or02 ix567 (.Y (enableRegister_281), .A0 (nx35823), .A1 (decoderOutput_281)
         ) ;
    or02 ix569 (.Y (enableRegister_282), .A0 (nx35823), .A1 (decoderOutput_282)
         ) ;
    or02 ix571 (.Y (enableRegister_283), .A0 (nx35823), .A1 (decoderOutput_283)
         ) ;
    or02 ix573 (.Y (enableRegister_284), .A0 (nx35823), .A1 (decoderOutput_284)
         ) ;
    or02 ix575 (.Y (enableRegister_285), .A0 (nx35823), .A1 (decoderOutput_285)
         ) ;
    or02 ix577 (.Y (enableRegister_286), .A0 (nx35825), .A1 (decoderOutput_286)
         ) ;
    or02 ix579 (.Y (enableRegister_287), .A0 (nx35825), .A1 (decoderOutput_287)
         ) ;
    or02 ix581 (.Y (enableRegister_288), .A0 (nx35825), .A1 (decoderOutput_288)
         ) ;
    or02 ix583 (.Y (enableRegister_289), .A0 (nx35825), .A1 (decoderOutput_289)
         ) ;
    or02 ix585 (.Y (enableRegister_290), .A0 (nx35825), .A1 (decoderOutput_290)
         ) ;
    or02 ix587 (.Y (enableRegister_291), .A0 (nx35825), .A1 (decoderOutput_291)
         ) ;
    or02 ix589 (.Y (enableRegister_292), .A0 (nx35825), .A1 (decoderOutput_292)
         ) ;
    or02 ix591 (.Y (enableRegister_293), .A0 (nx35827), .A1 (decoderOutput_293)
         ) ;
    or02 ix593 (.Y (enableRegister_294), .A0 (nx35827), .A1 (decoderOutput_294)
         ) ;
    or02 ix595 (.Y (enableRegister_295), .A0 (nx35827), .A1 (decoderOutput_295)
         ) ;
    or02 ix597 (.Y (enableRegister_296), .A0 (nx35827), .A1 (decoderOutput_296)
         ) ;
    or02 ix599 (.Y (enableRegister_297), .A0 (nx35827), .A1 (decoderOutput_297)
         ) ;
    or02 ix601 (.Y (enableRegister_298), .A0 (nx35827), .A1 (decoderOutput_298)
         ) ;
    or02 ix603 (.Y (enableRegister_299), .A0 (nx35827), .A1 (decoderOutput_299)
         ) ;
    or02 ix605 (.Y (enableRegister_300), .A0 (nx35829), .A1 (decoderOutput_300)
         ) ;
    or02 ix607 (.Y (enableRegister_301), .A0 (nx35829), .A1 (decoderOutput_301)
         ) ;
    or02 ix609 (.Y (enableRegister_302), .A0 (nx35829), .A1 (decoderOutput_302)
         ) ;
    or02 ix611 (.Y (enableRegister_303), .A0 (nx35829), .A1 (decoderOutput_303)
         ) ;
    or02 ix613 (.Y (enableRegister_304), .A0 (nx35829), .A1 (decoderOutput_304)
         ) ;
    or02 ix615 (.Y (enableRegister_305), .A0 (nx35829), .A1 (decoderOutput_305)
         ) ;
    or02 ix617 (.Y (enableRegister_306), .A0 (nx35829), .A1 (decoderOutput_306)
         ) ;
    or02 ix619 (.Y (enableRegister_307), .A0 (nx35831), .A1 (decoderOutput_307)
         ) ;
    or02 ix621 (.Y (enableRegister_308), .A0 (nx35831), .A1 (decoderOutput_308)
         ) ;
    or02 ix623 (.Y (enableRegister_309), .A0 (nx35831), .A1 (decoderOutput_309)
         ) ;
    or02 ix625 (.Y (enableRegister_310), .A0 (nx35831), .A1 (decoderOutput_310)
         ) ;
    or02 ix627 (.Y (enableRegister_311), .A0 (nx35831), .A1 (decoderOutput_311)
         ) ;
    or02 ix629 (.Y (enableRegister_312), .A0 (nx35831), .A1 (decoderOutput_312)
         ) ;
    or02 ix631 (.Y (enableRegister_313), .A0 (nx35831), .A1 (decoderOutput_313)
         ) ;
    or02 ix633 (.Y (enableRegister_314), .A0 (nx35833), .A1 (decoderOutput_314)
         ) ;
    or02 ix635 (.Y (enableRegister_315), .A0 (nx35833), .A1 (decoderOutput_315)
         ) ;
    or02 ix637 (.Y (enableRegister_316), .A0 (nx35833), .A1 (decoderOutput_316)
         ) ;
    or02 ix639 (.Y (enableRegister_317), .A0 (nx35833), .A1 (decoderOutput_317)
         ) ;
    or02 ix641 (.Y (enableRegister_318), .A0 (nx35833), .A1 (decoderOutput_318)
         ) ;
    or02 ix643 (.Y (enableRegister_319), .A0 (nx35833), .A1 (decoderOutput_319)
         ) ;
    or02 ix645 (.Y (enableRegister_320), .A0 (nx35833), .A1 (decoderOutput_320)
         ) ;
    or02 ix647 (.Y (enableRegister_321), .A0 (nx35835), .A1 (decoderOutput_321)
         ) ;
    or02 ix649 (.Y (enableRegister_322), .A0 (nx35835), .A1 (decoderOutput_322)
         ) ;
    or02 ix651 (.Y (enableRegister_323), .A0 (nx35835), .A1 (decoderOutput_323)
         ) ;
    or02 ix653 (.Y (enableRegister_324), .A0 (nx35835), .A1 (decoderOutput_324)
         ) ;
    or02 ix655 (.Y (enableRegister_325), .A0 (nx35835), .A1 (decoderOutput_325)
         ) ;
    or02 ix657 (.Y (enableRegister_326), .A0 (nx35835), .A1 (decoderOutput_326)
         ) ;
    or02 ix659 (.Y (enableRegister_327), .A0 (nx35835), .A1 (decoderOutput_327)
         ) ;
    or02 ix661 (.Y (enableRegister_328), .A0 (nx35837), .A1 (decoderOutput_328)
         ) ;
    or02 ix663 (.Y (enableRegister_329), .A0 (nx35837), .A1 (decoderOutput_329)
         ) ;
    or02 ix665 (.Y (enableRegister_330), .A0 (nx35837), .A1 (decoderOutput_330)
         ) ;
    or02 ix667 (.Y (enableRegister_331), .A0 (nx35837), .A1 (decoderOutput_331)
         ) ;
    or02 ix669 (.Y (enableRegister_332), .A0 (nx35837), .A1 (decoderOutput_332)
         ) ;
    or02 ix671 (.Y (enableRegister_333), .A0 (nx35837), .A1 (decoderOutput_333)
         ) ;
    or02 ix673 (.Y (enableRegister_334), .A0 (nx35837), .A1 (decoderOutput_334)
         ) ;
    or02 ix675 (.Y (enableRegister_335), .A0 (nx35839), .A1 (decoderOutput_335)
         ) ;
    or02 ix677 (.Y (enableRegister_336), .A0 (nx35839), .A1 (decoderOutput_336)
         ) ;
    or02 ix679 (.Y (enableRegister_337), .A0 (nx35839), .A1 (decoderOutput_337)
         ) ;
    or02 ix681 (.Y (enableRegister_338), .A0 (nx35839), .A1 (decoderOutput_338)
         ) ;
    or02 ix683 (.Y (enableRegister_339), .A0 (nx35839), .A1 (decoderOutput_339)
         ) ;
    or02 ix685 (.Y (enableRegister_340), .A0 (nx35839), .A1 (decoderOutput_340)
         ) ;
    or02 ix687 (.Y (enableRegister_341), .A0 (nx35839), .A1 (decoderOutput_341)
         ) ;
    or02 ix689 (.Y (enableRegister_342), .A0 (nx35841), .A1 (decoderOutput_342)
         ) ;
    or02 ix691 (.Y (enableRegister_343), .A0 (nx35841), .A1 (decoderOutput_343)
         ) ;
    or02 ix693 (.Y (enableRegister_344), .A0 (nx35841), .A1 (decoderOutput_344)
         ) ;
    or02 ix695 (.Y (enableRegister_345), .A0 (nx35841), .A1 (decoderOutput_345)
         ) ;
    or02 ix697 (.Y (enableRegister_346), .A0 (nx35841), .A1 (decoderOutput_346)
         ) ;
    or02 ix699 (.Y (enableRegister_347), .A0 (nx35841), .A1 (decoderOutput_347)
         ) ;
    or02 ix701 (.Y (enableRegister_348), .A0 (nx35841), .A1 (decoderOutput_348)
         ) ;
    or02 ix703 (.Y (enableRegister_349), .A0 (nx35843), .A1 (decoderOutput_349)
         ) ;
    or02 ix705 (.Y (enableRegister_350), .A0 (nx35843), .A1 (decoderOutput_350)
         ) ;
    or02 ix707 (.Y (enableRegister_351), .A0 (nx35843), .A1 (decoderOutput_351)
         ) ;
    or02 ix709 (.Y (enableRegister_352), .A0 (nx35843), .A1 (decoderOutput_352)
         ) ;
    or02 ix711 (.Y (enableRegister_353), .A0 (nx35843), .A1 (decoderOutput_353)
         ) ;
    or02 ix713 (.Y (enableRegister_354), .A0 (nx35843), .A1 (decoderOutput_354)
         ) ;
    or02 ix715 (.Y (enableRegister_355), .A0 (nx35843), .A1 (decoderOutput_355)
         ) ;
    or02 ix717 (.Y (enableRegister_356), .A0 (nx35845), .A1 (decoderOutput_356)
         ) ;
    or02 ix719 (.Y (enableRegister_357), .A0 (nx35845), .A1 (decoderOutput_357)
         ) ;
    or02 ix721 (.Y (enableRegister_358), .A0 (nx35845), .A1 (decoderOutput_358)
         ) ;
    or02 ix723 (.Y (enableRegister_359), .A0 (nx35845), .A1 (decoderOutput_359)
         ) ;
    or02 ix725 (.Y (enableRegister_360), .A0 (nx35845), .A1 (decoderOutput_360)
         ) ;
    or02 ix727 (.Y (enableRegister_361), .A0 (nx35845), .A1 (decoderOutput_361)
         ) ;
    or02 ix729 (.Y (enableRegister_362), .A0 (nx35845), .A1 (decoderOutput_362)
         ) ;
    or02 ix731 (.Y (enableRegister_363), .A0 (nx35847), .A1 (decoderOutput_363)
         ) ;
    or02 ix733 (.Y (enableRegister_364), .A0 (nx35847), .A1 (decoderOutput_364)
         ) ;
    or02 ix735 (.Y (enableRegister_365), .A0 (nx35847), .A1 (decoderOutput_365)
         ) ;
    or02 ix737 (.Y (enableRegister_366), .A0 (nx35847), .A1 (decoderOutput_366)
         ) ;
    or02 ix739 (.Y (enableRegister_367), .A0 (nx35847), .A1 (decoderOutput_367)
         ) ;
    or02 ix741 (.Y (enableRegister_368), .A0 (nx35847), .A1 (decoderOutput_368)
         ) ;
    or02 ix743 (.Y (enableRegister_369), .A0 (nx35847), .A1 (decoderOutput_369)
         ) ;
    or02 ix745 (.Y (enableRegister_370), .A0 (nx35849), .A1 (decoderOutput_370)
         ) ;
    or02 ix747 (.Y (enableRegister_371), .A0 (nx35849), .A1 (decoderOutput_371)
         ) ;
    or02 ix749 (.Y (enableRegister_372), .A0 (nx35849), .A1 (decoderOutput_372)
         ) ;
    or02 ix751 (.Y (enableRegister_373), .A0 (nx35849), .A1 (decoderOutput_373)
         ) ;
    or02 ix753 (.Y (enableRegister_374), .A0 (nx35849), .A1 (decoderOutput_374)
         ) ;
    or02 ix755 (.Y (enableRegister_375), .A0 (nx35849), .A1 (decoderOutput_375)
         ) ;
    or02 ix757 (.Y (enableRegister_376), .A0 (nx35849), .A1 (decoderOutput_376)
         ) ;
    or02 ix759 (.Y (enableRegister_377), .A0 (nx35851), .A1 (decoderOutput_377)
         ) ;
    or02 ix761 (.Y (enableRegister_378), .A0 (nx35851), .A1 (decoderOutput_378)
         ) ;
    or02 ix763 (.Y (enableRegister_379), .A0 (nx35851), .A1 (decoderOutput_379)
         ) ;
    or02 ix765 (.Y (enableRegister_380), .A0 (nx35851), .A1 (decoderOutput_380)
         ) ;
    or02 ix767 (.Y (enableRegister_381), .A0 (nx35851), .A1 (decoderOutput_381)
         ) ;
    or02 ix769 (.Y (enableRegister_382), .A0 (nx35851), .A1 (decoderOutput_382)
         ) ;
    or02 ix771 (.Y (enableRegister_383), .A0 (nx35851), .A1 (decoderOutput_383)
         ) ;
    or02 ix773 (.Y (enableRegister_384), .A0 (nx35853), .A1 (decoderOutput_384)
         ) ;
    or02 ix775 (.Y (enableRegister_385), .A0 (nx35853), .A1 (decoderOutput_385)
         ) ;
    or02 ix777 (.Y (enableRegister_386), .A0 (nx35853), .A1 (decoderOutput_386)
         ) ;
    or02 ix779 (.Y (enableRegister_387), .A0 (nx35853), .A1 (decoderOutput_387)
         ) ;
    or02 ix781 (.Y (enableRegister_388), .A0 (nx35853), .A1 (decoderOutput_388)
         ) ;
    or02 ix783 (.Y (enableRegister_389), .A0 (nx35853), .A1 (decoderOutput_389)
         ) ;
    or02 ix785 (.Y (enableRegister_390), .A0 (nx35853), .A1 (decoderOutput_390)
         ) ;
    or02 ix787 (.Y (enableRegister_391), .A0 (nx35855), .A1 (decoderOutput_391)
         ) ;
    or02 ix789 (.Y (enableRegister_392), .A0 (nx35855), .A1 (decoderOutput_392)
         ) ;
    or02 ix791 (.Y (enableRegister_393), .A0 (nx35855), .A1 (decoderOutput_393)
         ) ;
    or02 ix793 (.Y (enableRegister_394), .A0 (nx35855), .A1 (decoderOutput_394)
         ) ;
    or02 ix795 (.Y (enableRegister_395), .A0 (nx35855), .A1 (decoderOutput_395)
         ) ;
    or02 ix797 (.Y (enableRegister_396), .A0 (nx35855), .A1 (decoderOutput_396)
         ) ;
    or02 ix799 (.Y (enableRegister_397), .A0 (nx35855), .A1 (decoderOutput_397)
         ) ;
    or02 ix801 (.Y (enableRegister_398), .A0 (nx35857), .A1 (decoderOutput_398)
         ) ;
    or02 ix803 (.Y (enableRegister_399), .A0 (nx35857), .A1 (decoderOutput_399)
         ) ;
    or02 ix805 (.Y (enableRegister_400), .A0 (nx35857), .A1 (decoderOutput_400)
         ) ;
    or02 ix807 (.Y (enableRegister_401), .A0 (nx35857), .A1 (decoderOutput_401)
         ) ;
    or02 ix809 (.Y (enableRegister_402), .A0 (nx35857), .A1 (decoderOutput_402)
         ) ;
    or02 ix811 (.Y (enableRegister_403), .A0 (nx35857), .A1 (decoderOutput_403)
         ) ;
    or02 ix813 (.Y (enableRegister_404), .A0 (nx35857), .A1 (decoderOutput_404)
         ) ;
    or02 ix815 (.Y (enableRegister_405), .A0 (nx35859), .A1 (decoderOutput_405)
         ) ;
    or02 ix817 (.Y (enableRegister_406), .A0 (nx35859), .A1 (decoderOutput_406)
         ) ;
    or02 ix819 (.Y (enableRegister_407), .A0 (nx35859), .A1 (decoderOutput_407)
         ) ;
    or02 ix821 (.Y (enableRegister_408), .A0 (nx35859), .A1 (decoderOutput_408)
         ) ;
    or02 ix823 (.Y (enableRegister_409), .A0 (nx35859), .A1 (decoderOutput_409)
         ) ;
    or02 ix825 (.Y (enableRegister_410), .A0 (nx35859), .A1 (decoderOutput_410)
         ) ;
    or02 ix827 (.Y (enableRegister_411), .A0 (nx35859), .A1 (decoderOutput_411)
         ) ;
    or02 ix829 (.Y (enableRegister_412), .A0 (nx35861), .A1 (decoderOutput_412)
         ) ;
    or02 ix831 (.Y (enableRegister_413), .A0 (nx35861), .A1 (decoderOutput_413)
         ) ;
    or02 ix833 (.Y (enableRegister_414), .A0 (nx35861), .A1 (decoderOutput_414)
         ) ;
    or02 ix835 (.Y (enableRegister_415), .A0 (nx35861), .A1 (decoderOutput_415)
         ) ;
    or02 ix837 (.Y (enableRegister_416), .A0 (nx35861), .A1 (decoderOutput_416)
         ) ;
    or02 ix839 (.Y (enableRegister_417), .A0 (nx35861), .A1 (decoderOutput_417)
         ) ;
    or02 ix841 (.Y (enableRegister_418), .A0 (nx35861), .A1 (decoderOutput_418)
         ) ;
    or02 ix843 (.Y (enableRegister_419), .A0 (nx35863), .A1 (decoderOutput_419)
         ) ;
    or02 ix845 (.Y (enableRegister_420), .A0 (nx35863), .A1 (decoderOutput_420)
         ) ;
    or02 ix847 (.Y (enableRegister_421), .A0 (nx35863), .A1 (decoderOutput_421)
         ) ;
    or02 ix849 (.Y (enableRegister_422), .A0 (nx35863), .A1 (decoderOutput_422)
         ) ;
    or02 ix851 (.Y (enableRegister_423), .A0 (nx35863), .A1 (decoderOutput_423)
         ) ;
    or02 ix853 (.Y (enableRegister_424), .A0 (nx35863), .A1 (decoderOutput_424)
         ) ;
    or02 ix855 (.Y (enableRegister_425), .A0 (nx35863), .A1 (decoderOutput_425)
         ) ;
    or02 ix857 (.Y (enableRegister_426), .A0 (nx35865), .A1 (decoderOutput_426)
         ) ;
    or02 ix859 (.Y (enableRegister_427), .A0 (nx35865), .A1 (decoderOutput_427)
         ) ;
    or02 ix861 (.Y (enableRegister_428), .A0 (nx35865), .A1 (decoderOutput_428)
         ) ;
    or02 ix863 (.Y (enableRegister_429), .A0 (nx35865), .A1 (decoderOutput_429)
         ) ;
    or02 ix865 (.Y (enableRegister_430), .A0 (nx35865), .A1 (decoderOutput_430)
         ) ;
    or02 ix867 (.Y (enableRegister_431), .A0 (nx35865), .A1 (decoderOutput_431)
         ) ;
    or02 ix869 (.Y (enableRegister_432), .A0 (nx35865), .A1 (decoderOutput_432)
         ) ;
    or02 ix871 (.Y (enableRegister_433), .A0 (nx35867), .A1 (decoderOutput_433)
         ) ;
    or02 ix873 (.Y (enableRegister_434), .A0 (nx35867), .A1 (decoderOutput_434)
         ) ;
    or02 ix875 (.Y (enableRegister_435), .A0 (nx35867), .A1 (decoderOutput_435)
         ) ;
    or02 ix877 (.Y (enableRegister_436), .A0 (nx35867), .A1 (decoderOutput_436)
         ) ;
    or02 ix879 (.Y (enableRegister_437), .A0 (nx35867), .A1 (decoderOutput_437)
         ) ;
    or02 ix881 (.Y (enableRegister_438), .A0 (nx35867), .A1 (decoderOutput_438)
         ) ;
    or02 ix883 (.Y (enableRegister_439), .A0 (nx35867), .A1 (decoderOutput_439)
         ) ;
    or02 ix885 (.Y (enableRegister_440), .A0 (nx35869), .A1 (decoderOutput_440)
         ) ;
    or02 ix887 (.Y (enableRegister_441), .A0 (nx35869), .A1 (decoderOutput_441)
         ) ;
    or02 ix889 (.Y (enableRegister_442), .A0 (nx35869), .A1 (decoderOutput_442)
         ) ;
    or02 ix891 (.Y (enableRegister_443), .A0 (nx35869), .A1 (decoderOutput_443)
         ) ;
    or02 ix893 (.Y (enableRegister_444), .A0 (nx35869), .A1 (decoderOutput_444)
         ) ;
    or02 ix895 (.Y (enableRegister_445), .A0 (nx35869), .A1 (decoderOutput_445)
         ) ;
    or02 ix897 (.Y (enableRegister_446), .A0 (nx35869), .A1 (decoderOutput_446)
         ) ;
    or02 ix899 (.Y (enableRegister_447), .A0 (nx35871), .A1 (decoderOutput_447)
         ) ;
    or02 ix901 (.Y (enableRegister_448), .A0 (nx35871), .A1 (decoderOutput_448)
         ) ;
    or02 ix903 (.Y (enableRegister_449), .A0 (nx35871), .A1 (decoderOutput_449)
         ) ;
    or02 ix905 (.Y (enableRegister_450), .A0 (nx35871), .A1 (decoderOutput_450)
         ) ;
    or02 ix907 (.Y (enableRegister_451), .A0 (nx35871), .A1 (decoderOutput_451)
         ) ;
    or02 ix909 (.Y (enableRegister_452), .A0 (nx35871), .A1 (decoderOutput_452)
         ) ;
    or02 ix911 (.Y (enableRegister_453), .A0 (nx35871), .A1 (decoderOutput_453)
         ) ;
    or02 ix913 (.Y (enableRegister_454), .A0 (nx35873), .A1 (decoderOutput_454)
         ) ;
    or02 ix915 (.Y (enableRegister_455), .A0 (nx35873), .A1 (decoderOutput_455)
         ) ;
    or02 ix917 (.Y (enableRegister_456), .A0 (nx35873), .A1 (decoderOutput_456)
         ) ;
    or02 ix919 (.Y (enableRegister_457), .A0 (nx35873), .A1 (decoderOutput_457)
         ) ;
    or02 ix921 (.Y (enableRegister_458), .A0 (nx35873), .A1 (decoderOutput_458)
         ) ;
    or02 ix923 (.Y (enableRegister_459), .A0 (nx35873), .A1 (decoderOutput_459)
         ) ;
    or02 ix925 (.Y (enableRegister_460), .A0 (nx35873), .A1 (decoderOutput_460)
         ) ;
    or02 ix927 (.Y (enableRegister_461), .A0 (nx35875), .A1 (decoderOutput_461)
         ) ;
    or02 ix929 (.Y (enableRegister_462), .A0 (nx35875), .A1 (decoderOutput_462)
         ) ;
    or02 ix931 (.Y (enableRegister_463), .A0 (nx35875), .A1 (decoderOutput_463)
         ) ;
    or02 ix933 (.Y (enableRegister_464), .A0 (nx35875), .A1 (decoderOutput_464)
         ) ;
    or02 ix935 (.Y (enableRegister_465), .A0 (nx35875), .A1 (decoderOutput_465)
         ) ;
    or02 ix937 (.Y (enableRegister_466), .A0 (nx35875), .A1 (decoderOutput_466)
         ) ;
    or02 ix939 (.Y (enableRegister_467), .A0 (nx35875), .A1 (decoderOutput_467)
         ) ;
    or02 ix941 (.Y (enableRegister_468), .A0 (nx35877), .A1 (decoderOutput_468)
         ) ;
    or02 ix943 (.Y (enableRegister_469), .A0 (nx35877), .A1 (decoderOutput_469)
         ) ;
    or02 ix945 (.Y (enableRegister_470), .A0 (nx35877), .A1 (decoderOutput_470)
         ) ;
    or02 ix947 (.Y (enableRegister_471), .A0 (nx35877), .A1 (decoderOutput_471)
         ) ;
    or02 ix949 (.Y (enableRegister_472), .A0 (nx35877), .A1 (decoderOutput_472)
         ) ;
    or02 ix951 (.Y (enableRegister_473), .A0 (nx35877), .A1 (decoderOutput_473)
         ) ;
    or02 ix953 (.Y (enableRegister_474), .A0 (nx35877), .A1 (decoderOutput_474)
         ) ;
    or02 ix955 (.Y (enableRegister_475), .A0 (nx35879), .A1 (decoderOutput_475)
         ) ;
    or02 ix957 (.Y (enableRegister_476), .A0 (nx35879), .A1 (decoderOutput_476)
         ) ;
    or02 ix959 (.Y (enableRegister_477), .A0 (nx35879), .A1 (decoderOutput_477)
         ) ;
    or02 ix961 (.Y (enableRegister_478), .A0 (nx35879), .A1 (decoderOutput_478)
         ) ;
    or02 ix963 (.Y (enableRegister_479), .A0 (nx35879), .A1 (decoderOutput_479)
         ) ;
    or02 ix965 (.Y (enableRegister_480), .A0 (nx35879), .A1 (decoderOutput_480)
         ) ;
    or02 ix967 (.Y (enableRegister_481), .A0 (nx35879), .A1 (decoderOutput_481)
         ) ;
    or02 ix969 (.Y (enableRegister_482), .A0 (nx35881), .A1 (decoderOutput_482)
         ) ;
    or02 ix971 (.Y (enableRegister_483), .A0 (decoderOutput_483), .A1 (nx35881)
         ) ;
    buf02 ix33624 (.Y (nx33625), .A (registerSelector_8)) ;
    buf02 ix33626 (.Y (nx33627), .A (registerSelector_2)) ;
    buf02 ix33628 (.Y (nx33629), .A (registerSelector_2)) ;
    buf02 ix33630 (.Y (nx33631), .A (registerSelector_0)) ;
    buf02 ix33632 (.Y (nx33633), .A (registerSelector_0)) ;
    inv01 ix33638 (.Y (nx33639), .A (weightsBus[7])) ;
    inv01 ix33640 (.Y (nx33641), .A (nx38159)) ;
    inv01 ix33642 (.Y (nx33643), .A (nx38159)) ;
    inv01 ix33644 (.Y (nx33645), .A (nx38159)) ;
    inv01 ix33646 (.Y (nx33647), .A (nx38159)) ;
    inv01 ix33648 (.Y (nx33649), .A (nx38159)) ;
    inv01 ix33650 (.Y (nx33651), .A (nx38159)) ;
    inv01 ix33652 (.Y (nx33653), .A (nx38159)) ;
    inv01 ix33654 (.Y (nx33655), .A (nx38161)) ;
    inv01 ix33656 (.Y (nx33657), .A (nx38161)) ;
    inv01 ix33658 (.Y (nx33659), .A (nx38161)) ;
    inv01 ix33660 (.Y (nx33661), .A (nx38161)) ;
    inv01 ix33662 (.Y (nx33663), .A (nx38161)) ;
    inv01 ix33664 (.Y (nx33665), .A (nx38161)) ;
    inv01 ix33666 (.Y (nx33667), .A (nx38161)) ;
    inv01 ix33668 (.Y (nx33669), .A (nx38163)) ;
    inv01 ix33670 (.Y (nx33671), .A (nx38163)) ;
    inv01 ix33672 (.Y (nx33673), .A (nx38163)) ;
    inv01 ix33674 (.Y (nx33675), .A (nx38163)) ;
    inv01 ix33676 (.Y (nx33677), .A (nx38163)) ;
    inv01 ix33678 (.Y (nx33679), .A (nx38163)) ;
    inv01 ix33680 (.Y (nx33681), .A (nx38163)) ;
    inv01 ix33682 (.Y (nx33683), .A (nx38165)) ;
    inv01 ix33684 (.Y (nx33685), .A (nx38165)) ;
    inv01 ix33686 (.Y (nx33687), .A (nx38165)) ;
    inv01 ix33688 (.Y (nx33689), .A (nx38165)) ;
    inv01 ix33690 (.Y (nx33691), .A (nx38165)) ;
    inv01 ix33692 (.Y (nx33693), .A (nx38165)) ;
    inv01 ix33694 (.Y (nx33695), .A (nx38165)) ;
    inv01 ix33696 (.Y (nx33697), .A (nx38167)) ;
    inv01 ix33698 (.Y (nx33699), .A (nx38167)) ;
    inv01 ix33700 (.Y (nx33701), .A (nx38167)) ;
    inv01 ix33702 (.Y (nx33703), .A (nx38167)) ;
    inv01 ix33704 (.Y (nx33705), .A (nx38167)) ;
    inv01 ix33706 (.Y (nx33707), .A (nx38167)) ;
    inv01 ix33708 (.Y (nx33709), .A (nx38167)) ;
    inv01 ix33710 (.Y (nx33711), .A (nx38169)) ;
    inv01 ix33712 (.Y (nx33713), .A (nx38169)) ;
    inv01 ix33714 (.Y (nx33715), .A (nx38169)) ;
    inv01 ix33716 (.Y (nx33717), .A (nx38169)) ;
    inv01 ix33718 (.Y (nx33719), .A (nx38169)) ;
    inv01 ix33720 (.Y (nx33721), .A (nx38169)) ;
    inv01 ix33722 (.Y (nx33723), .A (nx38169)) ;
    inv01 ix33724 (.Y (nx33725), .A (nx38171)) ;
    inv01 ix33726 (.Y (nx33727), .A (nx38171)) ;
    inv01 ix33728 (.Y (nx33729), .A (nx38171)) ;
    inv01 ix33730 (.Y (nx33731), .A (nx38171)) ;
    inv01 ix33732 (.Y (nx33733), .A (nx38171)) ;
    inv01 ix33734 (.Y (nx33735), .A (nx38171)) ;
    inv01 ix33736 (.Y (nx33737), .A (nx38171)) ;
    inv01 ix33738 (.Y (nx33739), .A (nx38173)) ;
    inv01 ix33740 (.Y (nx33741), .A (nx38173)) ;
    inv01 ix33742 (.Y (nx33743), .A (nx38173)) ;
    inv01 ix33744 (.Y (nx33745), .A (nx38173)) ;
    inv01 ix33746 (.Y (nx33747), .A (nx38173)) ;
    inv01 ix33748 (.Y (nx33749), .A (nx38173)) ;
    inv01 ix33750 (.Y (nx33751), .A (nx38173)) ;
    inv01 ix33752 (.Y (nx33753), .A (nx38175)) ;
    inv01 ix33754 (.Y (nx33755), .A (nx38175)) ;
    inv01 ix33756 (.Y (nx33757), .A (nx38175)) ;
    inv01 ix33758 (.Y (nx33759), .A (nx38175)) ;
    inv01 ix33760 (.Y (nx33761), .A (nx38175)) ;
    inv01 ix33762 (.Y (nx33763), .A (nx38175)) ;
    inv01 ix33764 (.Y (nx33765), .A (nx38175)) ;
    inv01 ix33766 (.Y (nx33767), .A (nx38177)) ;
    inv01 ix33768 (.Y (nx33769), .A (nx38177)) ;
    inv01 ix33770 (.Y (nx33771), .A (nx38177)) ;
    inv01 ix33772 (.Y (nx33773), .A (nx38177)) ;
    inv01 ix33774 (.Y (nx33775), .A (nx38177)) ;
    inv01 ix33776 (.Y (nx33777), .A (nx38177)) ;
    inv01 ix33778 (.Y (nx33779), .A (nx38177)) ;
    inv01 ix33780 (.Y (nx33781), .A (nx38179)) ;
    inv01 ix33782 (.Y (nx33783), .A (nx38179)) ;
    inv01 ix33784 (.Y (nx33785), .A (nx38179)) ;
    inv01 ix33786 (.Y (nx33787), .A (nx38179)) ;
    inv01 ix33788 (.Y (nx33789), .A (nx38179)) ;
    inv01 ix33790 (.Y (nx33791), .A (nx38179)) ;
    inv01 ix33792 (.Y (nx33793), .A (nx38179)) ;
    inv01 ix33794 (.Y (nx33795), .A (nx38181)) ;
    inv01 ix33796 (.Y (nx33797), .A (nx38181)) ;
    inv01 ix33798 (.Y (nx33799), .A (nx38181)) ;
    inv01 ix33800 (.Y (nx33801), .A (nx38181)) ;
    inv01 ix33802 (.Y (nx33803), .A (nx38181)) ;
    inv01 ix33804 (.Y (nx33805), .A (nx38181)) ;
    inv01 ix33806 (.Y (nx33807), .A (nx38181)) ;
    inv01 ix33808 (.Y (nx33809), .A (nx38183)) ;
    inv01 ix33810 (.Y (nx33811), .A (nx38183)) ;
    inv01 ix33812 (.Y (nx33813), .A (nx38183)) ;
    inv01 ix33814 (.Y (nx33815), .A (nx38183)) ;
    inv01 ix33816 (.Y (nx33817), .A (nx38183)) ;
    inv01 ix33818 (.Y (nx33819), .A (nx38183)) ;
    inv01 ix33820 (.Y (nx33821), .A (nx38183)) ;
    inv01 ix33822 (.Y (nx33823), .A (nx38185)) ;
    inv01 ix33824 (.Y (nx33825), .A (nx38185)) ;
    inv01 ix33826 (.Y (nx33827), .A (nx38185)) ;
    inv01 ix33828 (.Y (nx33829), .A (nx38185)) ;
    inv01 ix33830 (.Y (nx33831), .A (nx38185)) ;
    inv01 ix33832 (.Y (nx33833), .A (nx38185)) ;
    inv01 ix33834 (.Y (nx33835), .A (nx38185)) ;
    inv01 ix33836 (.Y (nx33837), .A (nx38187)) ;
    inv01 ix33838 (.Y (nx33839), .A (nx38187)) ;
    inv01 ix33840 (.Y (nx33841), .A (nx38187)) ;
    inv01 ix33842 (.Y (nx33843), .A (nx38187)) ;
    inv01 ix33844 (.Y (nx33845), .A (nx38187)) ;
    inv01 ix33846 (.Y (nx33847), .A (nx38187)) ;
    inv01 ix33848 (.Y (nx33849), .A (nx38187)) ;
    inv01 ix33850 (.Y (nx33851), .A (nx38189)) ;
    inv01 ix33852 (.Y (nx33853), .A (nx38189)) ;
    inv01 ix33854 (.Y (nx33855), .A (nx38189)) ;
    inv01 ix33856 (.Y (nx33857), .A (nx38189)) ;
    inv01 ix33858 (.Y (nx33859), .A (nx38189)) ;
    inv01 ix33860 (.Y (nx33861), .A (nx38189)) ;
    inv01 ix33862 (.Y (nx33863), .A (nx38189)) ;
    inv01 ix33864 (.Y (nx33865), .A (nx38191)) ;
    inv01 ix33866 (.Y (nx33867), .A (nx38191)) ;
    inv01 ix33868 (.Y (nx33869), .A (nx38191)) ;
    inv01 ix33870 (.Y (nx33871), .A (nx38191)) ;
    inv01 ix33872 (.Y (nx33873), .A (nx38191)) ;
    inv01 ix33874 (.Y (nx33875), .A (nx38191)) ;
    inv01 ix33876 (.Y (nx33877), .A (nx38191)) ;
    inv01 ix33878 (.Y (nx33879), .A (nx38193)) ;
    inv01 ix33880 (.Y (nx33881), .A (nx38193)) ;
    inv01 ix33882 (.Y (nx33883), .A (nx38193)) ;
    inv01 ix33884 (.Y (nx33885), .A (nx38193)) ;
    inv01 ix33886 (.Y (nx33887), .A (nx38193)) ;
    inv01 ix33888 (.Y (nx33889), .A (nx38193)) ;
    inv01 ix33890 (.Y (nx33891), .A (nx38193)) ;
    inv01 ix33892 (.Y (nx33893), .A (nx38195)) ;
    inv01 ix33894 (.Y (nx33895), .A (nx38195)) ;
    inv01 ix33896 (.Y (nx33897), .A (nx38195)) ;
    inv01 ix33898 (.Y (nx33899), .A (nx38195)) ;
    inv01 ix33900 (.Y (nx33901), .A (nx38195)) ;
    inv01 ix33902 (.Y (nx33903), .A (nx38195)) ;
    inv01 ix33904 (.Y (nx33905), .A (nx38195)) ;
    inv01 ix33906 (.Y (nx33907), .A (nx38197)) ;
    inv01 ix33908 (.Y (nx33909), .A (nx38197)) ;
    inv01 ix33910 (.Y (nx33911), .A (nx38197)) ;
    inv01 ix33912 (.Y (nx33913), .A (nx38197)) ;
    inv01 ix33914 (.Y (nx33915), .A (nx38197)) ;
    inv01 ix33916 (.Y (nx33917), .A (nx38197)) ;
    inv01 ix33918 (.Y (nx33919), .A (nx38197)) ;
    inv01 ix33920 (.Y (nx33921), .A (nx38199)) ;
    inv01 ix33922 (.Y (nx33923), .A (nx38199)) ;
    inv01 ix33924 (.Y (nx33925), .A (nx38199)) ;
    inv01 ix33926 (.Y (nx33927), .A (nx38199)) ;
    inv01 ix33928 (.Y (nx33929), .A (nx38199)) ;
    inv01 ix33930 (.Y (nx33931), .A (nx38199)) ;
    inv01 ix33932 (.Y (nx33933), .A (nx38199)) ;
    inv01 ix33934 (.Y (nx33935), .A (nx38201)) ;
    inv01 ix33936 (.Y (nx33937), .A (nx38201)) ;
    inv01 ix33938 (.Y (nx33939), .A (nx38201)) ;
    inv01 ix33940 (.Y (nx33941), .A (nx38201)) ;
    inv01 ix33942 (.Y (nx33943), .A (nx38201)) ;
    inv01 ix33944 (.Y (nx33945), .A (nx38201)) ;
    inv01 ix33946 (.Y (nx33947), .A (nx38201)) ;
    inv01 ix33948 (.Y (nx33949), .A (nx38203)) ;
    inv01 ix33950 (.Y (nx33951), .A (nx38203)) ;
    inv01 ix33952 (.Y (nx33953), .A (nx38203)) ;
    inv01 ix33954 (.Y (nx33955), .A (nx38203)) ;
    inv01 ix33956 (.Y (nx33957), .A (nx38203)) ;
    inv01 ix33958 (.Y (nx33959), .A (nx38203)) ;
    inv01 ix33960 (.Y (nx33961), .A (nx38203)) ;
    inv01 ix33962 (.Y (nx33963), .A (nx38205)) ;
    inv01 ix33964 (.Y (nx33965), .A (nx38205)) ;
    inv01 ix33966 (.Y (nx33967), .A (nx38205)) ;
    inv01 ix33968 (.Y (nx33969), .A (nx38205)) ;
    inv01 ix33970 (.Y (nx33971), .A (nx38205)) ;
    inv01 ix33972 (.Y (nx33973), .A (nx38205)) ;
    inv01 ix33974 (.Y (nx33975), .A (nx38205)) ;
    inv01 ix33976 (.Y (nx33977), .A (nx38207)) ;
    inv01 ix33978 (.Y (nx33979), .A (nx38207)) ;
    inv01 ix33980 (.Y (nx33981), .A (nx38207)) ;
    inv01 ix33982 (.Y (nx33983), .A (nx38207)) ;
    inv01 ix33984 (.Y (nx33985), .A (nx38207)) ;
    inv01 ix33986 (.Y (nx33987), .A (nx38207)) ;
    inv01 ix33988 (.Y (nx33989), .A (nx38207)) ;
    inv01 ix33990 (.Y (nx33991), .A (nx38209)) ;
    inv01 ix33992 (.Y (nx33993), .A (nx38209)) ;
    inv01 ix33994 (.Y (nx33995), .A (nx38209)) ;
    inv01 ix33996 (.Y (nx33997), .A (nx38209)) ;
    inv01 ix33998 (.Y (nx33999), .A (nx38209)) ;
    inv01 ix34000 (.Y (nx34001), .A (nx38209)) ;
    inv01 ix34002 (.Y (nx34003), .A (nx38209)) ;
    inv01 ix34004 (.Y (nx34005), .A (nx38211)) ;
    inv01 ix34006 (.Y (nx34007), .A (nx38211)) ;
    inv01 ix34008 (.Y (nx34009), .A (nx38211)) ;
    inv01 ix34010 (.Y (nx34011), .A (nx38211)) ;
    inv01 ix34012 (.Y (nx34013), .A (nx38211)) ;
    inv01 ix34014 (.Y (nx34015), .A (nx38211)) ;
    inv01 ix34016 (.Y (nx34017), .A (nx38211)) ;
    inv01 ix34018 (.Y (nx34019), .A (nx38213)) ;
    inv01 ix34020 (.Y (nx34021), .A (nx38213)) ;
    inv01 ix34022 (.Y (nx34023), .A (nx38213)) ;
    inv01 ix34024 (.Y (nx34025), .A (nx38213)) ;
    inv01 ix34026 (.Y (nx34027), .A (nx38213)) ;
    inv01 ix34028 (.Y (nx34029), .A (nx38213)) ;
    inv01 ix34030 (.Y (nx34031), .A (nx38213)) ;
    inv01 ix34032 (.Y (nx34033), .A (nx38215)) ;
    inv01 ix34034 (.Y (nx34035), .A (nx38215)) ;
    inv01 ix34036 (.Y (nx34037), .A (nx38215)) ;
    inv01 ix34038 (.Y (nx34039), .A (nx38215)) ;
    inv01 ix34040 (.Y (nx34041), .A (nx38215)) ;
    inv01 ix34042 (.Y (nx34043), .A (nx38215)) ;
    inv01 ix34044 (.Y (nx34045), .A (nx38215)) ;
    inv01 ix34046 (.Y (nx34047), .A (nx38217)) ;
    inv01 ix34048 (.Y (nx34049), .A (nx38217)) ;
    inv01 ix34050 (.Y (nx34051), .A (nx38217)) ;
    inv01 ix34052 (.Y (nx34053), .A (nx38217)) ;
    inv01 ix34054 (.Y (nx34055), .A (nx38217)) ;
    inv01 ix34056 (.Y (nx34057), .A (nx38217)) ;
    inv01 ix34058 (.Y (nx34059), .A (nx38217)) ;
    inv01 ix34060 (.Y (nx34061), .A (nx38219)) ;
    inv01 ix34062 (.Y (nx34063), .A (nx38219)) ;
    inv01 ix34064 (.Y (nx34065), .A (nx38219)) ;
    inv01 ix34066 (.Y (nx34067), .A (nx38219)) ;
    inv01 ix34068 (.Y (nx34069), .A (nx38219)) ;
    inv01 ix34070 (.Y (nx34071), .A (nx38219)) ;
    inv01 ix34072 (.Y (nx34073), .A (nx38219)) ;
    inv01 ix34074 (.Y (nx34075), .A (nx38221)) ;
    inv01 ix34076 (.Y (nx34077), .A (nx38221)) ;
    inv01 ix34078 (.Y (nx34079), .A (nx38221)) ;
    inv01 ix34080 (.Y (nx34081), .A (nx38221)) ;
    inv01 ix34082 (.Y (nx34083), .A (nx38221)) ;
    inv01 ix34084 (.Y (nx34085), .A (nx38221)) ;
    inv01 ix34086 (.Y (nx34087), .A (nx38221)) ;
    inv01 ix34088 (.Y (nx34089), .A (nx38223)) ;
    inv01 ix34090 (.Y (nx34091), .A (nx38223)) ;
    inv01 ix34092 (.Y (nx34093), .A (nx38223)) ;
    inv01 ix34094 (.Y (nx34095), .A (nx38223)) ;
    inv01 ix34096 (.Y (nx34097), .A (nx38223)) ;
    inv01 ix34098 (.Y (nx34099), .A (nx38223)) ;
    inv01 ix34100 (.Y (nx34101), .A (nx38223)) ;
    inv01 ix34102 (.Y (nx34103), .A (nx38225)) ;
    inv01 ix34104 (.Y (nx34105), .A (nx38225)) ;
    inv01 ix34106 (.Y (nx34107), .A (nx38225)) ;
    inv01 ix34108 (.Y (nx34109), .A (nx38225)) ;
    inv01 ix34110 (.Y (nx34111), .A (nx38225)) ;
    inv01 ix34112 (.Y (nx34113), .A (nx38225)) ;
    inv01 ix34114 (.Y (nx34115), .A (nx38225)) ;
    inv01 ix34116 (.Y (nx34117), .A (nx38227)) ;
    inv01 ix34118 (.Y (nx34119), .A (nx38227)) ;
    inv01 ix34120 (.Y (nx34121), .A (nx38227)) ;
    inv01 ix34122 (.Y (nx34123), .A (nx38227)) ;
    inv01 ix34124 (.Y (nx34125), .A (nx38227)) ;
    inv01 ix34126 (.Y (nx34127), .A (nx38227)) ;
    inv01 ix34128 (.Y (nx34129), .A (nx38227)) ;
    inv01 ix34130 (.Y (nx34131), .A (nx38229)) ;
    inv01 ix34132 (.Y (nx34133), .A (nx38229)) ;
    inv01 ix34134 (.Y (nx34135), .A (nx38229)) ;
    inv01 ix34136 (.Y (nx34137), .A (nx38229)) ;
    inv01 ix34138 (.Y (nx34139), .A (nx38229)) ;
    inv01 ix34140 (.Y (nx34141), .A (nx38229)) ;
    inv01 ix34142 (.Y (nx34143), .A (nx38229)) ;
    inv01 ix34144 (.Y (nx34145), .A (nx38231)) ;
    inv01 ix34146 (.Y (nx34147), .A (nx38231)) ;
    inv01 ix34148 (.Y (nx34149), .A (nx38231)) ;
    inv01 ix34150 (.Y (nx34151), .A (nx38231)) ;
    inv01 ix34152 (.Y (nx34153), .A (nx38231)) ;
    inv01 ix34154 (.Y (nx34155), .A (nx38231)) ;
    inv01 ix34156 (.Y (nx34157), .A (nx38231)) ;
    inv01 ix34158 (.Y (nx34159), .A (nx38233)) ;
    inv01 ix34160 (.Y (nx34161), .A (nx38233)) ;
    inv01 ix34162 (.Y (nx34163), .A (nx38233)) ;
    inv01 ix34164 (.Y (nx34165), .A (nx38233)) ;
    inv01 ix34166 (.Y (nx34167), .A (nx38233)) ;
    inv01 ix34168 (.Y (nx34169), .A (nx38233)) ;
    inv01 ix34170 (.Y (nx34171), .A (nx38233)) ;
    inv01 ix34172 (.Y (nx34173), .A (nx38235)) ;
    inv01 ix34174 (.Y (nx34175), .A (nx38235)) ;
    inv01 ix34176 (.Y (nx34177), .A (nx38235)) ;
    inv01 ix34178 (.Y (nx34179), .A (nx38235)) ;
    inv01 ix34180 (.Y (nx34181), .A (nx38235)) ;
    inv01 ix34182 (.Y (nx34183), .A (nx38235)) ;
    inv01 ix34184 (.Y (nx34185), .A (nx38235)) ;
    inv01 ix34186 (.Y (nx34187), .A (nx38237)) ;
    inv01 ix34188 (.Y (nx34189), .A (nx38237)) ;
    inv01 ix34190 (.Y (nx34191), .A (nx38237)) ;
    inv01 ix34192 (.Y (nx34193), .A (nx38237)) ;
    inv01 ix34194 (.Y (nx34195), .A (nx38237)) ;
    inv01 ix34196 (.Y (nx34197), .A (nx38237)) ;
    inv01 ix34198 (.Y (nx34199), .A (nx38237)) ;
    inv01 ix34200 (.Y (nx34201), .A (nx38239)) ;
    inv01 ix34202 (.Y (nx34203), .A (nx38239)) ;
    inv01 ix34204 (.Y (nx34205), .A (nx38239)) ;
    inv01 ix34206 (.Y (nx34207), .A (nx38239)) ;
    inv01 ix34208 (.Y (nx34209), .A (nx38239)) ;
    inv01 ix34210 (.Y (nx34211), .A (nx38239)) ;
    inv01 ix34212 (.Y (nx34213), .A (nx38239)) ;
    inv01 ix34214 (.Y (nx34215), .A (nx38241)) ;
    inv01 ix34216 (.Y (nx34217), .A (nx38241)) ;
    inv01 ix34218 (.Y (nx34219), .A (nx38241)) ;
    inv01 ix34220 (.Y (nx34221), .A (nx38241)) ;
    inv01 ix34222 (.Y (nx34223), .A (nx38241)) ;
    inv01 ix34224 (.Y (nx34225), .A (nx38241)) ;
    inv01 ix34226 (.Y (nx34227), .A (nx38241)) ;
    inv01 ix34228 (.Y (nx34229), .A (nx38243)) ;
    inv01 ix34230 (.Y (nx34231), .A (nx38243)) ;
    inv01 ix34232 (.Y (nx34233), .A (nx38243)) ;
    inv01 ix34234 (.Y (nx34235), .A (nx38243)) ;
    inv01 ix34236 (.Y (nx34237), .A (nx38243)) ;
    inv01 ix34238 (.Y (nx34239), .A (nx38243)) ;
    inv01 ix34240 (.Y (nx34241), .A (nx38243)) ;
    inv01 ix34242 (.Y (nx34243), .A (nx38245)) ;
    inv01 ix34244 (.Y (nx34245), .A (nx38245)) ;
    inv01 ix34246 (.Y (nx34247), .A (nx38245)) ;
    inv01 ix34248 (.Y (nx34249), .A (nx38245)) ;
    inv01 ix34250 (.Y (nx34251), .A (nx38245)) ;
    inv01 ix34252 (.Y (nx34253), .A (nx38245)) ;
    inv01 ix34254 (.Y (nx34255), .A (nx38245)) ;
    inv01 ix34256 (.Y (nx34257), .A (nx38247)) ;
    inv01 ix34258 (.Y (nx34259), .A (nx38247)) ;
    inv01 ix34260 (.Y (nx34261), .A (nx38247)) ;
    inv01 ix34262 (.Y (nx34263), .A (nx38247)) ;
    inv01 ix34264 (.Y (nx34265), .A (nx38247)) ;
    inv01 ix34266 (.Y (nx34267), .A (nx38247)) ;
    inv01 ix34268 (.Y (nx34269), .A (nx38247)) ;
    inv01 ix34270 (.Y (nx34271), .A (nx38249)) ;
    inv01 ix34272 (.Y (nx34273), .A (nx38249)) ;
    inv01 ix34274 (.Y (nx34275), .A (nx38249)) ;
    inv01 ix34276 (.Y (nx34277), .A (nx38249)) ;
    inv01 ix34278 (.Y (nx34279), .A (nx38249)) ;
    inv01 ix34280 (.Y (nx34281), .A (nx38249)) ;
    inv01 ix34282 (.Y (nx34283), .A (nx38249)) ;
    inv01 ix34284 (.Y (nx34285), .A (nx38251)) ;
    inv01 ix34286 (.Y (nx34287), .A (nx38251)) ;
    inv01 ix34288 (.Y (nx34289), .A (nx38251)) ;
    inv01 ix34290 (.Y (nx34291), .A (nx38251)) ;
    inv01 ix34292 (.Y (nx34293), .A (nx38251)) ;
    inv01 ix34294 (.Y (nx34295), .A (nx38251)) ;
    inv01 ix34296 (.Y (nx34297), .A (nx38251)) ;
    inv01 ix34298 (.Y (nx34299), .A (nx38253)) ;
    inv01 ix34300 (.Y (nx34301), .A (nx38253)) ;
    inv01 ix34302 (.Y (nx34303), .A (nx38253)) ;
    inv01 ix34304 (.Y (nx34305), .A (nx38253)) ;
    inv01 ix34306 (.Y (nx34307), .A (nx38253)) ;
    inv01 ix34308 (.Y (nx34309), .A (nx38253)) ;
    inv01 ix34310 (.Y (nx34311), .A (nx38253)) ;
    inv01 ix34312 (.Y (nx34313), .A (nx38255)) ;
    inv01 ix34314 (.Y (nx34315), .A (nx38255)) ;
    inv01 ix34316 (.Y (nx34317), .A (nx38255)) ;
    inv01 ix34318 (.Y (nx34319), .A (nx38255)) ;
    inv01 ix34320 (.Y (nx34321), .A (nx38255)) ;
    inv01 ix34322 (.Y (nx34323), .A (nx38255)) ;
    inv01 ix34324 (.Y (nx34325), .A (nx38255)) ;
    inv01 ix34326 (.Y (nx34327), .A (nx38257)) ;
    inv01 ix34328 (.Y (nx34329), .A (nx38257)) ;
    inv01 ix34330 (.Y (nx34331), .A (nx38257)) ;
    inv01 ix34332 (.Y (nx34333), .A (nx38257)) ;
    inv01 ix34334 (.Y (nx34335), .A (nx38257)) ;
    inv01 ix34336 (.Y (nx34337), .A (nx38257)) ;
    inv01 ix34338 (.Y (nx34339), .A (nx38257)) ;
    inv01 ix34340 (.Y (nx34341), .A (nx38259)) ;
    inv01 ix34342 (.Y (nx34343), .A (nx38259)) ;
    inv01 ix34344 (.Y (nx34345), .A (nx38259)) ;
    inv01 ix34346 (.Y (nx34347), .A (nx38259)) ;
    inv01 ix34348 (.Y (nx34349), .A (nx38259)) ;
    inv01 ix34350 (.Y (nx34351), .A (nx38259)) ;
    inv01 ix34352 (.Y (nx34353), .A (nx38259)) ;
    inv01 ix34354 (.Y (nx34355), .A (nx38261)) ;
    inv01 ix34356 (.Y (nx34357), .A (nx38261)) ;
    inv01 ix34358 (.Y (nx34359), .A (nx38261)) ;
    inv01 ix34360 (.Y (nx34361), .A (nx38261)) ;
    inv01 ix34362 (.Y (nx34363), .A (nx38261)) ;
    inv01 ix34364 (.Y (nx34365), .A (nx38261)) ;
    inv01 ix34366 (.Y (nx34367), .A (nx38261)) ;
    inv01 ix34368 (.Y (nx34369), .A (nx38263)) ;
    inv01 ix34370 (.Y (nx34371), .A (nx38263)) ;
    inv01 ix34372 (.Y (nx34373), .A (nx38263)) ;
    inv01 ix34374 (.Y (nx34375), .A (nx38263)) ;
    inv01 ix34376 (.Y (nx34377), .A (nx38263)) ;
    inv01 ix34378 (.Y (nx34379), .A (nx38263)) ;
    inv01 ix34380 (.Y (nx34381), .A (nx38263)) ;
    inv01 ix34382 (.Y (nx34383), .A (nx38265)) ;
    inv01 ix34384 (.Y (nx34385), .A (nx38265)) ;
    inv01 ix34386 (.Y (nx34387), .A (nx38265)) ;
    inv01 ix34388 (.Y (nx34389), .A (nx38265)) ;
    inv01 ix34390 (.Y (nx34391), .A (nx38265)) ;
    inv01 ix34392 (.Y (nx34393), .A (nx38265)) ;
    inv01 ix34394 (.Y (nx34395), .A (nx38265)) ;
    inv01 ix34396 (.Y (nx34397), .A (nx38267)) ;
    inv01 ix34398 (.Y (nx34399), .A (nx38267)) ;
    inv01 ix34400 (.Y (nx34401), .A (nx38267)) ;
    inv01 ix34402 (.Y (nx34403), .A (nx38267)) ;
    inv01 ix34404 (.Y (nx34405), .A (nx38267)) ;
    inv01 ix34406 (.Y (nx34407), .A (nx38267)) ;
    inv01 ix34408 (.Y (nx34409), .A (nx38267)) ;
    inv01 ix34410 (.Y (nx34411), .A (nx38269)) ;
    inv01 ix34412 (.Y (nx34413), .A (nx38269)) ;
    inv01 ix34414 (.Y (nx34415), .A (nx38269)) ;
    inv01 ix34416 (.Y (nx34417), .A (nx38269)) ;
    inv01 ix34418 (.Y (nx34419), .A (nx38269)) ;
    inv01 ix34420 (.Y (nx34421), .A (nx38269)) ;
    inv01 ix34422 (.Y (nx34423), .A (nx38269)) ;
    inv01 ix34424 (.Y (nx34425), .A (nx38271)) ;
    inv01 ix34426 (.Y (nx34427), .A (nx38271)) ;
    inv01 ix34428 (.Y (nx34429), .A (nx38271)) ;
    inv01 ix34430 (.Y (nx34431), .A (nx38271)) ;
    inv01 ix34432 (.Y (nx34433), .A (nx38271)) ;
    inv01 ix34434 (.Y (nx34435), .A (nx38271)) ;
    inv01 ix34436 (.Y (nx34437), .A (nx38271)) ;
    inv01 ix34438 (.Y (nx34439), .A (nx38273)) ;
    inv01 ix34440 (.Y (nx34441), .A (nx38273)) ;
    inv01 ix34442 (.Y (nx34443), .A (nx38273)) ;
    inv01 ix34444 (.Y (nx34445), .A (nx38273)) ;
    inv01 ix34446 (.Y (nx34447), .A (nx38273)) ;
    inv01 ix34448 (.Y (nx34449), .A (nx38273)) ;
    inv01 ix34450 (.Y (nx34451), .A (nx38273)) ;
    inv01 ix34452 (.Y (nx34453), .A (nx38275)) ;
    inv01 ix34454 (.Y (nx34455), .A (nx38275)) ;
    inv01 ix34456 (.Y (nx34457), .A (nx38275)) ;
    inv01 ix34458 (.Y (nx34459), .A (nx38275)) ;
    inv01 ix34460 (.Y (nx34461), .A (nx38275)) ;
    inv01 ix34462 (.Y (nx34463), .A (nx38275)) ;
    inv01 ix34464 (.Y (nx34465), .A (nx38275)) ;
    inv01 ix34466 (.Y (nx34467), .A (nx38277)) ;
    inv01 ix34468 (.Y (nx34469), .A (nx38277)) ;
    inv01 ix34470 (.Y (nx34471), .A (nx38277)) ;
    inv01 ix34472 (.Y (nx34473), .A (nx38277)) ;
    inv01 ix34474 (.Y (nx34475), .A (nx38277)) ;
    inv01 ix34476 (.Y (nx34477), .A (nx38277)) ;
    inv01 ix34478 (.Y (nx34479), .A (nx38277)) ;
    inv01 ix34480 (.Y (nx34481), .A (nx38279)) ;
    inv01 ix34482 (.Y (nx34483), .A (nx38279)) ;
    inv01 ix34484 (.Y (nx34485), .A (nx38279)) ;
    inv01 ix34486 (.Y (nx34487), .A (nx38279)) ;
    inv01 ix34488 (.Y (nx34489), .A (nx38279)) ;
    inv01 ix34490 (.Y (nx34491), .A (nx38279)) ;
    inv01 ix34492 (.Y (nx34493), .A (nx38279)) ;
    inv01 ix34494 (.Y (nx34495), .A (nx38281)) ;
    inv01 ix34496 (.Y (nx34497), .A (nx38281)) ;
    inv01 ix34498 (.Y (nx34499), .A (nx38281)) ;
    inv01 ix34500 (.Y (nx34501), .A (nx38281)) ;
    inv01 ix34502 (.Y (nx34503), .A (nx38281)) ;
    inv01 ix34504 (.Y (nx34505), .A (nx38281)) ;
    inv01 ix34506 (.Y (nx34507), .A (nx38281)) ;
    inv01 ix34508 (.Y (nx34509), .A (nx38283)) ;
    inv01 ix34510 (.Y (nx34511), .A (nx38283)) ;
    inv01 ix34512 (.Y (nx34513), .A (nx38283)) ;
    inv01 ix34514 (.Y (nx34515), .A (nx38283)) ;
    inv01 ix34516 (.Y (nx34517), .A (nx38283)) ;
    inv01 ix34518 (.Y (nx34519), .A (nx38283)) ;
    inv01 ix34520 (.Y (nx34521), .A (nx38283)) ;
    inv01 ix34522 (.Y (nx34523), .A (nx38285)) ;
    inv01 ix34524 (.Y (nx34525), .A (nx38285)) ;
    inv01 ix34526 (.Y (nx34527), .A (nx38285)) ;
    inv01 ix34528 (.Y (nx34529), .A (nx38285)) ;
    inv01 ix34530 (.Y (nx34531), .A (nx38285)) ;
    inv01 ix34532 (.Y (nx34533), .A (nx38285)) ;
    inv01 ix34534 (.Y (nx34535), .A (nx38285)) ;
    inv01 ix34536 (.Y (nx34537), .A (nx38287)) ;
    inv01 ix34538 (.Y (nx34539), .A (nx38287)) ;
    inv01 ix34540 (.Y (nx34541), .A (nx38287)) ;
    inv01 ix34542 (.Y (nx34543), .A (nx38287)) ;
    inv01 ix34544 (.Y (nx34545), .A (nx38287)) ;
    inv01 ix34546 (.Y (nx34547), .A (nx38287)) ;
    inv01 ix34548 (.Y (nx34549), .A (nx38287)) ;
    inv01 ix34550 (.Y (nx34551), .A (nx38289)) ;
    inv01 ix34552 (.Y (nx34553), .A (nx38289)) ;
    inv01 ix34554 (.Y (nx34555), .A (nx38289)) ;
    inv01 ix34556 (.Y (nx34557), .A (nx38289)) ;
    inv01 ix34558 (.Y (nx34559), .A (nx38289)) ;
    inv01 ix34560 (.Y (nx34561), .A (nx38289)) ;
    inv01 ix34562 (.Y (nx34563), .A (nx38289)) ;
    inv01 ix34564 (.Y (nx34565), .A (nx38291)) ;
    inv01 ix34566 (.Y (nx34567), .A (nx38291)) ;
    inv01 ix34568 (.Y (nx34569), .A (nx38291)) ;
    inv01 ix34570 (.Y (nx34571), .A (nx38291)) ;
    inv01 ix34572 (.Y (nx34573), .A (nx38291)) ;
    inv01 ix34574 (.Y (nx34575), .A (nx38291)) ;
    inv01 ix34576 (.Y (nx34577), .A (nx38291)) ;
    inv01 ix34578 (.Y (nx34579), .A (nx38293)) ;
    inv01 ix34580 (.Y (nx34581), .A (nx38293)) ;
    inv01 ix34582 (.Y (nx34583), .A (nx38293)) ;
    inv01 ix34584 (.Y (nx34585), .A (nx38293)) ;
    inv01 ix34586 (.Y (nx34587), .A (nx38293)) ;
    inv01 ix34588 (.Y (nx34589), .A (nx38293)) ;
    inv01 ix34590 (.Y (nx34591), .A (nx38293)) ;
    inv01 ix34592 (.Y (nx34593), .A (nx38295)) ;
    inv01 ix34594 (.Y (nx34595), .A (nx38295)) ;
    inv01 ix34596 (.Y (nx34597), .A (nx38295)) ;
    inv01 ix34598 (.Y (nx34599), .A (nx38295)) ;
    inv01 ix34600 (.Y (nx34601), .A (nx38295)) ;
    inv01 ix34602 (.Y (nx34603), .A (nx38295)) ;
    inv01 ix34604 (.Y (nx34605), .A (nx38295)) ;
    inv01 ix34606 (.Y (nx34607), .A (nx33639)) ;
    inv01 ix34608 (.Y (nx34609), .A (weightsBus[6])) ;
    inv01 ix34610 (.Y (nx34611), .A (nx38297)) ;
    inv01 ix34612 (.Y (nx34613), .A (nx38297)) ;
    inv01 ix34614 (.Y (nx34615), .A (nx38297)) ;
    inv01 ix34616 (.Y (nx34617), .A (nx38297)) ;
    inv01 ix34618 (.Y (nx34619), .A (nx38297)) ;
    inv01 ix34620 (.Y (nx34621), .A (nx38297)) ;
    inv01 ix34622 (.Y (nx34623), .A (nx38297)) ;
    inv01 ix34624 (.Y (nx34625), .A (nx38299)) ;
    inv01 ix34626 (.Y (nx34627), .A (nx38299)) ;
    inv01 ix34628 (.Y (nx34629), .A (nx38299)) ;
    inv01 ix34630 (.Y (nx34631), .A (nx38299)) ;
    inv01 ix34632 (.Y (nx34633), .A (nx38299)) ;
    inv01 ix34634 (.Y (nx34635), .A (nx38299)) ;
    inv01 ix34636 (.Y (nx34637), .A (nx38299)) ;
    inv01 ix34638 (.Y (nx34639), .A (nx38301)) ;
    inv01 ix34640 (.Y (nx34641), .A (nx38301)) ;
    inv01 ix34642 (.Y (nx34643), .A (nx38301)) ;
    inv01 ix34644 (.Y (nx34645), .A (nx38301)) ;
    inv01 ix34646 (.Y (nx34647), .A (nx38301)) ;
    inv01 ix34648 (.Y (nx34649), .A (nx38301)) ;
    inv01 ix34650 (.Y (nx34651), .A (nx38301)) ;
    inv01 ix34652 (.Y (nx34653), .A (nx38303)) ;
    inv01 ix34654 (.Y (nx34655), .A (nx38303)) ;
    inv01 ix34656 (.Y (nx34657), .A (nx38303)) ;
    inv01 ix34658 (.Y (nx34659), .A (nx38303)) ;
    inv01 ix34660 (.Y (nx34661), .A (nx38303)) ;
    inv01 ix34662 (.Y (nx34663), .A (nx38303)) ;
    inv01 ix34664 (.Y (nx34665), .A (nx38303)) ;
    inv01 ix34666 (.Y (nx34667), .A (nx38305)) ;
    inv01 ix34668 (.Y (nx34669), .A (nx38305)) ;
    inv01 ix34670 (.Y (nx34671), .A (nx38305)) ;
    inv01 ix34672 (.Y (nx34673), .A (nx38305)) ;
    inv01 ix34674 (.Y (nx34675), .A (nx38305)) ;
    inv01 ix34676 (.Y (nx34677), .A (nx38305)) ;
    inv01 ix34678 (.Y (nx34679), .A (nx38305)) ;
    inv01 ix34680 (.Y (nx34681), .A (nx38307)) ;
    inv01 ix34682 (.Y (nx34683), .A (nx38307)) ;
    inv01 ix34684 (.Y (nx34685), .A (nx38307)) ;
    inv01 ix34686 (.Y (nx34687), .A (nx38307)) ;
    inv01 ix34688 (.Y (nx34689), .A (nx38307)) ;
    inv01 ix34690 (.Y (nx34691), .A (nx38307)) ;
    inv01 ix34692 (.Y (nx34693), .A (nx38307)) ;
    inv01 ix34694 (.Y (nx34695), .A (nx38309)) ;
    inv01 ix34696 (.Y (nx34697), .A (nx38309)) ;
    inv01 ix34698 (.Y (nx34699), .A (nx38309)) ;
    inv01 ix34700 (.Y (nx34701), .A (nx38309)) ;
    inv01 ix34702 (.Y (nx34703), .A (nx38309)) ;
    inv01 ix34704 (.Y (nx34705), .A (nx38309)) ;
    inv01 ix34706 (.Y (nx34707), .A (nx38309)) ;
    inv01 ix34708 (.Y (nx34709), .A (nx38311)) ;
    inv01 ix34710 (.Y (nx34711), .A (nx38311)) ;
    inv01 ix34712 (.Y (nx34713), .A (nx38311)) ;
    inv01 ix34714 (.Y (nx34715), .A (nx38311)) ;
    inv01 ix34716 (.Y (nx34717), .A (nx38311)) ;
    inv01 ix34718 (.Y (nx34719), .A (nx38311)) ;
    inv01 ix34720 (.Y (nx34721), .A (nx38311)) ;
    inv01 ix34722 (.Y (nx34723), .A (nx38313)) ;
    inv01 ix34724 (.Y (nx34725), .A (nx38313)) ;
    inv01 ix34726 (.Y (nx34727), .A (nx38313)) ;
    inv01 ix34728 (.Y (nx34729), .A (nx38313)) ;
    inv01 ix34730 (.Y (nx34731), .A (nx38313)) ;
    inv01 ix34732 (.Y (nx34733), .A (nx38313)) ;
    inv01 ix34734 (.Y (nx34735), .A (nx38313)) ;
    inv01 ix34736 (.Y (nx34737), .A (nx34609)) ;
    inv01 ix34738 (.Y (nx34739), .A (nx34609)) ;
    inv01 ix34740 (.Y (nx34741), .A (nx34609)) ;
    inv01 ix34742 (.Y (nx34743), .A (nx34609)) ;
    inv01 ix34744 (.Y (nx34745), .A (nx34609)) ;
    inv01 ix34746 (.Y (nx34747), .A (nx34609)) ;
    inv01 ix34748 (.Y (nx34749), .A (nx34609)) ;
    inv01 ix34750 (.Y (nx34751), .A (weightsBus[5])) ;
    inv01 ix34752 (.Y (nx34753), .A (nx38315)) ;
    inv01 ix34754 (.Y (nx34755), .A (nx38315)) ;
    inv01 ix34756 (.Y (nx34757), .A (nx38315)) ;
    inv01 ix34758 (.Y (nx34759), .A (nx38315)) ;
    inv01 ix34760 (.Y (nx34761), .A (nx38315)) ;
    inv01 ix34762 (.Y (nx34763), .A (nx38315)) ;
    inv01 ix34764 (.Y (nx34765), .A (nx38315)) ;
    inv01 ix34766 (.Y (nx34767), .A (nx38317)) ;
    inv01 ix34768 (.Y (nx34769), .A (nx38317)) ;
    inv01 ix34770 (.Y (nx34771), .A (nx38317)) ;
    inv01 ix34772 (.Y (nx34773), .A (nx38317)) ;
    inv01 ix34774 (.Y (nx34775), .A (nx38317)) ;
    inv01 ix34776 (.Y (nx34777), .A (nx38317)) ;
    inv01 ix34778 (.Y (nx34779), .A (nx38317)) ;
    inv01 ix34780 (.Y (nx34781), .A (nx38319)) ;
    inv01 ix34782 (.Y (nx34783), .A (nx38319)) ;
    inv01 ix34784 (.Y (nx34785), .A (nx38319)) ;
    inv01 ix34786 (.Y (nx34787), .A (nx38319)) ;
    inv01 ix34788 (.Y (nx34789), .A (nx38319)) ;
    inv01 ix34790 (.Y (nx34791), .A (nx38319)) ;
    inv01 ix34792 (.Y (nx34793), .A (nx38319)) ;
    inv01 ix34794 (.Y (nx34795), .A (nx38321)) ;
    inv01 ix34796 (.Y (nx34797), .A (nx38321)) ;
    inv01 ix34798 (.Y (nx34799), .A (nx38321)) ;
    inv01 ix34800 (.Y (nx34801), .A (nx38321)) ;
    inv01 ix34802 (.Y (nx34803), .A (nx38321)) ;
    inv01 ix34804 (.Y (nx34805), .A (nx38321)) ;
    inv01 ix34806 (.Y (nx34807), .A (nx38321)) ;
    inv01 ix34808 (.Y (nx34809), .A (nx38323)) ;
    inv01 ix34810 (.Y (nx34811), .A (nx38323)) ;
    inv01 ix34812 (.Y (nx34813), .A (nx38323)) ;
    inv01 ix34814 (.Y (nx34815), .A (nx38323)) ;
    inv01 ix34816 (.Y (nx34817), .A (nx38323)) ;
    inv01 ix34818 (.Y (nx34819), .A (nx38323)) ;
    inv01 ix34820 (.Y (nx34821), .A (nx38323)) ;
    inv01 ix34822 (.Y (nx34823), .A (nx38325)) ;
    inv01 ix34824 (.Y (nx34825), .A (nx38325)) ;
    inv01 ix34826 (.Y (nx34827), .A (nx38325)) ;
    inv01 ix34828 (.Y (nx34829), .A (nx38325)) ;
    inv01 ix34830 (.Y (nx34831), .A (nx38325)) ;
    inv01 ix34832 (.Y (nx34833), .A (nx38325)) ;
    inv01 ix34834 (.Y (nx34835), .A (nx38325)) ;
    inv01 ix34836 (.Y (nx34837), .A (nx38327)) ;
    inv01 ix34838 (.Y (nx34839), .A (nx38327)) ;
    inv01 ix34840 (.Y (nx34841), .A (nx38327)) ;
    inv01 ix34842 (.Y (nx34843), .A (nx38327)) ;
    inv01 ix34844 (.Y (nx34845), .A (nx38327)) ;
    inv01 ix34846 (.Y (nx34847), .A (nx38327)) ;
    inv01 ix34848 (.Y (nx34849), .A (nx38327)) ;
    inv01 ix34850 (.Y (nx34851), .A (nx38329)) ;
    inv01 ix34852 (.Y (nx34853), .A (nx38329)) ;
    inv01 ix34854 (.Y (nx34855), .A (nx38329)) ;
    inv01 ix34856 (.Y (nx34857), .A (nx38329)) ;
    inv01 ix34858 (.Y (nx34859), .A (nx38329)) ;
    inv01 ix34860 (.Y (nx34861), .A (nx38329)) ;
    inv01 ix34862 (.Y (nx34863), .A (nx38329)) ;
    inv01 ix34864 (.Y (nx34865), .A (nx38331)) ;
    inv01 ix34866 (.Y (nx34867), .A (nx38331)) ;
    inv01 ix34868 (.Y (nx34869), .A (nx38331)) ;
    inv01 ix34870 (.Y (nx34871), .A (nx38331)) ;
    inv01 ix34872 (.Y (nx34873), .A (nx38331)) ;
    inv01 ix34874 (.Y (nx34875), .A (nx38331)) ;
    inv01 ix34876 (.Y (nx34877), .A (nx38331)) ;
    inv01 ix34878 (.Y (nx34879), .A (nx34751)) ;
    inv01 ix34880 (.Y (nx34881), .A (nx34751)) ;
    inv01 ix34882 (.Y (nx34883), .A (nx34751)) ;
    inv01 ix34884 (.Y (nx34885), .A (nx34751)) ;
    inv01 ix34886 (.Y (nx34887), .A (nx34751)) ;
    inv01 ix34888 (.Y (nx34889), .A (nx34751)) ;
    inv01 ix34890 (.Y (nx34891), .A (nx34751)) ;
    inv01 ix34892 (.Y (nx34893), .A (weightsBus[4])) ;
    inv01 ix34894 (.Y (nx34895), .A (nx38333)) ;
    inv01 ix34896 (.Y (nx34897), .A (nx38333)) ;
    inv01 ix34898 (.Y (nx34899), .A (nx38333)) ;
    inv01 ix34900 (.Y (nx34901), .A (nx38333)) ;
    inv01 ix34902 (.Y (nx34903), .A (nx38333)) ;
    inv01 ix34904 (.Y (nx34905), .A (nx38333)) ;
    inv01 ix34906 (.Y (nx34907), .A (nx38333)) ;
    inv01 ix34908 (.Y (nx34909), .A (nx38335)) ;
    inv01 ix34910 (.Y (nx34911), .A (nx38335)) ;
    inv01 ix34912 (.Y (nx34913), .A (nx38335)) ;
    inv01 ix34914 (.Y (nx34915), .A (nx38335)) ;
    inv01 ix34916 (.Y (nx34917), .A (nx38335)) ;
    inv01 ix34918 (.Y (nx34919), .A (nx38335)) ;
    inv01 ix34920 (.Y (nx34921), .A (nx38335)) ;
    inv01 ix34922 (.Y (nx34923), .A (nx38337)) ;
    inv01 ix34924 (.Y (nx34925), .A (nx38337)) ;
    inv01 ix34926 (.Y (nx34927), .A (nx38337)) ;
    inv01 ix34928 (.Y (nx34929), .A (nx38337)) ;
    inv01 ix34930 (.Y (nx34931), .A (nx38337)) ;
    inv01 ix34932 (.Y (nx34933), .A (nx38337)) ;
    inv01 ix34934 (.Y (nx34935), .A (nx38337)) ;
    inv01 ix34936 (.Y (nx34937), .A (nx38339)) ;
    inv01 ix34938 (.Y (nx34939), .A (nx38339)) ;
    inv01 ix34940 (.Y (nx34941), .A (nx38339)) ;
    inv01 ix34942 (.Y (nx34943), .A (nx38339)) ;
    inv01 ix34944 (.Y (nx34945), .A (nx38339)) ;
    inv01 ix34946 (.Y (nx34947), .A (nx38339)) ;
    inv01 ix34948 (.Y (nx34949), .A (nx38339)) ;
    inv01 ix34950 (.Y (nx34951), .A (nx38341)) ;
    inv01 ix34952 (.Y (nx34953), .A (nx38341)) ;
    inv01 ix34954 (.Y (nx34955), .A (nx38341)) ;
    inv01 ix34956 (.Y (nx34957), .A (nx38341)) ;
    inv01 ix34958 (.Y (nx34959), .A (nx38341)) ;
    inv01 ix34960 (.Y (nx34961), .A (nx38341)) ;
    inv01 ix34962 (.Y (nx34963), .A (nx38341)) ;
    inv01 ix34964 (.Y (nx34965), .A (nx38343)) ;
    inv01 ix34966 (.Y (nx34967), .A (nx38343)) ;
    inv01 ix34968 (.Y (nx34969), .A (nx38343)) ;
    inv01 ix34970 (.Y (nx34971), .A (nx38343)) ;
    inv01 ix34972 (.Y (nx34973), .A (nx38343)) ;
    inv01 ix34974 (.Y (nx34975), .A (nx38343)) ;
    inv01 ix34976 (.Y (nx34977), .A (nx38343)) ;
    inv01 ix34978 (.Y (nx34979), .A (nx38345)) ;
    inv01 ix34980 (.Y (nx34981), .A (nx38345)) ;
    inv01 ix34982 (.Y (nx34983), .A (nx38345)) ;
    inv01 ix34984 (.Y (nx34985), .A (nx38345)) ;
    inv01 ix34986 (.Y (nx34987), .A (nx38345)) ;
    inv01 ix34988 (.Y (nx34989), .A (nx38345)) ;
    inv01 ix34990 (.Y (nx34991), .A (nx38345)) ;
    inv01 ix34992 (.Y (nx34993), .A (nx38347)) ;
    inv01 ix34994 (.Y (nx34995), .A (nx38347)) ;
    inv01 ix34996 (.Y (nx34997), .A (nx38347)) ;
    inv01 ix34998 (.Y (nx34999), .A (nx38347)) ;
    inv01 ix35000 (.Y (nx35001), .A (nx38347)) ;
    inv01 ix35002 (.Y (nx35003), .A (nx38347)) ;
    inv01 ix35004 (.Y (nx35005), .A (nx38347)) ;
    inv01 ix35006 (.Y (nx35007), .A (nx38349)) ;
    inv01 ix35008 (.Y (nx35009), .A (nx38349)) ;
    inv01 ix35010 (.Y (nx35011), .A (nx38349)) ;
    inv01 ix35012 (.Y (nx35013), .A (nx38349)) ;
    inv01 ix35014 (.Y (nx35015), .A (nx38349)) ;
    inv01 ix35016 (.Y (nx35017), .A (nx38349)) ;
    inv01 ix35018 (.Y (nx35019), .A (nx38349)) ;
    inv01 ix35020 (.Y (nx35021), .A (nx34893)) ;
    inv01 ix35022 (.Y (nx35023), .A (nx34893)) ;
    inv01 ix35024 (.Y (nx35025), .A (nx34893)) ;
    inv01 ix35026 (.Y (nx35027), .A (nx34893)) ;
    inv01 ix35028 (.Y (nx35029), .A (nx34893)) ;
    inv01 ix35030 (.Y (nx35031), .A (nx34893)) ;
    inv01 ix35032 (.Y (nx35033), .A (nx34893)) ;
    inv01 ix35034 (.Y (nx35035), .A (weightsBus[3])) ;
    inv01 ix35036 (.Y (nx35037), .A (nx38351)) ;
    inv01 ix35038 (.Y (nx35039), .A (nx38351)) ;
    inv01 ix35040 (.Y (nx35041), .A (nx38351)) ;
    inv01 ix35042 (.Y (nx35043), .A (nx38351)) ;
    inv01 ix35044 (.Y (nx35045), .A (nx38351)) ;
    inv01 ix35046 (.Y (nx35047), .A (nx38351)) ;
    inv01 ix35048 (.Y (nx35049), .A (nx38351)) ;
    inv01 ix35050 (.Y (nx35051), .A (nx38353)) ;
    inv01 ix35052 (.Y (nx35053), .A (nx38353)) ;
    inv01 ix35054 (.Y (nx35055), .A (nx38353)) ;
    inv01 ix35056 (.Y (nx35057), .A (nx38353)) ;
    inv01 ix35058 (.Y (nx35059), .A (nx38353)) ;
    inv01 ix35060 (.Y (nx35061), .A (nx38353)) ;
    inv01 ix35062 (.Y (nx35063), .A (nx38353)) ;
    inv01 ix35064 (.Y (nx35065), .A (nx38355)) ;
    inv01 ix35066 (.Y (nx35067), .A (nx38355)) ;
    inv01 ix35068 (.Y (nx35069), .A (nx38355)) ;
    inv01 ix35070 (.Y (nx35071), .A (nx38355)) ;
    inv01 ix35072 (.Y (nx35073), .A (nx38355)) ;
    inv01 ix35074 (.Y (nx35075), .A (nx38355)) ;
    inv01 ix35076 (.Y (nx35077), .A (nx38355)) ;
    inv01 ix35078 (.Y (nx35079), .A (nx38357)) ;
    inv01 ix35080 (.Y (nx35081), .A (nx38357)) ;
    inv01 ix35082 (.Y (nx35083), .A (nx38357)) ;
    inv01 ix35084 (.Y (nx35085), .A (nx38357)) ;
    inv01 ix35086 (.Y (nx35087), .A (nx38357)) ;
    inv01 ix35088 (.Y (nx35089), .A (nx38357)) ;
    inv01 ix35090 (.Y (nx35091), .A (nx38357)) ;
    inv01 ix35092 (.Y (nx35093), .A (nx38359)) ;
    inv01 ix35094 (.Y (nx35095), .A (nx38359)) ;
    inv01 ix35096 (.Y (nx35097), .A (nx38359)) ;
    inv01 ix35098 (.Y (nx35099), .A (nx38359)) ;
    inv01 ix35100 (.Y (nx35101), .A (nx38359)) ;
    inv01 ix35102 (.Y (nx35103), .A (nx38359)) ;
    inv01 ix35104 (.Y (nx35105), .A (nx38359)) ;
    inv01 ix35106 (.Y (nx35107), .A (nx38361)) ;
    inv01 ix35108 (.Y (nx35109), .A (nx38361)) ;
    inv01 ix35110 (.Y (nx35111), .A (nx38361)) ;
    inv01 ix35112 (.Y (nx35113), .A (nx38361)) ;
    inv01 ix35114 (.Y (nx35115), .A (nx38361)) ;
    inv01 ix35116 (.Y (nx35117), .A (nx38361)) ;
    inv01 ix35118 (.Y (nx35119), .A (nx38361)) ;
    inv01 ix35120 (.Y (nx35121), .A (nx38363)) ;
    inv01 ix35122 (.Y (nx35123), .A (nx38363)) ;
    inv01 ix35124 (.Y (nx35125), .A (nx38363)) ;
    inv01 ix35126 (.Y (nx35127), .A (nx38363)) ;
    inv01 ix35128 (.Y (nx35129), .A (nx38363)) ;
    inv01 ix35130 (.Y (nx35131), .A (nx38363)) ;
    inv01 ix35132 (.Y (nx35133), .A (nx38363)) ;
    inv01 ix35134 (.Y (nx35135), .A (nx38365)) ;
    inv01 ix35136 (.Y (nx35137), .A (nx38365)) ;
    inv01 ix35138 (.Y (nx35139), .A (nx38365)) ;
    inv01 ix35140 (.Y (nx35141), .A (nx38365)) ;
    inv01 ix35142 (.Y (nx35143), .A (nx38365)) ;
    inv01 ix35144 (.Y (nx35145), .A (nx38365)) ;
    inv01 ix35146 (.Y (nx35147), .A (nx38365)) ;
    inv01 ix35148 (.Y (nx35149), .A (nx38367)) ;
    inv01 ix35150 (.Y (nx35151), .A (nx38367)) ;
    inv01 ix35152 (.Y (nx35153), .A (nx38367)) ;
    inv01 ix35154 (.Y (nx35155), .A (nx38367)) ;
    inv01 ix35156 (.Y (nx35157), .A (nx38367)) ;
    inv01 ix35158 (.Y (nx35159), .A (nx38367)) ;
    inv01 ix35160 (.Y (nx35161), .A (nx38367)) ;
    inv01 ix35162 (.Y (nx35163), .A (nx35035)) ;
    inv01 ix35164 (.Y (nx35165), .A (nx35035)) ;
    inv01 ix35166 (.Y (nx35167), .A (nx35035)) ;
    inv01 ix35168 (.Y (nx35169), .A (nx35035)) ;
    inv01 ix35170 (.Y (nx35171), .A (nx35035)) ;
    inv01 ix35172 (.Y (nx35173), .A (nx35035)) ;
    inv01 ix35174 (.Y (nx35175), .A (nx35035)) ;
    inv01 ix35176 (.Y (nx35177), .A (weightsBus[2])) ;
    inv01 ix35178 (.Y (nx35179), .A (nx38369)) ;
    inv01 ix35180 (.Y (nx35181), .A (nx38369)) ;
    inv01 ix35182 (.Y (nx35183), .A (nx38369)) ;
    inv01 ix35184 (.Y (nx35185), .A (nx38369)) ;
    inv01 ix35186 (.Y (nx35187), .A (nx38369)) ;
    inv01 ix35188 (.Y (nx35189), .A (nx38369)) ;
    inv01 ix35190 (.Y (nx35191), .A (nx38369)) ;
    inv01 ix35192 (.Y (nx35193), .A (nx38371)) ;
    inv01 ix35194 (.Y (nx35195), .A (nx38371)) ;
    inv01 ix35196 (.Y (nx35197), .A (nx38371)) ;
    inv01 ix35198 (.Y (nx35199), .A (nx38371)) ;
    inv01 ix35200 (.Y (nx35201), .A (nx38371)) ;
    inv01 ix35202 (.Y (nx35203), .A (nx38371)) ;
    inv01 ix35204 (.Y (nx35205), .A (nx38371)) ;
    inv01 ix35206 (.Y (nx35207), .A (nx38373)) ;
    inv01 ix35208 (.Y (nx35209), .A (nx38373)) ;
    inv01 ix35210 (.Y (nx35211), .A (nx38373)) ;
    inv01 ix35212 (.Y (nx35213), .A (nx38373)) ;
    inv01 ix35214 (.Y (nx35215), .A (nx38373)) ;
    inv01 ix35216 (.Y (nx35217), .A (nx38373)) ;
    inv01 ix35218 (.Y (nx35219), .A (nx38373)) ;
    inv01 ix35220 (.Y (nx35221), .A (nx38375)) ;
    inv01 ix35222 (.Y (nx35223), .A (nx38375)) ;
    inv01 ix35224 (.Y (nx35225), .A (nx38375)) ;
    inv01 ix35226 (.Y (nx35227), .A (nx38375)) ;
    inv01 ix35228 (.Y (nx35229), .A (nx38375)) ;
    inv01 ix35230 (.Y (nx35231), .A (nx38375)) ;
    inv01 ix35232 (.Y (nx35233), .A (nx38375)) ;
    inv01 ix35234 (.Y (nx35235), .A (nx38377)) ;
    inv01 ix35236 (.Y (nx35237), .A (nx38377)) ;
    inv01 ix35238 (.Y (nx35239), .A (nx38377)) ;
    inv01 ix35240 (.Y (nx35241), .A (nx38377)) ;
    inv01 ix35242 (.Y (nx35243), .A (nx38377)) ;
    inv01 ix35244 (.Y (nx35245), .A (nx38377)) ;
    inv01 ix35246 (.Y (nx35247), .A (nx38377)) ;
    inv01 ix35248 (.Y (nx35249), .A (nx38379)) ;
    inv01 ix35250 (.Y (nx35251), .A (nx38379)) ;
    inv01 ix35252 (.Y (nx35253), .A (nx38379)) ;
    inv01 ix35254 (.Y (nx35255), .A (nx38379)) ;
    inv01 ix35256 (.Y (nx35257), .A (nx38379)) ;
    inv01 ix35258 (.Y (nx35259), .A (nx38379)) ;
    inv01 ix35260 (.Y (nx35261), .A (nx38379)) ;
    inv01 ix35262 (.Y (nx35263), .A (nx38381)) ;
    inv01 ix35264 (.Y (nx35265), .A (nx38381)) ;
    inv01 ix35266 (.Y (nx35267), .A (nx38381)) ;
    inv01 ix35268 (.Y (nx35269), .A (nx38381)) ;
    inv01 ix35270 (.Y (nx35271), .A (nx38381)) ;
    inv01 ix35272 (.Y (nx35273), .A (nx38381)) ;
    inv01 ix35274 (.Y (nx35275), .A (nx38381)) ;
    inv01 ix35276 (.Y (nx35277), .A (nx38383)) ;
    inv01 ix35278 (.Y (nx35279), .A (nx38383)) ;
    inv01 ix35280 (.Y (nx35281), .A (nx38383)) ;
    inv01 ix35282 (.Y (nx35283), .A (nx38383)) ;
    inv01 ix35284 (.Y (nx35285), .A (nx38383)) ;
    inv01 ix35286 (.Y (nx35287), .A (nx38383)) ;
    inv01 ix35288 (.Y (nx35289), .A (nx38383)) ;
    inv01 ix35290 (.Y (nx35291), .A (nx38385)) ;
    inv01 ix35292 (.Y (nx35293), .A (nx38385)) ;
    inv01 ix35294 (.Y (nx35295), .A (nx38385)) ;
    inv01 ix35296 (.Y (nx35297), .A (nx38385)) ;
    inv01 ix35298 (.Y (nx35299), .A (nx38385)) ;
    inv01 ix35300 (.Y (nx35301), .A (nx38385)) ;
    inv01 ix35302 (.Y (nx35303), .A (nx38385)) ;
    inv01 ix35304 (.Y (nx35305), .A (nx35177)) ;
    inv01 ix35306 (.Y (nx35307), .A (nx35177)) ;
    inv01 ix35308 (.Y (nx35309), .A (nx35177)) ;
    inv01 ix35310 (.Y (nx35311), .A (nx35177)) ;
    inv01 ix35312 (.Y (nx35313), .A (nx35177)) ;
    inv01 ix35314 (.Y (nx35315), .A (nx35177)) ;
    inv01 ix35316 (.Y (nx35317), .A (nx35177)) ;
    inv01 ix35318 (.Y (nx35319), .A (weightsBus[1])) ;
    inv01 ix35320 (.Y (nx35321), .A (nx38387)) ;
    inv01 ix35322 (.Y (nx35323), .A (nx38387)) ;
    inv01 ix35324 (.Y (nx35325), .A (nx38387)) ;
    inv01 ix35326 (.Y (nx35327), .A (nx38387)) ;
    inv01 ix35328 (.Y (nx35329), .A (nx38387)) ;
    inv01 ix35330 (.Y (nx35331), .A (nx38387)) ;
    inv01 ix35332 (.Y (nx35333), .A (nx38387)) ;
    inv01 ix35334 (.Y (nx35335), .A (nx38389)) ;
    inv01 ix35336 (.Y (nx35337), .A (nx38389)) ;
    inv01 ix35338 (.Y (nx35339), .A (nx38389)) ;
    inv01 ix35340 (.Y (nx35341), .A (nx38389)) ;
    inv01 ix35342 (.Y (nx35343), .A (nx38389)) ;
    inv01 ix35344 (.Y (nx35345), .A (nx38389)) ;
    inv01 ix35346 (.Y (nx35347), .A (nx38389)) ;
    inv01 ix35348 (.Y (nx35349), .A (nx38391)) ;
    inv01 ix35350 (.Y (nx35351), .A (nx38391)) ;
    inv01 ix35352 (.Y (nx35353), .A (nx38391)) ;
    inv01 ix35354 (.Y (nx35355), .A (nx38391)) ;
    inv01 ix35356 (.Y (nx35357), .A (nx38391)) ;
    inv01 ix35358 (.Y (nx35359), .A (nx38391)) ;
    inv01 ix35360 (.Y (nx35361), .A (nx38391)) ;
    inv01 ix35362 (.Y (nx35363), .A (nx38393)) ;
    inv01 ix35364 (.Y (nx35365), .A (nx38393)) ;
    inv01 ix35366 (.Y (nx35367), .A (nx38393)) ;
    inv01 ix35368 (.Y (nx35369), .A (nx38393)) ;
    inv01 ix35370 (.Y (nx35371), .A (nx38393)) ;
    inv01 ix35372 (.Y (nx35373), .A (nx38393)) ;
    inv01 ix35374 (.Y (nx35375), .A (nx38393)) ;
    inv01 ix35376 (.Y (nx35377), .A (nx38395)) ;
    inv01 ix35378 (.Y (nx35379), .A (nx38395)) ;
    inv01 ix35380 (.Y (nx35381), .A (nx38395)) ;
    inv01 ix35382 (.Y (nx35383), .A (nx38395)) ;
    inv01 ix35384 (.Y (nx35385), .A (nx38395)) ;
    inv01 ix35386 (.Y (nx35387), .A (nx38395)) ;
    inv01 ix35388 (.Y (nx35389), .A (nx38395)) ;
    inv01 ix35390 (.Y (nx35391), .A (nx38397)) ;
    inv01 ix35392 (.Y (nx35393), .A (nx38397)) ;
    inv01 ix35394 (.Y (nx35395), .A (nx38397)) ;
    inv01 ix35396 (.Y (nx35397), .A (nx38397)) ;
    inv01 ix35398 (.Y (nx35399), .A (nx38397)) ;
    inv01 ix35400 (.Y (nx35401), .A (nx38397)) ;
    inv01 ix35402 (.Y (nx35403), .A (nx38397)) ;
    inv01 ix35404 (.Y (nx35405), .A (nx38399)) ;
    inv01 ix35406 (.Y (nx35407), .A (nx38399)) ;
    inv01 ix35408 (.Y (nx35409), .A (nx38399)) ;
    inv01 ix35410 (.Y (nx35411), .A (nx38399)) ;
    inv01 ix35412 (.Y (nx35413), .A (nx38399)) ;
    inv01 ix35414 (.Y (nx35415), .A (nx38399)) ;
    inv01 ix35416 (.Y (nx35417), .A (nx38399)) ;
    inv01 ix35418 (.Y (nx35419), .A (nx38401)) ;
    inv01 ix35420 (.Y (nx35421), .A (nx38401)) ;
    inv01 ix35422 (.Y (nx35423), .A (nx38401)) ;
    inv01 ix35424 (.Y (nx35425), .A (nx38401)) ;
    inv01 ix35426 (.Y (nx35427), .A (nx38401)) ;
    inv01 ix35428 (.Y (nx35429), .A (nx38401)) ;
    inv01 ix35430 (.Y (nx35431), .A (nx38401)) ;
    inv01 ix35432 (.Y (nx35433), .A (nx38403)) ;
    inv01 ix35434 (.Y (nx35435), .A (nx38403)) ;
    inv01 ix35436 (.Y (nx35437), .A (nx38403)) ;
    inv01 ix35438 (.Y (nx35439), .A (nx38403)) ;
    inv01 ix35440 (.Y (nx35441), .A (nx38403)) ;
    inv01 ix35442 (.Y (nx35443), .A (nx38403)) ;
    inv01 ix35444 (.Y (nx35445), .A (nx38403)) ;
    inv01 ix35446 (.Y (nx35447), .A (nx35319)) ;
    inv01 ix35448 (.Y (nx35449), .A (nx35319)) ;
    inv01 ix35450 (.Y (nx35451), .A (nx35319)) ;
    inv01 ix35452 (.Y (nx35453), .A (nx35319)) ;
    inv01 ix35454 (.Y (nx35455), .A (nx35319)) ;
    inv01 ix35456 (.Y (nx35457), .A (nx35319)) ;
    inv01 ix35458 (.Y (nx35459), .A (nx35319)) ;
    inv01 ix35460 (.Y (nx35461), .A (weightsBus[0])) ;
    inv01 ix35462 (.Y (nx35463), .A (nx38405)) ;
    inv01 ix35464 (.Y (nx35465), .A (nx38405)) ;
    inv01 ix35466 (.Y (nx35467), .A (nx38405)) ;
    inv01 ix35468 (.Y (nx35469), .A (nx38405)) ;
    inv01 ix35470 (.Y (nx35471), .A (nx38405)) ;
    inv01 ix35472 (.Y (nx35473), .A (nx38405)) ;
    inv01 ix35474 (.Y (nx35475), .A (nx38405)) ;
    inv01 ix35476 (.Y (nx35477), .A (nx38407)) ;
    inv01 ix35478 (.Y (nx35479), .A (nx38407)) ;
    inv01 ix35480 (.Y (nx35481), .A (nx38407)) ;
    inv01 ix35482 (.Y (nx35483), .A (nx38407)) ;
    inv01 ix35484 (.Y (nx35485), .A (nx38407)) ;
    inv01 ix35486 (.Y (nx35487), .A (nx38407)) ;
    inv01 ix35488 (.Y (nx35489), .A (nx38407)) ;
    inv01 ix35490 (.Y (nx35491), .A (nx38409)) ;
    inv01 ix35492 (.Y (nx35493), .A (nx38409)) ;
    inv01 ix35494 (.Y (nx35495), .A (nx38409)) ;
    inv01 ix35496 (.Y (nx35497), .A (nx38409)) ;
    inv01 ix35498 (.Y (nx35499), .A (nx38409)) ;
    inv01 ix35500 (.Y (nx35501), .A (nx38409)) ;
    inv01 ix35502 (.Y (nx35503), .A (nx38409)) ;
    inv01 ix35504 (.Y (nx35505), .A (nx38411)) ;
    inv01 ix35506 (.Y (nx35507), .A (nx38411)) ;
    inv01 ix35508 (.Y (nx35509), .A (nx38411)) ;
    inv01 ix35510 (.Y (nx35511), .A (nx38411)) ;
    inv01 ix35512 (.Y (nx35513), .A (nx38411)) ;
    inv01 ix35514 (.Y (nx35515), .A (nx38411)) ;
    inv01 ix35516 (.Y (nx35517), .A (nx38411)) ;
    inv01 ix35518 (.Y (nx35519), .A (nx38413)) ;
    inv01 ix35520 (.Y (nx35521), .A (nx38413)) ;
    inv01 ix35522 (.Y (nx35523), .A (nx38413)) ;
    inv01 ix35524 (.Y (nx35525), .A (nx38413)) ;
    inv01 ix35526 (.Y (nx35527), .A (nx38413)) ;
    inv01 ix35528 (.Y (nx35529), .A (nx38413)) ;
    inv01 ix35530 (.Y (nx35531), .A (nx38413)) ;
    inv01 ix35532 (.Y (nx35533), .A (nx38415)) ;
    inv01 ix35534 (.Y (nx35535), .A (nx38415)) ;
    inv01 ix35536 (.Y (nx35537), .A (nx38415)) ;
    inv01 ix35538 (.Y (nx35539), .A (nx38415)) ;
    inv01 ix35540 (.Y (nx35541), .A (nx38415)) ;
    inv01 ix35542 (.Y (nx35543), .A (nx38415)) ;
    inv01 ix35544 (.Y (nx35545), .A (nx38415)) ;
    inv01 ix35546 (.Y (nx35547), .A (nx38417)) ;
    inv01 ix35548 (.Y (nx35549), .A (nx38417)) ;
    inv01 ix35550 (.Y (nx35551), .A (nx38417)) ;
    inv01 ix35552 (.Y (nx35553), .A (nx38417)) ;
    inv01 ix35554 (.Y (nx35555), .A (nx38417)) ;
    inv01 ix35556 (.Y (nx35557), .A (nx38417)) ;
    inv01 ix35558 (.Y (nx35559), .A (nx38417)) ;
    inv01 ix35560 (.Y (nx35561), .A (nx38419)) ;
    inv01 ix35562 (.Y (nx35563), .A (nx38419)) ;
    inv01 ix35564 (.Y (nx35565), .A (nx38419)) ;
    inv01 ix35566 (.Y (nx35567), .A (nx38419)) ;
    inv01 ix35568 (.Y (nx35569), .A (nx38419)) ;
    inv01 ix35570 (.Y (nx35571), .A (nx38419)) ;
    inv01 ix35572 (.Y (nx35573), .A (nx38419)) ;
    inv01 ix35574 (.Y (nx35575), .A (nx38421)) ;
    inv01 ix35576 (.Y (nx35577), .A (nx38421)) ;
    inv01 ix35578 (.Y (nx35579), .A (nx38421)) ;
    inv01 ix35580 (.Y (nx35581), .A (nx38421)) ;
    inv01 ix35582 (.Y (nx35583), .A (nx38421)) ;
    inv01 ix35584 (.Y (nx35585), .A (nx38421)) ;
    inv01 ix35586 (.Y (nx35587), .A (nx38421)) ;
    inv01 ix35588 (.Y (nx35589), .A (nx35461)) ;
    inv01 ix35590 (.Y (nx35591), .A (nx35461)) ;
    inv01 ix35592 (.Y (nx35593), .A (nx35461)) ;
    inv01 ix35594 (.Y (nx35595), .A (nx35461)) ;
    inv01 ix35596 (.Y (nx35597), .A (nx35461)) ;
    inv01 ix35598 (.Y (nx35599), .A (nx35461)) ;
    inv01 ix35600 (.Y (nx35601), .A (nx35461)) ;
    inv01 ix35602 (.Y (nx35603), .A (AllRead)) ;
    inv01 ix35604 (.Y (nx35605), .A (nx38423)) ;
    inv01 ix35606 (.Y (nx35607), .A (nx38423)) ;
    inv01 ix35608 (.Y (nx35609), .A (nx38423)) ;
    inv01 ix35610 (.Y (nx35611), .A (nx38423)) ;
    inv01 ix35612 (.Y (nx35613), .A (nx38423)) ;
    inv01 ix35614 (.Y (nx35615), .A (nx38423)) ;
    inv01 ix35616 (.Y (nx35617), .A (nx38423)) ;
    inv01 ix35618 (.Y (nx35619), .A (nx38425)) ;
    inv01 ix35620 (.Y (nx35621), .A (nx38425)) ;
    inv01 ix35622 (.Y (nx35623), .A (nx38425)) ;
    inv01 ix35624 (.Y (nx35625), .A (nx38425)) ;
    inv01 ix35626 (.Y (nx35627), .A (nx38425)) ;
    inv01 ix35628 (.Y (nx35629), .A (nx38425)) ;
    inv01 ix35630 (.Y (nx35631), .A (nx38425)) ;
    inv01 ix35632 (.Y (nx35633), .A (nx38427)) ;
    inv01 ix35634 (.Y (nx35635), .A (nx38427)) ;
    inv01 ix35636 (.Y (nx35637), .A (nx38427)) ;
    inv01 ix35638 (.Y (nx35639), .A (nx38427)) ;
    inv01 ix35640 (.Y (nx35641), .A (nx38427)) ;
    inv01 ix35642 (.Y (nx35643), .A (nx38427)) ;
    inv01 ix35644 (.Y (nx35645), .A (nx38427)) ;
    inv01 ix35646 (.Y (nx35647), .A (nx38429)) ;
    inv01 ix35648 (.Y (nx35649), .A (nx38429)) ;
    inv01 ix35650 (.Y (nx35651), .A (nx38429)) ;
    inv01 ix35652 (.Y (nx35653), .A (nx38429)) ;
    inv01 ix35654 (.Y (nx35655), .A (nx38429)) ;
    inv01 ix35656 (.Y (nx35657), .A (nx38429)) ;
    inv01 ix35658 (.Y (nx35659), .A (nx38429)) ;
    inv01 ix35660 (.Y (nx35661), .A (nx38431)) ;
    inv01 ix35662 (.Y (nx35663), .A (nx38431)) ;
    inv01 ix35664 (.Y (nx35665), .A (nx38431)) ;
    inv01 ix35666 (.Y (nx35667), .A (nx38431)) ;
    inv01 ix35668 (.Y (nx35669), .A (nx38431)) ;
    inv01 ix35670 (.Y (nx35671), .A (nx38431)) ;
    inv01 ix35672 (.Y (nx35673), .A (nx38431)) ;
    inv01 ix35674 (.Y (nx35675), .A (nx38433)) ;
    inv01 ix35676 (.Y (nx35677), .A (nx38433)) ;
    inv01 ix35678 (.Y (nx35679), .A (nx38433)) ;
    inv01 ix35680 (.Y (nx35681), .A (nx38433)) ;
    inv01 ix35682 (.Y (nx35683), .A (nx38433)) ;
    inv01 ix35684 (.Y (nx35685), .A (nx38433)) ;
    inv01 ix35686 (.Y (nx35687), .A (nx38433)) ;
    inv01 ix35688 (.Y (nx35689), .A (nx38435)) ;
    inv01 ix35690 (.Y (nx35691), .A (nx38435)) ;
    inv01 ix35692 (.Y (nx35693), .A (nx38435)) ;
    inv01 ix35694 (.Y (nx35695), .A (nx38435)) ;
    inv01 ix35696 (.Y (nx35697), .A (nx38435)) ;
    inv01 ix35698 (.Y (nx35699), .A (nx38435)) ;
    inv01 ix35700 (.Y (nx35701), .A (nx38435)) ;
    inv01 ix35702 (.Y (nx35703), .A (nx38437)) ;
    inv01 ix35704 (.Y (nx35705), .A (nx38437)) ;
    inv01 ix35706 (.Y (nx35707), .A (nx38437)) ;
    inv01 ix35708 (.Y (nx35709), .A (nx38437)) ;
    inv01 ix35710 (.Y (nx35711), .A (nx38437)) ;
    inv01 ix35712 (.Y (nx35713), .A (nx38437)) ;
    inv01 ix35714 (.Y (nx35715), .A (nx38437)) ;
    inv01 ix35716 (.Y (nx35717), .A (nx38439)) ;
    inv01 ix35718 (.Y (nx35719), .A (nx38439)) ;
    inv01 ix35720 (.Y (nx35721), .A (nx38439)) ;
    inv01 ix35722 (.Y (nx35723), .A (nx38439)) ;
    inv01 ix35724 (.Y (nx35725), .A (nx38439)) ;
    inv01 ix35726 (.Y (nx35727), .A (nx38439)) ;
    inv01 ix35728 (.Y (nx35729), .A (nx38439)) ;
    inv01 ix35730 (.Y (nx35731), .A (nx38441)) ;
    inv01 ix35732 (.Y (nx35733), .A (nx38441)) ;
    inv01 ix35734 (.Y (nx35735), .A (nx38441)) ;
    inv01 ix35736 (.Y (nx35737), .A (nx38441)) ;
    inv01 ix35738 (.Y (nx35739), .A (nx38441)) ;
    inv01 ix35740 (.Y (nx35741), .A (nx38441)) ;
    inv01 ix35742 (.Y (nx35743), .A (nx38441)) ;
    inv01 ix35744 (.Y (nx35745), .A (nx38443)) ;
    inv01 ix35746 (.Y (nx35747), .A (nx38443)) ;
    inv01 ix35748 (.Y (nx35749), .A (nx38443)) ;
    inv01 ix35750 (.Y (nx35751), .A (nx38443)) ;
    inv01 ix35752 (.Y (nx35753), .A (nx38443)) ;
    inv01 ix35754 (.Y (nx35755), .A (nx38443)) ;
    inv01 ix35756 (.Y (nx35757), .A (nx38443)) ;
    inv01 ix35758 (.Y (nx35759), .A (nx38445)) ;
    inv01 ix35760 (.Y (nx35761), .A (nx38445)) ;
    inv01 ix35762 (.Y (nx35763), .A (nx38445)) ;
    inv01 ix35764 (.Y (nx35765), .A (nx38445)) ;
    inv01 ix35766 (.Y (nx35767), .A (nx38445)) ;
    inv01 ix35768 (.Y (nx35769), .A (nx38445)) ;
    inv01 ix35770 (.Y (nx35771), .A (nx38445)) ;
    inv01 ix35772 (.Y (nx35773), .A (nx38447)) ;
    inv01 ix35774 (.Y (nx35775), .A (nx38447)) ;
    inv01 ix35776 (.Y (nx35777), .A (nx38447)) ;
    inv01 ix35778 (.Y (nx35779), .A (nx38447)) ;
    inv01 ix35780 (.Y (nx35781), .A (nx38447)) ;
    inv01 ix35782 (.Y (nx35783), .A (nx38447)) ;
    inv01 ix35784 (.Y (nx35785), .A (nx38447)) ;
    inv01 ix35786 (.Y (nx35787), .A (nx38449)) ;
    inv01 ix35788 (.Y (nx35789), .A (nx38449)) ;
    inv01 ix35790 (.Y (nx35791), .A (nx38449)) ;
    inv01 ix35792 (.Y (nx35793), .A (nx38449)) ;
    inv01 ix35794 (.Y (nx35795), .A (nx38449)) ;
    inv01 ix35796 (.Y (nx35797), .A (nx38449)) ;
    inv01 ix35798 (.Y (nx35799), .A (nx38449)) ;
    inv01 ix35800 (.Y (nx35801), .A (nx38451)) ;
    inv01 ix35802 (.Y (nx35803), .A (nx38451)) ;
    inv01 ix35804 (.Y (nx35805), .A (nx38451)) ;
    inv01 ix35806 (.Y (nx35807), .A (nx38451)) ;
    inv01 ix35808 (.Y (nx35809), .A (nx38451)) ;
    inv01 ix35810 (.Y (nx35811), .A (nx38451)) ;
    inv01 ix35812 (.Y (nx35813), .A (nx38451)) ;
    inv01 ix35814 (.Y (nx35815), .A (nx38453)) ;
    inv01 ix35816 (.Y (nx35817), .A (nx38453)) ;
    inv01 ix35818 (.Y (nx35819), .A (nx38453)) ;
    inv01 ix35820 (.Y (nx35821), .A (nx38453)) ;
    inv01 ix35822 (.Y (nx35823), .A (nx38453)) ;
    inv01 ix35824 (.Y (nx35825), .A (nx38453)) ;
    inv01 ix35826 (.Y (nx35827), .A (nx38453)) ;
    inv01 ix35828 (.Y (nx35829), .A (nx38455)) ;
    inv01 ix35830 (.Y (nx35831), .A (nx38455)) ;
    inv01 ix35832 (.Y (nx35833), .A (nx38455)) ;
    inv01 ix35834 (.Y (nx35835), .A (nx38455)) ;
    inv01 ix35836 (.Y (nx35837), .A (nx38455)) ;
    inv01 ix35838 (.Y (nx35839), .A (nx38455)) ;
    inv01 ix35840 (.Y (nx35841), .A (nx38455)) ;
    inv01 ix35842 (.Y (nx35843), .A (nx38457)) ;
    inv01 ix35844 (.Y (nx35845), .A (nx38457)) ;
    inv01 ix35846 (.Y (nx35847), .A (nx38457)) ;
    inv01 ix35848 (.Y (nx35849), .A (nx38457)) ;
    inv01 ix35850 (.Y (nx35851), .A (nx38457)) ;
    inv01 ix35852 (.Y (nx35853), .A (nx38457)) ;
    inv01 ix35854 (.Y (nx35855), .A (nx38457)) ;
    inv01 ix35856 (.Y (nx35857), .A (nx38459)) ;
    inv01 ix35858 (.Y (nx35859), .A (nx38459)) ;
    inv01 ix35860 (.Y (nx35861), .A (nx38459)) ;
    inv01 ix35862 (.Y (nx35863), .A (nx38459)) ;
    inv01 ix35864 (.Y (nx35865), .A (nx38459)) ;
    inv01 ix35866 (.Y (nx35867), .A (nx38459)) ;
    inv01 ix35868 (.Y (nx35869), .A (nx38459)) ;
    inv01 ix35870 (.Y (nx35871), .A (nx35603)) ;
    inv01 ix35872 (.Y (nx35873), .A (nx35603)) ;
    inv01 ix35874 (.Y (nx35875), .A (nx35603)) ;
    inv01 ix35876 (.Y (nx35877), .A (nx35603)) ;
    inv01 ix35878 (.Y (nx35879), .A (nx35603)) ;
    inv01 ix35880 (.Y (nx35881), .A (nx35603)) ;
    inv02 ix35884 (.Y (nx35885), .A (nx38461)) ;
    inv02 ix35886 (.Y (nx35887), .A (nx38461)) ;
    inv02 ix35888 (.Y (nx35889), .A (nx38461)) ;
    inv02 ix35890 (.Y (nx35891), .A (nx38461)) ;
    inv02 ix35892 (.Y (nx35893), .A (nx38461)) ;
    inv02 ix35894 (.Y (nx35895), .A (nx38461)) ;
    inv02 ix35896 (.Y (nx35897), .A (nx38461)) ;
    inv02 ix35898 (.Y (nx35899), .A (nx38463)) ;
    inv02 ix35900 (.Y (nx35901), .A (nx38463)) ;
    inv02 ix35902 (.Y (nx35903), .A (nx38463)) ;
    inv02 ix35904 (.Y (nx35905), .A (nx38463)) ;
    inv02 ix35906 (.Y (nx35907), .A (nx38463)) ;
    inv02 ix35908 (.Y (nx35909), .A (nx38463)) ;
    inv02 ix35910 (.Y (nx35911), .A (nx38463)) ;
    inv02 ix35912 (.Y (nx35913), .A (nx38465)) ;
    inv02 ix35914 (.Y (nx35915), .A (nx38465)) ;
    inv02 ix35916 (.Y (nx35917), .A (nx38465)) ;
    inv02 ix35918 (.Y (nx35919), .A (nx38465)) ;
    inv02 ix35920 (.Y (nx35921), .A (nx38465)) ;
    inv02 ix35922 (.Y (nx35923), .A (nx38465)) ;
    inv02 ix35924 (.Y (nx35925), .A (nx38465)) ;
    inv02 ix35926 (.Y (nx35927), .A (nx38467)) ;
    inv02 ix35928 (.Y (nx35929), .A (nx38467)) ;
    inv02 ix35930 (.Y (nx35931), .A (nx38467)) ;
    inv02 ix35932 (.Y (nx35933), .A (nx38467)) ;
    inv02 ix35934 (.Y (nx35935), .A (nx38467)) ;
    inv02 ix35936 (.Y (nx35937), .A (nx38467)) ;
    inv02 ix35938 (.Y (nx35939), .A (nx38467)) ;
    inv02 ix35940 (.Y (nx35941), .A (nx38469)) ;
    inv02 ix35942 (.Y (nx35943), .A (nx38469)) ;
    inv02 ix35944 (.Y (nx35945), .A (nx38469)) ;
    inv02 ix35946 (.Y (nx35947), .A (nx38469)) ;
    inv02 ix35948 (.Y (nx35949), .A (nx38469)) ;
    inv02 ix35950 (.Y (nx35951), .A (nx38469)) ;
    inv02 ix35952 (.Y (nx35953), .A (nx38469)) ;
    inv02 ix35954 (.Y (nx35955), .A (nx38471)) ;
    inv02 ix35956 (.Y (nx35957), .A (nx38471)) ;
    inv02 ix35958 (.Y (nx35959), .A (nx38471)) ;
    inv02 ix35960 (.Y (nx35961), .A (nx38471)) ;
    inv02 ix35962 (.Y (nx35963), .A (nx38471)) ;
    inv02 ix35964 (.Y (nx35965), .A (nx38471)) ;
    inv02 ix35966 (.Y (nx35967), .A (nx38471)) ;
    inv02 ix35968 (.Y (nx35969), .A (nx38473)) ;
    inv02 ix35970 (.Y (nx35971), .A (nx38473)) ;
    inv02 ix35972 (.Y (nx35973), .A (nx38473)) ;
    inv02 ix35974 (.Y (nx35975), .A (nx38473)) ;
    inv02 ix35976 (.Y (nx35977), .A (nx38473)) ;
    inv02 ix35978 (.Y (nx35979), .A (nx38473)) ;
    inv02 ix35980 (.Y (nx35981), .A (nx38473)) ;
    inv02 ix35982 (.Y (nx35983), .A (nx38475)) ;
    inv02 ix35984 (.Y (nx35985), .A (nx38475)) ;
    inv02 ix35986 (.Y (nx35987), .A (nx38475)) ;
    inv02 ix35988 (.Y (nx35989), .A (nx38475)) ;
    inv02 ix35990 (.Y (nx35991), .A (nx38475)) ;
    inv02 ix35992 (.Y (nx35993), .A (nx38475)) ;
    inv02 ix35994 (.Y (nx35995), .A (nx38475)) ;
    inv02 ix35996 (.Y (nx35997), .A (nx38477)) ;
    inv02 ix35998 (.Y (nx35999), .A (nx38477)) ;
    inv02 ix36000 (.Y (nx36001), .A (nx38477)) ;
    inv02 ix36002 (.Y (nx36003), .A (nx38477)) ;
    inv02 ix36004 (.Y (nx36005), .A (nx38477)) ;
    inv02 ix36006 (.Y (nx36007), .A (nx38477)) ;
    inv02 ix36008 (.Y (nx36009), .A (nx38477)) ;
    inv02 ix36010 (.Y (nx36011), .A (nx38479)) ;
    inv02 ix36012 (.Y (nx36013), .A (nx38479)) ;
    inv02 ix36014 (.Y (nx36015), .A (nx38479)) ;
    inv02 ix36016 (.Y (nx36017), .A (nx38479)) ;
    inv02 ix36018 (.Y (nx36019), .A (nx38479)) ;
    inv02 ix36020 (.Y (nx36021), .A (nx38479)) ;
    inv02 ix36022 (.Y (nx36023), .A (nx38479)) ;
    inv02 ix36026 (.Y (nx36027), .A (nx38481)) ;
    inv02 ix36028 (.Y (nx36029), .A (nx38481)) ;
    inv02 ix36030 (.Y (nx36031), .A (nx38481)) ;
    inv02 ix36032 (.Y (nx36033), .A (nx38481)) ;
    inv02 ix36034 (.Y (nx36035), .A (nx38481)) ;
    inv02 ix36036 (.Y (nx36037), .A (nx38481)) ;
    inv02 ix36038 (.Y (nx36039), .A (nx38481)) ;
    inv02 ix36040 (.Y (nx36041), .A (nx38483)) ;
    inv02 ix36042 (.Y (nx36043), .A (nx38483)) ;
    inv02 ix36044 (.Y (nx36045), .A (nx38483)) ;
    inv02 ix36046 (.Y (nx36047), .A (nx38483)) ;
    inv02 ix36048 (.Y (nx36049), .A (nx38483)) ;
    inv02 ix36050 (.Y (nx36051), .A (nx38483)) ;
    inv02 ix36052 (.Y (nx36053), .A (nx38483)) ;
    inv02 ix36054 (.Y (nx36055), .A (nx38485)) ;
    inv02 ix36056 (.Y (nx36057), .A (nx38485)) ;
    inv02 ix36058 (.Y (nx36059), .A (nx38485)) ;
    inv02 ix36060 (.Y (nx36061), .A (nx38485)) ;
    inv02 ix36062 (.Y (nx36063), .A (nx38485)) ;
    inv02 ix36064 (.Y (nx36065), .A (nx38485)) ;
    inv02 ix36066 (.Y (nx36067), .A (nx38485)) ;
    inv02 ix36068 (.Y (nx36069), .A (nx38487)) ;
    inv02 ix36070 (.Y (nx36071), .A (nx38487)) ;
    inv02 ix36072 (.Y (nx36073), .A (nx38487)) ;
    inv02 ix36074 (.Y (nx36075), .A (nx38487)) ;
    inv02 ix36076 (.Y (nx36077), .A (nx38487)) ;
    inv02 ix36078 (.Y (nx36079), .A (nx38487)) ;
    inv02 ix36080 (.Y (nx36081), .A (nx38487)) ;
    inv02 ix36082 (.Y (nx36083), .A (nx38489)) ;
    inv02 ix36084 (.Y (nx36085), .A (nx38489)) ;
    inv02 ix36086 (.Y (nx36087), .A (nx38489)) ;
    inv02 ix36088 (.Y (nx36089), .A (nx38489)) ;
    inv02 ix36090 (.Y (nx36091), .A (nx38489)) ;
    inv02 ix36092 (.Y (nx36093), .A (nx38489)) ;
    inv02 ix36094 (.Y (nx36095), .A (nx38489)) ;
    inv02 ix36096 (.Y (nx36097), .A (nx38491)) ;
    inv02 ix36098 (.Y (nx36099), .A (nx38491)) ;
    inv02 ix36100 (.Y (nx36101), .A (nx38491)) ;
    inv02 ix36102 (.Y (nx36103), .A (nx38491)) ;
    inv02 ix36104 (.Y (nx36105), .A (nx38491)) ;
    inv02 ix36106 (.Y (nx36107), .A (nx38491)) ;
    inv02 ix36108 (.Y (nx36109), .A (nx38491)) ;
    inv02 ix36110 (.Y (nx36111), .A (nx38493)) ;
    inv02 ix36112 (.Y (nx36113), .A (nx38493)) ;
    inv02 ix36114 (.Y (nx36115), .A (nx38493)) ;
    inv02 ix36116 (.Y (nx36117), .A (nx38493)) ;
    inv02 ix36118 (.Y (nx36119), .A (nx38493)) ;
    inv02 ix36120 (.Y (nx36121), .A (nx38493)) ;
    inv02 ix36122 (.Y (nx36123), .A (nx38493)) ;
    inv02 ix36124 (.Y (nx36125), .A (nx38495)) ;
    inv02 ix36126 (.Y (nx36127), .A (nx38495)) ;
    inv02 ix36128 (.Y (nx36129), .A (nx38495)) ;
    inv02 ix36130 (.Y (nx36131), .A (nx38495)) ;
    inv02 ix36132 (.Y (nx36133), .A (nx38495)) ;
    inv02 ix36134 (.Y (nx36135), .A (nx38495)) ;
    inv02 ix36136 (.Y (nx36137), .A (nx38495)) ;
    inv02 ix36138 (.Y (nx36139), .A (nx38497)) ;
    inv02 ix36140 (.Y (nx36141), .A (nx38497)) ;
    inv02 ix36142 (.Y (nx36143), .A (nx38497)) ;
    inv02 ix36144 (.Y (nx36145), .A (nx38497)) ;
    inv02 ix36146 (.Y (nx36147), .A (nx38497)) ;
    inv02 ix36148 (.Y (nx36149), .A (nx38497)) ;
    inv02 ix36150 (.Y (nx36151), .A (nx38497)) ;
    inv02 ix36152 (.Y (nx36153), .A (nx38499)) ;
    inv02 ix36154 (.Y (nx36155), .A (nx38499)) ;
    inv02 ix36156 (.Y (nx36157), .A (nx38499)) ;
    inv02 ix36158 (.Y (nx36159), .A (nx38499)) ;
    inv02 ix36160 (.Y (nx36161), .A (nx38499)) ;
    inv02 ix36162 (.Y (nx36163), .A (nx38499)) ;
    inv02 ix36164 (.Y (nx36165), .A (nx38499)) ;
    inv02 ix36168 (.Y (nx36169), .A (nx38501)) ;
    inv02 ix36170 (.Y (nx36171), .A (nx38501)) ;
    inv02 ix36172 (.Y (nx36173), .A (nx38501)) ;
    inv02 ix36174 (.Y (nx36175), .A (nx38501)) ;
    inv02 ix36176 (.Y (nx36177), .A (nx38501)) ;
    inv02 ix36178 (.Y (nx36179), .A (nx38501)) ;
    inv02 ix36180 (.Y (nx36181), .A (nx38501)) ;
    inv02 ix36182 (.Y (nx36183), .A (nx38503)) ;
    inv02 ix36184 (.Y (nx36185), .A (nx38503)) ;
    inv02 ix36186 (.Y (nx36187), .A (nx38503)) ;
    inv02 ix36188 (.Y (nx36189), .A (nx38503)) ;
    inv02 ix36190 (.Y (nx36191), .A (nx38503)) ;
    inv02 ix36192 (.Y (nx36193), .A (nx38503)) ;
    inv02 ix36194 (.Y (nx36195), .A (nx38503)) ;
    inv02 ix36196 (.Y (nx36197), .A (nx38505)) ;
    inv02 ix36198 (.Y (nx36199), .A (nx38505)) ;
    inv02 ix36200 (.Y (nx36201), .A (nx38505)) ;
    inv02 ix36202 (.Y (nx36203), .A (nx38505)) ;
    inv02 ix36204 (.Y (nx36205), .A (nx38505)) ;
    inv02 ix36206 (.Y (nx36207), .A (nx38505)) ;
    inv02 ix36208 (.Y (nx36209), .A (nx38505)) ;
    inv02 ix36210 (.Y (nx36211), .A (nx38507)) ;
    inv02 ix36212 (.Y (nx36213), .A (nx38507)) ;
    inv02 ix36214 (.Y (nx36215), .A (nx38507)) ;
    inv02 ix36216 (.Y (nx36217), .A (nx38507)) ;
    inv02 ix36218 (.Y (nx36219), .A (nx38507)) ;
    inv02 ix36220 (.Y (nx36221), .A (nx38507)) ;
    inv02 ix36222 (.Y (nx36223), .A (nx38507)) ;
    inv02 ix36224 (.Y (nx36225), .A (nx38509)) ;
    inv02 ix36226 (.Y (nx36227), .A (nx38509)) ;
    inv02 ix36228 (.Y (nx36229), .A (nx38509)) ;
    inv02 ix36230 (.Y (nx36231), .A (nx38509)) ;
    inv02 ix36232 (.Y (nx36233), .A (nx38509)) ;
    inv02 ix36234 (.Y (nx36235), .A (nx38509)) ;
    inv02 ix36236 (.Y (nx36237), .A (nx38509)) ;
    inv02 ix36238 (.Y (nx36239), .A (nx38511)) ;
    inv02 ix36240 (.Y (nx36241), .A (nx38511)) ;
    inv02 ix36242 (.Y (nx36243), .A (nx38511)) ;
    inv02 ix36244 (.Y (nx36245), .A (nx38511)) ;
    inv02 ix36246 (.Y (nx36247), .A (nx38511)) ;
    inv02 ix36248 (.Y (nx36249), .A (nx38511)) ;
    inv02 ix36250 (.Y (nx36251), .A (nx38511)) ;
    inv02 ix36252 (.Y (nx36253), .A (nx38513)) ;
    inv02 ix36254 (.Y (nx36255), .A (nx38513)) ;
    inv02 ix36256 (.Y (nx36257), .A (nx38513)) ;
    inv02 ix36258 (.Y (nx36259), .A (nx38513)) ;
    inv02 ix36260 (.Y (nx36261), .A (nx38513)) ;
    inv02 ix36262 (.Y (nx36263), .A (nx38513)) ;
    inv02 ix36264 (.Y (nx36265), .A (nx38513)) ;
    inv02 ix36266 (.Y (nx36267), .A (nx38515)) ;
    inv02 ix36268 (.Y (nx36269), .A (nx38515)) ;
    inv02 ix36270 (.Y (nx36271), .A (nx38515)) ;
    inv02 ix36272 (.Y (nx36273), .A (nx38515)) ;
    inv02 ix36274 (.Y (nx36275), .A (nx38515)) ;
    inv02 ix36276 (.Y (nx36277), .A (nx38515)) ;
    inv02 ix36278 (.Y (nx36279), .A (nx38515)) ;
    inv02 ix36280 (.Y (nx36281), .A (nx38517)) ;
    inv02 ix36282 (.Y (nx36283), .A (nx38517)) ;
    inv02 ix36284 (.Y (nx36285), .A (nx38517)) ;
    inv02 ix36286 (.Y (nx36287), .A (nx38517)) ;
    inv02 ix36288 (.Y (nx36289), .A (nx38517)) ;
    inv02 ix36290 (.Y (nx36291), .A (nx38517)) ;
    inv02 ix36292 (.Y (nx36293), .A (nx38517)) ;
    inv02 ix36294 (.Y (nx36295), .A (nx38519)) ;
    inv02 ix36296 (.Y (nx36297), .A (nx38519)) ;
    inv02 ix36298 (.Y (nx36299), .A (nx38519)) ;
    inv02 ix36300 (.Y (nx36301), .A (nx38519)) ;
    inv02 ix36302 (.Y (nx36303), .A (nx38519)) ;
    inv02 ix36304 (.Y (nx36305), .A (nx38519)) ;
    inv02 ix36306 (.Y (nx36307), .A (nx38519)) ;
    inv02 ix36310 (.Y (nx36311), .A (nx38521)) ;
    inv02 ix36312 (.Y (nx36313), .A (nx38521)) ;
    inv02 ix36314 (.Y (nx36315), .A (nx38521)) ;
    inv02 ix36316 (.Y (nx36317), .A (nx38521)) ;
    inv02 ix36318 (.Y (nx36319), .A (nx38521)) ;
    inv02 ix36320 (.Y (nx36321), .A (nx38521)) ;
    inv02 ix36322 (.Y (nx36323), .A (nx38521)) ;
    inv02 ix36324 (.Y (nx36325), .A (nx38523)) ;
    inv02 ix36326 (.Y (nx36327), .A (nx38523)) ;
    inv02 ix36328 (.Y (nx36329), .A (nx38523)) ;
    inv02 ix36330 (.Y (nx36331), .A (nx38523)) ;
    inv02 ix36332 (.Y (nx36333), .A (nx38523)) ;
    inv02 ix36334 (.Y (nx36335), .A (nx38523)) ;
    inv02 ix36336 (.Y (nx36337), .A (nx38523)) ;
    inv02 ix36338 (.Y (nx36339), .A (nx38525)) ;
    inv02 ix36340 (.Y (nx36341), .A (nx38525)) ;
    inv02 ix36342 (.Y (nx36343), .A (nx38525)) ;
    inv02 ix36344 (.Y (nx36345), .A (nx38525)) ;
    inv02 ix36346 (.Y (nx36347), .A (nx38525)) ;
    inv02 ix36348 (.Y (nx36349), .A (nx38525)) ;
    inv02 ix36350 (.Y (nx36351), .A (nx38525)) ;
    inv02 ix36352 (.Y (nx36353), .A (nx38527)) ;
    inv02 ix36354 (.Y (nx36355), .A (nx38527)) ;
    inv02 ix36356 (.Y (nx36357), .A (nx38527)) ;
    inv02 ix36358 (.Y (nx36359), .A (nx38527)) ;
    inv02 ix36360 (.Y (nx36361), .A (nx38527)) ;
    inv02 ix36362 (.Y (nx36363), .A (nx38527)) ;
    inv02 ix36364 (.Y (nx36365), .A (nx38527)) ;
    inv02 ix36366 (.Y (nx36367), .A (nx38529)) ;
    inv02 ix36368 (.Y (nx36369), .A (nx38529)) ;
    inv02 ix36370 (.Y (nx36371), .A (nx38529)) ;
    inv02 ix36372 (.Y (nx36373), .A (nx38529)) ;
    inv02 ix36374 (.Y (nx36375), .A (nx38529)) ;
    inv02 ix36376 (.Y (nx36377), .A (nx38529)) ;
    inv02 ix36378 (.Y (nx36379), .A (nx38529)) ;
    inv02 ix36380 (.Y (nx36381), .A (nx38531)) ;
    inv02 ix36382 (.Y (nx36383), .A (nx38531)) ;
    inv02 ix36384 (.Y (nx36385), .A (nx38531)) ;
    inv02 ix36386 (.Y (nx36387), .A (nx38531)) ;
    inv02 ix36388 (.Y (nx36389), .A (nx38531)) ;
    inv02 ix36390 (.Y (nx36391), .A (nx38531)) ;
    inv02 ix36392 (.Y (nx36393), .A (nx38531)) ;
    inv02 ix36394 (.Y (nx36395), .A (nx38533)) ;
    inv02 ix36396 (.Y (nx36397), .A (nx38533)) ;
    inv02 ix36398 (.Y (nx36399), .A (nx38533)) ;
    inv02 ix36400 (.Y (nx36401), .A (nx38533)) ;
    inv02 ix36402 (.Y (nx36403), .A (nx38533)) ;
    inv02 ix36404 (.Y (nx36405), .A (nx38533)) ;
    inv02 ix36406 (.Y (nx36407), .A (nx38533)) ;
    inv02 ix36408 (.Y (nx36409), .A (nx38535)) ;
    inv02 ix36410 (.Y (nx36411), .A (nx38535)) ;
    inv02 ix36412 (.Y (nx36413), .A (nx38535)) ;
    inv02 ix36414 (.Y (nx36415), .A (nx38535)) ;
    inv02 ix36416 (.Y (nx36417), .A (nx38535)) ;
    inv02 ix36418 (.Y (nx36419), .A (nx38535)) ;
    inv02 ix36420 (.Y (nx36421), .A (nx38535)) ;
    inv02 ix36422 (.Y (nx36423), .A (nx38537)) ;
    inv02 ix36424 (.Y (nx36425), .A (nx38537)) ;
    inv02 ix36426 (.Y (nx36427), .A (nx38537)) ;
    inv02 ix36428 (.Y (nx36429), .A (nx38537)) ;
    inv02 ix36430 (.Y (nx36431), .A (nx38537)) ;
    inv02 ix36432 (.Y (nx36433), .A (nx38537)) ;
    inv02 ix36434 (.Y (nx36435), .A (nx38537)) ;
    inv02 ix36436 (.Y (nx36437), .A (nx38539)) ;
    inv02 ix36438 (.Y (nx36439), .A (nx38539)) ;
    inv02 ix36440 (.Y (nx36441), .A (nx38539)) ;
    inv02 ix36442 (.Y (nx36443), .A (nx38539)) ;
    inv02 ix36444 (.Y (nx36445), .A (nx38539)) ;
    inv02 ix36446 (.Y (nx36447), .A (nx38539)) ;
    inv02 ix36448 (.Y (nx36449), .A (nx38539)) ;
    inv02 ix36452 (.Y (nx36453), .A (nx38541)) ;
    inv02 ix36454 (.Y (nx36455), .A (nx38541)) ;
    inv02 ix36456 (.Y (nx36457), .A (nx38541)) ;
    inv02 ix36458 (.Y (nx36459), .A (nx38541)) ;
    inv02 ix36460 (.Y (nx36461), .A (nx38541)) ;
    inv02 ix36462 (.Y (nx36463), .A (nx38541)) ;
    inv02 ix36464 (.Y (nx36465), .A (nx38541)) ;
    inv02 ix36466 (.Y (nx36467), .A (nx38543)) ;
    inv02 ix36468 (.Y (nx36469), .A (nx38543)) ;
    inv02 ix36470 (.Y (nx36471), .A (nx38543)) ;
    inv02 ix36472 (.Y (nx36473), .A (nx38543)) ;
    inv02 ix36474 (.Y (nx36475), .A (nx38543)) ;
    inv02 ix36476 (.Y (nx36477), .A (nx38543)) ;
    inv02 ix36478 (.Y (nx36479), .A (nx38543)) ;
    inv02 ix36480 (.Y (nx36481), .A (nx38545)) ;
    inv02 ix36482 (.Y (nx36483), .A (nx38545)) ;
    inv02 ix36484 (.Y (nx36485), .A (nx38545)) ;
    inv02 ix36486 (.Y (nx36487), .A (nx38545)) ;
    inv02 ix36488 (.Y (nx36489), .A (nx38545)) ;
    inv02 ix36490 (.Y (nx36491), .A (nx38545)) ;
    inv02 ix36492 (.Y (nx36493), .A (nx38545)) ;
    inv02 ix36494 (.Y (nx36495), .A (nx38547)) ;
    inv02 ix36496 (.Y (nx36497), .A (nx38547)) ;
    inv02 ix36498 (.Y (nx36499), .A (nx38547)) ;
    inv02 ix36500 (.Y (nx36501), .A (nx38547)) ;
    inv02 ix36502 (.Y (nx36503), .A (nx38547)) ;
    inv02 ix36504 (.Y (nx36505), .A (nx38547)) ;
    inv02 ix36506 (.Y (nx36507), .A (nx38547)) ;
    inv02 ix36508 (.Y (nx36509), .A (nx38549)) ;
    inv02 ix36510 (.Y (nx36511), .A (nx38549)) ;
    inv02 ix36512 (.Y (nx36513), .A (nx38549)) ;
    inv02 ix36514 (.Y (nx36515), .A (nx38549)) ;
    inv02 ix36516 (.Y (nx36517), .A (nx38549)) ;
    inv02 ix36518 (.Y (nx36519), .A (nx38549)) ;
    inv02 ix36520 (.Y (nx36521), .A (nx38549)) ;
    inv02 ix36522 (.Y (nx36523), .A (nx38551)) ;
    inv02 ix36524 (.Y (nx36525), .A (nx38551)) ;
    inv02 ix36526 (.Y (nx36527), .A (nx38551)) ;
    inv02 ix36528 (.Y (nx36529), .A (nx38551)) ;
    inv02 ix36530 (.Y (nx36531), .A (nx38551)) ;
    inv02 ix36532 (.Y (nx36533), .A (nx38551)) ;
    inv02 ix36534 (.Y (nx36535), .A (nx38551)) ;
    inv02 ix36536 (.Y (nx36537), .A (nx38553)) ;
    inv02 ix36538 (.Y (nx36539), .A (nx38553)) ;
    inv02 ix36540 (.Y (nx36541), .A (nx38553)) ;
    inv02 ix36542 (.Y (nx36543), .A (nx38553)) ;
    inv02 ix36544 (.Y (nx36545), .A (nx38553)) ;
    inv02 ix36546 (.Y (nx36547), .A (nx38553)) ;
    inv02 ix36548 (.Y (nx36549), .A (nx38553)) ;
    inv02 ix36550 (.Y (nx36551), .A (nx38555)) ;
    inv02 ix36552 (.Y (nx36553), .A (nx38555)) ;
    inv02 ix36554 (.Y (nx36555), .A (nx38555)) ;
    inv02 ix36556 (.Y (nx36557), .A (nx38555)) ;
    inv02 ix36558 (.Y (nx36559), .A (nx38555)) ;
    inv02 ix36560 (.Y (nx36561), .A (nx38555)) ;
    inv02 ix36562 (.Y (nx36563), .A (nx38555)) ;
    inv02 ix36564 (.Y (nx36565), .A (nx38557)) ;
    inv02 ix36566 (.Y (nx36567), .A (nx38557)) ;
    inv02 ix36568 (.Y (nx36569), .A (nx38557)) ;
    inv02 ix36570 (.Y (nx36571), .A (nx38557)) ;
    inv02 ix36572 (.Y (nx36573), .A (nx38557)) ;
    inv02 ix36574 (.Y (nx36575), .A (nx38557)) ;
    inv02 ix36576 (.Y (nx36577), .A (nx38557)) ;
    inv02 ix36578 (.Y (nx36579), .A (nx38559)) ;
    inv02 ix36580 (.Y (nx36581), .A (nx38559)) ;
    inv02 ix36582 (.Y (nx36583), .A (nx38559)) ;
    inv02 ix36584 (.Y (nx36585), .A (nx38559)) ;
    inv02 ix36586 (.Y (nx36587), .A (nx38559)) ;
    inv02 ix36588 (.Y (nx36589), .A (nx38559)) ;
    inv02 ix36590 (.Y (nx36591), .A (nx38559)) ;
    inv02 ix36594 (.Y (nx36595), .A (nx38561)) ;
    inv02 ix36596 (.Y (nx36597), .A (nx38561)) ;
    inv02 ix36598 (.Y (nx36599), .A (nx38561)) ;
    inv02 ix36600 (.Y (nx36601), .A (nx38561)) ;
    inv02 ix36602 (.Y (nx36603), .A (nx38561)) ;
    inv02 ix36604 (.Y (nx36605), .A (nx38561)) ;
    inv02 ix36606 (.Y (nx36607), .A (nx38561)) ;
    inv02 ix36608 (.Y (nx36609), .A (nx38563)) ;
    inv02 ix36610 (.Y (nx36611), .A (nx38563)) ;
    inv02 ix36612 (.Y (nx36613), .A (nx38563)) ;
    inv02 ix36614 (.Y (nx36615), .A (nx38563)) ;
    inv02 ix36616 (.Y (nx36617), .A (nx38563)) ;
    inv02 ix36618 (.Y (nx36619), .A (nx38563)) ;
    inv02 ix36620 (.Y (nx36621), .A (nx38563)) ;
    inv02 ix36622 (.Y (nx36623), .A (nx38565)) ;
    inv02 ix36624 (.Y (nx36625), .A (nx38565)) ;
    inv02 ix36626 (.Y (nx36627), .A (nx38565)) ;
    inv02 ix36628 (.Y (nx36629), .A (nx38565)) ;
    inv02 ix36630 (.Y (nx36631), .A (nx38565)) ;
    inv02 ix36632 (.Y (nx36633), .A (nx38565)) ;
    inv02 ix36634 (.Y (nx36635), .A (nx38565)) ;
    inv02 ix36636 (.Y (nx36637), .A (nx38567)) ;
    inv02 ix36638 (.Y (nx36639), .A (nx38567)) ;
    inv02 ix36640 (.Y (nx36641), .A (nx38567)) ;
    inv02 ix36642 (.Y (nx36643), .A (nx38567)) ;
    inv02 ix36644 (.Y (nx36645), .A (nx38567)) ;
    inv02 ix36646 (.Y (nx36647), .A (nx38567)) ;
    inv02 ix36648 (.Y (nx36649), .A (nx38567)) ;
    inv02 ix36650 (.Y (nx36651), .A (nx38569)) ;
    inv02 ix36652 (.Y (nx36653), .A (nx38569)) ;
    inv02 ix36654 (.Y (nx36655), .A (nx38569)) ;
    inv02 ix36656 (.Y (nx36657), .A (nx38569)) ;
    inv02 ix36658 (.Y (nx36659), .A (nx38569)) ;
    inv02 ix36660 (.Y (nx36661), .A (nx38569)) ;
    inv02 ix36662 (.Y (nx36663), .A (nx38569)) ;
    inv02 ix36664 (.Y (nx36665), .A (nx38571)) ;
    inv02 ix36666 (.Y (nx36667), .A (nx38571)) ;
    inv02 ix36668 (.Y (nx36669), .A (nx38571)) ;
    inv02 ix36670 (.Y (nx36671), .A (nx38571)) ;
    inv02 ix36672 (.Y (nx36673), .A (nx38571)) ;
    inv02 ix36674 (.Y (nx36675), .A (nx38571)) ;
    inv02 ix36676 (.Y (nx36677), .A (nx38571)) ;
    inv02 ix36678 (.Y (nx36679), .A (nx38573)) ;
    inv02 ix36680 (.Y (nx36681), .A (nx38573)) ;
    inv02 ix36682 (.Y (nx36683), .A (nx38573)) ;
    inv02 ix36684 (.Y (nx36685), .A (nx38573)) ;
    inv02 ix36686 (.Y (nx36687), .A (nx38573)) ;
    inv02 ix36688 (.Y (nx36689), .A (nx38573)) ;
    inv02 ix36690 (.Y (nx36691), .A (nx38573)) ;
    inv02 ix36692 (.Y (nx36693), .A (nx38575)) ;
    inv02 ix36694 (.Y (nx36695), .A (nx38575)) ;
    inv02 ix36696 (.Y (nx36697), .A (nx38575)) ;
    inv02 ix36698 (.Y (nx36699), .A (nx38575)) ;
    inv02 ix36700 (.Y (nx36701), .A (nx38575)) ;
    inv02 ix36702 (.Y (nx36703), .A (nx38575)) ;
    inv02 ix36704 (.Y (nx36705), .A (nx38575)) ;
    inv02 ix36706 (.Y (nx36707), .A (nx38577)) ;
    inv02 ix36708 (.Y (nx36709), .A (nx38577)) ;
    inv02 ix36710 (.Y (nx36711), .A (nx38577)) ;
    inv02 ix36712 (.Y (nx36713), .A (nx38577)) ;
    inv02 ix36714 (.Y (nx36715), .A (nx38577)) ;
    inv02 ix36716 (.Y (nx36717), .A (nx38577)) ;
    inv02 ix36718 (.Y (nx36719), .A (nx38577)) ;
    inv02 ix36720 (.Y (nx36721), .A (nx38579)) ;
    inv02 ix36722 (.Y (nx36723), .A (nx38579)) ;
    inv02 ix36724 (.Y (nx36725), .A (nx38579)) ;
    inv02 ix36726 (.Y (nx36727), .A (nx38579)) ;
    inv02 ix36728 (.Y (nx36729), .A (nx38579)) ;
    inv02 ix36730 (.Y (nx36731), .A (nx38579)) ;
    inv02 ix36732 (.Y (nx36733), .A (nx38579)) ;
    inv02 ix36736 (.Y (nx36737), .A (nx38581)) ;
    inv02 ix36738 (.Y (nx36739), .A (nx38581)) ;
    inv02 ix36740 (.Y (nx36741), .A (nx38581)) ;
    inv02 ix36742 (.Y (nx36743), .A (nx38581)) ;
    inv02 ix36744 (.Y (nx36745), .A (nx38581)) ;
    inv02 ix36746 (.Y (nx36747), .A (nx38581)) ;
    inv02 ix36748 (.Y (nx36749), .A (nx38581)) ;
    inv02 ix36750 (.Y (nx36751), .A (nx38583)) ;
    inv02 ix36752 (.Y (nx36753), .A (nx38583)) ;
    inv02 ix36754 (.Y (nx36755), .A (nx38583)) ;
    inv02 ix36756 (.Y (nx36757), .A (nx38583)) ;
    inv02 ix36758 (.Y (nx36759), .A (nx38583)) ;
    inv02 ix36760 (.Y (nx36761), .A (nx38583)) ;
    inv02 ix36762 (.Y (nx36763), .A (nx38583)) ;
    inv02 ix36764 (.Y (nx36765), .A (nx38585)) ;
    inv02 ix36766 (.Y (nx36767), .A (nx38585)) ;
    inv02 ix36768 (.Y (nx36769), .A (nx38585)) ;
    inv02 ix36770 (.Y (nx36771), .A (nx38585)) ;
    inv02 ix36772 (.Y (nx36773), .A (nx38585)) ;
    inv02 ix36774 (.Y (nx36775), .A (nx38585)) ;
    inv02 ix36776 (.Y (nx36777), .A (nx38585)) ;
    inv02 ix36778 (.Y (nx36779), .A (nx38587)) ;
    inv02 ix36780 (.Y (nx36781), .A (nx38587)) ;
    inv02 ix36782 (.Y (nx36783), .A (nx38587)) ;
    inv02 ix36784 (.Y (nx36785), .A (nx38587)) ;
    inv02 ix36786 (.Y (nx36787), .A (nx38587)) ;
    inv02 ix36788 (.Y (nx36789), .A (nx38587)) ;
    inv02 ix36790 (.Y (nx36791), .A (nx38587)) ;
    inv02 ix36792 (.Y (nx36793), .A (nx38589)) ;
    inv02 ix36794 (.Y (nx36795), .A (nx38589)) ;
    inv02 ix36796 (.Y (nx36797), .A (nx38589)) ;
    inv02 ix36798 (.Y (nx36799), .A (nx38589)) ;
    inv02 ix36800 (.Y (nx36801), .A (nx38589)) ;
    inv02 ix36802 (.Y (nx36803), .A (nx38589)) ;
    inv02 ix36804 (.Y (nx36805), .A (nx38589)) ;
    inv02 ix36806 (.Y (nx36807), .A (nx38591)) ;
    inv02 ix36808 (.Y (nx36809), .A (nx38591)) ;
    inv02 ix36810 (.Y (nx36811), .A (nx38591)) ;
    inv02 ix36812 (.Y (nx36813), .A (nx38591)) ;
    inv02 ix36814 (.Y (nx36815), .A (nx38591)) ;
    inv02 ix36816 (.Y (nx36817), .A (nx38591)) ;
    inv02 ix36818 (.Y (nx36819), .A (nx38591)) ;
    inv02 ix36820 (.Y (nx36821), .A (nx38593)) ;
    inv02 ix36822 (.Y (nx36823), .A (nx38593)) ;
    inv02 ix36824 (.Y (nx36825), .A (nx38593)) ;
    inv02 ix36826 (.Y (nx36827), .A (nx38593)) ;
    inv02 ix36828 (.Y (nx36829), .A (nx38593)) ;
    inv02 ix36830 (.Y (nx36831), .A (nx38593)) ;
    inv02 ix36832 (.Y (nx36833), .A (nx38593)) ;
    inv02 ix36834 (.Y (nx36835), .A (nx38595)) ;
    inv02 ix36836 (.Y (nx36837), .A (nx38595)) ;
    inv02 ix36838 (.Y (nx36839), .A (nx38595)) ;
    inv02 ix36840 (.Y (nx36841), .A (nx38595)) ;
    inv02 ix36842 (.Y (nx36843), .A (nx38595)) ;
    inv02 ix36844 (.Y (nx36845), .A (nx38595)) ;
    inv02 ix36846 (.Y (nx36847), .A (nx38595)) ;
    inv02 ix36848 (.Y (nx36849), .A (nx38597)) ;
    inv02 ix36850 (.Y (nx36851), .A (nx38597)) ;
    inv02 ix36852 (.Y (nx36853), .A (nx38597)) ;
    inv02 ix36854 (.Y (nx36855), .A (nx38597)) ;
    inv02 ix36856 (.Y (nx36857), .A (nx38597)) ;
    inv02 ix36858 (.Y (nx36859), .A (nx38597)) ;
    inv02 ix36860 (.Y (nx36861), .A (nx38597)) ;
    inv02 ix36862 (.Y (nx36863), .A (nx38599)) ;
    inv02 ix36864 (.Y (nx36865), .A (nx38599)) ;
    inv02 ix36866 (.Y (nx36867), .A (nx38599)) ;
    inv02 ix36868 (.Y (nx36869), .A (nx38599)) ;
    inv02 ix36870 (.Y (nx36871), .A (nx38599)) ;
    inv02 ix36872 (.Y (nx36873), .A (nx38599)) ;
    inv02 ix36874 (.Y (nx36875), .A (nx38599)) ;
    inv02 ix36878 (.Y (nx36879), .A (nx38601)) ;
    inv02 ix36880 (.Y (nx36881), .A (nx38601)) ;
    inv02 ix36882 (.Y (nx36883), .A (nx38601)) ;
    inv02 ix36884 (.Y (nx36885), .A (nx38601)) ;
    inv02 ix36886 (.Y (nx36887), .A (nx38601)) ;
    inv02 ix36888 (.Y (nx36889), .A (nx38601)) ;
    inv02 ix36890 (.Y (nx36891), .A (nx38601)) ;
    inv02 ix36892 (.Y (nx36893), .A (nx38603)) ;
    inv02 ix36894 (.Y (nx36895), .A (nx38603)) ;
    inv02 ix36896 (.Y (nx36897), .A (nx38603)) ;
    inv02 ix36898 (.Y (nx36899), .A (nx38603)) ;
    inv02 ix36900 (.Y (nx36901), .A (nx38603)) ;
    inv02 ix36902 (.Y (nx36903), .A (nx38603)) ;
    inv02 ix36904 (.Y (nx36905), .A (nx38603)) ;
    inv02 ix36906 (.Y (nx36907), .A (nx38605)) ;
    inv02 ix36908 (.Y (nx36909), .A (nx38605)) ;
    inv02 ix36910 (.Y (nx36911), .A (nx38605)) ;
    inv02 ix36912 (.Y (nx36913), .A (nx38605)) ;
    inv02 ix36914 (.Y (nx36915), .A (nx38605)) ;
    inv02 ix36916 (.Y (nx36917), .A (nx38605)) ;
    inv02 ix36918 (.Y (nx36919), .A (nx38605)) ;
    inv02 ix36920 (.Y (nx36921), .A (nx38607)) ;
    inv02 ix36922 (.Y (nx36923), .A (nx38607)) ;
    inv02 ix36924 (.Y (nx36925), .A (nx38607)) ;
    inv02 ix36926 (.Y (nx36927), .A (nx38607)) ;
    inv02 ix36928 (.Y (nx36929), .A (nx38607)) ;
    inv02 ix36930 (.Y (nx36931), .A (nx38607)) ;
    inv02 ix36932 (.Y (nx36933), .A (nx38607)) ;
    inv02 ix36934 (.Y (nx36935), .A (nx38609)) ;
    inv02 ix36936 (.Y (nx36937), .A (nx38609)) ;
    inv02 ix36938 (.Y (nx36939), .A (nx38609)) ;
    inv02 ix36940 (.Y (nx36941), .A (nx38609)) ;
    inv02 ix36942 (.Y (nx36943), .A (nx38609)) ;
    inv02 ix36944 (.Y (nx36945), .A (nx38609)) ;
    inv02 ix36946 (.Y (nx36947), .A (nx38609)) ;
    inv02 ix36948 (.Y (nx36949), .A (nx38611)) ;
    inv02 ix36950 (.Y (nx36951), .A (nx38611)) ;
    inv02 ix36952 (.Y (nx36953), .A (nx38611)) ;
    inv02 ix36954 (.Y (nx36955), .A (nx38611)) ;
    inv02 ix36956 (.Y (nx36957), .A (nx38611)) ;
    inv02 ix36958 (.Y (nx36959), .A (nx38611)) ;
    inv02 ix36960 (.Y (nx36961), .A (nx38611)) ;
    inv02 ix36962 (.Y (nx36963), .A (nx38613)) ;
    inv02 ix36964 (.Y (nx36965), .A (nx38613)) ;
    inv02 ix36966 (.Y (nx36967), .A (nx38613)) ;
    inv02 ix36968 (.Y (nx36969), .A (nx38613)) ;
    inv02 ix36970 (.Y (nx36971), .A (nx38613)) ;
    inv02 ix36972 (.Y (nx36973), .A (nx38613)) ;
    inv02 ix36974 (.Y (nx36975), .A (nx38613)) ;
    inv02 ix36976 (.Y (nx36977), .A (nx38615)) ;
    inv02 ix36978 (.Y (nx36979), .A (nx38615)) ;
    inv02 ix36980 (.Y (nx36981), .A (nx38615)) ;
    inv02 ix36982 (.Y (nx36983), .A (nx38615)) ;
    inv02 ix36984 (.Y (nx36985), .A (nx38615)) ;
    inv02 ix36986 (.Y (nx36987), .A (nx38615)) ;
    inv02 ix36988 (.Y (nx36989), .A (nx38615)) ;
    inv02 ix36990 (.Y (nx36991), .A (nx38617)) ;
    inv02 ix36992 (.Y (nx36993), .A (nx38617)) ;
    inv02 ix36994 (.Y (nx36995), .A (nx38617)) ;
    inv02 ix36996 (.Y (nx36997), .A (nx38617)) ;
    inv02 ix36998 (.Y (nx36999), .A (nx38617)) ;
    inv02 ix37000 (.Y (nx37001), .A (nx38617)) ;
    inv02 ix37002 (.Y (nx37003), .A (nx38617)) ;
    inv02 ix37004 (.Y (nx37005), .A (nx38619)) ;
    inv02 ix37006 (.Y (nx37007), .A (nx38619)) ;
    inv02 ix37008 (.Y (nx37009), .A (nx38619)) ;
    inv02 ix37010 (.Y (nx37011), .A (nx38619)) ;
    inv02 ix37012 (.Y (nx37013), .A (nx38619)) ;
    inv02 ix37014 (.Y (nx37015), .A (nx38619)) ;
    inv02 ix37016 (.Y (nx37017), .A (nx38619)) ;
    inv02 ix37020 (.Y (nx37021), .A (nx38621)) ;
    inv02 ix37022 (.Y (nx37023), .A (nx38621)) ;
    inv02 ix37024 (.Y (nx37025), .A (nx38621)) ;
    inv02 ix37026 (.Y (nx37027), .A (nx38621)) ;
    inv02 ix37028 (.Y (nx37029), .A (nx38621)) ;
    inv02 ix37030 (.Y (nx37031), .A (nx38621)) ;
    inv02 ix37032 (.Y (nx37033), .A (nx38621)) ;
    inv02 ix37034 (.Y (nx37035), .A (nx38623)) ;
    inv02 ix37036 (.Y (nx37037), .A (nx38623)) ;
    inv02 ix37038 (.Y (nx37039), .A (nx38623)) ;
    inv02 ix37040 (.Y (nx37041), .A (nx38623)) ;
    inv02 ix37042 (.Y (nx37043), .A (nx38623)) ;
    inv02 ix37044 (.Y (nx37045), .A (nx38623)) ;
    inv02 ix37046 (.Y (nx37047), .A (nx38623)) ;
    inv02 ix37048 (.Y (nx37049), .A (nx38625)) ;
    inv02 ix37050 (.Y (nx37051), .A (nx38625)) ;
    inv02 ix37052 (.Y (nx37053), .A (nx38625)) ;
    inv02 ix37054 (.Y (nx37055), .A (nx38625)) ;
    inv02 ix37056 (.Y (nx37057), .A (nx38625)) ;
    inv02 ix37058 (.Y (nx37059), .A (nx38625)) ;
    inv02 ix37060 (.Y (nx37061), .A (nx38625)) ;
    inv02 ix37062 (.Y (nx37063), .A (nx38627)) ;
    inv02 ix37064 (.Y (nx37065), .A (nx38627)) ;
    inv02 ix37066 (.Y (nx37067), .A (nx38627)) ;
    inv02 ix37068 (.Y (nx37069), .A (nx38627)) ;
    inv02 ix37070 (.Y (nx37071), .A (nx38627)) ;
    inv02 ix37072 (.Y (nx37073), .A (nx38627)) ;
    inv02 ix37074 (.Y (nx37075), .A (nx38627)) ;
    inv02 ix37076 (.Y (nx37077), .A (nx38629)) ;
    inv02 ix37078 (.Y (nx37079), .A (nx38629)) ;
    inv02 ix37080 (.Y (nx37081), .A (nx38629)) ;
    inv02 ix37082 (.Y (nx37083), .A (nx38629)) ;
    inv02 ix37084 (.Y (nx37085), .A (nx38629)) ;
    inv02 ix37086 (.Y (nx37087), .A (nx38629)) ;
    inv02 ix37088 (.Y (nx37089), .A (nx38629)) ;
    inv02 ix37090 (.Y (nx37091), .A (nx38631)) ;
    inv02 ix37092 (.Y (nx37093), .A (nx38631)) ;
    inv02 ix37094 (.Y (nx37095), .A (nx38631)) ;
    inv02 ix37096 (.Y (nx37097), .A (nx38631)) ;
    inv02 ix37098 (.Y (nx37099), .A (nx38631)) ;
    inv02 ix37100 (.Y (nx37101), .A (nx38631)) ;
    inv02 ix37102 (.Y (nx37103), .A (nx38631)) ;
    inv02 ix37104 (.Y (nx37105), .A (nx38633)) ;
    inv02 ix37106 (.Y (nx37107), .A (nx38633)) ;
    inv02 ix37108 (.Y (nx37109), .A (nx38633)) ;
    inv02 ix37110 (.Y (nx37111), .A (nx38633)) ;
    inv02 ix37112 (.Y (nx37113), .A (nx38633)) ;
    inv02 ix37114 (.Y (nx37115), .A (nx38633)) ;
    inv02 ix37116 (.Y (nx37117), .A (nx38633)) ;
    inv02 ix37118 (.Y (nx37119), .A (nx38635)) ;
    inv02 ix37120 (.Y (nx37121), .A (nx38635)) ;
    inv02 ix37122 (.Y (nx37123), .A (nx38635)) ;
    inv02 ix37124 (.Y (nx37125), .A (nx38635)) ;
    inv02 ix37126 (.Y (nx37127), .A (nx38635)) ;
    inv02 ix37128 (.Y (nx37129), .A (nx38635)) ;
    inv02 ix37130 (.Y (nx37131), .A (nx38635)) ;
    inv02 ix37132 (.Y (nx37133), .A (nx38637)) ;
    inv02 ix37134 (.Y (nx37135), .A (nx38637)) ;
    inv02 ix37136 (.Y (nx37137), .A (nx38637)) ;
    inv02 ix37138 (.Y (nx37139), .A (nx38637)) ;
    inv02 ix37140 (.Y (nx37141), .A (nx38637)) ;
    inv02 ix37142 (.Y (nx37143), .A (nx38637)) ;
    inv02 ix37144 (.Y (nx37145), .A (nx38637)) ;
    inv02 ix37146 (.Y (nx37147), .A (nx38639)) ;
    inv02 ix37148 (.Y (nx37149), .A (nx38639)) ;
    inv02 ix37150 (.Y (nx37151), .A (nx38639)) ;
    inv02 ix37152 (.Y (nx37153), .A (nx38639)) ;
    inv02 ix37154 (.Y (nx37155), .A (nx38639)) ;
    inv02 ix37156 (.Y (nx37157), .A (nx38639)) ;
    inv02 ix37158 (.Y (nx37159), .A (nx38639)) ;
    inv02 ix37162 (.Y (nx37163), .A (nx38641)) ;
    inv02 ix37164 (.Y (nx37165), .A (nx38641)) ;
    inv02 ix37166 (.Y (nx37167), .A (nx38641)) ;
    inv02 ix37168 (.Y (nx37169), .A (nx38641)) ;
    inv02 ix37170 (.Y (nx37171), .A (nx38641)) ;
    inv02 ix37172 (.Y (nx37173), .A (nx38641)) ;
    inv02 ix37174 (.Y (nx37175), .A (nx38641)) ;
    inv02 ix37176 (.Y (nx37177), .A (nx38643)) ;
    inv02 ix37178 (.Y (nx37179), .A (nx38643)) ;
    inv02 ix37180 (.Y (nx37181), .A (nx38643)) ;
    inv02 ix37182 (.Y (nx37183), .A (nx38643)) ;
    inv02 ix37184 (.Y (nx37185), .A (nx38643)) ;
    inv02 ix37186 (.Y (nx37187), .A (nx38643)) ;
    inv02 ix37188 (.Y (nx37189), .A (nx38643)) ;
    inv02 ix37190 (.Y (nx37191), .A (nx38645)) ;
    inv02 ix37192 (.Y (nx37193), .A (nx38645)) ;
    inv02 ix37194 (.Y (nx37195), .A (nx38645)) ;
    inv02 ix37196 (.Y (nx37197), .A (nx38645)) ;
    inv02 ix37198 (.Y (nx37199), .A (nx38645)) ;
    inv02 ix37200 (.Y (nx37201), .A (nx38645)) ;
    inv02 ix37202 (.Y (nx37203), .A (nx38645)) ;
    inv02 ix37204 (.Y (nx37205), .A (nx38647)) ;
    inv02 ix37206 (.Y (nx37207), .A (nx38647)) ;
    inv02 ix37208 (.Y (nx37209), .A (nx38647)) ;
    inv02 ix37210 (.Y (nx37211), .A (nx38647)) ;
    inv02 ix37212 (.Y (nx37213), .A (nx38647)) ;
    inv02 ix37214 (.Y (nx37215), .A (nx38647)) ;
    inv02 ix37216 (.Y (nx37217), .A (nx38647)) ;
    inv02 ix37218 (.Y (nx37219), .A (nx38649)) ;
    inv02 ix37220 (.Y (nx37221), .A (nx38649)) ;
    inv02 ix37222 (.Y (nx37223), .A (nx38649)) ;
    inv02 ix37224 (.Y (nx37225), .A (nx38649)) ;
    inv02 ix37226 (.Y (nx37227), .A (nx38649)) ;
    inv02 ix37228 (.Y (nx37229), .A (nx38649)) ;
    inv02 ix37230 (.Y (nx37231), .A (nx38649)) ;
    inv02 ix37232 (.Y (nx37233), .A (nx38651)) ;
    inv02 ix37234 (.Y (nx37235), .A (nx38651)) ;
    inv02 ix37236 (.Y (nx37237), .A (nx38651)) ;
    inv02 ix37238 (.Y (nx37239), .A (nx38651)) ;
    inv02 ix37240 (.Y (nx37241), .A (nx38651)) ;
    inv02 ix37242 (.Y (nx37243), .A (nx38651)) ;
    inv02 ix37244 (.Y (nx37245), .A (nx38651)) ;
    inv02 ix37246 (.Y (nx37247), .A (nx38653)) ;
    inv02 ix37248 (.Y (nx37249), .A (nx38653)) ;
    inv02 ix37250 (.Y (nx37251), .A (nx38653)) ;
    inv02 ix37252 (.Y (nx37253), .A (nx38653)) ;
    inv02 ix37254 (.Y (nx37255), .A (nx38653)) ;
    inv02 ix37256 (.Y (nx37257), .A (nx38653)) ;
    inv02 ix37258 (.Y (nx37259), .A (nx38653)) ;
    inv02 ix37260 (.Y (nx37261), .A (nx38655)) ;
    inv02 ix37262 (.Y (nx37263), .A (nx38655)) ;
    inv02 ix37264 (.Y (nx37265), .A (nx38655)) ;
    inv02 ix37266 (.Y (nx37267), .A (nx38655)) ;
    inv02 ix37268 (.Y (nx37269), .A (nx38655)) ;
    inv02 ix37270 (.Y (nx37271), .A (nx38655)) ;
    inv02 ix37272 (.Y (nx37273), .A (nx38655)) ;
    inv02 ix37274 (.Y (nx37275), .A (nx38657)) ;
    inv02 ix37276 (.Y (nx37277), .A (nx38657)) ;
    inv02 ix37278 (.Y (nx37279), .A (nx38657)) ;
    inv02 ix37280 (.Y (nx37281), .A (nx38657)) ;
    inv02 ix37282 (.Y (nx37283), .A (nx38657)) ;
    inv02 ix37284 (.Y (nx37285), .A (nx38657)) ;
    inv02 ix37286 (.Y (nx37287), .A (nx38657)) ;
    inv02 ix37288 (.Y (nx37289), .A (nx38659)) ;
    inv02 ix37290 (.Y (nx37291), .A (nx38659)) ;
    inv02 ix37292 (.Y (nx37293), .A (nx38659)) ;
    inv02 ix37294 (.Y (nx37295), .A (nx38659)) ;
    inv02 ix37296 (.Y (nx37297), .A (nx38659)) ;
    inv02 ix37298 (.Y (nx37299), .A (nx38659)) ;
    inv02 ix37300 (.Y (nx37301), .A (nx38659)) ;
    inv02 ix37304 (.Y (nx37305), .A (nx38661)) ;
    inv02 ix37306 (.Y (nx37307), .A (nx38661)) ;
    inv02 ix37308 (.Y (nx37309), .A (nx38661)) ;
    inv02 ix37310 (.Y (nx37311), .A (nx38661)) ;
    inv02 ix37312 (.Y (nx37313), .A (nx38661)) ;
    inv02 ix37314 (.Y (nx37315), .A (nx38661)) ;
    inv02 ix37316 (.Y (nx37317), .A (nx38661)) ;
    inv02 ix37318 (.Y (nx37319), .A (nx38663)) ;
    inv02 ix37320 (.Y (nx37321), .A (nx38663)) ;
    inv02 ix37322 (.Y (nx37323), .A (nx38663)) ;
    inv02 ix37324 (.Y (nx37325), .A (nx38663)) ;
    inv02 ix37326 (.Y (nx37327), .A (nx38663)) ;
    inv02 ix37328 (.Y (nx37329), .A (nx38663)) ;
    inv02 ix37330 (.Y (nx37331), .A (nx38663)) ;
    inv02 ix37332 (.Y (nx37333), .A (nx38665)) ;
    inv02 ix37334 (.Y (nx37335), .A (nx38665)) ;
    inv02 ix37336 (.Y (nx37337), .A (nx38665)) ;
    inv02 ix37338 (.Y (nx37339), .A (nx38665)) ;
    inv02 ix37340 (.Y (nx37341), .A (nx38665)) ;
    inv02 ix37342 (.Y (nx37343), .A (nx38665)) ;
    inv02 ix37344 (.Y (nx37345), .A (nx38665)) ;
    inv02 ix37346 (.Y (nx37347), .A (nx38667)) ;
    inv02 ix37348 (.Y (nx37349), .A (nx38667)) ;
    inv02 ix37350 (.Y (nx37351), .A (nx38667)) ;
    inv02 ix37352 (.Y (nx37353), .A (nx38667)) ;
    inv02 ix37354 (.Y (nx37355), .A (nx38667)) ;
    inv02 ix37356 (.Y (nx37357), .A (nx38667)) ;
    inv02 ix37358 (.Y (nx37359), .A (nx38667)) ;
    inv02 ix37360 (.Y (nx37361), .A (nx38669)) ;
    inv02 ix37362 (.Y (nx37363), .A (nx38669)) ;
    inv02 ix37364 (.Y (nx37365), .A (nx38669)) ;
    inv02 ix37366 (.Y (nx37367), .A (nx38669)) ;
    inv02 ix37368 (.Y (nx37369), .A (nx38669)) ;
    inv02 ix37370 (.Y (nx37371), .A (nx38669)) ;
    inv02 ix37372 (.Y (nx37373), .A (nx38669)) ;
    inv02 ix37374 (.Y (nx37375), .A (nx38671)) ;
    inv02 ix37376 (.Y (nx37377), .A (nx38671)) ;
    inv02 ix37378 (.Y (nx37379), .A (nx38671)) ;
    inv02 ix37380 (.Y (nx37381), .A (nx38671)) ;
    inv02 ix37382 (.Y (nx37383), .A (nx38671)) ;
    inv02 ix37384 (.Y (nx37385), .A (nx38671)) ;
    inv02 ix37386 (.Y (nx37387), .A (nx38671)) ;
    inv02 ix37388 (.Y (nx37389), .A (nx38673)) ;
    inv02 ix37390 (.Y (nx37391), .A (nx38673)) ;
    inv02 ix37392 (.Y (nx37393), .A (nx38673)) ;
    inv02 ix37394 (.Y (nx37395), .A (nx38673)) ;
    inv02 ix37396 (.Y (nx37397), .A (nx38673)) ;
    inv02 ix37398 (.Y (nx37399), .A (nx38673)) ;
    inv02 ix37400 (.Y (nx37401), .A (nx38673)) ;
    inv02 ix37402 (.Y (nx37403), .A (nx38675)) ;
    inv02 ix37404 (.Y (nx37405), .A (nx38675)) ;
    inv02 ix37406 (.Y (nx37407), .A (nx38675)) ;
    inv02 ix37408 (.Y (nx37409), .A (nx38675)) ;
    inv02 ix37410 (.Y (nx37411), .A (nx38675)) ;
    inv02 ix37412 (.Y (nx37413), .A (nx38675)) ;
    inv02 ix37414 (.Y (nx37415), .A (nx38675)) ;
    inv02 ix37416 (.Y (nx37417), .A (nx38677)) ;
    inv02 ix37418 (.Y (nx37419), .A (nx38677)) ;
    inv02 ix37420 (.Y (nx37421), .A (nx38677)) ;
    inv02 ix37422 (.Y (nx37423), .A (nx38677)) ;
    inv02 ix37424 (.Y (nx37425), .A (nx38677)) ;
    inv02 ix37426 (.Y (nx37427), .A (nx38677)) ;
    inv02 ix37428 (.Y (nx37429), .A (nx38677)) ;
    inv02 ix37430 (.Y (nx37431), .A (nx38679)) ;
    inv02 ix37432 (.Y (nx37433), .A (nx38679)) ;
    inv02 ix37434 (.Y (nx37435), .A (nx38679)) ;
    inv02 ix37436 (.Y (nx37437), .A (nx38679)) ;
    inv02 ix37438 (.Y (nx37439), .A (nx38679)) ;
    inv02 ix37440 (.Y (nx37441), .A (nx38679)) ;
    inv02 ix37442 (.Y (nx37443), .A (nx38679)) ;
    inv02 ix37446 (.Y (nx37447), .A (nx38681)) ;
    inv02 ix37448 (.Y (nx37449), .A (nx38681)) ;
    inv02 ix37450 (.Y (nx37451), .A (nx38681)) ;
    inv02 ix37452 (.Y (nx37453), .A (nx38681)) ;
    inv02 ix37454 (.Y (nx37455), .A (nx38681)) ;
    inv02 ix37456 (.Y (nx37457), .A (nx38681)) ;
    inv02 ix37458 (.Y (nx37459), .A (nx38681)) ;
    inv02 ix37460 (.Y (nx37461), .A (nx38683)) ;
    inv02 ix37462 (.Y (nx37463), .A (nx38683)) ;
    inv02 ix37464 (.Y (nx37465), .A (nx38683)) ;
    inv02 ix37466 (.Y (nx37467), .A (nx38683)) ;
    inv02 ix37468 (.Y (nx37469), .A (nx38683)) ;
    inv02 ix37470 (.Y (nx37471), .A (nx38683)) ;
    inv02 ix37472 (.Y (nx37473), .A (nx38683)) ;
    inv02 ix37474 (.Y (nx37475), .A (nx38685)) ;
    inv02 ix37476 (.Y (nx37477), .A (nx38685)) ;
    inv02 ix37478 (.Y (nx37479), .A (nx38685)) ;
    inv02 ix37480 (.Y (nx37481), .A (nx38685)) ;
    inv02 ix37482 (.Y (nx37483), .A (nx38685)) ;
    inv02 ix37484 (.Y (nx37485), .A (nx38685)) ;
    inv02 ix37486 (.Y (nx37487), .A (nx38685)) ;
    inv02 ix37488 (.Y (nx37489), .A (nx38687)) ;
    inv02 ix37490 (.Y (nx37491), .A (nx38687)) ;
    inv02 ix37492 (.Y (nx37493), .A (nx38687)) ;
    inv02 ix37494 (.Y (nx37495), .A (nx38687)) ;
    inv02 ix37496 (.Y (nx37497), .A (nx38687)) ;
    inv02 ix37498 (.Y (nx37499), .A (nx38687)) ;
    inv02 ix37500 (.Y (nx37501), .A (nx38687)) ;
    inv02 ix37502 (.Y (nx37503), .A (nx38689)) ;
    inv02 ix37504 (.Y (nx37505), .A (nx38689)) ;
    inv02 ix37506 (.Y (nx37507), .A (nx38689)) ;
    inv02 ix37508 (.Y (nx37509), .A (nx38689)) ;
    inv02 ix37510 (.Y (nx37511), .A (nx38689)) ;
    inv02 ix37512 (.Y (nx37513), .A (nx38689)) ;
    inv02 ix37514 (.Y (nx37515), .A (nx38689)) ;
    inv02 ix37516 (.Y (nx37517), .A (nx38691)) ;
    inv02 ix37518 (.Y (nx37519), .A (nx38691)) ;
    inv02 ix37520 (.Y (nx37521), .A (nx38691)) ;
    inv02 ix37522 (.Y (nx37523), .A (nx38691)) ;
    inv02 ix37524 (.Y (nx37525), .A (nx38691)) ;
    inv02 ix37526 (.Y (nx37527), .A (nx38691)) ;
    inv02 ix37528 (.Y (nx37529), .A (nx38691)) ;
    inv02 ix37530 (.Y (nx37531), .A (nx38693)) ;
    inv02 ix37532 (.Y (nx37533), .A (nx38693)) ;
    inv02 ix37534 (.Y (nx37535), .A (nx38693)) ;
    inv02 ix37536 (.Y (nx37537), .A (nx38693)) ;
    inv02 ix37538 (.Y (nx37539), .A (nx38693)) ;
    inv02 ix37540 (.Y (nx37541), .A (nx38693)) ;
    inv02 ix37542 (.Y (nx37543), .A (nx38693)) ;
    inv02 ix37544 (.Y (nx37545), .A (nx38695)) ;
    inv02 ix37546 (.Y (nx37547), .A (nx38695)) ;
    inv02 ix37548 (.Y (nx37549), .A (nx38695)) ;
    inv02 ix37550 (.Y (nx37551), .A (nx38695)) ;
    inv02 ix37552 (.Y (nx37553), .A (nx38695)) ;
    inv02 ix37554 (.Y (nx37555), .A (nx38695)) ;
    inv02 ix37556 (.Y (nx37557), .A (nx38695)) ;
    inv02 ix37558 (.Y (nx37559), .A (nx38697)) ;
    inv02 ix37560 (.Y (nx37561), .A (nx38697)) ;
    inv02 ix37562 (.Y (nx37563), .A (nx38697)) ;
    inv02 ix37564 (.Y (nx37565), .A (nx38697)) ;
    inv02 ix37566 (.Y (nx37567), .A (nx38697)) ;
    inv02 ix37568 (.Y (nx37569), .A (nx38697)) ;
    inv02 ix37570 (.Y (nx37571), .A (nx38697)) ;
    inv02 ix37572 (.Y (nx37573), .A (nx38699)) ;
    inv02 ix37574 (.Y (nx37575), .A (nx38699)) ;
    inv02 ix37576 (.Y (nx37577), .A (nx38699)) ;
    inv02 ix37578 (.Y (nx37579), .A (nx38699)) ;
    inv02 ix37580 (.Y (nx37581), .A (nx38699)) ;
    inv02 ix37582 (.Y (nx37583), .A (nx38699)) ;
    inv02 ix37584 (.Y (nx37585), .A (nx38699)) ;
    inv02 ix37588 (.Y (nx37589), .A (nx38701)) ;
    inv02 ix37590 (.Y (nx37591), .A (nx38701)) ;
    inv02 ix37592 (.Y (nx37593), .A (nx38701)) ;
    inv02 ix37594 (.Y (nx37595), .A (nx38701)) ;
    inv02 ix37596 (.Y (nx37597), .A (nx38701)) ;
    inv02 ix37598 (.Y (nx37599), .A (nx38701)) ;
    inv02 ix37600 (.Y (nx37601), .A (nx38701)) ;
    inv02 ix37602 (.Y (nx37603), .A (nx38703)) ;
    inv02 ix37604 (.Y (nx37605), .A (nx38703)) ;
    inv02 ix37606 (.Y (nx37607), .A (nx38703)) ;
    inv02 ix37608 (.Y (nx37609), .A (nx38703)) ;
    inv02 ix37610 (.Y (nx37611), .A (nx38703)) ;
    inv02 ix37612 (.Y (nx37613), .A (nx38703)) ;
    inv02 ix37614 (.Y (nx37615), .A (nx38703)) ;
    inv02 ix37616 (.Y (nx37617), .A (nx38705)) ;
    inv02 ix37618 (.Y (nx37619), .A (nx38705)) ;
    inv02 ix37620 (.Y (nx37621), .A (nx38705)) ;
    inv02 ix37622 (.Y (nx37623), .A (nx38705)) ;
    inv02 ix37624 (.Y (nx37625), .A (nx38705)) ;
    inv02 ix37626 (.Y (nx37627), .A (nx38705)) ;
    inv02 ix37628 (.Y (nx37629), .A (nx38705)) ;
    inv02 ix37630 (.Y (nx37631), .A (nx38707)) ;
    inv02 ix37632 (.Y (nx37633), .A (nx38707)) ;
    inv02 ix37634 (.Y (nx37635), .A (nx38707)) ;
    inv02 ix37636 (.Y (nx37637), .A (nx38707)) ;
    inv02 ix37638 (.Y (nx37639), .A (nx38707)) ;
    inv02 ix37640 (.Y (nx37641), .A (nx38707)) ;
    inv02 ix37642 (.Y (nx37643), .A (nx38707)) ;
    inv02 ix37644 (.Y (nx37645), .A (nx38709)) ;
    inv02 ix37646 (.Y (nx37647), .A (nx38709)) ;
    inv02 ix37648 (.Y (nx37649), .A (nx38709)) ;
    inv02 ix37650 (.Y (nx37651), .A (nx38709)) ;
    inv02 ix37652 (.Y (nx37653), .A (nx38709)) ;
    inv02 ix37654 (.Y (nx37655), .A (nx38709)) ;
    inv02 ix37656 (.Y (nx37657), .A (nx38709)) ;
    inv02 ix37658 (.Y (nx37659), .A (nx38711)) ;
    inv02 ix37660 (.Y (nx37661), .A (nx38711)) ;
    inv02 ix37662 (.Y (nx37663), .A (nx38711)) ;
    inv02 ix37664 (.Y (nx37665), .A (nx38711)) ;
    inv02 ix37666 (.Y (nx37667), .A (nx38711)) ;
    inv02 ix37668 (.Y (nx37669), .A (nx38711)) ;
    inv02 ix37670 (.Y (nx37671), .A (nx38711)) ;
    inv02 ix37672 (.Y (nx37673), .A (nx38713)) ;
    inv02 ix37674 (.Y (nx37675), .A (nx38713)) ;
    inv02 ix37676 (.Y (nx37677), .A (nx38713)) ;
    inv02 ix37678 (.Y (nx37679), .A (nx38713)) ;
    inv02 ix37680 (.Y (nx37681), .A (nx38713)) ;
    inv02 ix37682 (.Y (nx37683), .A (nx38713)) ;
    inv02 ix37684 (.Y (nx37685), .A (nx38713)) ;
    inv02 ix37686 (.Y (nx37687), .A (nx38715)) ;
    inv02 ix37688 (.Y (nx37689), .A (nx38715)) ;
    inv02 ix37690 (.Y (nx37691), .A (nx38715)) ;
    inv02 ix37692 (.Y (nx37693), .A (nx38715)) ;
    inv02 ix37694 (.Y (nx37695), .A (nx38715)) ;
    inv02 ix37696 (.Y (nx37697), .A (nx38715)) ;
    inv02 ix37698 (.Y (nx37699), .A (nx38715)) ;
    inv02 ix37700 (.Y (nx37701), .A (nx38717)) ;
    inv02 ix37702 (.Y (nx37703), .A (nx38717)) ;
    inv02 ix37704 (.Y (nx37705), .A (nx38717)) ;
    inv02 ix37706 (.Y (nx37707), .A (nx38717)) ;
    inv02 ix37708 (.Y (nx37709), .A (nx38717)) ;
    inv02 ix37710 (.Y (nx37711), .A (nx38717)) ;
    inv02 ix37712 (.Y (nx37713), .A (nx38717)) ;
    inv02 ix37714 (.Y (nx37715), .A (nx38719)) ;
    inv02 ix37716 (.Y (nx37717), .A (nx38719)) ;
    inv02 ix37718 (.Y (nx37719), .A (nx38719)) ;
    inv02 ix37720 (.Y (nx37721), .A (nx38719)) ;
    inv02 ix37722 (.Y (nx37723), .A (nx38719)) ;
    inv02 ix37724 (.Y (nx37725), .A (nx38719)) ;
    inv02 ix37726 (.Y (nx37727), .A (nx38719)) ;
    inv02 ix37730 (.Y (nx37731), .A (nx38721)) ;
    inv02 ix37732 (.Y (nx37733), .A (nx38721)) ;
    inv02 ix37734 (.Y (nx37735), .A (nx38721)) ;
    inv02 ix37736 (.Y (nx37737), .A (nx38721)) ;
    inv02 ix37738 (.Y (nx37739), .A (nx38721)) ;
    inv02 ix37740 (.Y (nx37741), .A (nx38721)) ;
    inv02 ix37742 (.Y (nx37743), .A (nx38721)) ;
    inv02 ix37744 (.Y (nx37745), .A (nx38723)) ;
    inv02 ix37746 (.Y (nx37747), .A (nx38723)) ;
    inv02 ix37748 (.Y (nx37749), .A (nx38723)) ;
    inv02 ix37750 (.Y (nx37751), .A (nx38723)) ;
    inv02 ix37752 (.Y (nx37753), .A (nx38723)) ;
    inv02 ix37754 (.Y (nx37755), .A (nx38723)) ;
    inv02 ix37756 (.Y (nx37757), .A (nx38723)) ;
    inv02 ix37758 (.Y (nx37759), .A (nx38725)) ;
    inv02 ix37760 (.Y (nx37761), .A (nx38725)) ;
    inv02 ix37762 (.Y (nx37763), .A (nx38725)) ;
    inv02 ix37764 (.Y (nx37765), .A (nx38725)) ;
    inv02 ix37766 (.Y (nx37767), .A (nx38725)) ;
    inv02 ix37768 (.Y (nx37769), .A (nx38725)) ;
    inv02 ix37770 (.Y (nx37771), .A (nx38725)) ;
    inv02 ix37772 (.Y (nx37773), .A (nx38727)) ;
    inv02 ix37774 (.Y (nx37775), .A (nx38727)) ;
    inv02 ix37776 (.Y (nx37777), .A (nx38727)) ;
    inv02 ix37778 (.Y (nx37779), .A (nx38727)) ;
    inv02 ix37780 (.Y (nx37781), .A (nx38727)) ;
    inv02 ix37782 (.Y (nx37783), .A (nx38727)) ;
    inv02 ix37784 (.Y (nx37785), .A (nx38727)) ;
    inv02 ix37786 (.Y (nx37787), .A (nx38729)) ;
    inv02 ix37788 (.Y (nx37789), .A (nx38729)) ;
    inv02 ix37790 (.Y (nx37791), .A (nx38729)) ;
    inv02 ix37792 (.Y (nx37793), .A (nx38729)) ;
    inv02 ix37794 (.Y (nx37795), .A (nx38729)) ;
    inv02 ix37796 (.Y (nx37797), .A (nx38729)) ;
    inv02 ix37798 (.Y (nx37799), .A (nx38729)) ;
    inv02 ix37800 (.Y (nx37801), .A (nx38731)) ;
    inv02 ix37802 (.Y (nx37803), .A (nx38731)) ;
    inv02 ix37804 (.Y (nx37805), .A (nx38731)) ;
    inv02 ix37806 (.Y (nx37807), .A (nx38731)) ;
    inv02 ix37808 (.Y (nx37809), .A (nx38731)) ;
    inv02 ix37810 (.Y (nx37811), .A (nx38731)) ;
    inv02 ix37812 (.Y (nx37813), .A (nx38731)) ;
    inv02 ix37814 (.Y (nx37815), .A (nx38733)) ;
    inv02 ix37816 (.Y (nx37817), .A (nx38733)) ;
    inv02 ix37818 (.Y (nx37819), .A (nx38733)) ;
    inv02 ix37820 (.Y (nx37821), .A (nx38733)) ;
    inv02 ix37822 (.Y (nx37823), .A (nx38733)) ;
    inv02 ix37824 (.Y (nx37825), .A (nx38733)) ;
    inv02 ix37826 (.Y (nx37827), .A (nx38733)) ;
    inv02 ix37828 (.Y (nx37829), .A (nx38735)) ;
    inv02 ix37830 (.Y (nx37831), .A (nx38735)) ;
    inv02 ix37832 (.Y (nx37833), .A (nx38735)) ;
    inv02 ix37834 (.Y (nx37835), .A (nx38735)) ;
    inv02 ix37836 (.Y (nx37837), .A (nx38735)) ;
    inv02 ix37838 (.Y (nx37839), .A (nx38735)) ;
    inv02 ix37840 (.Y (nx37841), .A (nx38735)) ;
    inv02 ix37842 (.Y (nx37843), .A (nx38737)) ;
    inv02 ix37844 (.Y (nx37845), .A (nx38737)) ;
    inv02 ix37846 (.Y (nx37847), .A (nx38737)) ;
    inv02 ix37848 (.Y (nx37849), .A (nx38737)) ;
    inv02 ix37850 (.Y (nx37851), .A (nx38737)) ;
    inv02 ix37852 (.Y (nx37853), .A (nx38737)) ;
    inv02 ix37854 (.Y (nx37855), .A (nx38737)) ;
    inv02 ix37856 (.Y (nx37857), .A (nx38739)) ;
    inv02 ix37858 (.Y (nx37859), .A (nx38739)) ;
    inv02 ix37860 (.Y (nx37861), .A (nx38739)) ;
    inv02 ix37862 (.Y (nx37863), .A (nx38739)) ;
    inv02 ix37864 (.Y (nx37865), .A (nx38739)) ;
    inv02 ix37866 (.Y (nx37867), .A (nx38739)) ;
    inv02 ix37868 (.Y (nx37869), .A (nx38739)) ;
    inv02 ix37872 (.Y (nx37873), .A (nx38741)) ;
    inv02 ix37874 (.Y (nx37875), .A (nx38741)) ;
    inv02 ix37876 (.Y (nx37877), .A (nx38741)) ;
    inv02 ix37878 (.Y (nx37879), .A (nx38741)) ;
    inv02 ix37880 (.Y (nx37881), .A (nx38741)) ;
    inv02 ix37882 (.Y (nx37883), .A (nx38741)) ;
    inv02 ix37884 (.Y (nx37885), .A (nx38741)) ;
    inv02 ix37886 (.Y (nx37887), .A (nx38743)) ;
    inv02 ix37888 (.Y (nx37889), .A (nx38743)) ;
    inv02 ix37890 (.Y (nx37891), .A (nx38743)) ;
    inv02 ix37892 (.Y (nx37893), .A (nx38743)) ;
    inv02 ix37894 (.Y (nx37895), .A (nx38743)) ;
    inv02 ix37896 (.Y (nx37897), .A (nx38743)) ;
    inv02 ix37898 (.Y (nx37899), .A (nx38743)) ;
    inv02 ix37900 (.Y (nx37901), .A (nx38745)) ;
    inv02 ix37902 (.Y (nx37903), .A (nx38745)) ;
    inv02 ix37904 (.Y (nx37905), .A (nx38745)) ;
    inv02 ix37906 (.Y (nx37907), .A (nx38745)) ;
    inv02 ix37908 (.Y (nx37909), .A (nx38745)) ;
    inv02 ix37910 (.Y (nx37911), .A (nx38745)) ;
    inv02 ix37912 (.Y (nx37913), .A (nx38745)) ;
    inv02 ix37914 (.Y (nx37915), .A (nx38747)) ;
    inv02 ix37916 (.Y (nx37917), .A (nx38747)) ;
    inv02 ix37918 (.Y (nx37919), .A (nx38747)) ;
    inv02 ix37920 (.Y (nx37921), .A (nx38747)) ;
    inv02 ix37922 (.Y (nx37923), .A (nx38747)) ;
    inv02 ix37924 (.Y (nx37925), .A (nx38747)) ;
    inv02 ix37926 (.Y (nx37927), .A (nx38747)) ;
    inv02 ix37928 (.Y (nx37929), .A (nx38749)) ;
    inv02 ix37930 (.Y (nx37931), .A (nx38749)) ;
    inv02 ix37932 (.Y (nx37933), .A (nx38749)) ;
    inv02 ix37934 (.Y (nx37935), .A (nx38749)) ;
    inv02 ix37936 (.Y (nx37937), .A (nx38749)) ;
    inv02 ix37938 (.Y (nx37939), .A (nx38749)) ;
    inv02 ix37940 (.Y (nx37941), .A (nx38749)) ;
    inv02 ix37942 (.Y (nx37943), .A (nx38751)) ;
    inv02 ix37944 (.Y (nx37945), .A (nx38751)) ;
    inv02 ix37946 (.Y (nx37947), .A (nx38751)) ;
    inv02 ix37948 (.Y (nx37949), .A (nx38751)) ;
    inv02 ix37950 (.Y (nx37951), .A (nx38751)) ;
    inv02 ix37952 (.Y (nx37953), .A (nx38751)) ;
    inv02 ix37954 (.Y (nx37955), .A (nx38751)) ;
    inv02 ix37956 (.Y (nx37957), .A (nx38753)) ;
    inv02 ix37958 (.Y (nx37959), .A (nx38753)) ;
    inv02 ix37960 (.Y (nx37961), .A (nx38753)) ;
    inv02 ix37962 (.Y (nx37963), .A (nx38753)) ;
    inv02 ix37964 (.Y (nx37965), .A (nx38753)) ;
    inv02 ix37966 (.Y (nx37967), .A (nx38753)) ;
    inv02 ix37968 (.Y (nx37969), .A (nx38753)) ;
    inv02 ix37970 (.Y (nx37971), .A (nx38755)) ;
    inv02 ix37972 (.Y (nx37973), .A (nx38755)) ;
    inv02 ix37974 (.Y (nx37975), .A (nx38755)) ;
    inv02 ix37976 (.Y (nx37977), .A (nx38755)) ;
    inv02 ix37978 (.Y (nx37979), .A (nx38755)) ;
    inv02 ix37980 (.Y (nx37981), .A (nx38755)) ;
    inv02 ix37982 (.Y (nx37983), .A (nx38755)) ;
    inv02 ix37984 (.Y (nx37985), .A (nx38757)) ;
    inv02 ix37986 (.Y (nx37987), .A (nx38757)) ;
    inv02 ix37988 (.Y (nx37989), .A (nx38757)) ;
    inv02 ix37990 (.Y (nx37991), .A (nx38757)) ;
    inv02 ix37992 (.Y (nx37993), .A (nx38757)) ;
    inv02 ix37994 (.Y (nx37995), .A (nx38757)) ;
    inv02 ix37996 (.Y (nx37997), .A (nx38757)) ;
    inv02 ix37998 (.Y (nx37999), .A (nx38759)) ;
    inv02 ix38000 (.Y (nx38001), .A (nx38759)) ;
    inv02 ix38002 (.Y (nx38003), .A (nx38759)) ;
    inv02 ix38004 (.Y (nx38005), .A (nx38759)) ;
    inv02 ix38006 (.Y (nx38007), .A (nx38759)) ;
    inv02 ix38008 (.Y (nx38009), .A (nx38759)) ;
    inv02 ix38010 (.Y (nx38011), .A (nx38759)) ;
    inv02 ix38014 (.Y (nx38015), .A (nx38761)) ;
    inv02 ix38016 (.Y (nx38017), .A (nx38761)) ;
    inv02 ix38018 (.Y (nx38019), .A (nx38761)) ;
    inv02 ix38020 (.Y (nx38021), .A (nx38761)) ;
    inv02 ix38022 (.Y (nx38023), .A (nx38761)) ;
    inv02 ix38024 (.Y (nx38025), .A (nx38761)) ;
    inv02 ix38026 (.Y (nx38027), .A (nx38761)) ;
    inv02 ix38028 (.Y (nx38029), .A (nx38763)) ;
    inv02 ix38030 (.Y (nx38031), .A (nx38763)) ;
    inv02 ix38032 (.Y (nx38033), .A (nx38763)) ;
    inv02 ix38034 (.Y (nx38035), .A (nx38763)) ;
    inv02 ix38036 (.Y (nx38037), .A (nx38763)) ;
    inv02 ix38038 (.Y (nx38039), .A (nx38763)) ;
    inv02 ix38040 (.Y (nx38041), .A (nx38763)) ;
    inv02 ix38042 (.Y (nx38043), .A (nx38765)) ;
    inv02 ix38044 (.Y (nx38045), .A (nx38765)) ;
    inv02 ix38046 (.Y (nx38047), .A (nx38765)) ;
    inv02 ix38048 (.Y (nx38049), .A (nx38765)) ;
    inv02 ix38050 (.Y (nx38051), .A (nx38765)) ;
    inv02 ix38052 (.Y (nx38053), .A (nx38765)) ;
    inv02 ix38054 (.Y (nx38055), .A (nx38765)) ;
    inv02 ix38056 (.Y (nx38057), .A (nx38767)) ;
    inv02 ix38058 (.Y (nx38059), .A (nx38767)) ;
    inv02 ix38060 (.Y (nx38061), .A (nx38767)) ;
    inv02 ix38062 (.Y (nx38063), .A (nx38767)) ;
    inv02 ix38064 (.Y (nx38065), .A (nx38767)) ;
    inv02 ix38066 (.Y (nx38067), .A (nx38767)) ;
    inv02 ix38068 (.Y (nx38069), .A (nx38767)) ;
    inv02 ix38070 (.Y (nx38071), .A (nx38769)) ;
    inv02 ix38072 (.Y (nx38073), .A (nx38769)) ;
    inv02 ix38074 (.Y (nx38075), .A (nx38769)) ;
    inv02 ix38076 (.Y (nx38077), .A (nx38769)) ;
    inv02 ix38078 (.Y (nx38079), .A (nx38769)) ;
    inv02 ix38080 (.Y (nx38081), .A (nx38769)) ;
    inv02 ix38082 (.Y (nx38083), .A (nx38769)) ;
    inv02 ix38084 (.Y (nx38085), .A (nx38771)) ;
    inv02 ix38086 (.Y (nx38087), .A (nx38771)) ;
    inv02 ix38088 (.Y (nx38089), .A (nx38771)) ;
    inv02 ix38090 (.Y (nx38091), .A (nx38771)) ;
    inv02 ix38092 (.Y (nx38093), .A (nx38771)) ;
    inv02 ix38094 (.Y (nx38095), .A (nx38771)) ;
    inv02 ix38096 (.Y (nx38097), .A (nx38771)) ;
    inv02 ix38098 (.Y (nx38099), .A (nx38773)) ;
    inv02 ix38100 (.Y (nx38101), .A (nx38773)) ;
    inv02 ix38102 (.Y (nx38103), .A (nx38773)) ;
    inv02 ix38104 (.Y (nx38105), .A (nx38773)) ;
    inv02 ix38106 (.Y (nx38107), .A (nx38773)) ;
    inv02 ix38108 (.Y (nx38109), .A (nx38773)) ;
    inv02 ix38110 (.Y (nx38111), .A (nx38773)) ;
    inv02 ix38112 (.Y (nx38113), .A (nx38775)) ;
    inv02 ix38114 (.Y (nx38115), .A (nx38775)) ;
    inv02 ix38116 (.Y (nx38117), .A (nx38775)) ;
    inv02 ix38118 (.Y (nx38119), .A (nx38775)) ;
    inv02 ix38120 (.Y (nx38121), .A (nx38775)) ;
    inv02 ix38122 (.Y (nx38123), .A (nx38775)) ;
    inv02 ix38124 (.Y (nx38125), .A (nx38775)) ;
    inv02 ix38126 (.Y (nx38127), .A (nx38777)) ;
    inv02 ix38128 (.Y (nx38129), .A (nx38777)) ;
    inv02 ix38130 (.Y (nx38131), .A (nx38777)) ;
    inv02 ix38132 (.Y (nx38133), .A (nx38777)) ;
    inv02 ix38134 (.Y (nx38135), .A (nx38777)) ;
    inv02 ix38136 (.Y (nx38137), .A (nx38777)) ;
    inv02 ix38138 (.Y (nx38139), .A (nx38777)) ;
    inv02 ix38140 (.Y (nx38141), .A (nx38779)) ;
    inv02 ix38142 (.Y (nx38143), .A (nx38779)) ;
    inv02 ix38144 (.Y (nx38145), .A (nx38779)) ;
    inv02 ix38146 (.Y (nx38147), .A (nx38779)) ;
    inv02 ix38148 (.Y (nx38149), .A (nx38779)) ;
    inv02 ix38150 (.Y (nx38151), .A (nx38779)) ;
    inv02 ix38152 (.Y (nx38153), .A (nx38779)) ;
    buf02 ix38154 (.Y (nx38155), .A (registerSelector_6)) ;
    buf02 ix38156 (.Y (nx38157), .A (registerSelector_3)) ;
    inv01 ix38158 (.Y (nx38159), .A (nx38879)) ;
    inv01 ix38160 (.Y (nx38161), .A (nx38879)) ;
    inv01 ix38162 (.Y (nx38163), .A (nx38879)) ;
    inv01 ix38164 (.Y (nx38165), .A (nx38879)) ;
    inv01 ix38166 (.Y (nx38167), .A (nx38879)) ;
    inv01 ix38168 (.Y (nx38169), .A (nx38879)) ;
    inv01 ix38170 (.Y (nx38171), .A (nx38879)) ;
    inv01 ix38172 (.Y (nx38173), .A (nx38881)) ;
    inv01 ix38174 (.Y (nx38175), .A (nx38881)) ;
    inv01 ix38176 (.Y (nx38177), .A (nx38881)) ;
    inv01 ix38178 (.Y (nx38179), .A (nx38881)) ;
    inv01 ix38180 (.Y (nx38181), .A (nx38881)) ;
    inv01 ix38182 (.Y (nx38183), .A (nx38881)) ;
    inv01 ix38184 (.Y (nx38185), .A (nx38881)) ;
    inv01 ix38186 (.Y (nx38187), .A (nx38883)) ;
    inv01 ix38188 (.Y (nx38189), .A (nx38883)) ;
    inv01 ix38190 (.Y (nx38191), .A (nx38883)) ;
    inv01 ix38192 (.Y (nx38193), .A (nx38883)) ;
    inv01 ix38194 (.Y (nx38195), .A (nx38883)) ;
    inv01 ix38196 (.Y (nx38197), .A (nx38883)) ;
    inv01 ix38198 (.Y (nx38199), .A (nx38883)) ;
    inv01 ix38200 (.Y (nx38201), .A (nx38885)) ;
    inv01 ix38202 (.Y (nx38203), .A (nx38885)) ;
    inv01 ix38204 (.Y (nx38205), .A (nx38885)) ;
    inv01 ix38206 (.Y (nx38207), .A (nx38885)) ;
    inv01 ix38208 (.Y (nx38209), .A (nx38885)) ;
    inv01 ix38210 (.Y (nx38211), .A (nx38885)) ;
    inv01 ix38212 (.Y (nx38213), .A (nx38885)) ;
    inv01 ix38214 (.Y (nx38215), .A (nx38887)) ;
    inv01 ix38216 (.Y (nx38217), .A (nx38887)) ;
    inv01 ix38218 (.Y (nx38219), .A (nx38887)) ;
    inv01 ix38220 (.Y (nx38221), .A (nx38887)) ;
    inv01 ix38222 (.Y (nx38223), .A (nx38887)) ;
    inv01 ix38224 (.Y (nx38225), .A (nx38887)) ;
    inv01 ix38226 (.Y (nx38227), .A (nx38887)) ;
    inv01 ix38228 (.Y (nx38229), .A (nx38889)) ;
    inv01 ix38230 (.Y (nx38231), .A (nx38889)) ;
    inv01 ix38232 (.Y (nx38233), .A (nx38889)) ;
    inv01 ix38234 (.Y (nx38235), .A (nx38889)) ;
    inv01 ix38236 (.Y (nx38237), .A (nx38889)) ;
    inv01 ix38238 (.Y (nx38239), .A (nx38889)) ;
    inv01 ix38240 (.Y (nx38241), .A (nx38889)) ;
    inv01 ix38242 (.Y (nx38243), .A (nx38891)) ;
    inv01 ix38244 (.Y (nx38245), .A (nx38891)) ;
    inv01 ix38246 (.Y (nx38247), .A (nx38891)) ;
    inv01 ix38248 (.Y (nx38249), .A (nx38891)) ;
    inv01 ix38250 (.Y (nx38251), .A (nx38891)) ;
    inv01 ix38252 (.Y (nx38253), .A (nx38891)) ;
    inv01 ix38254 (.Y (nx38255), .A (nx38891)) ;
    inv01 ix38256 (.Y (nx38257), .A (nx38893)) ;
    inv01 ix38258 (.Y (nx38259), .A (nx38893)) ;
    inv01 ix38260 (.Y (nx38261), .A (nx38893)) ;
    inv01 ix38262 (.Y (nx38263), .A (nx38893)) ;
    inv01 ix38264 (.Y (nx38265), .A (nx38893)) ;
    inv01 ix38266 (.Y (nx38267), .A (nx38893)) ;
    inv01 ix38268 (.Y (nx38269), .A (nx38893)) ;
    inv01 ix38270 (.Y (nx38271), .A (nx38895)) ;
    inv01 ix38272 (.Y (nx38273), .A (nx38895)) ;
    inv01 ix38274 (.Y (nx38275), .A (nx38895)) ;
    inv01 ix38276 (.Y (nx38277), .A (nx38895)) ;
    inv01 ix38278 (.Y (nx38279), .A (nx38895)) ;
    inv01 ix38280 (.Y (nx38281), .A (nx38895)) ;
    inv01 ix38282 (.Y (nx38283), .A (nx38895)) ;
    inv01 ix38284 (.Y (nx38285), .A (nx38897)) ;
    inv01 ix38286 (.Y (nx38287), .A (nx38897)) ;
    inv01 ix38288 (.Y (nx38289), .A (nx38897)) ;
    inv01 ix38290 (.Y (nx38291), .A (nx38897)) ;
    inv01 ix38292 (.Y (nx38293), .A (nx38897)) ;
    inv01 ix38294 (.Y (nx38295), .A (nx38897)) ;
    inv01 ix38296 (.Y (nx38297), .A (nx38899)) ;
    inv01 ix38298 (.Y (nx38299), .A (nx38899)) ;
    inv01 ix38300 (.Y (nx38301), .A (nx38899)) ;
    inv01 ix38302 (.Y (nx38303), .A (nx38899)) ;
    inv01 ix38304 (.Y (nx38305), .A (nx38899)) ;
    inv01 ix38306 (.Y (nx38307), .A (nx38899)) ;
    inv01 ix38308 (.Y (nx38309), .A (nx38899)) ;
    inv01 ix38310 (.Y (nx38311), .A (nx38901)) ;
    inv01 ix38312 (.Y (nx38313), .A (nx38901)) ;
    inv01 ix38314 (.Y (nx38315), .A (nx38785)) ;
    inv01 ix38316 (.Y (nx38317), .A (nx38785)) ;
    inv01 ix38318 (.Y (nx38319), .A (nx38785)) ;
    inv01 ix38320 (.Y (nx38321), .A (nx38785)) ;
    inv01 ix38322 (.Y (nx38323), .A (nx38785)) ;
    inv01 ix38324 (.Y (nx38325), .A (nx38785)) ;
    inv01 ix38326 (.Y (nx38327), .A (nx38785)) ;
    inv01 ix38328 (.Y (nx38329), .A (nx38787)) ;
    inv01 ix38330 (.Y (nx38331), .A (nx38787)) ;
    inv01 ix38332 (.Y (nx38333), .A (nx38789)) ;
    inv01 ix38334 (.Y (nx38335), .A (nx38789)) ;
    inv01 ix38336 (.Y (nx38337), .A (nx38789)) ;
    inv01 ix38338 (.Y (nx38339), .A (nx38789)) ;
    inv01 ix38340 (.Y (nx38341), .A (nx38789)) ;
    inv01 ix38342 (.Y (nx38343), .A (nx38789)) ;
    inv01 ix38344 (.Y (nx38345), .A (nx38789)) ;
    inv01 ix38346 (.Y (nx38347), .A (nx38791)) ;
    inv01 ix38348 (.Y (nx38349), .A (nx38791)) ;
    inv01 ix38350 (.Y (nx38351), .A (nx38793)) ;
    inv01 ix38352 (.Y (nx38353), .A (nx38793)) ;
    inv01 ix38354 (.Y (nx38355), .A (nx38793)) ;
    inv01 ix38356 (.Y (nx38357), .A (nx38793)) ;
    inv01 ix38358 (.Y (nx38359), .A (nx38793)) ;
    inv01 ix38360 (.Y (nx38361), .A (nx38793)) ;
    inv01 ix38362 (.Y (nx38363), .A (nx38793)) ;
    inv01 ix38364 (.Y (nx38365), .A (nx38795)) ;
    inv01 ix38366 (.Y (nx38367), .A (nx38795)) ;
    inv01 ix38368 (.Y (nx38369), .A (nx38797)) ;
    inv01 ix38370 (.Y (nx38371), .A (nx38797)) ;
    inv01 ix38372 (.Y (nx38373), .A (nx38797)) ;
    inv01 ix38374 (.Y (nx38375), .A (nx38797)) ;
    inv01 ix38376 (.Y (nx38377), .A (nx38797)) ;
    inv01 ix38378 (.Y (nx38379), .A (nx38797)) ;
    inv01 ix38380 (.Y (nx38381), .A (nx38797)) ;
    inv01 ix38382 (.Y (nx38383), .A (nx38799)) ;
    inv01 ix38384 (.Y (nx38385), .A (nx38799)) ;
    inv01 ix38386 (.Y (nx38387), .A (nx38801)) ;
    inv01 ix38388 (.Y (nx38389), .A (nx38801)) ;
    inv01 ix38390 (.Y (nx38391), .A (nx38801)) ;
    inv01 ix38392 (.Y (nx38393), .A (nx38801)) ;
    inv01 ix38394 (.Y (nx38395), .A (nx38801)) ;
    inv01 ix38396 (.Y (nx38397), .A (nx38801)) ;
    inv01 ix38398 (.Y (nx38399), .A (nx38801)) ;
    inv01 ix38400 (.Y (nx38401), .A (nx38803)) ;
    inv01 ix38402 (.Y (nx38403), .A (nx38803)) ;
    inv01 ix38404 (.Y (nx38405), .A (nx38805)) ;
    inv01 ix38406 (.Y (nx38407), .A (nx38805)) ;
    inv01 ix38408 (.Y (nx38409), .A (nx38805)) ;
    inv01 ix38410 (.Y (nx38411), .A (nx38805)) ;
    inv01 ix38412 (.Y (nx38413), .A (nx38805)) ;
    inv01 ix38414 (.Y (nx38415), .A (nx38805)) ;
    inv01 ix38416 (.Y (nx38417), .A (nx38805)) ;
    inv01 ix38418 (.Y (nx38419), .A (nx38807)) ;
    inv01 ix38420 (.Y (nx38421), .A (nx38807)) ;
    inv01 ix38422 (.Y (nx38423), .A (nx38809)) ;
    inv01 ix38424 (.Y (nx38425), .A (nx38809)) ;
    inv01 ix38426 (.Y (nx38427), .A (nx38809)) ;
    inv01 ix38428 (.Y (nx38429), .A (nx38809)) ;
    inv01 ix38430 (.Y (nx38431), .A (nx38809)) ;
    inv01 ix38432 (.Y (nx38433), .A (nx38809)) ;
    inv01 ix38434 (.Y (nx38435), .A (nx38809)) ;
    inv01 ix38436 (.Y (nx38437), .A (nx38811)) ;
    inv01 ix38438 (.Y (nx38439), .A (nx38811)) ;
    inv01 ix38440 (.Y (nx38441), .A (nx38811)) ;
    inv01 ix38442 (.Y (nx38443), .A (nx38811)) ;
    inv01 ix38444 (.Y (nx38445), .A (nx38811)) ;
    inv01 ix38446 (.Y (nx38447), .A (nx38811)) ;
    inv01 ix38448 (.Y (nx38449), .A (nx38811)) ;
    inv01 ix38450 (.Y (nx38451), .A (nx38813)) ;
    inv01 ix38452 (.Y (nx38453), .A (nx38813)) ;
    inv01 ix38454 (.Y (nx38455), .A (nx38813)) ;
    inv01 ix38456 (.Y (nx38457), .A (nx38813)) ;
    inv01 ix38458 (.Y (nx38459), .A (nx38813)) ;
    inv02 ix38460 (.Y (nx38461), .A (sumInput[15])) ;
    inv02 ix38462 (.Y (nx38463), .A (nx38815)) ;
    inv02 ix38464 (.Y (nx38465), .A (nx38815)) ;
    inv02 ix38466 (.Y (nx38467), .A (nx38815)) ;
    inv02 ix38468 (.Y (nx38469), .A (nx38815)) ;
    inv02 ix38470 (.Y (nx38471), .A (nx38815)) ;
    inv02 ix38472 (.Y (nx38473), .A (nx38817)) ;
    inv02 ix38474 (.Y (nx38475), .A (nx38817)) ;
    inv02 ix38476 (.Y (nx38477), .A (nx38817)) ;
    inv02 ix38478 (.Y (nx38479), .A (nx38817)) ;
    inv02 ix38480 (.Y (nx38481), .A (sumInput[14])) ;
    inv02 ix38482 (.Y (nx38483), .A (nx38819)) ;
    inv02 ix38484 (.Y (nx38485), .A (nx38819)) ;
    inv02 ix38486 (.Y (nx38487), .A (nx38819)) ;
    inv02 ix38488 (.Y (nx38489), .A (nx38819)) ;
    inv02 ix38490 (.Y (nx38491), .A (nx38819)) ;
    inv02 ix38492 (.Y (nx38493), .A (nx38821)) ;
    inv02 ix38494 (.Y (nx38495), .A (nx38821)) ;
    inv02 ix38496 (.Y (nx38497), .A (nx38821)) ;
    inv02 ix38498 (.Y (nx38499), .A (nx38821)) ;
    inv02 ix38500 (.Y (nx38501), .A (sumInput[13])) ;
    inv02 ix38502 (.Y (nx38503), .A (nx38823)) ;
    inv02 ix38504 (.Y (nx38505), .A (nx38823)) ;
    inv02 ix38506 (.Y (nx38507), .A (nx38823)) ;
    inv02 ix38508 (.Y (nx38509), .A (nx38823)) ;
    inv02 ix38510 (.Y (nx38511), .A (nx38823)) ;
    inv02 ix38512 (.Y (nx38513), .A (nx38825)) ;
    inv02 ix38514 (.Y (nx38515), .A (nx38825)) ;
    inv02 ix38516 (.Y (nx38517), .A (nx38825)) ;
    inv02 ix38518 (.Y (nx38519), .A (nx38825)) ;
    inv02 ix38520 (.Y (nx38521), .A (sumInput[12])) ;
    inv02 ix38522 (.Y (nx38523), .A (nx38827)) ;
    inv02 ix38524 (.Y (nx38525), .A (nx38827)) ;
    inv02 ix38526 (.Y (nx38527), .A (nx38827)) ;
    inv02 ix38528 (.Y (nx38529), .A (nx38827)) ;
    inv02 ix38530 (.Y (nx38531), .A (nx38827)) ;
    inv02 ix38532 (.Y (nx38533), .A (nx38829)) ;
    inv02 ix38534 (.Y (nx38535), .A (nx38829)) ;
    inv02 ix38536 (.Y (nx38537), .A (nx38829)) ;
    inv02 ix38538 (.Y (nx38539), .A (nx38829)) ;
    inv02 ix38540 (.Y (nx38541), .A (sumInput[11])) ;
    inv02 ix38542 (.Y (nx38543), .A (nx38831)) ;
    inv02 ix38544 (.Y (nx38545), .A (nx38831)) ;
    inv02 ix38546 (.Y (nx38547), .A (nx38831)) ;
    inv02 ix38548 (.Y (nx38549), .A (nx38831)) ;
    inv02 ix38550 (.Y (nx38551), .A (nx38831)) ;
    inv02 ix38552 (.Y (nx38553), .A (nx38833)) ;
    inv02 ix38554 (.Y (nx38555), .A (nx38833)) ;
    inv02 ix38556 (.Y (nx38557), .A (nx38833)) ;
    inv02 ix38558 (.Y (nx38559), .A (nx38833)) ;
    inv02 ix38560 (.Y (nx38561), .A (sumInput[10])) ;
    inv02 ix38562 (.Y (nx38563), .A (nx38835)) ;
    inv02 ix38564 (.Y (nx38565), .A (nx38835)) ;
    inv02 ix38566 (.Y (nx38567), .A (nx38835)) ;
    inv02 ix38568 (.Y (nx38569), .A (nx38835)) ;
    inv02 ix38570 (.Y (nx38571), .A (nx38835)) ;
    inv02 ix38572 (.Y (nx38573), .A (nx38837)) ;
    inv02 ix38574 (.Y (nx38575), .A (nx38837)) ;
    inv02 ix38576 (.Y (nx38577), .A (nx38837)) ;
    inv02 ix38578 (.Y (nx38579), .A (nx38837)) ;
    inv02 ix38580 (.Y (nx38581), .A (sumInput[9])) ;
    inv02 ix38582 (.Y (nx38583), .A (nx38839)) ;
    inv02 ix38584 (.Y (nx38585), .A (nx38839)) ;
    inv02 ix38586 (.Y (nx38587), .A (nx38839)) ;
    inv02 ix38588 (.Y (nx38589), .A (nx38839)) ;
    inv02 ix38590 (.Y (nx38591), .A (nx38839)) ;
    inv02 ix38592 (.Y (nx38593), .A (nx38841)) ;
    inv02 ix38594 (.Y (nx38595), .A (nx38841)) ;
    inv02 ix38596 (.Y (nx38597), .A (nx38841)) ;
    inv02 ix38598 (.Y (nx38599), .A (nx38841)) ;
    inv02 ix38600 (.Y (nx38601), .A (sumInput[8])) ;
    inv02 ix38602 (.Y (nx38603), .A (nx38843)) ;
    inv02 ix38604 (.Y (nx38605), .A (nx38843)) ;
    inv02 ix38606 (.Y (nx38607), .A (nx38843)) ;
    inv02 ix38608 (.Y (nx38609), .A (nx38843)) ;
    inv02 ix38610 (.Y (nx38611), .A (nx38843)) ;
    inv02 ix38612 (.Y (nx38613), .A (nx38845)) ;
    inv02 ix38614 (.Y (nx38615), .A (nx38845)) ;
    inv02 ix38616 (.Y (nx38617), .A (nx38845)) ;
    inv02 ix38618 (.Y (nx38619), .A (nx38845)) ;
    inv02 ix38620 (.Y (nx38621), .A (sumInput[7])) ;
    inv02 ix38622 (.Y (nx38623), .A (nx38847)) ;
    inv02 ix38624 (.Y (nx38625), .A (nx38847)) ;
    inv02 ix38626 (.Y (nx38627), .A (nx38847)) ;
    inv02 ix38628 (.Y (nx38629), .A (nx38847)) ;
    inv02 ix38630 (.Y (nx38631), .A (nx38847)) ;
    inv02 ix38632 (.Y (nx38633), .A (nx38849)) ;
    inv02 ix38634 (.Y (nx38635), .A (nx38849)) ;
    inv02 ix38636 (.Y (nx38637), .A (nx38849)) ;
    inv02 ix38638 (.Y (nx38639), .A (nx38849)) ;
    inv02 ix38640 (.Y (nx38641), .A (sumInput[6])) ;
    inv02 ix38642 (.Y (nx38643), .A (nx38851)) ;
    inv02 ix38644 (.Y (nx38645), .A (nx38851)) ;
    inv02 ix38646 (.Y (nx38647), .A (nx38851)) ;
    inv02 ix38648 (.Y (nx38649), .A (nx38851)) ;
    inv02 ix38650 (.Y (nx38651), .A (nx38851)) ;
    inv02 ix38652 (.Y (nx38653), .A (nx38853)) ;
    inv02 ix38654 (.Y (nx38655), .A (nx38853)) ;
    inv02 ix38656 (.Y (nx38657), .A (nx38853)) ;
    inv02 ix38658 (.Y (nx38659), .A (nx38853)) ;
    inv02 ix38660 (.Y (nx38661), .A (sumInput[5])) ;
    inv02 ix38662 (.Y (nx38663), .A (nx38855)) ;
    inv02 ix38664 (.Y (nx38665), .A (nx38855)) ;
    inv02 ix38666 (.Y (nx38667), .A (nx38855)) ;
    inv02 ix38668 (.Y (nx38669), .A (nx38855)) ;
    inv02 ix38670 (.Y (nx38671), .A (nx38855)) ;
    inv02 ix38672 (.Y (nx38673), .A (nx38857)) ;
    inv02 ix38674 (.Y (nx38675), .A (nx38857)) ;
    inv02 ix38676 (.Y (nx38677), .A (nx38857)) ;
    inv02 ix38678 (.Y (nx38679), .A (nx38857)) ;
    inv02 ix38680 (.Y (nx38681), .A (sumInput[4])) ;
    inv02 ix38682 (.Y (nx38683), .A (nx38859)) ;
    inv02 ix38684 (.Y (nx38685), .A (nx38859)) ;
    inv02 ix38686 (.Y (nx38687), .A (nx38859)) ;
    inv02 ix38688 (.Y (nx38689), .A (nx38859)) ;
    inv02 ix38690 (.Y (nx38691), .A (nx38859)) ;
    inv02 ix38692 (.Y (nx38693), .A (nx38861)) ;
    inv02 ix38694 (.Y (nx38695), .A (nx38861)) ;
    inv02 ix38696 (.Y (nx38697), .A (nx38861)) ;
    inv02 ix38698 (.Y (nx38699), .A (nx38861)) ;
    inv02 ix38700 (.Y (nx38701), .A (sumInput[3])) ;
    inv02 ix38702 (.Y (nx38703), .A (nx38863)) ;
    inv02 ix38704 (.Y (nx38705), .A (nx38863)) ;
    inv02 ix38706 (.Y (nx38707), .A (nx38863)) ;
    inv02 ix38708 (.Y (nx38709), .A (nx38863)) ;
    inv02 ix38710 (.Y (nx38711), .A (nx38863)) ;
    inv02 ix38712 (.Y (nx38713), .A (nx38865)) ;
    inv02 ix38714 (.Y (nx38715), .A (nx38865)) ;
    inv02 ix38716 (.Y (nx38717), .A (nx38865)) ;
    inv02 ix38718 (.Y (nx38719), .A (nx38865)) ;
    inv02 ix38720 (.Y (nx38721), .A (sumInput[2])) ;
    inv02 ix38722 (.Y (nx38723), .A (nx38867)) ;
    inv02 ix38724 (.Y (nx38725), .A (nx38867)) ;
    inv02 ix38726 (.Y (nx38727), .A (nx38867)) ;
    inv02 ix38728 (.Y (nx38729), .A (nx38867)) ;
    inv02 ix38730 (.Y (nx38731), .A (nx38867)) ;
    inv02 ix38732 (.Y (nx38733), .A (nx38869)) ;
    inv02 ix38734 (.Y (nx38735), .A (nx38869)) ;
    inv02 ix38736 (.Y (nx38737), .A (nx38869)) ;
    inv02 ix38738 (.Y (nx38739), .A (nx38869)) ;
    inv02 ix38740 (.Y (nx38741), .A (sumInput[1])) ;
    inv02 ix38742 (.Y (nx38743), .A (nx38871)) ;
    inv02 ix38744 (.Y (nx38745), .A (nx38871)) ;
    inv02 ix38746 (.Y (nx38747), .A (nx38871)) ;
    inv02 ix38748 (.Y (nx38749), .A (nx38871)) ;
    inv02 ix38750 (.Y (nx38751), .A (nx38871)) ;
    inv02 ix38752 (.Y (nx38753), .A (nx38873)) ;
    inv02 ix38754 (.Y (nx38755), .A (nx38873)) ;
    inv02 ix38756 (.Y (nx38757), .A (nx38873)) ;
    inv02 ix38758 (.Y (nx38759), .A (nx38873)) ;
    inv02 ix38760 (.Y (nx38761), .A (sumInput[0])) ;
    inv02 ix38762 (.Y (nx38763), .A (nx38875)) ;
    inv02 ix38764 (.Y (nx38765), .A (nx38875)) ;
    inv02 ix38766 (.Y (nx38767), .A (nx38875)) ;
    inv02 ix38768 (.Y (nx38769), .A (nx38875)) ;
    inv02 ix38770 (.Y (nx38771), .A (nx38875)) ;
    inv02 ix38772 (.Y (nx38773), .A (nx38877)) ;
    inv02 ix38774 (.Y (nx38775), .A (nx38877)) ;
    inv02 ix38776 (.Y (nx38777), .A (nx38877)) ;
    inv02 ix38778 (.Y (nx38779), .A (nx38877)) ;
    inv01 ix38784 (.Y (nx38785), .A (nx34751)) ;
    inv01 ix38786 (.Y (nx38787), .A (nx34751)) ;
    inv01 ix38788 (.Y (nx38789), .A (nx34893)) ;
    inv01 ix38790 (.Y (nx38791), .A (nx34893)) ;
    inv01 ix38792 (.Y (nx38793), .A (nx35035)) ;
    inv01 ix38794 (.Y (nx38795), .A (nx35035)) ;
    inv01 ix38796 (.Y (nx38797), .A (nx35177)) ;
    inv01 ix38798 (.Y (nx38799), .A (nx35177)) ;
    inv01 ix38800 (.Y (nx38801), .A (nx35319)) ;
    inv01 ix38802 (.Y (nx38803), .A (nx35319)) ;
    inv01 ix38804 (.Y (nx38805), .A (nx35461)) ;
    inv01 ix38806 (.Y (nx38807), .A (nx35461)) ;
    inv01 ix38808 (.Y (nx38809), .A (nx35603)) ;
    inv01 ix38810 (.Y (nx38811), .A (nx35603)) ;
    inv01 ix38812 (.Y (nx38813), .A (nx35603)) ;
    inv01 ix38814 (.Y (nx38815), .A (nx38461)) ;
    inv01 ix38816 (.Y (nx38817), .A (nx38461)) ;
    inv01 ix38818 (.Y (nx38819), .A (nx38481)) ;
    inv01 ix38820 (.Y (nx38821), .A (nx38481)) ;
    inv01 ix38822 (.Y (nx38823), .A (nx38501)) ;
    inv01 ix38824 (.Y (nx38825), .A (nx38501)) ;
    inv01 ix38826 (.Y (nx38827), .A (nx38521)) ;
    inv01 ix38828 (.Y (nx38829), .A (nx38521)) ;
    inv01 ix38830 (.Y (nx38831), .A (nx38541)) ;
    inv01 ix38832 (.Y (nx38833), .A (nx38541)) ;
    inv01 ix38834 (.Y (nx38835), .A (nx38561)) ;
    inv01 ix38836 (.Y (nx38837), .A (nx38561)) ;
    inv01 ix38838 (.Y (nx38839), .A (nx38581)) ;
    inv01 ix38840 (.Y (nx38841), .A (nx38581)) ;
    inv01 ix38842 (.Y (nx38843), .A (nx38601)) ;
    inv01 ix38844 (.Y (nx38845), .A (nx38601)) ;
    inv01 ix38846 (.Y (nx38847), .A (nx38621)) ;
    inv01 ix38848 (.Y (nx38849), .A (nx38621)) ;
    inv01 ix38850 (.Y (nx38851), .A (nx38641)) ;
    inv01 ix38852 (.Y (nx38853), .A (nx38641)) ;
    inv01 ix38854 (.Y (nx38855), .A (nx38661)) ;
    inv01 ix38856 (.Y (nx38857), .A (nx38661)) ;
    inv01 ix38858 (.Y (nx38859), .A (nx38681)) ;
    inv01 ix38860 (.Y (nx38861), .A (nx38681)) ;
    inv01 ix38862 (.Y (nx38863), .A (nx38701)) ;
    inv01 ix38864 (.Y (nx38865), .A (nx38701)) ;
    inv01 ix38866 (.Y (nx38867), .A (nx38721)) ;
    inv01 ix38868 (.Y (nx38869), .A (nx38721)) ;
    inv01 ix38870 (.Y (nx38871), .A (nx38741)) ;
    inv01 ix38872 (.Y (nx38873), .A (nx38741)) ;
    inv01 ix38874 (.Y (nx38875), .A (nx38761)) ;
    inv01 ix38876 (.Y (nx38877), .A (nx38761)) ;
    inv01 ix38878 (.Y (nx38879), .A (nx33639)) ;
    inv01 ix38880 (.Y (nx38881), .A (nx33639)) ;
    inv01 ix38882 (.Y (nx38883), .A (nx33639)) ;
    inv01 ix38884 (.Y (nx38885), .A (nx33639)) ;
    inv01 ix38886 (.Y (nx38887), .A (nx33639)) ;
    inv01 ix38888 (.Y (nx38889), .A (nx33639)) ;
    inv01 ix38890 (.Y (nx38891), .A (nx33639)) ;
    inv01 ix38892 (.Y (nx38893), .A (nx33639)) ;
    inv01 ix38894 (.Y (nx38895), .A (nx33639)) ;
    inv01 ix38896 (.Y (nx38897), .A (nx33639)) ;
    inv01 ix38898 (.Y (nx38899), .A (nx34609)) ;
    inv01 ix38900 (.Y (nx38901), .A (nx34609)) ;
endmodule


module Counter_9 ( en, reset, clk, count ) ;

    input en ;
    input reset ;
    input clk ;
    output [8:0]count ;

    wire addedOne_8, addedOne_7, addedOne_6, addedOne_5, addedOne_4, addedOne_3, 
         addedOne_2, addedOne_1, addedOne_0, finalReset, oneSignal_8, PWR;
    wire [0:0] \$dummy ;




    Reg_9 counterReg (.D ({addedOne_8,addedOne_7,addedOne_6,addedOne_5,
          addedOne_4,addedOne_3,addedOne_2,addedOne_1,addedOne_0}), .en (en), .clk (
          clk), .rst (finalReset), .Q ({count[8],count[7],count[6],count[5],
          count[4],count[3],count[2],count[1],count[0]})) ;
    NBitAdder_9 nextCount (.a ({count[8],count[7],count[6],count[5],count[4],
                count[3],count[2],count[1],count[0]}), .b ({oneSignal_8,
                oneSignal_8,oneSignal_8,oneSignal_8,oneSignal_8,oneSignal_8,
                oneSignal_8,oneSignal_8,oneSignal_8}), .carryIn (PWR), .sum ({
                addedOne_8,addedOne_7,addedOne_6,addedOne_5,addedOne_4,
                addedOne_3,addedOne_2,addedOne_1,addedOne_0}), .carryOut (
                \$dummy [0])) ;
    fake_vcc ix29 (.Y (PWR)) ;
    fake_gnd ix27 (.Y (oneSignal_8)) ;
    and02 ix1 (.Y (finalReset), .A0 (reset), .A1 (clk)) ;
endmodule


module NBitAdder_9 ( a, b, carryIn, sum, carryOut ) ;

    input [8:0]a ;
    input [8:0]b ;
    input carryIn ;
    output [8:0]sum ;
    output carryOut ;

    wire temp_7, temp_6, temp_5, temp_4, temp_3, temp_2, temp_1, temp_0;



    FullAdder f0 (.a (a[0]), .b (b[0]), .cin (carryIn), .s (sum[0]), .cout (
              temp_0)) ;
    FullAdder loop1_1_fx (.a (a[1]), .b (b[1]), .cin (temp_0), .s (sum[1]), .cout (
              temp_1)) ;
    FullAdder loop1_2_fx (.a (a[2]), .b (b[2]), .cin (temp_1), .s (sum[2]), .cout (
              temp_2)) ;
    FullAdder loop1_3_fx (.a (a[3]), .b (b[3]), .cin (temp_2), .s (sum[3]), .cout (
              temp_3)) ;
    FullAdder loop1_4_fx (.a (a[4]), .b (b[4]), .cin (temp_3), .s (sum[4]), .cout (
              temp_4)) ;
    FullAdder loop1_5_fx (.a (a[5]), .b (b[5]), .cin (temp_4), .s (sum[5]), .cout (
              temp_5)) ;
    FullAdder loop1_6_fx (.a (a[6]), .b (b[6]), .cin (temp_5), .s (sum[6]), .cout (
              temp_6)) ;
    FullAdder loop1_7_fx (.a (a[7]), .b (b[7]), .cin (temp_6), .s (sum[7]), .cout (
              temp_7)) ;
    FullAdder loop1_8_fx (.a (a[8]), .b (b[8]), .cin (temp_7), .s (sum[8]), .cout (
              carryOut)) ;
endmodule


module Reg_9 ( D, en, clk, rst, Q ) ;

    input [8:0]D ;
    input en ;
    input clk ;
    input rst ;
    output [8:0]Q ;

    wire nx144, nx154, nx164, nx174, nx184, nx194, nx204, nx214, nx224, nx266, 
         nx268, nx270, nx272, nx274, nx276;
    wire [8:0] \$dummy ;




    dffr reg_Q_0 (.Q (Q[0]), .QB (\$dummy [0]), .D (nx144), .CLK (nx270), .R (
         nx266)) ;
    mux21_ni ix145 (.Y (nx144), .A0 (Q[0]), .A1 (D[0]), .S0 (nx274)) ;
    dffr reg_Q_1 (.Q (Q[1]), .QB (\$dummy [1]), .D (nx154), .CLK (nx270), .R (
         nx266)) ;
    mux21_ni ix155 (.Y (nx154), .A0 (Q[1]), .A1 (D[1]), .S0 (nx274)) ;
    dffr reg_Q_2 (.Q (Q[2]), .QB (\$dummy [2]), .D (nx164), .CLK (nx270), .R (
         nx266)) ;
    mux21_ni ix165 (.Y (nx164), .A0 (Q[2]), .A1 (D[2]), .S0 (nx274)) ;
    dffr reg_Q_3 (.Q (Q[3]), .QB (\$dummy [3]), .D (nx174), .CLK (nx270), .R (
         nx266)) ;
    mux21_ni ix175 (.Y (nx174), .A0 (Q[3]), .A1 (D[3]), .S0 (nx274)) ;
    dffr reg_Q_4 (.Q (Q[4]), .QB (\$dummy [4]), .D (nx184), .CLK (nx270), .R (
         nx266)) ;
    mux21_ni ix185 (.Y (nx184), .A0 (Q[4]), .A1 (D[4]), .S0 (nx274)) ;
    dffr reg_Q_5 (.Q (Q[5]), .QB (\$dummy [5]), .D (nx194), .CLK (nx270), .R (
         nx266)) ;
    mux21_ni ix195 (.Y (nx194), .A0 (Q[5]), .A1 (D[5]), .S0 (nx274)) ;
    dffr reg_Q_6 (.Q (Q[6]), .QB (\$dummy [6]), .D (nx204), .CLK (nx270), .R (
         nx266)) ;
    mux21_ni ix205 (.Y (nx204), .A0 (Q[6]), .A1 (D[6]), .S0 (nx274)) ;
    dffr reg_Q_7 (.Q (Q[7]), .QB (\$dummy [7]), .D (nx214), .CLK (nx272), .R (
         nx268)) ;
    mux21_ni ix215 (.Y (nx214), .A0 (Q[7]), .A1 (D[7]), .S0 (nx276)) ;
    dffr reg_Q_8 (.Q (Q[8]), .QB (\$dummy [8]), .D (nx224), .CLK (nx272), .R (
         nx268)) ;
    mux21_ni ix225 (.Y (nx224), .A0 (Q[8]), .A1 (D[8]), .S0 (nx276)) ;
    buf02 ix265 (.Y (nx266), .A (rst)) ;
    buf02 ix267 (.Y (nx268), .A (rst)) ;
    buf02 ix269 (.Y (nx270), .A (clk)) ;
    buf02 ix271 (.Y (nx272), .A (clk)) ;
    buf02 ix273 (.Y (nx274), .A (en)) ;
    buf02 ix275 (.Y (nx276), .A (en)) ;
endmodule


module Mux_512 ( inputs_0__15, inputs_0__14, inputs_0__13, inputs_0__12, 
                 inputs_0__11, inputs_0__10, inputs_0__9, inputs_0__8, 
                 inputs_0__7, inputs_0__6, inputs_0__5, inputs_0__4, inputs_0__3, 
                 inputs_0__2, inputs_0__1, inputs_0__0, inputs_1__15, 
                 inputs_1__14, inputs_1__13, inputs_1__12, inputs_1__11, 
                 inputs_1__10, inputs_1__9, inputs_1__8, inputs_1__7, 
                 inputs_1__6, inputs_1__5, inputs_1__4, inputs_1__3, inputs_1__2, 
                 inputs_1__1, inputs_1__0, inputs_2__15, inputs_2__14, 
                 inputs_2__13, inputs_2__12, inputs_2__11, inputs_2__10, 
                 inputs_2__9, inputs_2__8, inputs_2__7, inputs_2__6, inputs_2__5, 
                 inputs_2__4, inputs_2__3, inputs_2__2, inputs_2__1, inputs_2__0, 
                 inputs_3__15, inputs_3__14, inputs_3__13, inputs_3__12, 
                 inputs_3__11, inputs_3__10, inputs_3__9, inputs_3__8, 
                 inputs_3__7, inputs_3__6, inputs_3__5, inputs_3__4, inputs_3__3, 
                 inputs_3__2, inputs_3__1, inputs_3__0, inputs_4__15, 
                 inputs_4__14, inputs_4__13, inputs_4__12, inputs_4__11, 
                 inputs_4__10, inputs_4__9, inputs_4__8, inputs_4__7, 
                 inputs_4__6, inputs_4__5, inputs_4__4, inputs_4__3, inputs_4__2, 
                 inputs_4__1, inputs_4__0, inputs_5__15, inputs_5__14, 
                 inputs_5__13, inputs_5__12, inputs_5__11, inputs_5__10, 
                 inputs_5__9, inputs_5__8, inputs_5__7, inputs_5__6, inputs_5__5, 
                 inputs_5__4, inputs_5__3, inputs_5__2, inputs_5__1, inputs_5__0, 
                 inputs_6__15, inputs_6__14, inputs_6__13, inputs_6__12, 
                 inputs_6__11, inputs_6__10, inputs_6__9, inputs_6__8, 
                 inputs_6__7, inputs_6__6, inputs_6__5, inputs_6__4, inputs_6__3, 
                 inputs_6__2, inputs_6__1, inputs_6__0, inputs_7__15, 
                 inputs_7__14, inputs_7__13, inputs_7__12, inputs_7__11, 
                 inputs_7__10, inputs_7__9, inputs_7__8, inputs_7__7, 
                 inputs_7__6, inputs_7__5, inputs_7__4, inputs_7__3, inputs_7__2, 
                 inputs_7__1, inputs_7__0, inputs_8__15, inputs_8__14, 
                 inputs_8__13, inputs_8__12, inputs_8__11, inputs_8__10, 
                 inputs_8__9, inputs_8__8, inputs_8__7, inputs_8__6, inputs_8__5, 
                 inputs_8__4, inputs_8__3, inputs_8__2, inputs_8__1, inputs_8__0, 
                 inputs_9__15, inputs_9__14, inputs_9__13, inputs_9__12, 
                 inputs_9__11, inputs_9__10, inputs_9__9, inputs_9__8, 
                 inputs_9__7, inputs_9__6, inputs_9__5, inputs_9__4, inputs_9__3, 
                 inputs_9__2, inputs_9__1, inputs_9__0, inputs_10__15, 
                 inputs_10__14, inputs_10__13, inputs_10__12, inputs_10__11, 
                 inputs_10__10, inputs_10__9, inputs_10__8, inputs_10__7, 
                 inputs_10__6, inputs_10__5, inputs_10__4, inputs_10__3, 
                 inputs_10__2, inputs_10__1, inputs_10__0, inputs_11__15, 
                 inputs_11__14, inputs_11__13, inputs_11__12, inputs_11__11, 
                 inputs_11__10, inputs_11__9, inputs_11__8, inputs_11__7, 
                 inputs_11__6, inputs_11__5, inputs_11__4, inputs_11__3, 
                 inputs_11__2, inputs_11__1, inputs_11__0, inputs_12__15, 
                 inputs_12__14, inputs_12__13, inputs_12__12, inputs_12__11, 
                 inputs_12__10, inputs_12__9, inputs_12__8, inputs_12__7, 
                 inputs_12__6, inputs_12__5, inputs_12__4, inputs_12__3, 
                 inputs_12__2, inputs_12__1, inputs_12__0, inputs_13__15, 
                 inputs_13__14, inputs_13__13, inputs_13__12, inputs_13__11, 
                 inputs_13__10, inputs_13__9, inputs_13__8, inputs_13__7, 
                 inputs_13__6, inputs_13__5, inputs_13__4, inputs_13__3, 
                 inputs_13__2, inputs_13__1, inputs_13__0, inputs_14__15, 
                 inputs_14__14, inputs_14__13, inputs_14__12, inputs_14__11, 
                 inputs_14__10, inputs_14__9, inputs_14__8, inputs_14__7, 
                 inputs_14__6, inputs_14__5, inputs_14__4, inputs_14__3, 
                 inputs_14__2, inputs_14__1, inputs_14__0, inputs_15__15, 
                 inputs_15__14, inputs_15__13, inputs_15__12, inputs_15__11, 
                 inputs_15__10, inputs_15__9, inputs_15__8, inputs_15__7, 
                 inputs_15__6, inputs_15__5, inputs_15__4, inputs_15__3, 
                 inputs_15__2, inputs_15__1, inputs_15__0, inputs_16__15, 
                 inputs_16__14, inputs_16__13, inputs_16__12, inputs_16__11, 
                 inputs_16__10, inputs_16__9, inputs_16__8, inputs_16__7, 
                 inputs_16__6, inputs_16__5, inputs_16__4, inputs_16__3, 
                 inputs_16__2, inputs_16__1, inputs_16__0, inputs_17__15, 
                 inputs_17__14, inputs_17__13, inputs_17__12, inputs_17__11, 
                 inputs_17__10, inputs_17__9, inputs_17__8, inputs_17__7, 
                 inputs_17__6, inputs_17__5, inputs_17__4, inputs_17__3, 
                 inputs_17__2, inputs_17__1, inputs_17__0, inputs_18__15, 
                 inputs_18__14, inputs_18__13, inputs_18__12, inputs_18__11, 
                 inputs_18__10, inputs_18__9, inputs_18__8, inputs_18__7, 
                 inputs_18__6, inputs_18__5, inputs_18__4, inputs_18__3, 
                 inputs_18__2, inputs_18__1, inputs_18__0, inputs_19__15, 
                 inputs_19__14, inputs_19__13, inputs_19__12, inputs_19__11, 
                 inputs_19__10, inputs_19__9, inputs_19__8, inputs_19__7, 
                 inputs_19__6, inputs_19__5, inputs_19__4, inputs_19__3, 
                 inputs_19__2, inputs_19__1, inputs_19__0, inputs_20__15, 
                 inputs_20__14, inputs_20__13, inputs_20__12, inputs_20__11, 
                 inputs_20__10, inputs_20__9, inputs_20__8, inputs_20__7, 
                 inputs_20__6, inputs_20__5, inputs_20__4, inputs_20__3, 
                 inputs_20__2, inputs_20__1, inputs_20__0, inputs_21__15, 
                 inputs_21__14, inputs_21__13, inputs_21__12, inputs_21__11, 
                 inputs_21__10, inputs_21__9, inputs_21__8, inputs_21__7, 
                 inputs_21__6, inputs_21__5, inputs_21__4, inputs_21__3, 
                 inputs_21__2, inputs_21__1, inputs_21__0, inputs_22__15, 
                 inputs_22__14, inputs_22__13, inputs_22__12, inputs_22__11, 
                 inputs_22__10, inputs_22__9, inputs_22__8, inputs_22__7, 
                 inputs_22__6, inputs_22__5, inputs_22__4, inputs_22__3, 
                 inputs_22__2, inputs_22__1, inputs_22__0, inputs_23__15, 
                 inputs_23__14, inputs_23__13, inputs_23__12, inputs_23__11, 
                 inputs_23__10, inputs_23__9, inputs_23__8, inputs_23__7, 
                 inputs_23__6, inputs_23__5, inputs_23__4, inputs_23__3, 
                 inputs_23__2, inputs_23__1, inputs_23__0, inputs_24__15, 
                 inputs_24__14, inputs_24__13, inputs_24__12, inputs_24__11, 
                 inputs_24__10, inputs_24__9, inputs_24__8, inputs_24__7, 
                 inputs_24__6, inputs_24__5, inputs_24__4, inputs_24__3, 
                 inputs_24__2, inputs_24__1, inputs_24__0, inputs_25__15, 
                 inputs_25__14, inputs_25__13, inputs_25__12, inputs_25__11, 
                 inputs_25__10, inputs_25__9, inputs_25__8, inputs_25__7, 
                 inputs_25__6, inputs_25__5, inputs_25__4, inputs_25__3, 
                 inputs_25__2, inputs_25__1, inputs_25__0, inputs_26__15, 
                 inputs_26__14, inputs_26__13, inputs_26__12, inputs_26__11, 
                 inputs_26__10, inputs_26__9, inputs_26__8, inputs_26__7, 
                 inputs_26__6, inputs_26__5, inputs_26__4, inputs_26__3, 
                 inputs_26__2, inputs_26__1, inputs_26__0, inputs_27__15, 
                 inputs_27__14, inputs_27__13, inputs_27__12, inputs_27__11, 
                 inputs_27__10, inputs_27__9, inputs_27__8, inputs_27__7, 
                 inputs_27__6, inputs_27__5, inputs_27__4, inputs_27__3, 
                 inputs_27__2, inputs_27__1, inputs_27__0, inputs_28__15, 
                 inputs_28__14, inputs_28__13, inputs_28__12, inputs_28__11, 
                 inputs_28__10, inputs_28__9, inputs_28__8, inputs_28__7, 
                 inputs_28__6, inputs_28__5, inputs_28__4, inputs_28__3, 
                 inputs_28__2, inputs_28__1, inputs_28__0, inputs_29__15, 
                 inputs_29__14, inputs_29__13, inputs_29__12, inputs_29__11, 
                 inputs_29__10, inputs_29__9, inputs_29__8, inputs_29__7, 
                 inputs_29__6, inputs_29__5, inputs_29__4, inputs_29__3, 
                 inputs_29__2, inputs_29__1, inputs_29__0, inputs_30__15, 
                 inputs_30__14, inputs_30__13, inputs_30__12, inputs_30__11, 
                 inputs_30__10, inputs_30__9, inputs_30__8, inputs_30__7, 
                 inputs_30__6, inputs_30__5, inputs_30__4, inputs_30__3, 
                 inputs_30__2, inputs_30__1, inputs_30__0, inputs_31__15, 
                 inputs_31__14, inputs_31__13, inputs_31__12, inputs_31__11, 
                 inputs_31__10, inputs_31__9, inputs_31__8, inputs_31__7, 
                 inputs_31__6, inputs_31__5, inputs_31__4, inputs_31__3, 
                 inputs_31__2, inputs_31__1, inputs_31__0, inputs_32__15, 
                 inputs_32__14, inputs_32__13, inputs_32__12, inputs_32__11, 
                 inputs_32__10, inputs_32__9, inputs_32__8, inputs_32__7, 
                 inputs_32__6, inputs_32__5, inputs_32__4, inputs_32__3, 
                 inputs_32__2, inputs_32__1, inputs_32__0, inputs_33__15, 
                 inputs_33__14, inputs_33__13, inputs_33__12, inputs_33__11, 
                 inputs_33__10, inputs_33__9, inputs_33__8, inputs_33__7, 
                 inputs_33__6, inputs_33__5, inputs_33__4, inputs_33__3, 
                 inputs_33__2, inputs_33__1, inputs_33__0, inputs_34__15, 
                 inputs_34__14, inputs_34__13, inputs_34__12, inputs_34__11, 
                 inputs_34__10, inputs_34__9, inputs_34__8, inputs_34__7, 
                 inputs_34__6, inputs_34__5, inputs_34__4, inputs_34__3, 
                 inputs_34__2, inputs_34__1, inputs_34__0, inputs_35__15, 
                 inputs_35__14, inputs_35__13, inputs_35__12, inputs_35__11, 
                 inputs_35__10, inputs_35__9, inputs_35__8, inputs_35__7, 
                 inputs_35__6, inputs_35__5, inputs_35__4, inputs_35__3, 
                 inputs_35__2, inputs_35__1, inputs_35__0, inputs_36__15, 
                 inputs_36__14, inputs_36__13, inputs_36__12, inputs_36__11, 
                 inputs_36__10, inputs_36__9, inputs_36__8, inputs_36__7, 
                 inputs_36__6, inputs_36__5, inputs_36__4, inputs_36__3, 
                 inputs_36__2, inputs_36__1, inputs_36__0, inputs_37__15, 
                 inputs_37__14, inputs_37__13, inputs_37__12, inputs_37__11, 
                 inputs_37__10, inputs_37__9, inputs_37__8, inputs_37__7, 
                 inputs_37__6, inputs_37__5, inputs_37__4, inputs_37__3, 
                 inputs_37__2, inputs_37__1, inputs_37__0, inputs_38__15, 
                 inputs_38__14, inputs_38__13, inputs_38__12, inputs_38__11, 
                 inputs_38__10, inputs_38__9, inputs_38__8, inputs_38__7, 
                 inputs_38__6, inputs_38__5, inputs_38__4, inputs_38__3, 
                 inputs_38__2, inputs_38__1, inputs_38__0, inputs_39__15, 
                 inputs_39__14, inputs_39__13, inputs_39__12, inputs_39__11, 
                 inputs_39__10, inputs_39__9, inputs_39__8, inputs_39__7, 
                 inputs_39__6, inputs_39__5, inputs_39__4, inputs_39__3, 
                 inputs_39__2, inputs_39__1, inputs_39__0, inputs_40__15, 
                 inputs_40__14, inputs_40__13, inputs_40__12, inputs_40__11, 
                 inputs_40__10, inputs_40__9, inputs_40__8, inputs_40__7, 
                 inputs_40__6, inputs_40__5, inputs_40__4, inputs_40__3, 
                 inputs_40__2, inputs_40__1, inputs_40__0, inputs_41__15, 
                 inputs_41__14, inputs_41__13, inputs_41__12, inputs_41__11, 
                 inputs_41__10, inputs_41__9, inputs_41__8, inputs_41__7, 
                 inputs_41__6, inputs_41__5, inputs_41__4, inputs_41__3, 
                 inputs_41__2, inputs_41__1, inputs_41__0, inputs_42__15, 
                 inputs_42__14, inputs_42__13, inputs_42__12, inputs_42__11, 
                 inputs_42__10, inputs_42__9, inputs_42__8, inputs_42__7, 
                 inputs_42__6, inputs_42__5, inputs_42__4, inputs_42__3, 
                 inputs_42__2, inputs_42__1, inputs_42__0, inputs_43__15, 
                 inputs_43__14, inputs_43__13, inputs_43__12, inputs_43__11, 
                 inputs_43__10, inputs_43__9, inputs_43__8, inputs_43__7, 
                 inputs_43__6, inputs_43__5, inputs_43__4, inputs_43__3, 
                 inputs_43__2, inputs_43__1, inputs_43__0, inputs_44__15, 
                 inputs_44__14, inputs_44__13, inputs_44__12, inputs_44__11, 
                 inputs_44__10, inputs_44__9, inputs_44__8, inputs_44__7, 
                 inputs_44__6, inputs_44__5, inputs_44__4, inputs_44__3, 
                 inputs_44__2, inputs_44__1, inputs_44__0, inputs_45__15, 
                 inputs_45__14, inputs_45__13, inputs_45__12, inputs_45__11, 
                 inputs_45__10, inputs_45__9, inputs_45__8, inputs_45__7, 
                 inputs_45__6, inputs_45__5, inputs_45__4, inputs_45__3, 
                 inputs_45__2, inputs_45__1, inputs_45__0, inputs_46__15, 
                 inputs_46__14, inputs_46__13, inputs_46__12, inputs_46__11, 
                 inputs_46__10, inputs_46__9, inputs_46__8, inputs_46__7, 
                 inputs_46__6, inputs_46__5, inputs_46__4, inputs_46__3, 
                 inputs_46__2, inputs_46__1, inputs_46__0, inputs_47__15, 
                 inputs_47__14, inputs_47__13, inputs_47__12, inputs_47__11, 
                 inputs_47__10, inputs_47__9, inputs_47__8, inputs_47__7, 
                 inputs_47__6, inputs_47__5, inputs_47__4, inputs_47__3, 
                 inputs_47__2, inputs_47__1, inputs_47__0, inputs_48__15, 
                 inputs_48__14, inputs_48__13, inputs_48__12, inputs_48__11, 
                 inputs_48__10, inputs_48__9, inputs_48__8, inputs_48__7, 
                 inputs_48__6, inputs_48__5, inputs_48__4, inputs_48__3, 
                 inputs_48__2, inputs_48__1, inputs_48__0, inputs_49__15, 
                 inputs_49__14, inputs_49__13, inputs_49__12, inputs_49__11, 
                 inputs_49__10, inputs_49__9, inputs_49__8, inputs_49__7, 
                 inputs_49__6, inputs_49__5, inputs_49__4, inputs_49__3, 
                 inputs_49__2, inputs_49__1, inputs_49__0, inputs_50__15, 
                 inputs_50__14, inputs_50__13, inputs_50__12, inputs_50__11, 
                 inputs_50__10, inputs_50__9, inputs_50__8, inputs_50__7, 
                 inputs_50__6, inputs_50__5, inputs_50__4, inputs_50__3, 
                 inputs_50__2, inputs_50__1, inputs_50__0, inputs_51__15, 
                 inputs_51__14, inputs_51__13, inputs_51__12, inputs_51__11, 
                 inputs_51__10, inputs_51__9, inputs_51__8, inputs_51__7, 
                 inputs_51__6, inputs_51__5, inputs_51__4, inputs_51__3, 
                 inputs_51__2, inputs_51__1, inputs_51__0, inputs_52__15, 
                 inputs_52__14, inputs_52__13, inputs_52__12, inputs_52__11, 
                 inputs_52__10, inputs_52__9, inputs_52__8, inputs_52__7, 
                 inputs_52__6, inputs_52__5, inputs_52__4, inputs_52__3, 
                 inputs_52__2, inputs_52__1, inputs_52__0, inputs_53__15, 
                 inputs_53__14, inputs_53__13, inputs_53__12, inputs_53__11, 
                 inputs_53__10, inputs_53__9, inputs_53__8, inputs_53__7, 
                 inputs_53__6, inputs_53__5, inputs_53__4, inputs_53__3, 
                 inputs_53__2, inputs_53__1, inputs_53__0, inputs_54__15, 
                 inputs_54__14, inputs_54__13, inputs_54__12, inputs_54__11, 
                 inputs_54__10, inputs_54__9, inputs_54__8, inputs_54__7, 
                 inputs_54__6, inputs_54__5, inputs_54__4, inputs_54__3, 
                 inputs_54__2, inputs_54__1, inputs_54__0, inputs_55__15, 
                 inputs_55__14, inputs_55__13, inputs_55__12, inputs_55__11, 
                 inputs_55__10, inputs_55__9, inputs_55__8, inputs_55__7, 
                 inputs_55__6, inputs_55__5, inputs_55__4, inputs_55__3, 
                 inputs_55__2, inputs_55__1, inputs_55__0, inputs_56__15, 
                 inputs_56__14, inputs_56__13, inputs_56__12, inputs_56__11, 
                 inputs_56__10, inputs_56__9, inputs_56__8, inputs_56__7, 
                 inputs_56__6, inputs_56__5, inputs_56__4, inputs_56__3, 
                 inputs_56__2, inputs_56__1, inputs_56__0, inputs_57__15, 
                 inputs_57__14, inputs_57__13, inputs_57__12, inputs_57__11, 
                 inputs_57__10, inputs_57__9, inputs_57__8, inputs_57__7, 
                 inputs_57__6, inputs_57__5, inputs_57__4, inputs_57__3, 
                 inputs_57__2, inputs_57__1, inputs_57__0, inputs_58__15, 
                 inputs_58__14, inputs_58__13, inputs_58__12, inputs_58__11, 
                 inputs_58__10, inputs_58__9, inputs_58__8, inputs_58__7, 
                 inputs_58__6, inputs_58__5, inputs_58__4, inputs_58__3, 
                 inputs_58__2, inputs_58__1, inputs_58__0, inputs_59__15, 
                 inputs_59__14, inputs_59__13, inputs_59__12, inputs_59__11, 
                 inputs_59__10, inputs_59__9, inputs_59__8, inputs_59__7, 
                 inputs_59__6, inputs_59__5, inputs_59__4, inputs_59__3, 
                 inputs_59__2, inputs_59__1, inputs_59__0, inputs_60__15, 
                 inputs_60__14, inputs_60__13, inputs_60__12, inputs_60__11, 
                 inputs_60__10, inputs_60__9, inputs_60__8, inputs_60__7, 
                 inputs_60__6, inputs_60__5, inputs_60__4, inputs_60__3, 
                 inputs_60__2, inputs_60__1, inputs_60__0, inputs_61__15, 
                 inputs_61__14, inputs_61__13, inputs_61__12, inputs_61__11, 
                 inputs_61__10, inputs_61__9, inputs_61__8, inputs_61__7, 
                 inputs_61__6, inputs_61__5, inputs_61__4, inputs_61__3, 
                 inputs_61__2, inputs_61__1, inputs_61__0, inputs_62__15, 
                 inputs_62__14, inputs_62__13, inputs_62__12, inputs_62__11, 
                 inputs_62__10, inputs_62__9, inputs_62__8, inputs_62__7, 
                 inputs_62__6, inputs_62__5, inputs_62__4, inputs_62__3, 
                 inputs_62__2, inputs_62__1, inputs_62__0, inputs_63__15, 
                 inputs_63__14, inputs_63__13, inputs_63__12, inputs_63__11, 
                 inputs_63__10, inputs_63__9, inputs_63__8, inputs_63__7, 
                 inputs_63__6, inputs_63__5, inputs_63__4, inputs_63__3, 
                 inputs_63__2, inputs_63__1, inputs_63__0, inputs_64__15, 
                 inputs_64__14, inputs_64__13, inputs_64__12, inputs_64__11, 
                 inputs_64__10, inputs_64__9, inputs_64__8, inputs_64__7, 
                 inputs_64__6, inputs_64__5, inputs_64__4, inputs_64__3, 
                 inputs_64__2, inputs_64__1, inputs_64__0, inputs_65__15, 
                 inputs_65__14, inputs_65__13, inputs_65__12, inputs_65__11, 
                 inputs_65__10, inputs_65__9, inputs_65__8, inputs_65__7, 
                 inputs_65__6, inputs_65__5, inputs_65__4, inputs_65__3, 
                 inputs_65__2, inputs_65__1, inputs_65__0, inputs_66__15, 
                 inputs_66__14, inputs_66__13, inputs_66__12, inputs_66__11, 
                 inputs_66__10, inputs_66__9, inputs_66__8, inputs_66__7, 
                 inputs_66__6, inputs_66__5, inputs_66__4, inputs_66__3, 
                 inputs_66__2, inputs_66__1, inputs_66__0, inputs_67__15, 
                 inputs_67__14, inputs_67__13, inputs_67__12, inputs_67__11, 
                 inputs_67__10, inputs_67__9, inputs_67__8, inputs_67__7, 
                 inputs_67__6, inputs_67__5, inputs_67__4, inputs_67__3, 
                 inputs_67__2, inputs_67__1, inputs_67__0, inputs_68__15, 
                 inputs_68__14, inputs_68__13, inputs_68__12, inputs_68__11, 
                 inputs_68__10, inputs_68__9, inputs_68__8, inputs_68__7, 
                 inputs_68__6, inputs_68__5, inputs_68__4, inputs_68__3, 
                 inputs_68__2, inputs_68__1, inputs_68__0, inputs_69__15, 
                 inputs_69__14, inputs_69__13, inputs_69__12, inputs_69__11, 
                 inputs_69__10, inputs_69__9, inputs_69__8, inputs_69__7, 
                 inputs_69__6, inputs_69__5, inputs_69__4, inputs_69__3, 
                 inputs_69__2, inputs_69__1, inputs_69__0, inputs_70__15, 
                 inputs_70__14, inputs_70__13, inputs_70__12, inputs_70__11, 
                 inputs_70__10, inputs_70__9, inputs_70__8, inputs_70__7, 
                 inputs_70__6, inputs_70__5, inputs_70__4, inputs_70__3, 
                 inputs_70__2, inputs_70__1, inputs_70__0, inputs_71__15, 
                 inputs_71__14, inputs_71__13, inputs_71__12, inputs_71__11, 
                 inputs_71__10, inputs_71__9, inputs_71__8, inputs_71__7, 
                 inputs_71__6, inputs_71__5, inputs_71__4, inputs_71__3, 
                 inputs_71__2, inputs_71__1, inputs_71__0, inputs_72__15, 
                 inputs_72__14, inputs_72__13, inputs_72__12, inputs_72__11, 
                 inputs_72__10, inputs_72__9, inputs_72__8, inputs_72__7, 
                 inputs_72__6, inputs_72__5, inputs_72__4, inputs_72__3, 
                 inputs_72__2, inputs_72__1, inputs_72__0, inputs_73__15, 
                 inputs_73__14, inputs_73__13, inputs_73__12, inputs_73__11, 
                 inputs_73__10, inputs_73__9, inputs_73__8, inputs_73__7, 
                 inputs_73__6, inputs_73__5, inputs_73__4, inputs_73__3, 
                 inputs_73__2, inputs_73__1, inputs_73__0, inputs_74__15, 
                 inputs_74__14, inputs_74__13, inputs_74__12, inputs_74__11, 
                 inputs_74__10, inputs_74__9, inputs_74__8, inputs_74__7, 
                 inputs_74__6, inputs_74__5, inputs_74__4, inputs_74__3, 
                 inputs_74__2, inputs_74__1, inputs_74__0, inputs_75__15, 
                 inputs_75__14, inputs_75__13, inputs_75__12, inputs_75__11, 
                 inputs_75__10, inputs_75__9, inputs_75__8, inputs_75__7, 
                 inputs_75__6, inputs_75__5, inputs_75__4, inputs_75__3, 
                 inputs_75__2, inputs_75__1, inputs_75__0, inputs_76__15, 
                 inputs_76__14, inputs_76__13, inputs_76__12, inputs_76__11, 
                 inputs_76__10, inputs_76__9, inputs_76__8, inputs_76__7, 
                 inputs_76__6, inputs_76__5, inputs_76__4, inputs_76__3, 
                 inputs_76__2, inputs_76__1, inputs_76__0, inputs_77__15, 
                 inputs_77__14, inputs_77__13, inputs_77__12, inputs_77__11, 
                 inputs_77__10, inputs_77__9, inputs_77__8, inputs_77__7, 
                 inputs_77__6, inputs_77__5, inputs_77__4, inputs_77__3, 
                 inputs_77__2, inputs_77__1, inputs_77__0, inputs_78__15, 
                 inputs_78__14, inputs_78__13, inputs_78__12, inputs_78__11, 
                 inputs_78__10, inputs_78__9, inputs_78__8, inputs_78__7, 
                 inputs_78__6, inputs_78__5, inputs_78__4, inputs_78__3, 
                 inputs_78__2, inputs_78__1, inputs_78__0, inputs_79__15, 
                 inputs_79__14, inputs_79__13, inputs_79__12, inputs_79__11, 
                 inputs_79__10, inputs_79__9, inputs_79__8, inputs_79__7, 
                 inputs_79__6, inputs_79__5, inputs_79__4, inputs_79__3, 
                 inputs_79__2, inputs_79__1, inputs_79__0, inputs_80__15, 
                 inputs_80__14, inputs_80__13, inputs_80__12, inputs_80__11, 
                 inputs_80__10, inputs_80__9, inputs_80__8, inputs_80__7, 
                 inputs_80__6, inputs_80__5, inputs_80__4, inputs_80__3, 
                 inputs_80__2, inputs_80__1, inputs_80__0, inputs_81__15, 
                 inputs_81__14, inputs_81__13, inputs_81__12, inputs_81__11, 
                 inputs_81__10, inputs_81__9, inputs_81__8, inputs_81__7, 
                 inputs_81__6, inputs_81__5, inputs_81__4, inputs_81__3, 
                 inputs_81__2, inputs_81__1, inputs_81__0, inputs_82__15, 
                 inputs_82__14, inputs_82__13, inputs_82__12, inputs_82__11, 
                 inputs_82__10, inputs_82__9, inputs_82__8, inputs_82__7, 
                 inputs_82__6, inputs_82__5, inputs_82__4, inputs_82__3, 
                 inputs_82__2, inputs_82__1, inputs_82__0, inputs_83__15, 
                 inputs_83__14, inputs_83__13, inputs_83__12, inputs_83__11, 
                 inputs_83__10, inputs_83__9, inputs_83__8, inputs_83__7, 
                 inputs_83__6, inputs_83__5, inputs_83__4, inputs_83__3, 
                 inputs_83__2, inputs_83__1, inputs_83__0, inputs_84__15, 
                 inputs_84__14, inputs_84__13, inputs_84__12, inputs_84__11, 
                 inputs_84__10, inputs_84__9, inputs_84__8, inputs_84__7, 
                 inputs_84__6, inputs_84__5, inputs_84__4, inputs_84__3, 
                 inputs_84__2, inputs_84__1, inputs_84__0, inputs_85__15, 
                 inputs_85__14, inputs_85__13, inputs_85__12, inputs_85__11, 
                 inputs_85__10, inputs_85__9, inputs_85__8, inputs_85__7, 
                 inputs_85__6, inputs_85__5, inputs_85__4, inputs_85__3, 
                 inputs_85__2, inputs_85__1, inputs_85__0, inputs_86__15, 
                 inputs_86__14, inputs_86__13, inputs_86__12, inputs_86__11, 
                 inputs_86__10, inputs_86__9, inputs_86__8, inputs_86__7, 
                 inputs_86__6, inputs_86__5, inputs_86__4, inputs_86__3, 
                 inputs_86__2, inputs_86__1, inputs_86__0, inputs_87__15, 
                 inputs_87__14, inputs_87__13, inputs_87__12, inputs_87__11, 
                 inputs_87__10, inputs_87__9, inputs_87__8, inputs_87__7, 
                 inputs_87__6, inputs_87__5, inputs_87__4, inputs_87__3, 
                 inputs_87__2, inputs_87__1, inputs_87__0, inputs_88__15, 
                 inputs_88__14, inputs_88__13, inputs_88__12, inputs_88__11, 
                 inputs_88__10, inputs_88__9, inputs_88__8, inputs_88__7, 
                 inputs_88__6, inputs_88__5, inputs_88__4, inputs_88__3, 
                 inputs_88__2, inputs_88__1, inputs_88__0, inputs_89__15, 
                 inputs_89__14, inputs_89__13, inputs_89__12, inputs_89__11, 
                 inputs_89__10, inputs_89__9, inputs_89__8, inputs_89__7, 
                 inputs_89__6, inputs_89__5, inputs_89__4, inputs_89__3, 
                 inputs_89__2, inputs_89__1, inputs_89__0, inputs_90__15, 
                 inputs_90__14, inputs_90__13, inputs_90__12, inputs_90__11, 
                 inputs_90__10, inputs_90__9, inputs_90__8, inputs_90__7, 
                 inputs_90__6, inputs_90__5, inputs_90__4, inputs_90__3, 
                 inputs_90__2, inputs_90__1, inputs_90__0, inputs_91__15, 
                 inputs_91__14, inputs_91__13, inputs_91__12, inputs_91__11, 
                 inputs_91__10, inputs_91__9, inputs_91__8, inputs_91__7, 
                 inputs_91__6, inputs_91__5, inputs_91__4, inputs_91__3, 
                 inputs_91__2, inputs_91__1, inputs_91__0, inputs_92__15, 
                 inputs_92__14, inputs_92__13, inputs_92__12, inputs_92__11, 
                 inputs_92__10, inputs_92__9, inputs_92__8, inputs_92__7, 
                 inputs_92__6, inputs_92__5, inputs_92__4, inputs_92__3, 
                 inputs_92__2, inputs_92__1, inputs_92__0, inputs_93__15, 
                 inputs_93__14, inputs_93__13, inputs_93__12, inputs_93__11, 
                 inputs_93__10, inputs_93__9, inputs_93__8, inputs_93__7, 
                 inputs_93__6, inputs_93__5, inputs_93__4, inputs_93__3, 
                 inputs_93__2, inputs_93__1, inputs_93__0, inputs_94__15, 
                 inputs_94__14, inputs_94__13, inputs_94__12, inputs_94__11, 
                 inputs_94__10, inputs_94__9, inputs_94__8, inputs_94__7, 
                 inputs_94__6, inputs_94__5, inputs_94__4, inputs_94__3, 
                 inputs_94__2, inputs_94__1, inputs_94__0, inputs_95__15, 
                 inputs_95__14, inputs_95__13, inputs_95__12, inputs_95__11, 
                 inputs_95__10, inputs_95__9, inputs_95__8, inputs_95__7, 
                 inputs_95__6, inputs_95__5, inputs_95__4, inputs_95__3, 
                 inputs_95__2, inputs_95__1, inputs_95__0, inputs_96__15, 
                 inputs_96__14, inputs_96__13, inputs_96__12, inputs_96__11, 
                 inputs_96__10, inputs_96__9, inputs_96__8, inputs_96__7, 
                 inputs_96__6, inputs_96__5, inputs_96__4, inputs_96__3, 
                 inputs_96__2, inputs_96__1, inputs_96__0, inputs_97__15, 
                 inputs_97__14, inputs_97__13, inputs_97__12, inputs_97__11, 
                 inputs_97__10, inputs_97__9, inputs_97__8, inputs_97__7, 
                 inputs_97__6, inputs_97__5, inputs_97__4, inputs_97__3, 
                 inputs_97__2, inputs_97__1, inputs_97__0, inputs_98__15, 
                 inputs_98__14, inputs_98__13, inputs_98__12, inputs_98__11, 
                 inputs_98__10, inputs_98__9, inputs_98__8, inputs_98__7, 
                 inputs_98__6, inputs_98__5, inputs_98__4, inputs_98__3, 
                 inputs_98__2, inputs_98__1, inputs_98__0, inputs_99__15, 
                 inputs_99__14, inputs_99__13, inputs_99__12, inputs_99__11, 
                 inputs_99__10, inputs_99__9, inputs_99__8, inputs_99__7, 
                 inputs_99__6, inputs_99__5, inputs_99__4, inputs_99__3, 
                 inputs_99__2, inputs_99__1, inputs_99__0, inputs_100__15, 
                 inputs_100__14, inputs_100__13, inputs_100__12, inputs_100__11, 
                 inputs_100__10, inputs_100__9, inputs_100__8, inputs_100__7, 
                 inputs_100__6, inputs_100__5, inputs_100__4, inputs_100__3, 
                 inputs_100__2, inputs_100__1, inputs_100__0, inputs_101__15, 
                 inputs_101__14, inputs_101__13, inputs_101__12, inputs_101__11, 
                 inputs_101__10, inputs_101__9, inputs_101__8, inputs_101__7, 
                 inputs_101__6, inputs_101__5, inputs_101__4, inputs_101__3, 
                 inputs_101__2, inputs_101__1, inputs_101__0, inputs_102__15, 
                 inputs_102__14, inputs_102__13, inputs_102__12, inputs_102__11, 
                 inputs_102__10, inputs_102__9, inputs_102__8, inputs_102__7, 
                 inputs_102__6, inputs_102__5, inputs_102__4, inputs_102__3, 
                 inputs_102__2, inputs_102__1, inputs_102__0, inputs_103__15, 
                 inputs_103__14, inputs_103__13, inputs_103__12, inputs_103__11, 
                 inputs_103__10, inputs_103__9, inputs_103__8, inputs_103__7, 
                 inputs_103__6, inputs_103__5, inputs_103__4, inputs_103__3, 
                 inputs_103__2, inputs_103__1, inputs_103__0, inputs_104__15, 
                 inputs_104__14, inputs_104__13, inputs_104__12, inputs_104__11, 
                 inputs_104__10, inputs_104__9, inputs_104__8, inputs_104__7, 
                 inputs_104__6, inputs_104__5, inputs_104__4, inputs_104__3, 
                 inputs_104__2, inputs_104__1, inputs_104__0, inputs_105__15, 
                 inputs_105__14, inputs_105__13, inputs_105__12, inputs_105__11, 
                 inputs_105__10, inputs_105__9, inputs_105__8, inputs_105__7, 
                 inputs_105__6, inputs_105__5, inputs_105__4, inputs_105__3, 
                 inputs_105__2, inputs_105__1, inputs_105__0, inputs_106__15, 
                 inputs_106__14, inputs_106__13, inputs_106__12, inputs_106__11, 
                 inputs_106__10, inputs_106__9, inputs_106__8, inputs_106__7, 
                 inputs_106__6, inputs_106__5, inputs_106__4, inputs_106__3, 
                 inputs_106__2, inputs_106__1, inputs_106__0, inputs_107__15, 
                 inputs_107__14, inputs_107__13, inputs_107__12, inputs_107__11, 
                 inputs_107__10, inputs_107__9, inputs_107__8, inputs_107__7, 
                 inputs_107__6, inputs_107__5, inputs_107__4, inputs_107__3, 
                 inputs_107__2, inputs_107__1, inputs_107__0, inputs_108__15, 
                 inputs_108__14, inputs_108__13, inputs_108__12, inputs_108__11, 
                 inputs_108__10, inputs_108__9, inputs_108__8, inputs_108__7, 
                 inputs_108__6, inputs_108__5, inputs_108__4, inputs_108__3, 
                 inputs_108__2, inputs_108__1, inputs_108__0, inputs_109__15, 
                 inputs_109__14, inputs_109__13, inputs_109__12, inputs_109__11, 
                 inputs_109__10, inputs_109__9, inputs_109__8, inputs_109__7, 
                 inputs_109__6, inputs_109__5, inputs_109__4, inputs_109__3, 
                 inputs_109__2, inputs_109__1, inputs_109__0, inputs_110__15, 
                 inputs_110__14, inputs_110__13, inputs_110__12, inputs_110__11, 
                 inputs_110__10, inputs_110__9, inputs_110__8, inputs_110__7, 
                 inputs_110__6, inputs_110__5, inputs_110__4, inputs_110__3, 
                 inputs_110__2, inputs_110__1, inputs_110__0, inputs_111__15, 
                 inputs_111__14, inputs_111__13, inputs_111__12, inputs_111__11, 
                 inputs_111__10, inputs_111__9, inputs_111__8, inputs_111__7, 
                 inputs_111__6, inputs_111__5, inputs_111__4, inputs_111__3, 
                 inputs_111__2, inputs_111__1, inputs_111__0, inputs_112__15, 
                 inputs_112__14, inputs_112__13, inputs_112__12, inputs_112__11, 
                 inputs_112__10, inputs_112__9, inputs_112__8, inputs_112__7, 
                 inputs_112__6, inputs_112__5, inputs_112__4, inputs_112__3, 
                 inputs_112__2, inputs_112__1, inputs_112__0, inputs_113__15, 
                 inputs_113__14, inputs_113__13, inputs_113__12, inputs_113__11, 
                 inputs_113__10, inputs_113__9, inputs_113__8, inputs_113__7, 
                 inputs_113__6, inputs_113__5, inputs_113__4, inputs_113__3, 
                 inputs_113__2, inputs_113__1, inputs_113__0, inputs_114__15, 
                 inputs_114__14, inputs_114__13, inputs_114__12, inputs_114__11, 
                 inputs_114__10, inputs_114__9, inputs_114__8, inputs_114__7, 
                 inputs_114__6, inputs_114__5, inputs_114__4, inputs_114__3, 
                 inputs_114__2, inputs_114__1, inputs_114__0, inputs_115__15, 
                 inputs_115__14, inputs_115__13, inputs_115__12, inputs_115__11, 
                 inputs_115__10, inputs_115__9, inputs_115__8, inputs_115__7, 
                 inputs_115__6, inputs_115__5, inputs_115__4, inputs_115__3, 
                 inputs_115__2, inputs_115__1, inputs_115__0, inputs_116__15, 
                 inputs_116__14, inputs_116__13, inputs_116__12, inputs_116__11, 
                 inputs_116__10, inputs_116__9, inputs_116__8, inputs_116__7, 
                 inputs_116__6, inputs_116__5, inputs_116__4, inputs_116__3, 
                 inputs_116__2, inputs_116__1, inputs_116__0, inputs_117__15, 
                 inputs_117__14, inputs_117__13, inputs_117__12, inputs_117__11, 
                 inputs_117__10, inputs_117__9, inputs_117__8, inputs_117__7, 
                 inputs_117__6, inputs_117__5, inputs_117__4, inputs_117__3, 
                 inputs_117__2, inputs_117__1, inputs_117__0, inputs_118__15, 
                 inputs_118__14, inputs_118__13, inputs_118__12, inputs_118__11, 
                 inputs_118__10, inputs_118__9, inputs_118__8, inputs_118__7, 
                 inputs_118__6, inputs_118__5, inputs_118__4, inputs_118__3, 
                 inputs_118__2, inputs_118__1, inputs_118__0, inputs_119__15, 
                 inputs_119__14, inputs_119__13, inputs_119__12, inputs_119__11, 
                 inputs_119__10, inputs_119__9, inputs_119__8, inputs_119__7, 
                 inputs_119__6, inputs_119__5, inputs_119__4, inputs_119__3, 
                 inputs_119__2, inputs_119__1, inputs_119__0, inputs_120__15, 
                 inputs_120__14, inputs_120__13, inputs_120__12, inputs_120__11, 
                 inputs_120__10, inputs_120__9, inputs_120__8, inputs_120__7, 
                 inputs_120__6, inputs_120__5, inputs_120__4, inputs_120__3, 
                 inputs_120__2, inputs_120__1, inputs_120__0, inputs_121__15, 
                 inputs_121__14, inputs_121__13, inputs_121__12, inputs_121__11, 
                 inputs_121__10, inputs_121__9, inputs_121__8, inputs_121__7, 
                 inputs_121__6, inputs_121__5, inputs_121__4, inputs_121__3, 
                 inputs_121__2, inputs_121__1, inputs_121__0, inputs_122__15, 
                 inputs_122__14, inputs_122__13, inputs_122__12, inputs_122__11, 
                 inputs_122__10, inputs_122__9, inputs_122__8, inputs_122__7, 
                 inputs_122__6, inputs_122__5, inputs_122__4, inputs_122__3, 
                 inputs_122__2, inputs_122__1, inputs_122__0, inputs_123__15, 
                 inputs_123__14, inputs_123__13, inputs_123__12, inputs_123__11, 
                 inputs_123__10, inputs_123__9, inputs_123__8, inputs_123__7, 
                 inputs_123__6, inputs_123__5, inputs_123__4, inputs_123__3, 
                 inputs_123__2, inputs_123__1, inputs_123__0, inputs_124__15, 
                 inputs_124__14, inputs_124__13, inputs_124__12, inputs_124__11, 
                 inputs_124__10, inputs_124__9, inputs_124__8, inputs_124__7, 
                 inputs_124__6, inputs_124__5, inputs_124__4, inputs_124__3, 
                 inputs_124__2, inputs_124__1, inputs_124__0, inputs_125__15, 
                 inputs_125__14, inputs_125__13, inputs_125__12, inputs_125__11, 
                 inputs_125__10, inputs_125__9, inputs_125__8, inputs_125__7, 
                 inputs_125__6, inputs_125__5, inputs_125__4, inputs_125__3, 
                 inputs_125__2, inputs_125__1, inputs_125__0, inputs_126__15, 
                 inputs_126__14, inputs_126__13, inputs_126__12, inputs_126__11, 
                 inputs_126__10, inputs_126__9, inputs_126__8, inputs_126__7, 
                 inputs_126__6, inputs_126__5, inputs_126__4, inputs_126__3, 
                 inputs_126__2, inputs_126__1, inputs_126__0, inputs_127__15, 
                 inputs_127__14, inputs_127__13, inputs_127__12, inputs_127__11, 
                 inputs_127__10, inputs_127__9, inputs_127__8, inputs_127__7, 
                 inputs_127__6, inputs_127__5, inputs_127__4, inputs_127__3, 
                 inputs_127__2, inputs_127__1, inputs_127__0, inputs_128__15, 
                 inputs_128__14, inputs_128__13, inputs_128__12, inputs_128__11, 
                 inputs_128__10, inputs_128__9, inputs_128__8, inputs_128__7, 
                 inputs_128__6, inputs_128__5, inputs_128__4, inputs_128__3, 
                 inputs_128__2, inputs_128__1, inputs_128__0, inputs_129__15, 
                 inputs_129__14, inputs_129__13, inputs_129__12, inputs_129__11, 
                 inputs_129__10, inputs_129__9, inputs_129__8, inputs_129__7, 
                 inputs_129__6, inputs_129__5, inputs_129__4, inputs_129__3, 
                 inputs_129__2, inputs_129__1, inputs_129__0, inputs_130__15, 
                 inputs_130__14, inputs_130__13, inputs_130__12, inputs_130__11, 
                 inputs_130__10, inputs_130__9, inputs_130__8, inputs_130__7, 
                 inputs_130__6, inputs_130__5, inputs_130__4, inputs_130__3, 
                 inputs_130__2, inputs_130__1, inputs_130__0, inputs_131__15, 
                 inputs_131__14, inputs_131__13, inputs_131__12, inputs_131__11, 
                 inputs_131__10, inputs_131__9, inputs_131__8, inputs_131__7, 
                 inputs_131__6, inputs_131__5, inputs_131__4, inputs_131__3, 
                 inputs_131__2, inputs_131__1, inputs_131__0, inputs_132__15, 
                 inputs_132__14, inputs_132__13, inputs_132__12, inputs_132__11, 
                 inputs_132__10, inputs_132__9, inputs_132__8, inputs_132__7, 
                 inputs_132__6, inputs_132__5, inputs_132__4, inputs_132__3, 
                 inputs_132__2, inputs_132__1, inputs_132__0, inputs_133__15, 
                 inputs_133__14, inputs_133__13, inputs_133__12, inputs_133__11, 
                 inputs_133__10, inputs_133__9, inputs_133__8, inputs_133__7, 
                 inputs_133__6, inputs_133__5, inputs_133__4, inputs_133__3, 
                 inputs_133__2, inputs_133__1, inputs_133__0, inputs_134__15, 
                 inputs_134__14, inputs_134__13, inputs_134__12, inputs_134__11, 
                 inputs_134__10, inputs_134__9, inputs_134__8, inputs_134__7, 
                 inputs_134__6, inputs_134__5, inputs_134__4, inputs_134__3, 
                 inputs_134__2, inputs_134__1, inputs_134__0, inputs_135__15, 
                 inputs_135__14, inputs_135__13, inputs_135__12, inputs_135__11, 
                 inputs_135__10, inputs_135__9, inputs_135__8, inputs_135__7, 
                 inputs_135__6, inputs_135__5, inputs_135__4, inputs_135__3, 
                 inputs_135__2, inputs_135__1, inputs_135__0, inputs_136__15, 
                 inputs_136__14, inputs_136__13, inputs_136__12, inputs_136__11, 
                 inputs_136__10, inputs_136__9, inputs_136__8, inputs_136__7, 
                 inputs_136__6, inputs_136__5, inputs_136__4, inputs_136__3, 
                 inputs_136__2, inputs_136__1, inputs_136__0, inputs_137__15, 
                 inputs_137__14, inputs_137__13, inputs_137__12, inputs_137__11, 
                 inputs_137__10, inputs_137__9, inputs_137__8, inputs_137__7, 
                 inputs_137__6, inputs_137__5, inputs_137__4, inputs_137__3, 
                 inputs_137__2, inputs_137__1, inputs_137__0, inputs_138__15, 
                 inputs_138__14, inputs_138__13, inputs_138__12, inputs_138__11, 
                 inputs_138__10, inputs_138__9, inputs_138__8, inputs_138__7, 
                 inputs_138__6, inputs_138__5, inputs_138__4, inputs_138__3, 
                 inputs_138__2, inputs_138__1, inputs_138__0, inputs_139__15, 
                 inputs_139__14, inputs_139__13, inputs_139__12, inputs_139__11, 
                 inputs_139__10, inputs_139__9, inputs_139__8, inputs_139__7, 
                 inputs_139__6, inputs_139__5, inputs_139__4, inputs_139__3, 
                 inputs_139__2, inputs_139__1, inputs_139__0, inputs_140__15, 
                 inputs_140__14, inputs_140__13, inputs_140__12, inputs_140__11, 
                 inputs_140__10, inputs_140__9, inputs_140__8, inputs_140__7, 
                 inputs_140__6, inputs_140__5, inputs_140__4, inputs_140__3, 
                 inputs_140__2, inputs_140__1, inputs_140__0, inputs_141__15, 
                 inputs_141__14, inputs_141__13, inputs_141__12, inputs_141__11, 
                 inputs_141__10, inputs_141__9, inputs_141__8, inputs_141__7, 
                 inputs_141__6, inputs_141__5, inputs_141__4, inputs_141__3, 
                 inputs_141__2, inputs_141__1, inputs_141__0, inputs_142__15, 
                 inputs_142__14, inputs_142__13, inputs_142__12, inputs_142__11, 
                 inputs_142__10, inputs_142__9, inputs_142__8, inputs_142__7, 
                 inputs_142__6, inputs_142__5, inputs_142__4, inputs_142__3, 
                 inputs_142__2, inputs_142__1, inputs_142__0, inputs_143__15, 
                 inputs_143__14, inputs_143__13, inputs_143__12, inputs_143__11, 
                 inputs_143__10, inputs_143__9, inputs_143__8, inputs_143__7, 
                 inputs_143__6, inputs_143__5, inputs_143__4, inputs_143__3, 
                 inputs_143__2, inputs_143__1, inputs_143__0, inputs_144__15, 
                 inputs_144__14, inputs_144__13, inputs_144__12, inputs_144__11, 
                 inputs_144__10, inputs_144__9, inputs_144__8, inputs_144__7, 
                 inputs_144__6, inputs_144__5, inputs_144__4, inputs_144__3, 
                 inputs_144__2, inputs_144__1, inputs_144__0, inputs_145__15, 
                 inputs_145__14, inputs_145__13, inputs_145__12, inputs_145__11, 
                 inputs_145__10, inputs_145__9, inputs_145__8, inputs_145__7, 
                 inputs_145__6, inputs_145__5, inputs_145__4, inputs_145__3, 
                 inputs_145__2, inputs_145__1, inputs_145__0, inputs_146__15, 
                 inputs_146__14, inputs_146__13, inputs_146__12, inputs_146__11, 
                 inputs_146__10, inputs_146__9, inputs_146__8, inputs_146__7, 
                 inputs_146__6, inputs_146__5, inputs_146__4, inputs_146__3, 
                 inputs_146__2, inputs_146__1, inputs_146__0, inputs_147__15, 
                 inputs_147__14, inputs_147__13, inputs_147__12, inputs_147__11, 
                 inputs_147__10, inputs_147__9, inputs_147__8, inputs_147__7, 
                 inputs_147__6, inputs_147__5, inputs_147__4, inputs_147__3, 
                 inputs_147__2, inputs_147__1, inputs_147__0, inputs_148__15, 
                 inputs_148__14, inputs_148__13, inputs_148__12, inputs_148__11, 
                 inputs_148__10, inputs_148__9, inputs_148__8, inputs_148__7, 
                 inputs_148__6, inputs_148__5, inputs_148__4, inputs_148__3, 
                 inputs_148__2, inputs_148__1, inputs_148__0, inputs_149__15, 
                 inputs_149__14, inputs_149__13, inputs_149__12, inputs_149__11, 
                 inputs_149__10, inputs_149__9, inputs_149__8, inputs_149__7, 
                 inputs_149__6, inputs_149__5, inputs_149__4, inputs_149__3, 
                 inputs_149__2, inputs_149__1, inputs_149__0, inputs_150__15, 
                 inputs_150__14, inputs_150__13, inputs_150__12, inputs_150__11, 
                 inputs_150__10, inputs_150__9, inputs_150__8, inputs_150__7, 
                 inputs_150__6, inputs_150__5, inputs_150__4, inputs_150__3, 
                 inputs_150__2, inputs_150__1, inputs_150__0, inputs_151__15, 
                 inputs_151__14, inputs_151__13, inputs_151__12, inputs_151__11, 
                 inputs_151__10, inputs_151__9, inputs_151__8, inputs_151__7, 
                 inputs_151__6, inputs_151__5, inputs_151__4, inputs_151__3, 
                 inputs_151__2, inputs_151__1, inputs_151__0, inputs_152__15, 
                 inputs_152__14, inputs_152__13, inputs_152__12, inputs_152__11, 
                 inputs_152__10, inputs_152__9, inputs_152__8, inputs_152__7, 
                 inputs_152__6, inputs_152__5, inputs_152__4, inputs_152__3, 
                 inputs_152__2, inputs_152__1, inputs_152__0, inputs_153__15, 
                 inputs_153__14, inputs_153__13, inputs_153__12, inputs_153__11, 
                 inputs_153__10, inputs_153__9, inputs_153__8, inputs_153__7, 
                 inputs_153__6, inputs_153__5, inputs_153__4, inputs_153__3, 
                 inputs_153__2, inputs_153__1, inputs_153__0, inputs_154__15, 
                 inputs_154__14, inputs_154__13, inputs_154__12, inputs_154__11, 
                 inputs_154__10, inputs_154__9, inputs_154__8, inputs_154__7, 
                 inputs_154__6, inputs_154__5, inputs_154__4, inputs_154__3, 
                 inputs_154__2, inputs_154__1, inputs_154__0, inputs_155__15, 
                 inputs_155__14, inputs_155__13, inputs_155__12, inputs_155__11, 
                 inputs_155__10, inputs_155__9, inputs_155__8, inputs_155__7, 
                 inputs_155__6, inputs_155__5, inputs_155__4, inputs_155__3, 
                 inputs_155__2, inputs_155__1, inputs_155__0, inputs_156__15, 
                 inputs_156__14, inputs_156__13, inputs_156__12, inputs_156__11, 
                 inputs_156__10, inputs_156__9, inputs_156__8, inputs_156__7, 
                 inputs_156__6, inputs_156__5, inputs_156__4, inputs_156__3, 
                 inputs_156__2, inputs_156__1, inputs_156__0, inputs_157__15, 
                 inputs_157__14, inputs_157__13, inputs_157__12, inputs_157__11, 
                 inputs_157__10, inputs_157__9, inputs_157__8, inputs_157__7, 
                 inputs_157__6, inputs_157__5, inputs_157__4, inputs_157__3, 
                 inputs_157__2, inputs_157__1, inputs_157__0, inputs_158__15, 
                 inputs_158__14, inputs_158__13, inputs_158__12, inputs_158__11, 
                 inputs_158__10, inputs_158__9, inputs_158__8, inputs_158__7, 
                 inputs_158__6, inputs_158__5, inputs_158__4, inputs_158__3, 
                 inputs_158__2, inputs_158__1, inputs_158__0, inputs_159__15, 
                 inputs_159__14, inputs_159__13, inputs_159__12, inputs_159__11, 
                 inputs_159__10, inputs_159__9, inputs_159__8, inputs_159__7, 
                 inputs_159__6, inputs_159__5, inputs_159__4, inputs_159__3, 
                 inputs_159__2, inputs_159__1, inputs_159__0, inputs_160__15, 
                 inputs_160__14, inputs_160__13, inputs_160__12, inputs_160__11, 
                 inputs_160__10, inputs_160__9, inputs_160__8, inputs_160__7, 
                 inputs_160__6, inputs_160__5, inputs_160__4, inputs_160__3, 
                 inputs_160__2, inputs_160__1, inputs_160__0, inputs_161__15, 
                 inputs_161__14, inputs_161__13, inputs_161__12, inputs_161__11, 
                 inputs_161__10, inputs_161__9, inputs_161__8, inputs_161__7, 
                 inputs_161__6, inputs_161__5, inputs_161__4, inputs_161__3, 
                 inputs_161__2, inputs_161__1, inputs_161__0, inputs_162__15, 
                 inputs_162__14, inputs_162__13, inputs_162__12, inputs_162__11, 
                 inputs_162__10, inputs_162__9, inputs_162__8, inputs_162__7, 
                 inputs_162__6, inputs_162__5, inputs_162__4, inputs_162__3, 
                 inputs_162__2, inputs_162__1, inputs_162__0, inputs_163__15, 
                 inputs_163__14, inputs_163__13, inputs_163__12, inputs_163__11, 
                 inputs_163__10, inputs_163__9, inputs_163__8, inputs_163__7, 
                 inputs_163__6, inputs_163__5, inputs_163__4, inputs_163__3, 
                 inputs_163__2, inputs_163__1, inputs_163__0, inputs_164__15, 
                 inputs_164__14, inputs_164__13, inputs_164__12, inputs_164__11, 
                 inputs_164__10, inputs_164__9, inputs_164__8, inputs_164__7, 
                 inputs_164__6, inputs_164__5, inputs_164__4, inputs_164__3, 
                 inputs_164__2, inputs_164__1, inputs_164__0, inputs_165__15, 
                 inputs_165__14, inputs_165__13, inputs_165__12, inputs_165__11, 
                 inputs_165__10, inputs_165__9, inputs_165__8, inputs_165__7, 
                 inputs_165__6, inputs_165__5, inputs_165__4, inputs_165__3, 
                 inputs_165__2, inputs_165__1, inputs_165__0, inputs_166__15, 
                 inputs_166__14, inputs_166__13, inputs_166__12, inputs_166__11, 
                 inputs_166__10, inputs_166__9, inputs_166__8, inputs_166__7, 
                 inputs_166__6, inputs_166__5, inputs_166__4, inputs_166__3, 
                 inputs_166__2, inputs_166__1, inputs_166__0, inputs_167__15, 
                 inputs_167__14, inputs_167__13, inputs_167__12, inputs_167__11, 
                 inputs_167__10, inputs_167__9, inputs_167__8, inputs_167__7, 
                 inputs_167__6, inputs_167__5, inputs_167__4, inputs_167__3, 
                 inputs_167__2, inputs_167__1, inputs_167__0, inputs_168__15, 
                 inputs_168__14, inputs_168__13, inputs_168__12, inputs_168__11, 
                 inputs_168__10, inputs_168__9, inputs_168__8, inputs_168__7, 
                 inputs_168__6, inputs_168__5, inputs_168__4, inputs_168__3, 
                 inputs_168__2, inputs_168__1, inputs_168__0, inputs_169__15, 
                 inputs_169__14, inputs_169__13, inputs_169__12, inputs_169__11, 
                 inputs_169__10, inputs_169__9, inputs_169__8, inputs_169__7, 
                 inputs_169__6, inputs_169__5, inputs_169__4, inputs_169__3, 
                 inputs_169__2, inputs_169__1, inputs_169__0, inputs_170__15, 
                 inputs_170__14, inputs_170__13, inputs_170__12, inputs_170__11, 
                 inputs_170__10, inputs_170__9, inputs_170__8, inputs_170__7, 
                 inputs_170__6, inputs_170__5, inputs_170__4, inputs_170__3, 
                 inputs_170__2, inputs_170__1, inputs_170__0, inputs_171__15, 
                 inputs_171__14, inputs_171__13, inputs_171__12, inputs_171__11, 
                 inputs_171__10, inputs_171__9, inputs_171__8, inputs_171__7, 
                 inputs_171__6, inputs_171__5, inputs_171__4, inputs_171__3, 
                 inputs_171__2, inputs_171__1, inputs_171__0, inputs_172__15, 
                 inputs_172__14, inputs_172__13, inputs_172__12, inputs_172__11, 
                 inputs_172__10, inputs_172__9, inputs_172__8, inputs_172__7, 
                 inputs_172__6, inputs_172__5, inputs_172__4, inputs_172__3, 
                 inputs_172__2, inputs_172__1, inputs_172__0, inputs_173__15, 
                 inputs_173__14, inputs_173__13, inputs_173__12, inputs_173__11, 
                 inputs_173__10, inputs_173__9, inputs_173__8, inputs_173__7, 
                 inputs_173__6, inputs_173__5, inputs_173__4, inputs_173__3, 
                 inputs_173__2, inputs_173__1, inputs_173__0, inputs_174__15, 
                 inputs_174__14, inputs_174__13, inputs_174__12, inputs_174__11, 
                 inputs_174__10, inputs_174__9, inputs_174__8, inputs_174__7, 
                 inputs_174__6, inputs_174__5, inputs_174__4, inputs_174__3, 
                 inputs_174__2, inputs_174__1, inputs_174__0, inputs_175__15, 
                 inputs_175__14, inputs_175__13, inputs_175__12, inputs_175__11, 
                 inputs_175__10, inputs_175__9, inputs_175__8, inputs_175__7, 
                 inputs_175__6, inputs_175__5, inputs_175__4, inputs_175__3, 
                 inputs_175__2, inputs_175__1, inputs_175__0, inputs_176__15, 
                 inputs_176__14, inputs_176__13, inputs_176__12, inputs_176__11, 
                 inputs_176__10, inputs_176__9, inputs_176__8, inputs_176__7, 
                 inputs_176__6, inputs_176__5, inputs_176__4, inputs_176__3, 
                 inputs_176__2, inputs_176__1, inputs_176__0, inputs_177__15, 
                 inputs_177__14, inputs_177__13, inputs_177__12, inputs_177__11, 
                 inputs_177__10, inputs_177__9, inputs_177__8, inputs_177__7, 
                 inputs_177__6, inputs_177__5, inputs_177__4, inputs_177__3, 
                 inputs_177__2, inputs_177__1, inputs_177__0, inputs_178__15, 
                 inputs_178__14, inputs_178__13, inputs_178__12, inputs_178__11, 
                 inputs_178__10, inputs_178__9, inputs_178__8, inputs_178__7, 
                 inputs_178__6, inputs_178__5, inputs_178__4, inputs_178__3, 
                 inputs_178__2, inputs_178__1, inputs_178__0, inputs_179__15, 
                 inputs_179__14, inputs_179__13, inputs_179__12, inputs_179__11, 
                 inputs_179__10, inputs_179__9, inputs_179__8, inputs_179__7, 
                 inputs_179__6, inputs_179__5, inputs_179__4, inputs_179__3, 
                 inputs_179__2, inputs_179__1, inputs_179__0, inputs_180__15, 
                 inputs_180__14, inputs_180__13, inputs_180__12, inputs_180__11, 
                 inputs_180__10, inputs_180__9, inputs_180__8, inputs_180__7, 
                 inputs_180__6, inputs_180__5, inputs_180__4, inputs_180__3, 
                 inputs_180__2, inputs_180__1, inputs_180__0, inputs_181__15, 
                 inputs_181__14, inputs_181__13, inputs_181__12, inputs_181__11, 
                 inputs_181__10, inputs_181__9, inputs_181__8, inputs_181__7, 
                 inputs_181__6, inputs_181__5, inputs_181__4, inputs_181__3, 
                 inputs_181__2, inputs_181__1, inputs_181__0, inputs_182__15, 
                 inputs_182__14, inputs_182__13, inputs_182__12, inputs_182__11, 
                 inputs_182__10, inputs_182__9, inputs_182__8, inputs_182__7, 
                 inputs_182__6, inputs_182__5, inputs_182__4, inputs_182__3, 
                 inputs_182__2, inputs_182__1, inputs_182__0, inputs_183__15, 
                 inputs_183__14, inputs_183__13, inputs_183__12, inputs_183__11, 
                 inputs_183__10, inputs_183__9, inputs_183__8, inputs_183__7, 
                 inputs_183__6, inputs_183__5, inputs_183__4, inputs_183__3, 
                 inputs_183__2, inputs_183__1, inputs_183__0, inputs_184__15, 
                 inputs_184__14, inputs_184__13, inputs_184__12, inputs_184__11, 
                 inputs_184__10, inputs_184__9, inputs_184__8, inputs_184__7, 
                 inputs_184__6, inputs_184__5, inputs_184__4, inputs_184__3, 
                 inputs_184__2, inputs_184__1, inputs_184__0, inputs_185__15, 
                 inputs_185__14, inputs_185__13, inputs_185__12, inputs_185__11, 
                 inputs_185__10, inputs_185__9, inputs_185__8, inputs_185__7, 
                 inputs_185__6, inputs_185__5, inputs_185__4, inputs_185__3, 
                 inputs_185__2, inputs_185__1, inputs_185__0, inputs_186__15, 
                 inputs_186__14, inputs_186__13, inputs_186__12, inputs_186__11, 
                 inputs_186__10, inputs_186__9, inputs_186__8, inputs_186__7, 
                 inputs_186__6, inputs_186__5, inputs_186__4, inputs_186__3, 
                 inputs_186__2, inputs_186__1, inputs_186__0, inputs_187__15, 
                 inputs_187__14, inputs_187__13, inputs_187__12, inputs_187__11, 
                 inputs_187__10, inputs_187__9, inputs_187__8, inputs_187__7, 
                 inputs_187__6, inputs_187__5, inputs_187__4, inputs_187__3, 
                 inputs_187__2, inputs_187__1, inputs_187__0, inputs_188__15, 
                 inputs_188__14, inputs_188__13, inputs_188__12, inputs_188__11, 
                 inputs_188__10, inputs_188__9, inputs_188__8, inputs_188__7, 
                 inputs_188__6, inputs_188__5, inputs_188__4, inputs_188__3, 
                 inputs_188__2, inputs_188__1, inputs_188__0, inputs_189__15, 
                 inputs_189__14, inputs_189__13, inputs_189__12, inputs_189__11, 
                 inputs_189__10, inputs_189__9, inputs_189__8, inputs_189__7, 
                 inputs_189__6, inputs_189__5, inputs_189__4, inputs_189__3, 
                 inputs_189__2, inputs_189__1, inputs_189__0, inputs_190__15, 
                 inputs_190__14, inputs_190__13, inputs_190__12, inputs_190__11, 
                 inputs_190__10, inputs_190__9, inputs_190__8, inputs_190__7, 
                 inputs_190__6, inputs_190__5, inputs_190__4, inputs_190__3, 
                 inputs_190__2, inputs_190__1, inputs_190__0, inputs_191__15, 
                 inputs_191__14, inputs_191__13, inputs_191__12, inputs_191__11, 
                 inputs_191__10, inputs_191__9, inputs_191__8, inputs_191__7, 
                 inputs_191__6, inputs_191__5, inputs_191__4, inputs_191__3, 
                 inputs_191__2, inputs_191__1, inputs_191__0, inputs_192__15, 
                 inputs_192__14, inputs_192__13, inputs_192__12, inputs_192__11, 
                 inputs_192__10, inputs_192__9, inputs_192__8, inputs_192__7, 
                 inputs_192__6, inputs_192__5, inputs_192__4, inputs_192__3, 
                 inputs_192__2, inputs_192__1, inputs_192__0, inputs_193__15, 
                 inputs_193__14, inputs_193__13, inputs_193__12, inputs_193__11, 
                 inputs_193__10, inputs_193__9, inputs_193__8, inputs_193__7, 
                 inputs_193__6, inputs_193__5, inputs_193__4, inputs_193__3, 
                 inputs_193__2, inputs_193__1, inputs_193__0, inputs_194__15, 
                 inputs_194__14, inputs_194__13, inputs_194__12, inputs_194__11, 
                 inputs_194__10, inputs_194__9, inputs_194__8, inputs_194__7, 
                 inputs_194__6, inputs_194__5, inputs_194__4, inputs_194__3, 
                 inputs_194__2, inputs_194__1, inputs_194__0, inputs_195__15, 
                 inputs_195__14, inputs_195__13, inputs_195__12, inputs_195__11, 
                 inputs_195__10, inputs_195__9, inputs_195__8, inputs_195__7, 
                 inputs_195__6, inputs_195__5, inputs_195__4, inputs_195__3, 
                 inputs_195__2, inputs_195__1, inputs_195__0, inputs_196__15, 
                 inputs_196__14, inputs_196__13, inputs_196__12, inputs_196__11, 
                 inputs_196__10, inputs_196__9, inputs_196__8, inputs_196__7, 
                 inputs_196__6, inputs_196__5, inputs_196__4, inputs_196__3, 
                 inputs_196__2, inputs_196__1, inputs_196__0, inputs_197__15, 
                 inputs_197__14, inputs_197__13, inputs_197__12, inputs_197__11, 
                 inputs_197__10, inputs_197__9, inputs_197__8, inputs_197__7, 
                 inputs_197__6, inputs_197__5, inputs_197__4, inputs_197__3, 
                 inputs_197__2, inputs_197__1, inputs_197__0, inputs_198__15, 
                 inputs_198__14, inputs_198__13, inputs_198__12, inputs_198__11, 
                 inputs_198__10, inputs_198__9, inputs_198__8, inputs_198__7, 
                 inputs_198__6, inputs_198__5, inputs_198__4, inputs_198__3, 
                 inputs_198__2, inputs_198__1, inputs_198__0, inputs_199__15, 
                 inputs_199__14, inputs_199__13, inputs_199__12, inputs_199__11, 
                 inputs_199__10, inputs_199__9, inputs_199__8, inputs_199__7, 
                 inputs_199__6, inputs_199__5, inputs_199__4, inputs_199__3, 
                 inputs_199__2, inputs_199__1, inputs_199__0, inputs_200__15, 
                 inputs_200__14, inputs_200__13, inputs_200__12, inputs_200__11, 
                 inputs_200__10, inputs_200__9, inputs_200__8, inputs_200__7, 
                 inputs_200__6, inputs_200__5, inputs_200__4, inputs_200__3, 
                 inputs_200__2, inputs_200__1, inputs_200__0, inputs_201__15, 
                 inputs_201__14, inputs_201__13, inputs_201__12, inputs_201__11, 
                 inputs_201__10, inputs_201__9, inputs_201__8, inputs_201__7, 
                 inputs_201__6, inputs_201__5, inputs_201__4, inputs_201__3, 
                 inputs_201__2, inputs_201__1, inputs_201__0, inputs_202__15, 
                 inputs_202__14, inputs_202__13, inputs_202__12, inputs_202__11, 
                 inputs_202__10, inputs_202__9, inputs_202__8, inputs_202__7, 
                 inputs_202__6, inputs_202__5, inputs_202__4, inputs_202__3, 
                 inputs_202__2, inputs_202__1, inputs_202__0, inputs_203__15, 
                 inputs_203__14, inputs_203__13, inputs_203__12, inputs_203__11, 
                 inputs_203__10, inputs_203__9, inputs_203__8, inputs_203__7, 
                 inputs_203__6, inputs_203__5, inputs_203__4, inputs_203__3, 
                 inputs_203__2, inputs_203__1, inputs_203__0, inputs_204__15, 
                 inputs_204__14, inputs_204__13, inputs_204__12, inputs_204__11, 
                 inputs_204__10, inputs_204__9, inputs_204__8, inputs_204__7, 
                 inputs_204__6, inputs_204__5, inputs_204__4, inputs_204__3, 
                 inputs_204__2, inputs_204__1, inputs_204__0, inputs_205__15, 
                 inputs_205__14, inputs_205__13, inputs_205__12, inputs_205__11, 
                 inputs_205__10, inputs_205__9, inputs_205__8, inputs_205__7, 
                 inputs_205__6, inputs_205__5, inputs_205__4, inputs_205__3, 
                 inputs_205__2, inputs_205__1, inputs_205__0, inputs_206__15, 
                 inputs_206__14, inputs_206__13, inputs_206__12, inputs_206__11, 
                 inputs_206__10, inputs_206__9, inputs_206__8, inputs_206__7, 
                 inputs_206__6, inputs_206__5, inputs_206__4, inputs_206__3, 
                 inputs_206__2, inputs_206__1, inputs_206__0, inputs_207__15, 
                 inputs_207__14, inputs_207__13, inputs_207__12, inputs_207__11, 
                 inputs_207__10, inputs_207__9, inputs_207__8, inputs_207__7, 
                 inputs_207__6, inputs_207__5, inputs_207__4, inputs_207__3, 
                 inputs_207__2, inputs_207__1, inputs_207__0, inputs_208__15, 
                 inputs_208__14, inputs_208__13, inputs_208__12, inputs_208__11, 
                 inputs_208__10, inputs_208__9, inputs_208__8, inputs_208__7, 
                 inputs_208__6, inputs_208__5, inputs_208__4, inputs_208__3, 
                 inputs_208__2, inputs_208__1, inputs_208__0, inputs_209__15, 
                 inputs_209__14, inputs_209__13, inputs_209__12, inputs_209__11, 
                 inputs_209__10, inputs_209__9, inputs_209__8, inputs_209__7, 
                 inputs_209__6, inputs_209__5, inputs_209__4, inputs_209__3, 
                 inputs_209__2, inputs_209__1, inputs_209__0, inputs_210__15, 
                 inputs_210__14, inputs_210__13, inputs_210__12, inputs_210__11, 
                 inputs_210__10, inputs_210__9, inputs_210__8, inputs_210__7, 
                 inputs_210__6, inputs_210__5, inputs_210__4, inputs_210__3, 
                 inputs_210__2, inputs_210__1, inputs_210__0, inputs_211__15, 
                 inputs_211__14, inputs_211__13, inputs_211__12, inputs_211__11, 
                 inputs_211__10, inputs_211__9, inputs_211__8, inputs_211__7, 
                 inputs_211__6, inputs_211__5, inputs_211__4, inputs_211__3, 
                 inputs_211__2, inputs_211__1, inputs_211__0, inputs_212__15, 
                 inputs_212__14, inputs_212__13, inputs_212__12, inputs_212__11, 
                 inputs_212__10, inputs_212__9, inputs_212__8, inputs_212__7, 
                 inputs_212__6, inputs_212__5, inputs_212__4, inputs_212__3, 
                 inputs_212__2, inputs_212__1, inputs_212__0, inputs_213__15, 
                 inputs_213__14, inputs_213__13, inputs_213__12, inputs_213__11, 
                 inputs_213__10, inputs_213__9, inputs_213__8, inputs_213__7, 
                 inputs_213__6, inputs_213__5, inputs_213__4, inputs_213__3, 
                 inputs_213__2, inputs_213__1, inputs_213__0, inputs_214__15, 
                 inputs_214__14, inputs_214__13, inputs_214__12, inputs_214__11, 
                 inputs_214__10, inputs_214__9, inputs_214__8, inputs_214__7, 
                 inputs_214__6, inputs_214__5, inputs_214__4, inputs_214__3, 
                 inputs_214__2, inputs_214__1, inputs_214__0, inputs_215__15, 
                 inputs_215__14, inputs_215__13, inputs_215__12, inputs_215__11, 
                 inputs_215__10, inputs_215__9, inputs_215__8, inputs_215__7, 
                 inputs_215__6, inputs_215__5, inputs_215__4, inputs_215__3, 
                 inputs_215__2, inputs_215__1, inputs_215__0, inputs_216__15, 
                 inputs_216__14, inputs_216__13, inputs_216__12, inputs_216__11, 
                 inputs_216__10, inputs_216__9, inputs_216__8, inputs_216__7, 
                 inputs_216__6, inputs_216__5, inputs_216__4, inputs_216__3, 
                 inputs_216__2, inputs_216__1, inputs_216__0, inputs_217__15, 
                 inputs_217__14, inputs_217__13, inputs_217__12, inputs_217__11, 
                 inputs_217__10, inputs_217__9, inputs_217__8, inputs_217__7, 
                 inputs_217__6, inputs_217__5, inputs_217__4, inputs_217__3, 
                 inputs_217__2, inputs_217__1, inputs_217__0, inputs_218__15, 
                 inputs_218__14, inputs_218__13, inputs_218__12, inputs_218__11, 
                 inputs_218__10, inputs_218__9, inputs_218__8, inputs_218__7, 
                 inputs_218__6, inputs_218__5, inputs_218__4, inputs_218__3, 
                 inputs_218__2, inputs_218__1, inputs_218__0, inputs_219__15, 
                 inputs_219__14, inputs_219__13, inputs_219__12, inputs_219__11, 
                 inputs_219__10, inputs_219__9, inputs_219__8, inputs_219__7, 
                 inputs_219__6, inputs_219__5, inputs_219__4, inputs_219__3, 
                 inputs_219__2, inputs_219__1, inputs_219__0, inputs_220__15, 
                 inputs_220__14, inputs_220__13, inputs_220__12, inputs_220__11, 
                 inputs_220__10, inputs_220__9, inputs_220__8, inputs_220__7, 
                 inputs_220__6, inputs_220__5, inputs_220__4, inputs_220__3, 
                 inputs_220__2, inputs_220__1, inputs_220__0, inputs_221__15, 
                 inputs_221__14, inputs_221__13, inputs_221__12, inputs_221__11, 
                 inputs_221__10, inputs_221__9, inputs_221__8, inputs_221__7, 
                 inputs_221__6, inputs_221__5, inputs_221__4, inputs_221__3, 
                 inputs_221__2, inputs_221__1, inputs_221__0, inputs_222__15, 
                 inputs_222__14, inputs_222__13, inputs_222__12, inputs_222__11, 
                 inputs_222__10, inputs_222__9, inputs_222__8, inputs_222__7, 
                 inputs_222__6, inputs_222__5, inputs_222__4, inputs_222__3, 
                 inputs_222__2, inputs_222__1, inputs_222__0, inputs_223__15, 
                 inputs_223__14, inputs_223__13, inputs_223__12, inputs_223__11, 
                 inputs_223__10, inputs_223__9, inputs_223__8, inputs_223__7, 
                 inputs_223__6, inputs_223__5, inputs_223__4, inputs_223__3, 
                 inputs_223__2, inputs_223__1, inputs_223__0, inputs_224__15, 
                 inputs_224__14, inputs_224__13, inputs_224__12, inputs_224__11, 
                 inputs_224__10, inputs_224__9, inputs_224__8, inputs_224__7, 
                 inputs_224__6, inputs_224__5, inputs_224__4, inputs_224__3, 
                 inputs_224__2, inputs_224__1, inputs_224__0, inputs_225__15, 
                 inputs_225__14, inputs_225__13, inputs_225__12, inputs_225__11, 
                 inputs_225__10, inputs_225__9, inputs_225__8, inputs_225__7, 
                 inputs_225__6, inputs_225__5, inputs_225__4, inputs_225__3, 
                 inputs_225__2, inputs_225__1, inputs_225__0, inputs_226__15, 
                 inputs_226__14, inputs_226__13, inputs_226__12, inputs_226__11, 
                 inputs_226__10, inputs_226__9, inputs_226__8, inputs_226__7, 
                 inputs_226__6, inputs_226__5, inputs_226__4, inputs_226__3, 
                 inputs_226__2, inputs_226__1, inputs_226__0, inputs_227__15, 
                 inputs_227__14, inputs_227__13, inputs_227__12, inputs_227__11, 
                 inputs_227__10, inputs_227__9, inputs_227__8, inputs_227__7, 
                 inputs_227__6, inputs_227__5, inputs_227__4, inputs_227__3, 
                 inputs_227__2, inputs_227__1, inputs_227__0, inputs_228__15, 
                 inputs_228__14, inputs_228__13, inputs_228__12, inputs_228__11, 
                 inputs_228__10, inputs_228__9, inputs_228__8, inputs_228__7, 
                 inputs_228__6, inputs_228__5, inputs_228__4, inputs_228__3, 
                 inputs_228__2, inputs_228__1, inputs_228__0, inputs_229__15, 
                 inputs_229__14, inputs_229__13, inputs_229__12, inputs_229__11, 
                 inputs_229__10, inputs_229__9, inputs_229__8, inputs_229__7, 
                 inputs_229__6, inputs_229__5, inputs_229__4, inputs_229__3, 
                 inputs_229__2, inputs_229__1, inputs_229__0, inputs_230__15, 
                 inputs_230__14, inputs_230__13, inputs_230__12, inputs_230__11, 
                 inputs_230__10, inputs_230__9, inputs_230__8, inputs_230__7, 
                 inputs_230__6, inputs_230__5, inputs_230__4, inputs_230__3, 
                 inputs_230__2, inputs_230__1, inputs_230__0, inputs_231__15, 
                 inputs_231__14, inputs_231__13, inputs_231__12, inputs_231__11, 
                 inputs_231__10, inputs_231__9, inputs_231__8, inputs_231__7, 
                 inputs_231__6, inputs_231__5, inputs_231__4, inputs_231__3, 
                 inputs_231__2, inputs_231__1, inputs_231__0, inputs_232__15, 
                 inputs_232__14, inputs_232__13, inputs_232__12, inputs_232__11, 
                 inputs_232__10, inputs_232__9, inputs_232__8, inputs_232__7, 
                 inputs_232__6, inputs_232__5, inputs_232__4, inputs_232__3, 
                 inputs_232__2, inputs_232__1, inputs_232__0, inputs_233__15, 
                 inputs_233__14, inputs_233__13, inputs_233__12, inputs_233__11, 
                 inputs_233__10, inputs_233__9, inputs_233__8, inputs_233__7, 
                 inputs_233__6, inputs_233__5, inputs_233__4, inputs_233__3, 
                 inputs_233__2, inputs_233__1, inputs_233__0, inputs_234__15, 
                 inputs_234__14, inputs_234__13, inputs_234__12, inputs_234__11, 
                 inputs_234__10, inputs_234__9, inputs_234__8, inputs_234__7, 
                 inputs_234__6, inputs_234__5, inputs_234__4, inputs_234__3, 
                 inputs_234__2, inputs_234__1, inputs_234__0, inputs_235__15, 
                 inputs_235__14, inputs_235__13, inputs_235__12, inputs_235__11, 
                 inputs_235__10, inputs_235__9, inputs_235__8, inputs_235__7, 
                 inputs_235__6, inputs_235__5, inputs_235__4, inputs_235__3, 
                 inputs_235__2, inputs_235__1, inputs_235__0, inputs_236__15, 
                 inputs_236__14, inputs_236__13, inputs_236__12, inputs_236__11, 
                 inputs_236__10, inputs_236__9, inputs_236__8, inputs_236__7, 
                 inputs_236__6, inputs_236__5, inputs_236__4, inputs_236__3, 
                 inputs_236__2, inputs_236__1, inputs_236__0, inputs_237__15, 
                 inputs_237__14, inputs_237__13, inputs_237__12, inputs_237__11, 
                 inputs_237__10, inputs_237__9, inputs_237__8, inputs_237__7, 
                 inputs_237__6, inputs_237__5, inputs_237__4, inputs_237__3, 
                 inputs_237__2, inputs_237__1, inputs_237__0, inputs_238__15, 
                 inputs_238__14, inputs_238__13, inputs_238__12, inputs_238__11, 
                 inputs_238__10, inputs_238__9, inputs_238__8, inputs_238__7, 
                 inputs_238__6, inputs_238__5, inputs_238__4, inputs_238__3, 
                 inputs_238__2, inputs_238__1, inputs_238__0, inputs_239__15, 
                 inputs_239__14, inputs_239__13, inputs_239__12, inputs_239__11, 
                 inputs_239__10, inputs_239__9, inputs_239__8, inputs_239__7, 
                 inputs_239__6, inputs_239__5, inputs_239__4, inputs_239__3, 
                 inputs_239__2, inputs_239__1, inputs_239__0, inputs_240__15, 
                 inputs_240__14, inputs_240__13, inputs_240__12, inputs_240__11, 
                 inputs_240__10, inputs_240__9, inputs_240__8, inputs_240__7, 
                 inputs_240__6, inputs_240__5, inputs_240__4, inputs_240__3, 
                 inputs_240__2, inputs_240__1, inputs_240__0, inputs_241__15, 
                 inputs_241__14, inputs_241__13, inputs_241__12, inputs_241__11, 
                 inputs_241__10, inputs_241__9, inputs_241__8, inputs_241__7, 
                 inputs_241__6, inputs_241__5, inputs_241__4, inputs_241__3, 
                 inputs_241__2, inputs_241__1, inputs_241__0, inputs_242__15, 
                 inputs_242__14, inputs_242__13, inputs_242__12, inputs_242__11, 
                 inputs_242__10, inputs_242__9, inputs_242__8, inputs_242__7, 
                 inputs_242__6, inputs_242__5, inputs_242__4, inputs_242__3, 
                 inputs_242__2, inputs_242__1, inputs_242__0, inputs_243__15, 
                 inputs_243__14, inputs_243__13, inputs_243__12, inputs_243__11, 
                 inputs_243__10, inputs_243__9, inputs_243__8, inputs_243__7, 
                 inputs_243__6, inputs_243__5, inputs_243__4, inputs_243__3, 
                 inputs_243__2, inputs_243__1, inputs_243__0, inputs_244__15, 
                 inputs_244__14, inputs_244__13, inputs_244__12, inputs_244__11, 
                 inputs_244__10, inputs_244__9, inputs_244__8, inputs_244__7, 
                 inputs_244__6, inputs_244__5, inputs_244__4, inputs_244__3, 
                 inputs_244__2, inputs_244__1, inputs_244__0, inputs_245__15, 
                 inputs_245__14, inputs_245__13, inputs_245__12, inputs_245__11, 
                 inputs_245__10, inputs_245__9, inputs_245__8, inputs_245__7, 
                 inputs_245__6, inputs_245__5, inputs_245__4, inputs_245__3, 
                 inputs_245__2, inputs_245__1, inputs_245__0, inputs_246__15, 
                 inputs_246__14, inputs_246__13, inputs_246__12, inputs_246__11, 
                 inputs_246__10, inputs_246__9, inputs_246__8, inputs_246__7, 
                 inputs_246__6, inputs_246__5, inputs_246__4, inputs_246__3, 
                 inputs_246__2, inputs_246__1, inputs_246__0, inputs_247__15, 
                 inputs_247__14, inputs_247__13, inputs_247__12, inputs_247__11, 
                 inputs_247__10, inputs_247__9, inputs_247__8, inputs_247__7, 
                 inputs_247__6, inputs_247__5, inputs_247__4, inputs_247__3, 
                 inputs_247__2, inputs_247__1, inputs_247__0, inputs_248__15, 
                 inputs_248__14, inputs_248__13, inputs_248__12, inputs_248__11, 
                 inputs_248__10, inputs_248__9, inputs_248__8, inputs_248__7, 
                 inputs_248__6, inputs_248__5, inputs_248__4, inputs_248__3, 
                 inputs_248__2, inputs_248__1, inputs_248__0, inputs_249__15, 
                 inputs_249__14, inputs_249__13, inputs_249__12, inputs_249__11, 
                 inputs_249__10, inputs_249__9, inputs_249__8, inputs_249__7, 
                 inputs_249__6, inputs_249__5, inputs_249__4, inputs_249__3, 
                 inputs_249__2, inputs_249__1, inputs_249__0, inputs_250__15, 
                 inputs_250__14, inputs_250__13, inputs_250__12, inputs_250__11, 
                 inputs_250__10, inputs_250__9, inputs_250__8, inputs_250__7, 
                 inputs_250__6, inputs_250__5, inputs_250__4, inputs_250__3, 
                 inputs_250__2, inputs_250__1, inputs_250__0, inputs_251__15, 
                 inputs_251__14, inputs_251__13, inputs_251__12, inputs_251__11, 
                 inputs_251__10, inputs_251__9, inputs_251__8, inputs_251__7, 
                 inputs_251__6, inputs_251__5, inputs_251__4, inputs_251__3, 
                 inputs_251__2, inputs_251__1, inputs_251__0, inputs_252__15, 
                 inputs_252__14, inputs_252__13, inputs_252__12, inputs_252__11, 
                 inputs_252__10, inputs_252__9, inputs_252__8, inputs_252__7, 
                 inputs_252__6, inputs_252__5, inputs_252__4, inputs_252__3, 
                 inputs_252__2, inputs_252__1, inputs_252__0, inputs_253__15, 
                 inputs_253__14, inputs_253__13, inputs_253__12, inputs_253__11, 
                 inputs_253__10, inputs_253__9, inputs_253__8, inputs_253__7, 
                 inputs_253__6, inputs_253__5, inputs_253__4, inputs_253__3, 
                 inputs_253__2, inputs_253__1, inputs_253__0, inputs_254__15, 
                 inputs_254__14, inputs_254__13, inputs_254__12, inputs_254__11, 
                 inputs_254__10, inputs_254__9, inputs_254__8, inputs_254__7, 
                 inputs_254__6, inputs_254__5, inputs_254__4, inputs_254__3, 
                 inputs_254__2, inputs_254__1, inputs_254__0, inputs_255__15, 
                 inputs_255__14, inputs_255__13, inputs_255__12, inputs_255__11, 
                 inputs_255__10, inputs_255__9, inputs_255__8, inputs_255__7, 
                 inputs_255__6, inputs_255__5, inputs_255__4, inputs_255__3, 
                 inputs_255__2, inputs_255__1, inputs_255__0, inputs_256__15, 
                 inputs_256__14, inputs_256__13, inputs_256__12, inputs_256__11, 
                 inputs_256__10, inputs_256__9, inputs_256__8, inputs_256__7, 
                 inputs_256__6, inputs_256__5, inputs_256__4, inputs_256__3, 
                 inputs_256__2, inputs_256__1, inputs_256__0, inputs_257__15, 
                 inputs_257__14, inputs_257__13, inputs_257__12, inputs_257__11, 
                 inputs_257__10, inputs_257__9, inputs_257__8, inputs_257__7, 
                 inputs_257__6, inputs_257__5, inputs_257__4, inputs_257__3, 
                 inputs_257__2, inputs_257__1, inputs_257__0, inputs_258__15, 
                 inputs_258__14, inputs_258__13, inputs_258__12, inputs_258__11, 
                 inputs_258__10, inputs_258__9, inputs_258__8, inputs_258__7, 
                 inputs_258__6, inputs_258__5, inputs_258__4, inputs_258__3, 
                 inputs_258__2, inputs_258__1, inputs_258__0, inputs_259__15, 
                 inputs_259__14, inputs_259__13, inputs_259__12, inputs_259__11, 
                 inputs_259__10, inputs_259__9, inputs_259__8, inputs_259__7, 
                 inputs_259__6, inputs_259__5, inputs_259__4, inputs_259__3, 
                 inputs_259__2, inputs_259__1, inputs_259__0, inputs_260__15, 
                 inputs_260__14, inputs_260__13, inputs_260__12, inputs_260__11, 
                 inputs_260__10, inputs_260__9, inputs_260__8, inputs_260__7, 
                 inputs_260__6, inputs_260__5, inputs_260__4, inputs_260__3, 
                 inputs_260__2, inputs_260__1, inputs_260__0, inputs_261__15, 
                 inputs_261__14, inputs_261__13, inputs_261__12, inputs_261__11, 
                 inputs_261__10, inputs_261__9, inputs_261__8, inputs_261__7, 
                 inputs_261__6, inputs_261__5, inputs_261__4, inputs_261__3, 
                 inputs_261__2, inputs_261__1, inputs_261__0, inputs_262__15, 
                 inputs_262__14, inputs_262__13, inputs_262__12, inputs_262__11, 
                 inputs_262__10, inputs_262__9, inputs_262__8, inputs_262__7, 
                 inputs_262__6, inputs_262__5, inputs_262__4, inputs_262__3, 
                 inputs_262__2, inputs_262__1, inputs_262__0, inputs_263__15, 
                 inputs_263__14, inputs_263__13, inputs_263__12, inputs_263__11, 
                 inputs_263__10, inputs_263__9, inputs_263__8, inputs_263__7, 
                 inputs_263__6, inputs_263__5, inputs_263__4, inputs_263__3, 
                 inputs_263__2, inputs_263__1, inputs_263__0, inputs_264__15, 
                 inputs_264__14, inputs_264__13, inputs_264__12, inputs_264__11, 
                 inputs_264__10, inputs_264__9, inputs_264__8, inputs_264__7, 
                 inputs_264__6, inputs_264__5, inputs_264__4, inputs_264__3, 
                 inputs_264__2, inputs_264__1, inputs_264__0, inputs_265__15, 
                 inputs_265__14, inputs_265__13, inputs_265__12, inputs_265__11, 
                 inputs_265__10, inputs_265__9, inputs_265__8, inputs_265__7, 
                 inputs_265__6, inputs_265__5, inputs_265__4, inputs_265__3, 
                 inputs_265__2, inputs_265__1, inputs_265__0, inputs_266__15, 
                 inputs_266__14, inputs_266__13, inputs_266__12, inputs_266__11, 
                 inputs_266__10, inputs_266__9, inputs_266__8, inputs_266__7, 
                 inputs_266__6, inputs_266__5, inputs_266__4, inputs_266__3, 
                 inputs_266__2, inputs_266__1, inputs_266__0, inputs_267__15, 
                 inputs_267__14, inputs_267__13, inputs_267__12, inputs_267__11, 
                 inputs_267__10, inputs_267__9, inputs_267__8, inputs_267__7, 
                 inputs_267__6, inputs_267__5, inputs_267__4, inputs_267__3, 
                 inputs_267__2, inputs_267__1, inputs_267__0, inputs_268__15, 
                 inputs_268__14, inputs_268__13, inputs_268__12, inputs_268__11, 
                 inputs_268__10, inputs_268__9, inputs_268__8, inputs_268__7, 
                 inputs_268__6, inputs_268__5, inputs_268__4, inputs_268__3, 
                 inputs_268__2, inputs_268__1, inputs_268__0, inputs_269__15, 
                 inputs_269__14, inputs_269__13, inputs_269__12, inputs_269__11, 
                 inputs_269__10, inputs_269__9, inputs_269__8, inputs_269__7, 
                 inputs_269__6, inputs_269__5, inputs_269__4, inputs_269__3, 
                 inputs_269__2, inputs_269__1, inputs_269__0, inputs_270__15, 
                 inputs_270__14, inputs_270__13, inputs_270__12, inputs_270__11, 
                 inputs_270__10, inputs_270__9, inputs_270__8, inputs_270__7, 
                 inputs_270__6, inputs_270__5, inputs_270__4, inputs_270__3, 
                 inputs_270__2, inputs_270__1, inputs_270__0, inputs_271__15, 
                 inputs_271__14, inputs_271__13, inputs_271__12, inputs_271__11, 
                 inputs_271__10, inputs_271__9, inputs_271__8, inputs_271__7, 
                 inputs_271__6, inputs_271__5, inputs_271__4, inputs_271__3, 
                 inputs_271__2, inputs_271__1, inputs_271__0, inputs_272__15, 
                 inputs_272__14, inputs_272__13, inputs_272__12, inputs_272__11, 
                 inputs_272__10, inputs_272__9, inputs_272__8, inputs_272__7, 
                 inputs_272__6, inputs_272__5, inputs_272__4, inputs_272__3, 
                 inputs_272__2, inputs_272__1, inputs_272__0, inputs_273__15, 
                 inputs_273__14, inputs_273__13, inputs_273__12, inputs_273__11, 
                 inputs_273__10, inputs_273__9, inputs_273__8, inputs_273__7, 
                 inputs_273__6, inputs_273__5, inputs_273__4, inputs_273__3, 
                 inputs_273__2, inputs_273__1, inputs_273__0, inputs_274__15, 
                 inputs_274__14, inputs_274__13, inputs_274__12, inputs_274__11, 
                 inputs_274__10, inputs_274__9, inputs_274__8, inputs_274__7, 
                 inputs_274__6, inputs_274__5, inputs_274__4, inputs_274__3, 
                 inputs_274__2, inputs_274__1, inputs_274__0, inputs_275__15, 
                 inputs_275__14, inputs_275__13, inputs_275__12, inputs_275__11, 
                 inputs_275__10, inputs_275__9, inputs_275__8, inputs_275__7, 
                 inputs_275__6, inputs_275__5, inputs_275__4, inputs_275__3, 
                 inputs_275__2, inputs_275__1, inputs_275__0, inputs_276__15, 
                 inputs_276__14, inputs_276__13, inputs_276__12, inputs_276__11, 
                 inputs_276__10, inputs_276__9, inputs_276__8, inputs_276__7, 
                 inputs_276__6, inputs_276__5, inputs_276__4, inputs_276__3, 
                 inputs_276__2, inputs_276__1, inputs_276__0, inputs_277__15, 
                 inputs_277__14, inputs_277__13, inputs_277__12, inputs_277__11, 
                 inputs_277__10, inputs_277__9, inputs_277__8, inputs_277__7, 
                 inputs_277__6, inputs_277__5, inputs_277__4, inputs_277__3, 
                 inputs_277__2, inputs_277__1, inputs_277__0, inputs_278__15, 
                 inputs_278__14, inputs_278__13, inputs_278__12, inputs_278__11, 
                 inputs_278__10, inputs_278__9, inputs_278__8, inputs_278__7, 
                 inputs_278__6, inputs_278__5, inputs_278__4, inputs_278__3, 
                 inputs_278__2, inputs_278__1, inputs_278__0, inputs_279__15, 
                 inputs_279__14, inputs_279__13, inputs_279__12, inputs_279__11, 
                 inputs_279__10, inputs_279__9, inputs_279__8, inputs_279__7, 
                 inputs_279__6, inputs_279__5, inputs_279__4, inputs_279__3, 
                 inputs_279__2, inputs_279__1, inputs_279__0, inputs_280__15, 
                 inputs_280__14, inputs_280__13, inputs_280__12, inputs_280__11, 
                 inputs_280__10, inputs_280__9, inputs_280__8, inputs_280__7, 
                 inputs_280__6, inputs_280__5, inputs_280__4, inputs_280__3, 
                 inputs_280__2, inputs_280__1, inputs_280__0, inputs_281__15, 
                 inputs_281__14, inputs_281__13, inputs_281__12, inputs_281__11, 
                 inputs_281__10, inputs_281__9, inputs_281__8, inputs_281__7, 
                 inputs_281__6, inputs_281__5, inputs_281__4, inputs_281__3, 
                 inputs_281__2, inputs_281__1, inputs_281__0, inputs_282__15, 
                 inputs_282__14, inputs_282__13, inputs_282__12, inputs_282__11, 
                 inputs_282__10, inputs_282__9, inputs_282__8, inputs_282__7, 
                 inputs_282__6, inputs_282__5, inputs_282__4, inputs_282__3, 
                 inputs_282__2, inputs_282__1, inputs_282__0, inputs_283__15, 
                 inputs_283__14, inputs_283__13, inputs_283__12, inputs_283__11, 
                 inputs_283__10, inputs_283__9, inputs_283__8, inputs_283__7, 
                 inputs_283__6, inputs_283__5, inputs_283__4, inputs_283__3, 
                 inputs_283__2, inputs_283__1, inputs_283__0, inputs_284__15, 
                 inputs_284__14, inputs_284__13, inputs_284__12, inputs_284__11, 
                 inputs_284__10, inputs_284__9, inputs_284__8, inputs_284__7, 
                 inputs_284__6, inputs_284__5, inputs_284__4, inputs_284__3, 
                 inputs_284__2, inputs_284__1, inputs_284__0, inputs_285__15, 
                 inputs_285__14, inputs_285__13, inputs_285__12, inputs_285__11, 
                 inputs_285__10, inputs_285__9, inputs_285__8, inputs_285__7, 
                 inputs_285__6, inputs_285__5, inputs_285__4, inputs_285__3, 
                 inputs_285__2, inputs_285__1, inputs_285__0, inputs_286__15, 
                 inputs_286__14, inputs_286__13, inputs_286__12, inputs_286__11, 
                 inputs_286__10, inputs_286__9, inputs_286__8, inputs_286__7, 
                 inputs_286__6, inputs_286__5, inputs_286__4, inputs_286__3, 
                 inputs_286__2, inputs_286__1, inputs_286__0, inputs_287__15, 
                 inputs_287__14, inputs_287__13, inputs_287__12, inputs_287__11, 
                 inputs_287__10, inputs_287__9, inputs_287__8, inputs_287__7, 
                 inputs_287__6, inputs_287__5, inputs_287__4, inputs_287__3, 
                 inputs_287__2, inputs_287__1, inputs_287__0, inputs_288__15, 
                 inputs_288__14, inputs_288__13, inputs_288__12, inputs_288__11, 
                 inputs_288__10, inputs_288__9, inputs_288__8, inputs_288__7, 
                 inputs_288__6, inputs_288__5, inputs_288__4, inputs_288__3, 
                 inputs_288__2, inputs_288__1, inputs_288__0, inputs_289__15, 
                 inputs_289__14, inputs_289__13, inputs_289__12, inputs_289__11, 
                 inputs_289__10, inputs_289__9, inputs_289__8, inputs_289__7, 
                 inputs_289__6, inputs_289__5, inputs_289__4, inputs_289__3, 
                 inputs_289__2, inputs_289__1, inputs_289__0, inputs_290__15, 
                 inputs_290__14, inputs_290__13, inputs_290__12, inputs_290__11, 
                 inputs_290__10, inputs_290__9, inputs_290__8, inputs_290__7, 
                 inputs_290__6, inputs_290__5, inputs_290__4, inputs_290__3, 
                 inputs_290__2, inputs_290__1, inputs_290__0, inputs_291__15, 
                 inputs_291__14, inputs_291__13, inputs_291__12, inputs_291__11, 
                 inputs_291__10, inputs_291__9, inputs_291__8, inputs_291__7, 
                 inputs_291__6, inputs_291__5, inputs_291__4, inputs_291__3, 
                 inputs_291__2, inputs_291__1, inputs_291__0, inputs_292__15, 
                 inputs_292__14, inputs_292__13, inputs_292__12, inputs_292__11, 
                 inputs_292__10, inputs_292__9, inputs_292__8, inputs_292__7, 
                 inputs_292__6, inputs_292__5, inputs_292__4, inputs_292__3, 
                 inputs_292__2, inputs_292__1, inputs_292__0, inputs_293__15, 
                 inputs_293__14, inputs_293__13, inputs_293__12, inputs_293__11, 
                 inputs_293__10, inputs_293__9, inputs_293__8, inputs_293__7, 
                 inputs_293__6, inputs_293__5, inputs_293__4, inputs_293__3, 
                 inputs_293__2, inputs_293__1, inputs_293__0, inputs_294__15, 
                 inputs_294__14, inputs_294__13, inputs_294__12, inputs_294__11, 
                 inputs_294__10, inputs_294__9, inputs_294__8, inputs_294__7, 
                 inputs_294__6, inputs_294__5, inputs_294__4, inputs_294__3, 
                 inputs_294__2, inputs_294__1, inputs_294__0, inputs_295__15, 
                 inputs_295__14, inputs_295__13, inputs_295__12, inputs_295__11, 
                 inputs_295__10, inputs_295__9, inputs_295__8, inputs_295__7, 
                 inputs_295__6, inputs_295__5, inputs_295__4, inputs_295__3, 
                 inputs_295__2, inputs_295__1, inputs_295__0, inputs_296__15, 
                 inputs_296__14, inputs_296__13, inputs_296__12, inputs_296__11, 
                 inputs_296__10, inputs_296__9, inputs_296__8, inputs_296__7, 
                 inputs_296__6, inputs_296__5, inputs_296__4, inputs_296__3, 
                 inputs_296__2, inputs_296__1, inputs_296__0, inputs_297__15, 
                 inputs_297__14, inputs_297__13, inputs_297__12, inputs_297__11, 
                 inputs_297__10, inputs_297__9, inputs_297__8, inputs_297__7, 
                 inputs_297__6, inputs_297__5, inputs_297__4, inputs_297__3, 
                 inputs_297__2, inputs_297__1, inputs_297__0, inputs_298__15, 
                 inputs_298__14, inputs_298__13, inputs_298__12, inputs_298__11, 
                 inputs_298__10, inputs_298__9, inputs_298__8, inputs_298__7, 
                 inputs_298__6, inputs_298__5, inputs_298__4, inputs_298__3, 
                 inputs_298__2, inputs_298__1, inputs_298__0, inputs_299__15, 
                 inputs_299__14, inputs_299__13, inputs_299__12, inputs_299__11, 
                 inputs_299__10, inputs_299__9, inputs_299__8, inputs_299__7, 
                 inputs_299__6, inputs_299__5, inputs_299__4, inputs_299__3, 
                 inputs_299__2, inputs_299__1, inputs_299__0, inputs_300__15, 
                 inputs_300__14, inputs_300__13, inputs_300__12, inputs_300__11, 
                 inputs_300__10, inputs_300__9, inputs_300__8, inputs_300__7, 
                 inputs_300__6, inputs_300__5, inputs_300__4, inputs_300__3, 
                 inputs_300__2, inputs_300__1, inputs_300__0, inputs_301__15, 
                 inputs_301__14, inputs_301__13, inputs_301__12, inputs_301__11, 
                 inputs_301__10, inputs_301__9, inputs_301__8, inputs_301__7, 
                 inputs_301__6, inputs_301__5, inputs_301__4, inputs_301__3, 
                 inputs_301__2, inputs_301__1, inputs_301__0, inputs_302__15, 
                 inputs_302__14, inputs_302__13, inputs_302__12, inputs_302__11, 
                 inputs_302__10, inputs_302__9, inputs_302__8, inputs_302__7, 
                 inputs_302__6, inputs_302__5, inputs_302__4, inputs_302__3, 
                 inputs_302__2, inputs_302__1, inputs_302__0, inputs_303__15, 
                 inputs_303__14, inputs_303__13, inputs_303__12, inputs_303__11, 
                 inputs_303__10, inputs_303__9, inputs_303__8, inputs_303__7, 
                 inputs_303__6, inputs_303__5, inputs_303__4, inputs_303__3, 
                 inputs_303__2, inputs_303__1, inputs_303__0, inputs_304__15, 
                 inputs_304__14, inputs_304__13, inputs_304__12, inputs_304__11, 
                 inputs_304__10, inputs_304__9, inputs_304__8, inputs_304__7, 
                 inputs_304__6, inputs_304__5, inputs_304__4, inputs_304__3, 
                 inputs_304__2, inputs_304__1, inputs_304__0, inputs_305__15, 
                 inputs_305__14, inputs_305__13, inputs_305__12, inputs_305__11, 
                 inputs_305__10, inputs_305__9, inputs_305__8, inputs_305__7, 
                 inputs_305__6, inputs_305__5, inputs_305__4, inputs_305__3, 
                 inputs_305__2, inputs_305__1, inputs_305__0, inputs_306__15, 
                 inputs_306__14, inputs_306__13, inputs_306__12, inputs_306__11, 
                 inputs_306__10, inputs_306__9, inputs_306__8, inputs_306__7, 
                 inputs_306__6, inputs_306__5, inputs_306__4, inputs_306__3, 
                 inputs_306__2, inputs_306__1, inputs_306__0, inputs_307__15, 
                 inputs_307__14, inputs_307__13, inputs_307__12, inputs_307__11, 
                 inputs_307__10, inputs_307__9, inputs_307__8, inputs_307__7, 
                 inputs_307__6, inputs_307__5, inputs_307__4, inputs_307__3, 
                 inputs_307__2, inputs_307__1, inputs_307__0, inputs_308__15, 
                 inputs_308__14, inputs_308__13, inputs_308__12, inputs_308__11, 
                 inputs_308__10, inputs_308__9, inputs_308__8, inputs_308__7, 
                 inputs_308__6, inputs_308__5, inputs_308__4, inputs_308__3, 
                 inputs_308__2, inputs_308__1, inputs_308__0, inputs_309__15, 
                 inputs_309__14, inputs_309__13, inputs_309__12, inputs_309__11, 
                 inputs_309__10, inputs_309__9, inputs_309__8, inputs_309__7, 
                 inputs_309__6, inputs_309__5, inputs_309__4, inputs_309__3, 
                 inputs_309__2, inputs_309__1, inputs_309__0, inputs_310__15, 
                 inputs_310__14, inputs_310__13, inputs_310__12, inputs_310__11, 
                 inputs_310__10, inputs_310__9, inputs_310__8, inputs_310__7, 
                 inputs_310__6, inputs_310__5, inputs_310__4, inputs_310__3, 
                 inputs_310__2, inputs_310__1, inputs_310__0, inputs_311__15, 
                 inputs_311__14, inputs_311__13, inputs_311__12, inputs_311__11, 
                 inputs_311__10, inputs_311__9, inputs_311__8, inputs_311__7, 
                 inputs_311__6, inputs_311__5, inputs_311__4, inputs_311__3, 
                 inputs_311__2, inputs_311__1, inputs_311__0, inputs_312__15, 
                 inputs_312__14, inputs_312__13, inputs_312__12, inputs_312__11, 
                 inputs_312__10, inputs_312__9, inputs_312__8, inputs_312__7, 
                 inputs_312__6, inputs_312__5, inputs_312__4, inputs_312__3, 
                 inputs_312__2, inputs_312__1, inputs_312__0, inputs_313__15, 
                 inputs_313__14, inputs_313__13, inputs_313__12, inputs_313__11, 
                 inputs_313__10, inputs_313__9, inputs_313__8, inputs_313__7, 
                 inputs_313__6, inputs_313__5, inputs_313__4, inputs_313__3, 
                 inputs_313__2, inputs_313__1, inputs_313__0, inputs_314__15, 
                 inputs_314__14, inputs_314__13, inputs_314__12, inputs_314__11, 
                 inputs_314__10, inputs_314__9, inputs_314__8, inputs_314__7, 
                 inputs_314__6, inputs_314__5, inputs_314__4, inputs_314__3, 
                 inputs_314__2, inputs_314__1, inputs_314__0, inputs_315__15, 
                 inputs_315__14, inputs_315__13, inputs_315__12, inputs_315__11, 
                 inputs_315__10, inputs_315__9, inputs_315__8, inputs_315__7, 
                 inputs_315__6, inputs_315__5, inputs_315__4, inputs_315__3, 
                 inputs_315__2, inputs_315__1, inputs_315__0, inputs_316__15, 
                 inputs_316__14, inputs_316__13, inputs_316__12, inputs_316__11, 
                 inputs_316__10, inputs_316__9, inputs_316__8, inputs_316__7, 
                 inputs_316__6, inputs_316__5, inputs_316__4, inputs_316__3, 
                 inputs_316__2, inputs_316__1, inputs_316__0, inputs_317__15, 
                 inputs_317__14, inputs_317__13, inputs_317__12, inputs_317__11, 
                 inputs_317__10, inputs_317__9, inputs_317__8, inputs_317__7, 
                 inputs_317__6, inputs_317__5, inputs_317__4, inputs_317__3, 
                 inputs_317__2, inputs_317__1, inputs_317__0, inputs_318__15, 
                 inputs_318__14, inputs_318__13, inputs_318__12, inputs_318__11, 
                 inputs_318__10, inputs_318__9, inputs_318__8, inputs_318__7, 
                 inputs_318__6, inputs_318__5, inputs_318__4, inputs_318__3, 
                 inputs_318__2, inputs_318__1, inputs_318__0, inputs_319__15, 
                 inputs_319__14, inputs_319__13, inputs_319__12, inputs_319__11, 
                 inputs_319__10, inputs_319__9, inputs_319__8, inputs_319__7, 
                 inputs_319__6, inputs_319__5, inputs_319__4, inputs_319__3, 
                 inputs_319__2, inputs_319__1, inputs_319__0, inputs_320__15, 
                 inputs_320__14, inputs_320__13, inputs_320__12, inputs_320__11, 
                 inputs_320__10, inputs_320__9, inputs_320__8, inputs_320__7, 
                 inputs_320__6, inputs_320__5, inputs_320__4, inputs_320__3, 
                 inputs_320__2, inputs_320__1, inputs_320__0, inputs_321__15, 
                 inputs_321__14, inputs_321__13, inputs_321__12, inputs_321__11, 
                 inputs_321__10, inputs_321__9, inputs_321__8, inputs_321__7, 
                 inputs_321__6, inputs_321__5, inputs_321__4, inputs_321__3, 
                 inputs_321__2, inputs_321__1, inputs_321__0, inputs_322__15, 
                 inputs_322__14, inputs_322__13, inputs_322__12, inputs_322__11, 
                 inputs_322__10, inputs_322__9, inputs_322__8, inputs_322__7, 
                 inputs_322__6, inputs_322__5, inputs_322__4, inputs_322__3, 
                 inputs_322__2, inputs_322__1, inputs_322__0, inputs_323__15, 
                 inputs_323__14, inputs_323__13, inputs_323__12, inputs_323__11, 
                 inputs_323__10, inputs_323__9, inputs_323__8, inputs_323__7, 
                 inputs_323__6, inputs_323__5, inputs_323__4, inputs_323__3, 
                 inputs_323__2, inputs_323__1, inputs_323__0, inputs_324__15, 
                 inputs_324__14, inputs_324__13, inputs_324__12, inputs_324__11, 
                 inputs_324__10, inputs_324__9, inputs_324__8, inputs_324__7, 
                 inputs_324__6, inputs_324__5, inputs_324__4, inputs_324__3, 
                 inputs_324__2, inputs_324__1, inputs_324__0, inputs_325__15, 
                 inputs_325__14, inputs_325__13, inputs_325__12, inputs_325__11, 
                 inputs_325__10, inputs_325__9, inputs_325__8, inputs_325__7, 
                 inputs_325__6, inputs_325__5, inputs_325__4, inputs_325__3, 
                 inputs_325__2, inputs_325__1, inputs_325__0, inputs_326__15, 
                 inputs_326__14, inputs_326__13, inputs_326__12, inputs_326__11, 
                 inputs_326__10, inputs_326__9, inputs_326__8, inputs_326__7, 
                 inputs_326__6, inputs_326__5, inputs_326__4, inputs_326__3, 
                 inputs_326__2, inputs_326__1, inputs_326__0, inputs_327__15, 
                 inputs_327__14, inputs_327__13, inputs_327__12, inputs_327__11, 
                 inputs_327__10, inputs_327__9, inputs_327__8, inputs_327__7, 
                 inputs_327__6, inputs_327__5, inputs_327__4, inputs_327__3, 
                 inputs_327__2, inputs_327__1, inputs_327__0, inputs_328__15, 
                 inputs_328__14, inputs_328__13, inputs_328__12, inputs_328__11, 
                 inputs_328__10, inputs_328__9, inputs_328__8, inputs_328__7, 
                 inputs_328__6, inputs_328__5, inputs_328__4, inputs_328__3, 
                 inputs_328__2, inputs_328__1, inputs_328__0, inputs_329__15, 
                 inputs_329__14, inputs_329__13, inputs_329__12, inputs_329__11, 
                 inputs_329__10, inputs_329__9, inputs_329__8, inputs_329__7, 
                 inputs_329__6, inputs_329__5, inputs_329__4, inputs_329__3, 
                 inputs_329__2, inputs_329__1, inputs_329__0, inputs_330__15, 
                 inputs_330__14, inputs_330__13, inputs_330__12, inputs_330__11, 
                 inputs_330__10, inputs_330__9, inputs_330__8, inputs_330__7, 
                 inputs_330__6, inputs_330__5, inputs_330__4, inputs_330__3, 
                 inputs_330__2, inputs_330__1, inputs_330__0, inputs_331__15, 
                 inputs_331__14, inputs_331__13, inputs_331__12, inputs_331__11, 
                 inputs_331__10, inputs_331__9, inputs_331__8, inputs_331__7, 
                 inputs_331__6, inputs_331__5, inputs_331__4, inputs_331__3, 
                 inputs_331__2, inputs_331__1, inputs_331__0, inputs_332__15, 
                 inputs_332__14, inputs_332__13, inputs_332__12, inputs_332__11, 
                 inputs_332__10, inputs_332__9, inputs_332__8, inputs_332__7, 
                 inputs_332__6, inputs_332__5, inputs_332__4, inputs_332__3, 
                 inputs_332__2, inputs_332__1, inputs_332__0, inputs_333__15, 
                 inputs_333__14, inputs_333__13, inputs_333__12, inputs_333__11, 
                 inputs_333__10, inputs_333__9, inputs_333__8, inputs_333__7, 
                 inputs_333__6, inputs_333__5, inputs_333__4, inputs_333__3, 
                 inputs_333__2, inputs_333__1, inputs_333__0, inputs_334__15, 
                 inputs_334__14, inputs_334__13, inputs_334__12, inputs_334__11, 
                 inputs_334__10, inputs_334__9, inputs_334__8, inputs_334__7, 
                 inputs_334__6, inputs_334__5, inputs_334__4, inputs_334__3, 
                 inputs_334__2, inputs_334__1, inputs_334__0, inputs_335__15, 
                 inputs_335__14, inputs_335__13, inputs_335__12, inputs_335__11, 
                 inputs_335__10, inputs_335__9, inputs_335__8, inputs_335__7, 
                 inputs_335__6, inputs_335__5, inputs_335__4, inputs_335__3, 
                 inputs_335__2, inputs_335__1, inputs_335__0, inputs_336__15, 
                 inputs_336__14, inputs_336__13, inputs_336__12, inputs_336__11, 
                 inputs_336__10, inputs_336__9, inputs_336__8, inputs_336__7, 
                 inputs_336__6, inputs_336__5, inputs_336__4, inputs_336__3, 
                 inputs_336__2, inputs_336__1, inputs_336__0, inputs_337__15, 
                 inputs_337__14, inputs_337__13, inputs_337__12, inputs_337__11, 
                 inputs_337__10, inputs_337__9, inputs_337__8, inputs_337__7, 
                 inputs_337__6, inputs_337__5, inputs_337__4, inputs_337__3, 
                 inputs_337__2, inputs_337__1, inputs_337__0, inputs_338__15, 
                 inputs_338__14, inputs_338__13, inputs_338__12, inputs_338__11, 
                 inputs_338__10, inputs_338__9, inputs_338__8, inputs_338__7, 
                 inputs_338__6, inputs_338__5, inputs_338__4, inputs_338__3, 
                 inputs_338__2, inputs_338__1, inputs_338__0, inputs_339__15, 
                 inputs_339__14, inputs_339__13, inputs_339__12, inputs_339__11, 
                 inputs_339__10, inputs_339__9, inputs_339__8, inputs_339__7, 
                 inputs_339__6, inputs_339__5, inputs_339__4, inputs_339__3, 
                 inputs_339__2, inputs_339__1, inputs_339__0, inputs_340__15, 
                 inputs_340__14, inputs_340__13, inputs_340__12, inputs_340__11, 
                 inputs_340__10, inputs_340__9, inputs_340__8, inputs_340__7, 
                 inputs_340__6, inputs_340__5, inputs_340__4, inputs_340__3, 
                 inputs_340__2, inputs_340__1, inputs_340__0, inputs_341__15, 
                 inputs_341__14, inputs_341__13, inputs_341__12, inputs_341__11, 
                 inputs_341__10, inputs_341__9, inputs_341__8, inputs_341__7, 
                 inputs_341__6, inputs_341__5, inputs_341__4, inputs_341__3, 
                 inputs_341__2, inputs_341__1, inputs_341__0, inputs_342__15, 
                 inputs_342__14, inputs_342__13, inputs_342__12, inputs_342__11, 
                 inputs_342__10, inputs_342__9, inputs_342__8, inputs_342__7, 
                 inputs_342__6, inputs_342__5, inputs_342__4, inputs_342__3, 
                 inputs_342__2, inputs_342__1, inputs_342__0, inputs_343__15, 
                 inputs_343__14, inputs_343__13, inputs_343__12, inputs_343__11, 
                 inputs_343__10, inputs_343__9, inputs_343__8, inputs_343__7, 
                 inputs_343__6, inputs_343__5, inputs_343__4, inputs_343__3, 
                 inputs_343__2, inputs_343__1, inputs_343__0, inputs_344__15, 
                 inputs_344__14, inputs_344__13, inputs_344__12, inputs_344__11, 
                 inputs_344__10, inputs_344__9, inputs_344__8, inputs_344__7, 
                 inputs_344__6, inputs_344__5, inputs_344__4, inputs_344__3, 
                 inputs_344__2, inputs_344__1, inputs_344__0, inputs_345__15, 
                 inputs_345__14, inputs_345__13, inputs_345__12, inputs_345__11, 
                 inputs_345__10, inputs_345__9, inputs_345__8, inputs_345__7, 
                 inputs_345__6, inputs_345__5, inputs_345__4, inputs_345__3, 
                 inputs_345__2, inputs_345__1, inputs_345__0, inputs_346__15, 
                 inputs_346__14, inputs_346__13, inputs_346__12, inputs_346__11, 
                 inputs_346__10, inputs_346__9, inputs_346__8, inputs_346__7, 
                 inputs_346__6, inputs_346__5, inputs_346__4, inputs_346__3, 
                 inputs_346__2, inputs_346__1, inputs_346__0, inputs_347__15, 
                 inputs_347__14, inputs_347__13, inputs_347__12, inputs_347__11, 
                 inputs_347__10, inputs_347__9, inputs_347__8, inputs_347__7, 
                 inputs_347__6, inputs_347__5, inputs_347__4, inputs_347__3, 
                 inputs_347__2, inputs_347__1, inputs_347__0, inputs_348__15, 
                 inputs_348__14, inputs_348__13, inputs_348__12, inputs_348__11, 
                 inputs_348__10, inputs_348__9, inputs_348__8, inputs_348__7, 
                 inputs_348__6, inputs_348__5, inputs_348__4, inputs_348__3, 
                 inputs_348__2, inputs_348__1, inputs_348__0, inputs_349__15, 
                 inputs_349__14, inputs_349__13, inputs_349__12, inputs_349__11, 
                 inputs_349__10, inputs_349__9, inputs_349__8, inputs_349__7, 
                 inputs_349__6, inputs_349__5, inputs_349__4, inputs_349__3, 
                 inputs_349__2, inputs_349__1, inputs_349__0, inputs_350__15, 
                 inputs_350__14, inputs_350__13, inputs_350__12, inputs_350__11, 
                 inputs_350__10, inputs_350__9, inputs_350__8, inputs_350__7, 
                 inputs_350__6, inputs_350__5, inputs_350__4, inputs_350__3, 
                 inputs_350__2, inputs_350__1, inputs_350__0, inputs_351__15, 
                 inputs_351__14, inputs_351__13, inputs_351__12, inputs_351__11, 
                 inputs_351__10, inputs_351__9, inputs_351__8, inputs_351__7, 
                 inputs_351__6, inputs_351__5, inputs_351__4, inputs_351__3, 
                 inputs_351__2, inputs_351__1, inputs_351__0, inputs_352__15, 
                 inputs_352__14, inputs_352__13, inputs_352__12, inputs_352__11, 
                 inputs_352__10, inputs_352__9, inputs_352__8, inputs_352__7, 
                 inputs_352__6, inputs_352__5, inputs_352__4, inputs_352__3, 
                 inputs_352__2, inputs_352__1, inputs_352__0, inputs_353__15, 
                 inputs_353__14, inputs_353__13, inputs_353__12, inputs_353__11, 
                 inputs_353__10, inputs_353__9, inputs_353__8, inputs_353__7, 
                 inputs_353__6, inputs_353__5, inputs_353__4, inputs_353__3, 
                 inputs_353__2, inputs_353__1, inputs_353__0, inputs_354__15, 
                 inputs_354__14, inputs_354__13, inputs_354__12, inputs_354__11, 
                 inputs_354__10, inputs_354__9, inputs_354__8, inputs_354__7, 
                 inputs_354__6, inputs_354__5, inputs_354__4, inputs_354__3, 
                 inputs_354__2, inputs_354__1, inputs_354__0, inputs_355__15, 
                 inputs_355__14, inputs_355__13, inputs_355__12, inputs_355__11, 
                 inputs_355__10, inputs_355__9, inputs_355__8, inputs_355__7, 
                 inputs_355__6, inputs_355__5, inputs_355__4, inputs_355__3, 
                 inputs_355__2, inputs_355__1, inputs_355__0, inputs_356__15, 
                 inputs_356__14, inputs_356__13, inputs_356__12, inputs_356__11, 
                 inputs_356__10, inputs_356__9, inputs_356__8, inputs_356__7, 
                 inputs_356__6, inputs_356__5, inputs_356__4, inputs_356__3, 
                 inputs_356__2, inputs_356__1, inputs_356__0, inputs_357__15, 
                 inputs_357__14, inputs_357__13, inputs_357__12, inputs_357__11, 
                 inputs_357__10, inputs_357__9, inputs_357__8, inputs_357__7, 
                 inputs_357__6, inputs_357__5, inputs_357__4, inputs_357__3, 
                 inputs_357__2, inputs_357__1, inputs_357__0, inputs_358__15, 
                 inputs_358__14, inputs_358__13, inputs_358__12, inputs_358__11, 
                 inputs_358__10, inputs_358__9, inputs_358__8, inputs_358__7, 
                 inputs_358__6, inputs_358__5, inputs_358__4, inputs_358__3, 
                 inputs_358__2, inputs_358__1, inputs_358__0, inputs_359__15, 
                 inputs_359__14, inputs_359__13, inputs_359__12, inputs_359__11, 
                 inputs_359__10, inputs_359__9, inputs_359__8, inputs_359__7, 
                 inputs_359__6, inputs_359__5, inputs_359__4, inputs_359__3, 
                 inputs_359__2, inputs_359__1, inputs_359__0, inputs_360__15, 
                 inputs_360__14, inputs_360__13, inputs_360__12, inputs_360__11, 
                 inputs_360__10, inputs_360__9, inputs_360__8, inputs_360__7, 
                 inputs_360__6, inputs_360__5, inputs_360__4, inputs_360__3, 
                 inputs_360__2, inputs_360__1, inputs_360__0, inputs_361__15, 
                 inputs_361__14, inputs_361__13, inputs_361__12, inputs_361__11, 
                 inputs_361__10, inputs_361__9, inputs_361__8, inputs_361__7, 
                 inputs_361__6, inputs_361__5, inputs_361__4, inputs_361__3, 
                 inputs_361__2, inputs_361__1, inputs_361__0, inputs_362__15, 
                 inputs_362__14, inputs_362__13, inputs_362__12, inputs_362__11, 
                 inputs_362__10, inputs_362__9, inputs_362__8, inputs_362__7, 
                 inputs_362__6, inputs_362__5, inputs_362__4, inputs_362__3, 
                 inputs_362__2, inputs_362__1, inputs_362__0, inputs_363__15, 
                 inputs_363__14, inputs_363__13, inputs_363__12, inputs_363__11, 
                 inputs_363__10, inputs_363__9, inputs_363__8, inputs_363__7, 
                 inputs_363__6, inputs_363__5, inputs_363__4, inputs_363__3, 
                 inputs_363__2, inputs_363__1, inputs_363__0, inputs_364__15, 
                 inputs_364__14, inputs_364__13, inputs_364__12, inputs_364__11, 
                 inputs_364__10, inputs_364__9, inputs_364__8, inputs_364__7, 
                 inputs_364__6, inputs_364__5, inputs_364__4, inputs_364__3, 
                 inputs_364__2, inputs_364__1, inputs_364__0, inputs_365__15, 
                 inputs_365__14, inputs_365__13, inputs_365__12, inputs_365__11, 
                 inputs_365__10, inputs_365__9, inputs_365__8, inputs_365__7, 
                 inputs_365__6, inputs_365__5, inputs_365__4, inputs_365__3, 
                 inputs_365__2, inputs_365__1, inputs_365__0, inputs_366__15, 
                 inputs_366__14, inputs_366__13, inputs_366__12, inputs_366__11, 
                 inputs_366__10, inputs_366__9, inputs_366__8, inputs_366__7, 
                 inputs_366__6, inputs_366__5, inputs_366__4, inputs_366__3, 
                 inputs_366__2, inputs_366__1, inputs_366__0, inputs_367__15, 
                 inputs_367__14, inputs_367__13, inputs_367__12, inputs_367__11, 
                 inputs_367__10, inputs_367__9, inputs_367__8, inputs_367__7, 
                 inputs_367__6, inputs_367__5, inputs_367__4, inputs_367__3, 
                 inputs_367__2, inputs_367__1, inputs_367__0, inputs_368__15, 
                 inputs_368__14, inputs_368__13, inputs_368__12, inputs_368__11, 
                 inputs_368__10, inputs_368__9, inputs_368__8, inputs_368__7, 
                 inputs_368__6, inputs_368__5, inputs_368__4, inputs_368__3, 
                 inputs_368__2, inputs_368__1, inputs_368__0, inputs_369__15, 
                 inputs_369__14, inputs_369__13, inputs_369__12, inputs_369__11, 
                 inputs_369__10, inputs_369__9, inputs_369__8, inputs_369__7, 
                 inputs_369__6, inputs_369__5, inputs_369__4, inputs_369__3, 
                 inputs_369__2, inputs_369__1, inputs_369__0, inputs_370__15, 
                 inputs_370__14, inputs_370__13, inputs_370__12, inputs_370__11, 
                 inputs_370__10, inputs_370__9, inputs_370__8, inputs_370__7, 
                 inputs_370__6, inputs_370__5, inputs_370__4, inputs_370__3, 
                 inputs_370__2, inputs_370__1, inputs_370__0, inputs_371__15, 
                 inputs_371__14, inputs_371__13, inputs_371__12, inputs_371__11, 
                 inputs_371__10, inputs_371__9, inputs_371__8, inputs_371__7, 
                 inputs_371__6, inputs_371__5, inputs_371__4, inputs_371__3, 
                 inputs_371__2, inputs_371__1, inputs_371__0, inputs_372__15, 
                 inputs_372__14, inputs_372__13, inputs_372__12, inputs_372__11, 
                 inputs_372__10, inputs_372__9, inputs_372__8, inputs_372__7, 
                 inputs_372__6, inputs_372__5, inputs_372__4, inputs_372__3, 
                 inputs_372__2, inputs_372__1, inputs_372__0, inputs_373__15, 
                 inputs_373__14, inputs_373__13, inputs_373__12, inputs_373__11, 
                 inputs_373__10, inputs_373__9, inputs_373__8, inputs_373__7, 
                 inputs_373__6, inputs_373__5, inputs_373__4, inputs_373__3, 
                 inputs_373__2, inputs_373__1, inputs_373__0, inputs_374__15, 
                 inputs_374__14, inputs_374__13, inputs_374__12, inputs_374__11, 
                 inputs_374__10, inputs_374__9, inputs_374__8, inputs_374__7, 
                 inputs_374__6, inputs_374__5, inputs_374__4, inputs_374__3, 
                 inputs_374__2, inputs_374__1, inputs_374__0, inputs_375__15, 
                 inputs_375__14, inputs_375__13, inputs_375__12, inputs_375__11, 
                 inputs_375__10, inputs_375__9, inputs_375__8, inputs_375__7, 
                 inputs_375__6, inputs_375__5, inputs_375__4, inputs_375__3, 
                 inputs_375__2, inputs_375__1, inputs_375__0, inputs_376__15, 
                 inputs_376__14, inputs_376__13, inputs_376__12, inputs_376__11, 
                 inputs_376__10, inputs_376__9, inputs_376__8, inputs_376__7, 
                 inputs_376__6, inputs_376__5, inputs_376__4, inputs_376__3, 
                 inputs_376__2, inputs_376__1, inputs_376__0, inputs_377__15, 
                 inputs_377__14, inputs_377__13, inputs_377__12, inputs_377__11, 
                 inputs_377__10, inputs_377__9, inputs_377__8, inputs_377__7, 
                 inputs_377__6, inputs_377__5, inputs_377__4, inputs_377__3, 
                 inputs_377__2, inputs_377__1, inputs_377__0, inputs_378__15, 
                 inputs_378__14, inputs_378__13, inputs_378__12, inputs_378__11, 
                 inputs_378__10, inputs_378__9, inputs_378__8, inputs_378__7, 
                 inputs_378__6, inputs_378__5, inputs_378__4, inputs_378__3, 
                 inputs_378__2, inputs_378__1, inputs_378__0, inputs_379__15, 
                 inputs_379__14, inputs_379__13, inputs_379__12, inputs_379__11, 
                 inputs_379__10, inputs_379__9, inputs_379__8, inputs_379__7, 
                 inputs_379__6, inputs_379__5, inputs_379__4, inputs_379__3, 
                 inputs_379__2, inputs_379__1, inputs_379__0, inputs_380__15, 
                 inputs_380__14, inputs_380__13, inputs_380__12, inputs_380__11, 
                 inputs_380__10, inputs_380__9, inputs_380__8, inputs_380__7, 
                 inputs_380__6, inputs_380__5, inputs_380__4, inputs_380__3, 
                 inputs_380__2, inputs_380__1, inputs_380__0, inputs_381__15, 
                 inputs_381__14, inputs_381__13, inputs_381__12, inputs_381__11, 
                 inputs_381__10, inputs_381__9, inputs_381__8, inputs_381__7, 
                 inputs_381__6, inputs_381__5, inputs_381__4, inputs_381__3, 
                 inputs_381__2, inputs_381__1, inputs_381__0, inputs_382__15, 
                 inputs_382__14, inputs_382__13, inputs_382__12, inputs_382__11, 
                 inputs_382__10, inputs_382__9, inputs_382__8, inputs_382__7, 
                 inputs_382__6, inputs_382__5, inputs_382__4, inputs_382__3, 
                 inputs_382__2, inputs_382__1, inputs_382__0, inputs_383__15, 
                 inputs_383__14, inputs_383__13, inputs_383__12, inputs_383__11, 
                 inputs_383__10, inputs_383__9, inputs_383__8, inputs_383__7, 
                 inputs_383__6, inputs_383__5, inputs_383__4, inputs_383__3, 
                 inputs_383__2, inputs_383__1, inputs_383__0, inputs_384__15, 
                 inputs_384__14, inputs_384__13, inputs_384__12, inputs_384__11, 
                 inputs_384__10, inputs_384__9, inputs_384__8, inputs_384__7, 
                 inputs_384__6, inputs_384__5, inputs_384__4, inputs_384__3, 
                 inputs_384__2, inputs_384__1, inputs_384__0, inputs_385__15, 
                 inputs_385__14, inputs_385__13, inputs_385__12, inputs_385__11, 
                 inputs_385__10, inputs_385__9, inputs_385__8, inputs_385__7, 
                 inputs_385__6, inputs_385__5, inputs_385__4, inputs_385__3, 
                 inputs_385__2, inputs_385__1, inputs_385__0, inputs_386__15, 
                 inputs_386__14, inputs_386__13, inputs_386__12, inputs_386__11, 
                 inputs_386__10, inputs_386__9, inputs_386__8, inputs_386__7, 
                 inputs_386__6, inputs_386__5, inputs_386__4, inputs_386__3, 
                 inputs_386__2, inputs_386__1, inputs_386__0, inputs_387__15, 
                 inputs_387__14, inputs_387__13, inputs_387__12, inputs_387__11, 
                 inputs_387__10, inputs_387__9, inputs_387__8, inputs_387__7, 
                 inputs_387__6, inputs_387__5, inputs_387__4, inputs_387__3, 
                 inputs_387__2, inputs_387__1, inputs_387__0, inputs_388__15, 
                 inputs_388__14, inputs_388__13, inputs_388__12, inputs_388__11, 
                 inputs_388__10, inputs_388__9, inputs_388__8, inputs_388__7, 
                 inputs_388__6, inputs_388__5, inputs_388__4, inputs_388__3, 
                 inputs_388__2, inputs_388__1, inputs_388__0, inputs_389__15, 
                 inputs_389__14, inputs_389__13, inputs_389__12, inputs_389__11, 
                 inputs_389__10, inputs_389__9, inputs_389__8, inputs_389__7, 
                 inputs_389__6, inputs_389__5, inputs_389__4, inputs_389__3, 
                 inputs_389__2, inputs_389__1, inputs_389__0, inputs_390__15, 
                 inputs_390__14, inputs_390__13, inputs_390__12, inputs_390__11, 
                 inputs_390__10, inputs_390__9, inputs_390__8, inputs_390__7, 
                 inputs_390__6, inputs_390__5, inputs_390__4, inputs_390__3, 
                 inputs_390__2, inputs_390__1, inputs_390__0, inputs_391__15, 
                 inputs_391__14, inputs_391__13, inputs_391__12, inputs_391__11, 
                 inputs_391__10, inputs_391__9, inputs_391__8, inputs_391__7, 
                 inputs_391__6, inputs_391__5, inputs_391__4, inputs_391__3, 
                 inputs_391__2, inputs_391__1, inputs_391__0, inputs_392__15, 
                 inputs_392__14, inputs_392__13, inputs_392__12, inputs_392__11, 
                 inputs_392__10, inputs_392__9, inputs_392__8, inputs_392__7, 
                 inputs_392__6, inputs_392__5, inputs_392__4, inputs_392__3, 
                 inputs_392__2, inputs_392__1, inputs_392__0, inputs_393__15, 
                 inputs_393__14, inputs_393__13, inputs_393__12, inputs_393__11, 
                 inputs_393__10, inputs_393__9, inputs_393__8, inputs_393__7, 
                 inputs_393__6, inputs_393__5, inputs_393__4, inputs_393__3, 
                 inputs_393__2, inputs_393__1, inputs_393__0, inputs_394__15, 
                 inputs_394__14, inputs_394__13, inputs_394__12, inputs_394__11, 
                 inputs_394__10, inputs_394__9, inputs_394__8, inputs_394__7, 
                 inputs_394__6, inputs_394__5, inputs_394__4, inputs_394__3, 
                 inputs_394__2, inputs_394__1, inputs_394__0, inputs_395__15, 
                 inputs_395__14, inputs_395__13, inputs_395__12, inputs_395__11, 
                 inputs_395__10, inputs_395__9, inputs_395__8, inputs_395__7, 
                 inputs_395__6, inputs_395__5, inputs_395__4, inputs_395__3, 
                 inputs_395__2, inputs_395__1, inputs_395__0, inputs_396__15, 
                 inputs_396__14, inputs_396__13, inputs_396__12, inputs_396__11, 
                 inputs_396__10, inputs_396__9, inputs_396__8, inputs_396__7, 
                 inputs_396__6, inputs_396__5, inputs_396__4, inputs_396__3, 
                 inputs_396__2, inputs_396__1, inputs_396__0, inputs_397__15, 
                 inputs_397__14, inputs_397__13, inputs_397__12, inputs_397__11, 
                 inputs_397__10, inputs_397__9, inputs_397__8, inputs_397__7, 
                 inputs_397__6, inputs_397__5, inputs_397__4, inputs_397__3, 
                 inputs_397__2, inputs_397__1, inputs_397__0, inputs_398__15, 
                 inputs_398__14, inputs_398__13, inputs_398__12, inputs_398__11, 
                 inputs_398__10, inputs_398__9, inputs_398__8, inputs_398__7, 
                 inputs_398__6, inputs_398__5, inputs_398__4, inputs_398__3, 
                 inputs_398__2, inputs_398__1, inputs_398__0, inputs_399__15, 
                 inputs_399__14, inputs_399__13, inputs_399__12, inputs_399__11, 
                 inputs_399__10, inputs_399__9, inputs_399__8, inputs_399__7, 
                 inputs_399__6, inputs_399__5, inputs_399__4, inputs_399__3, 
                 inputs_399__2, inputs_399__1, inputs_399__0, inputs_400__15, 
                 inputs_400__14, inputs_400__13, inputs_400__12, inputs_400__11, 
                 inputs_400__10, inputs_400__9, inputs_400__8, inputs_400__7, 
                 inputs_400__6, inputs_400__5, inputs_400__4, inputs_400__3, 
                 inputs_400__2, inputs_400__1, inputs_400__0, inputs_401__15, 
                 inputs_401__14, inputs_401__13, inputs_401__12, inputs_401__11, 
                 inputs_401__10, inputs_401__9, inputs_401__8, inputs_401__7, 
                 inputs_401__6, inputs_401__5, inputs_401__4, inputs_401__3, 
                 inputs_401__2, inputs_401__1, inputs_401__0, inputs_402__15, 
                 inputs_402__14, inputs_402__13, inputs_402__12, inputs_402__11, 
                 inputs_402__10, inputs_402__9, inputs_402__8, inputs_402__7, 
                 inputs_402__6, inputs_402__5, inputs_402__4, inputs_402__3, 
                 inputs_402__2, inputs_402__1, inputs_402__0, inputs_403__15, 
                 inputs_403__14, inputs_403__13, inputs_403__12, inputs_403__11, 
                 inputs_403__10, inputs_403__9, inputs_403__8, inputs_403__7, 
                 inputs_403__6, inputs_403__5, inputs_403__4, inputs_403__3, 
                 inputs_403__2, inputs_403__1, inputs_403__0, inputs_404__15, 
                 inputs_404__14, inputs_404__13, inputs_404__12, inputs_404__11, 
                 inputs_404__10, inputs_404__9, inputs_404__8, inputs_404__7, 
                 inputs_404__6, inputs_404__5, inputs_404__4, inputs_404__3, 
                 inputs_404__2, inputs_404__1, inputs_404__0, inputs_405__15, 
                 inputs_405__14, inputs_405__13, inputs_405__12, inputs_405__11, 
                 inputs_405__10, inputs_405__9, inputs_405__8, inputs_405__7, 
                 inputs_405__6, inputs_405__5, inputs_405__4, inputs_405__3, 
                 inputs_405__2, inputs_405__1, inputs_405__0, inputs_406__15, 
                 inputs_406__14, inputs_406__13, inputs_406__12, inputs_406__11, 
                 inputs_406__10, inputs_406__9, inputs_406__8, inputs_406__7, 
                 inputs_406__6, inputs_406__5, inputs_406__4, inputs_406__3, 
                 inputs_406__2, inputs_406__1, inputs_406__0, inputs_407__15, 
                 inputs_407__14, inputs_407__13, inputs_407__12, inputs_407__11, 
                 inputs_407__10, inputs_407__9, inputs_407__8, inputs_407__7, 
                 inputs_407__6, inputs_407__5, inputs_407__4, inputs_407__3, 
                 inputs_407__2, inputs_407__1, inputs_407__0, inputs_408__15, 
                 inputs_408__14, inputs_408__13, inputs_408__12, inputs_408__11, 
                 inputs_408__10, inputs_408__9, inputs_408__8, inputs_408__7, 
                 inputs_408__6, inputs_408__5, inputs_408__4, inputs_408__3, 
                 inputs_408__2, inputs_408__1, inputs_408__0, inputs_409__15, 
                 inputs_409__14, inputs_409__13, inputs_409__12, inputs_409__11, 
                 inputs_409__10, inputs_409__9, inputs_409__8, inputs_409__7, 
                 inputs_409__6, inputs_409__5, inputs_409__4, inputs_409__3, 
                 inputs_409__2, inputs_409__1, inputs_409__0, inputs_410__15, 
                 inputs_410__14, inputs_410__13, inputs_410__12, inputs_410__11, 
                 inputs_410__10, inputs_410__9, inputs_410__8, inputs_410__7, 
                 inputs_410__6, inputs_410__5, inputs_410__4, inputs_410__3, 
                 inputs_410__2, inputs_410__1, inputs_410__0, inputs_411__15, 
                 inputs_411__14, inputs_411__13, inputs_411__12, inputs_411__11, 
                 inputs_411__10, inputs_411__9, inputs_411__8, inputs_411__7, 
                 inputs_411__6, inputs_411__5, inputs_411__4, inputs_411__3, 
                 inputs_411__2, inputs_411__1, inputs_411__0, inputs_412__15, 
                 inputs_412__14, inputs_412__13, inputs_412__12, inputs_412__11, 
                 inputs_412__10, inputs_412__9, inputs_412__8, inputs_412__7, 
                 inputs_412__6, inputs_412__5, inputs_412__4, inputs_412__3, 
                 inputs_412__2, inputs_412__1, inputs_412__0, inputs_413__15, 
                 inputs_413__14, inputs_413__13, inputs_413__12, inputs_413__11, 
                 inputs_413__10, inputs_413__9, inputs_413__8, inputs_413__7, 
                 inputs_413__6, inputs_413__5, inputs_413__4, inputs_413__3, 
                 inputs_413__2, inputs_413__1, inputs_413__0, inputs_414__15, 
                 inputs_414__14, inputs_414__13, inputs_414__12, inputs_414__11, 
                 inputs_414__10, inputs_414__9, inputs_414__8, inputs_414__7, 
                 inputs_414__6, inputs_414__5, inputs_414__4, inputs_414__3, 
                 inputs_414__2, inputs_414__1, inputs_414__0, inputs_415__15, 
                 inputs_415__14, inputs_415__13, inputs_415__12, inputs_415__11, 
                 inputs_415__10, inputs_415__9, inputs_415__8, inputs_415__7, 
                 inputs_415__6, inputs_415__5, inputs_415__4, inputs_415__3, 
                 inputs_415__2, inputs_415__1, inputs_415__0, inputs_416__15, 
                 inputs_416__14, inputs_416__13, inputs_416__12, inputs_416__11, 
                 inputs_416__10, inputs_416__9, inputs_416__8, inputs_416__7, 
                 inputs_416__6, inputs_416__5, inputs_416__4, inputs_416__3, 
                 inputs_416__2, inputs_416__1, inputs_416__0, inputs_417__15, 
                 inputs_417__14, inputs_417__13, inputs_417__12, inputs_417__11, 
                 inputs_417__10, inputs_417__9, inputs_417__8, inputs_417__7, 
                 inputs_417__6, inputs_417__5, inputs_417__4, inputs_417__3, 
                 inputs_417__2, inputs_417__1, inputs_417__0, inputs_418__15, 
                 inputs_418__14, inputs_418__13, inputs_418__12, inputs_418__11, 
                 inputs_418__10, inputs_418__9, inputs_418__8, inputs_418__7, 
                 inputs_418__6, inputs_418__5, inputs_418__4, inputs_418__3, 
                 inputs_418__2, inputs_418__1, inputs_418__0, inputs_419__15, 
                 inputs_419__14, inputs_419__13, inputs_419__12, inputs_419__11, 
                 inputs_419__10, inputs_419__9, inputs_419__8, inputs_419__7, 
                 inputs_419__6, inputs_419__5, inputs_419__4, inputs_419__3, 
                 inputs_419__2, inputs_419__1, inputs_419__0, inputs_420__15, 
                 inputs_420__14, inputs_420__13, inputs_420__12, inputs_420__11, 
                 inputs_420__10, inputs_420__9, inputs_420__8, inputs_420__7, 
                 inputs_420__6, inputs_420__5, inputs_420__4, inputs_420__3, 
                 inputs_420__2, inputs_420__1, inputs_420__0, inputs_421__15, 
                 inputs_421__14, inputs_421__13, inputs_421__12, inputs_421__11, 
                 inputs_421__10, inputs_421__9, inputs_421__8, inputs_421__7, 
                 inputs_421__6, inputs_421__5, inputs_421__4, inputs_421__3, 
                 inputs_421__2, inputs_421__1, inputs_421__0, inputs_422__15, 
                 inputs_422__14, inputs_422__13, inputs_422__12, inputs_422__11, 
                 inputs_422__10, inputs_422__9, inputs_422__8, inputs_422__7, 
                 inputs_422__6, inputs_422__5, inputs_422__4, inputs_422__3, 
                 inputs_422__2, inputs_422__1, inputs_422__0, inputs_423__15, 
                 inputs_423__14, inputs_423__13, inputs_423__12, inputs_423__11, 
                 inputs_423__10, inputs_423__9, inputs_423__8, inputs_423__7, 
                 inputs_423__6, inputs_423__5, inputs_423__4, inputs_423__3, 
                 inputs_423__2, inputs_423__1, inputs_423__0, inputs_424__15, 
                 inputs_424__14, inputs_424__13, inputs_424__12, inputs_424__11, 
                 inputs_424__10, inputs_424__9, inputs_424__8, inputs_424__7, 
                 inputs_424__6, inputs_424__5, inputs_424__4, inputs_424__3, 
                 inputs_424__2, inputs_424__1, inputs_424__0, inputs_425__15, 
                 inputs_425__14, inputs_425__13, inputs_425__12, inputs_425__11, 
                 inputs_425__10, inputs_425__9, inputs_425__8, inputs_425__7, 
                 inputs_425__6, inputs_425__5, inputs_425__4, inputs_425__3, 
                 inputs_425__2, inputs_425__1, inputs_425__0, inputs_426__15, 
                 inputs_426__14, inputs_426__13, inputs_426__12, inputs_426__11, 
                 inputs_426__10, inputs_426__9, inputs_426__8, inputs_426__7, 
                 inputs_426__6, inputs_426__5, inputs_426__4, inputs_426__3, 
                 inputs_426__2, inputs_426__1, inputs_426__0, inputs_427__15, 
                 inputs_427__14, inputs_427__13, inputs_427__12, inputs_427__11, 
                 inputs_427__10, inputs_427__9, inputs_427__8, inputs_427__7, 
                 inputs_427__6, inputs_427__5, inputs_427__4, inputs_427__3, 
                 inputs_427__2, inputs_427__1, inputs_427__0, inputs_428__15, 
                 inputs_428__14, inputs_428__13, inputs_428__12, inputs_428__11, 
                 inputs_428__10, inputs_428__9, inputs_428__8, inputs_428__7, 
                 inputs_428__6, inputs_428__5, inputs_428__4, inputs_428__3, 
                 inputs_428__2, inputs_428__1, inputs_428__0, inputs_429__15, 
                 inputs_429__14, inputs_429__13, inputs_429__12, inputs_429__11, 
                 inputs_429__10, inputs_429__9, inputs_429__8, inputs_429__7, 
                 inputs_429__6, inputs_429__5, inputs_429__4, inputs_429__3, 
                 inputs_429__2, inputs_429__1, inputs_429__0, inputs_430__15, 
                 inputs_430__14, inputs_430__13, inputs_430__12, inputs_430__11, 
                 inputs_430__10, inputs_430__9, inputs_430__8, inputs_430__7, 
                 inputs_430__6, inputs_430__5, inputs_430__4, inputs_430__3, 
                 inputs_430__2, inputs_430__1, inputs_430__0, inputs_431__15, 
                 inputs_431__14, inputs_431__13, inputs_431__12, inputs_431__11, 
                 inputs_431__10, inputs_431__9, inputs_431__8, inputs_431__7, 
                 inputs_431__6, inputs_431__5, inputs_431__4, inputs_431__3, 
                 inputs_431__2, inputs_431__1, inputs_431__0, inputs_432__15, 
                 inputs_432__14, inputs_432__13, inputs_432__12, inputs_432__11, 
                 inputs_432__10, inputs_432__9, inputs_432__8, inputs_432__7, 
                 inputs_432__6, inputs_432__5, inputs_432__4, inputs_432__3, 
                 inputs_432__2, inputs_432__1, inputs_432__0, inputs_433__15, 
                 inputs_433__14, inputs_433__13, inputs_433__12, inputs_433__11, 
                 inputs_433__10, inputs_433__9, inputs_433__8, inputs_433__7, 
                 inputs_433__6, inputs_433__5, inputs_433__4, inputs_433__3, 
                 inputs_433__2, inputs_433__1, inputs_433__0, inputs_434__15, 
                 inputs_434__14, inputs_434__13, inputs_434__12, inputs_434__11, 
                 inputs_434__10, inputs_434__9, inputs_434__8, inputs_434__7, 
                 inputs_434__6, inputs_434__5, inputs_434__4, inputs_434__3, 
                 inputs_434__2, inputs_434__1, inputs_434__0, inputs_435__15, 
                 inputs_435__14, inputs_435__13, inputs_435__12, inputs_435__11, 
                 inputs_435__10, inputs_435__9, inputs_435__8, inputs_435__7, 
                 inputs_435__6, inputs_435__5, inputs_435__4, inputs_435__3, 
                 inputs_435__2, inputs_435__1, inputs_435__0, inputs_436__15, 
                 inputs_436__14, inputs_436__13, inputs_436__12, inputs_436__11, 
                 inputs_436__10, inputs_436__9, inputs_436__8, inputs_436__7, 
                 inputs_436__6, inputs_436__5, inputs_436__4, inputs_436__3, 
                 inputs_436__2, inputs_436__1, inputs_436__0, inputs_437__15, 
                 inputs_437__14, inputs_437__13, inputs_437__12, inputs_437__11, 
                 inputs_437__10, inputs_437__9, inputs_437__8, inputs_437__7, 
                 inputs_437__6, inputs_437__5, inputs_437__4, inputs_437__3, 
                 inputs_437__2, inputs_437__1, inputs_437__0, inputs_438__15, 
                 inputs_438__14, inputs_438__13, inputs_438__12, inputs_438__11, 
                 inputs_438__10, inputs_438__9, inputs_438__8, inputs_438__7, 
                 inputs_438__6, inputs_438__5, inputs_438__4, inputs_438__3, 
                 inputs_438__2, inputs_438__1, inputs_438__0, inputs_439__15, 
                 inputs_439__14, inputs_439__13, inputs_439__12, inputs_439__11, 
                 inputs_439__10, inputs_439__9, inputs_439__8, inputs_439__7, 
                 inputs_439__6, inputs_439__5, inputs_439__4, inputs_439__3, 
                 inputs_439__2, inputs_439__1, inputs_439__0, inputs_440__15, 
                 inputs_440__14, inputs_440__13, inputs_440__12, inputs_440__11, 
                 inputs_440__10, inputs_440__9, inputs_440__8, inputs_440__7, 
                 inputs_440__6, inputs_440__5, inputs_440__4, inputs_440__3, 
                 inputs_440__2, inputs_440__1, inputs_440__0, inputs_441__15, 
                 inputs_441__14, inputs_441__13, inputs_441__12, inputs_441__11, 
                 inputs_441__10, inputs_441__9, inputs_441__8, inputs_441__7, 
                 inputs_441__6, inputs_441__5, inputs_441__4, inputs_441__3, 
                 inputs_441__2, inputs_441__1, inputs_441__0, inputs_442__15, 
                 inputs_442__14, inputs_442__13, inputs_442__12, inputs_442__11, 
                 inputs_442__10, inputs_442__9, inputs_442__8, inputs_442__7, 
                 inputs_442__6, inputs_442__5, inputs_442__4, inputs_442__3, 
                 inputs_442__2, inputs_442__1, inputs_442__0, inputs_443__15, 
                 inputs_443__14, inputs_443__13, inputs_443__12, inputs_443__11, 
                 inputs_443__10, inputs_443__9, inputs_443__8, inputs_443__7, 
                 inputs_443__6, inputs_443__5, inputs_443__4, inputs_443__3, 
                 inputs_443__2, inputs_443__1, inputs_443__0, inputs_444__15, 
                 inputs_444__14, inputs_444__13, inputs_444__12, inputs_444__11, 
                 inputs_444__10, inputs_444__9, inputs_444__8, inputs_444__7, 
                 inputs_444__6, inputs_444__5, inputs_444__4, inputs_444__3, 
                 inputs_444__2, inputs_444__1, inputs_444__0, inputs_445__15, 
                 inputs_445__14, inputs_445__13, inputs_445__12, inputs_445__11, 
                 inputs_445__10, inputs_445__9, inputs_445__8, inputs_445__7, 
                 inputs_445__6, inputs_445__5, inputs_445__4, inputs_445__3, 
                 inputs_445__2, inputs_445__1, inputs_445__0, inputs_446__15, 
                 inputs_446__14, inputs_446__13, inputs_446__12, inputs_446__11, 
                 inputs_446__10, inputs_446__9, inputs_446__8, inputs_446__7, 
                 inputs_446__6, inputs_446__5, inputs_446__4, inputs_446__3, 
                 inputs_446__2, inputs_446__1, inputs_446__0, inputs_447__15, 
                 inputs_447__14, inputs_447__13, inputs_447__12, inputs_447__11, 
                 inputs_447__10, inputs_447__9, inputs_447__8, inputs_447__7, 
                 inputs_447__6, inputs_447__5, inputs_447__4, inputs_447__3, 
                 inputs_447__2, inputs_447__1, inputs_447__0, inputs_448__15, 
                 inputs_448__14, inputs_448__13, inputs_448__12, inputs_448__11, 
                 inputs_448__10, inputs_448__9, inputs_448__8, inputs_448__7, 
                 inputs_448__6, inputs_448__5, inputs_448__4, inputs_448__3, 
                 inputs_448__2, inputs_448__1, inputs_448__0, inputs_449__15, 
                 inputs_449__14, inputs_449__13, inputs_449__12, inputs_449__11, 
                 inputs_449__10, inputs_449__9, inputs_449__8, inputs_449__7, 
                 inputs_449__6, inputs_449__5, inputs_449__4, inputs_449__3, 
                 inputs_449__2, inputs_449__1, inputs_449__0, inputs_450__15, 
                 inputs_450__14, inputs_450__13, inputs_450__12, inputs_450__11, 
                 inputs_450__10, inputs_450__9, inputs_450__8, inputs_450__7, 
                 inputs_450__6, inputs_450__5, inputs_450__4, inputs_450__3, 
                 inputs_450__2, inputs_450__1, inputs_450__0, inputs_451__15, 
                 inputs_451__14, inputs_451__13, inputs_451__12, inputs_451__11, 
                 inputs_451__10, inputs_451__9, inputs_451__8, inputs_451__7, 
                 inputs_451__6, inputs_451__5, inputs_451__4, inputs_451__3, 
                 inputs_451__2, inputs_451__1, inputs_451__0, inputs_452__15, 
                 inputs_452__14, inputs_452__13, inputs_452__12, inputs_452__11, 
                 inputs_452__10, inputs_452__9, inputs_452__8, inputs_452__7, 
                 inputs_452__6, inputs_452__5, inputs_452__4, inputs_452__3, 
                 inputs_452__2, inputs_452__1, inputs_452__0, inputs_453__15, 
                 inputs_453__14, inputs_453__13, inputs_453__12, inputs_453__11, 
                 inputs_453__10, inputs_453__9, inputs_453__8, inputs_453__7, 
                 inputs_453__6, inputs_453__5, inputs_453__4, inputs_453__3, 
                 inputs_453__2, inputs_453__1, inputs_453__0, inputs_454__15, 
                 inputs_454__14, inputs_454__13, inputs_454__12, inputs_454__11, 
                 inputs_454__10, inputs_454__9, inputs_454__8, inputs_454__7, 
                 inputs_454__6, inputs_454__5, inputs_454__4, inputs_454__3, 
                 inputs_454__2, inputs_454__1, inputs_454__0, inputs_455__15, 
                 inputs_455__14, inputs_455__13, inputs_455__12, inputs_455__11, 
                 inputs_455__10, inputs_455__9, inputs_455__8, inputs_455__7, 
                 inputs_455__6, inputs_455__5, inputs_455__4, inputs_455__3, 
                 inputs_455__2, inputs_455__1, inputs_455__0, inputs_456__15, 
                 inputs_456__14, inputs_456__13, inputs_456__12, inputs_456__11, 
                 inputs_456__10, inputs_456__9, inputs_456__8, inputs_456__7, 
                 inputs_456__6, inputs_456__5, inputs_456__4, inputs_456__3, 
                 inputs_456__2, inputs_456__1, inputs_456__0, inputs_457__15, 
                 inputs_457__14, inputs_457__13, inputs_457__12, inputs_457__11, 
                 inputs_457__10, inputs_457__9, inputs_457__8, inputs_457__7, 
                 inputs_457__6, inputs_457__5, inputs_457__4, inputs_457__3, 
                 inputs_457__2, inputs_457__1, inputs_457__0, inputs_458__15, 
                 inputs_458__14, inputs_458__13, inputs_458__12, inputs_458__11, 
                 inputs_458__10, inputs_458__9, inputs_458__8, inputs_458__7, 
                 inputs_458__6, inputs_458__5, inputs_458__4, inputs_458__3, 
                 inputs_458__2, inputs_458__1, inputs_458__0, inputs_459__15, 
                 inputs_459__14, inputs_459__13, inputs_459__12, inputs_459__11, 
                 inputs_459__10, inputs_459__9, inputs_459__8, inputs_459__7, 
                 inputs_459__6, inputs_459__5, inputs_459__4, inputs_459__3, 
                 inputs_459__2, inputs_459__1, inputs_459__0, inputs_460__15, 
                 inputs_460__14, inputs_460__13, inputs_460__12, inputs_460__11, 
                 inputs_460__10, inputs_460__9, inputs_460__8, inputs_460__7, 
                 inputs_460__6, inputs_460__5, inputs_460__4, inputs_460__3, 
                 inputs_460__2, inputs_460__1, inputs_460__0, inputs_461__15, 
                 inputs_461__14, inputs_461__13, inputs_461__12, inputs_461__11, 
                 inputs_461__10, inputs_461__9, inputs_461__8, inputs_461__7, 
                 inputs_461__6, inputs_461__5, inputs_461__4, inputs_461__3, 
                 inputs_461__2, inputs_461__1, inputs_461__0, inputs_462__15, 
                 inputs_462__14, inputs_462__13, inputs_462__12, inputs_462__11, 
                 inputs_462__10, inputs_462__9, inputs_462__8, inputs_462__7, 
                 inputs_462__6, inputs_462__5, inputs_462__4, inputs_462__3, 
                 inputs_462__2, inputs_462__1, inputs_462__0, inputs_463__15, 
                 inputs_463__14, inputs_463__13, inputs_463__12, inputs_463__11, 
                 inputs_463__10, inputs_463__9, inputs_463__8, inputs_463__7, 
                 inputs_463__6, inputs_463__5, inputs_463__4, inputs_463__3, 
                 inputs_463__2, inputs_463__1, inputs_463__0, inputs_464__15, 
                 inputs_464__14, inputs_464__13, inputs_464__12, inputs_464__11, 
                 inputs_464__10, inputs_464__9, inputs_464__8, inputs_464__7, 
                 inputs_464__6, inputs_464__5, inputs_464__4, inputs_464__3, 
                 inputs_464__2, inputs_464__1, inputs_464__0, inputs_465__15, 
                 inputs_465__14, inputs_465__13, inputs_465__12, inputs_465__11, 
                 inputs_465__10, inputs_465__9, inputs_465__8, inputs_465__7, 
                 inputs_465__6, inputs_465__5, inputs_465__4, inputs_465__3, 
                 inputs_465__2, inputs_465__1, inputs_465__0, inputs_466__15, 
                 inputs_466__14, inputs_466__13, inputs_466__12, inputs_466__11, 
                 inputs_466__10, inputs_466__9, inputs_466__8, inputs_466__7, 
                 inputs_466__6, inputs_466__5, inputs_466__4, inputs_466__3, 
                 inputs_466__2, inputs_466__1, inputs_466__0, inputs_467__15, 
                 inputs_467__14, inputs_467__13, inputs_467__12, inputs_467__11, 
                 inputs_467__10, inputs_467__9, inputs_467__8, inputs_467__7, 
                 inputs_467__6, inputs_467__5, inputs_467__4, inputs_467__3, 
                 inputs_467__2, inputs_467__1, inputs_467__0, inputs_468__15, 
                 inputs_468__14, inputs_468__13, inputs_468__12, inputs_468__11, 
                 inputs_468__10, inputs_468__9, inputs_468__8, inputs_468__7, 
                 inputs_468__6, inputs_468__5, inputs_468__4, inputs_468__3, 
                 inputs_468__2, inputs_468__1, inputs_468__0, inputs_469__15, 
                 inputs_469__14, inputs_469__13, inputs_469__12, inputs_469__11, 
                 inputs_469__10, inputs_469__9, inputs_469__8, inputs_469__7, 
                 inputs_469__6, inputs_469__5, inputs_469__4, inputs_469__3, 
                 inputs_469__2, inputs_469__1, inputs_469__0, inputs_470__15, 
                 inputs_470__14, inputs_470__13, inputs_470__12, inputs_470__11, 
                 inputs_470__10, inputs_470__9, inputs_470__8, inputs_470__7, 
                 inputs_470__6, inputs_470__5, inputs_470__4, inputs_470__3, 
                 inputs_470__2, inputs_470__1, inputs_470__0, inputs_471__15, 
                 inputs_471__14, inputs_471__13, inputs_471__12, inputs_471__11, 
                 inputs_471__10, inputs_471__9, inputs_471__8, inputs_471__7, 
                 inputs_471__6, inputs_471__5, inputs_471__4, inputs_471__3, 
                 inputs_471__2, inputs_471__1, inputs_471__0, inputs_472__15, 
                 inputs_472__14, inputs_472__13, inputs_472__12, inputs_472__11, 
                 inputs_472__10, inputs_472__9, inputs_472__8, inputs_472__7, 
                 inputs_472__6, inputs_472__5, inputs_472__4, inputs_472__3, 
                 inputs_472__2, inputs_472__1, inputs_472__0, inputs_473__15, 
                 inputs_473__14, inputs_473__13, inputs_473__12, inputs_473__11, 
                 inputs_473__10, inputs_473__9, inputs_473__8, inputs_473__7, 
                 inputs_473__6, inputs_473__5, inputs_473__4, inputs_473__3, 
                 inputs_473__2, inputs_473__1, inputs_473__0, inputs_474__15, 
                 inputs_474__14, inputs_474__13, inputs_474__12, inputs_474__11, 
                 inputs_474__10, inputs_474__9, inputs_474__8, inputs_474__7, 
                 inputs_474__6, inputs_474__5, inputs_474__4, inputs_474__3, 
                 inputs_474__2, inputs_474__1, inputs_474__0, inputs_475__15, 
                 inputs_475__14, inputs_475__13, inputs_475__12, inputs_475__11, 
                 inputs_475__10, inputs_475__9, inputs_475__8, inputs_475__7, 
                 inputs_475__6, inputs_475__5, inputs_475__4, inputs_475__3, 
                 inputs_475__2, inputs_475__1, inputs_475__0, inputs_476__15, 
                 inputs_476__14, inputs_476__13, inputs_476__12, inputs_476__11, 
                 inputs_476__10, inputs_476__9, inputs_476__8, inputs_476__7, 
                 inputs_476__6, inputs_476__5, inputs_476__4, inputs_476__3, 
                 inputs_476__2, inputs_476__1, inputs_476__0, inputs_477__15, 
                 inputs_477__14, inputs_477__13, inputs_477__12, inputs_477__11, 
                 inputs_477__10, inputs_477__9, inputs_477__8, inputs_477__7, 
                 inputs_477__6, inputs_477__5, inputs_477__4, inputs_477__3, 
                 inputs_477__2, inputs_477__1, inputs_477__0, inputs_478__15, 
                 inputs_478__14, inputs_478__13, inputs_478__12, inputs_478__11, 
                 inputs_478__10, inputs_478__9, inputs_478__8, inputs_478__7, 
                 inputs_478__6, inputs_478__5, inputs_478__4, inputs_478__3, 
                 inputs_478__2, inputs_478__1, inputs_478__0, inputs_479__15, 
                 inputs_479__14, inputs_479__13, inputs_479__12, inputs_479__11, 
                 inputs_479__10, inputs_479__9, inputs_479__8, inputs_479__7, 
                 inputs_479__6, inputs_479__5, inputs_479__4, inputs_479__3, 
                 inputs_479__2, inputs_479__1, inputs_479__0, inputs_480__15, 
                 inputs_480__14, inputs_480__13, inputs_480__12, inputs_480__11, 
                 inputs_480__10, inputs_480__9, inputs_480__8, inputs_480__7, 
                 inputs_480__6, inputs_480__5, inputs_480__4, inputs_480__3, 
                 inputs_480__2, inputs_480__1, inputs_480__0, inputs_481__15, 
                 inputs_481__14, inputs_481__13, inputs_481__12, inputs_481__11, 
                 inputs_481__10, inputs_481__9, inputs_481__8, inputs_481__7, 
                 inputs_481__6, inputs_481__5, inputs_481__4, inputs_481__3, 
                 inputs_481__2, inputs_481__1, inputs_481__0, inputs_482__15, 
                 inputs_482__14, inputs_482__13, inputs_482__12, inputs_482__11, 
                 inputs_482__10, inputs_482__9, inputs_482__8, inputs_482__7, 
                 inputs_482__6, inputs_482__5, inputs_482__4, inputs_482__3, 
                 inputs_482__2, inputs_482__1, inputs_482__0, inputs_483__15, 
                 inputs_483__14, inputs_483__13, inputs_483__12, inputs_483__11, 
                 inputs_483__10, inputs_483__9, inputs_483__8, inputs_483__7, 
                 inputs_483__6, inputs_483__5, inputs_483__4, inputs_483__3, 
                 inputs_483__2, inputs_483__1, inputs_483__0, inputs_484__15, 
                 inputs_484__14, inputs_484__13, inputs_484__12, inputs_484__11, 
                 inputs_484__10, inputs_484__9, inputs_484__8, inputs_484__7, 
                 inputs_484__6, inputs_484__5, inputs_484__4, inputs_484__3, 
                 inputs_484__2, inputs_484__1, inputs_484__0, inputs_485__15, 
                 inputs_485__14, inputs_485__13, inputs_485__12, inputs_485__11, 
                 inputs_485__10, inputs_485__9, inputs_485__8, inputs_485__7, 
                 inputs_485__6, inputs_485__5, inputs_485__4, inputs_485__3, 
                 inputs_485__2, inputs_485__1, inputs_485__0, inputs_486__15, 
                 inputs_486__14, inputs_486__13, inputs_486__12, inputs_486__11, 
                 inputs_486__10, inputs_486__9, inputs_486__8, inputs_486__7, 
                 inputs_486__6, inputs_486__5, inputs_486__4, inputs_486__3, 
                 inputs_486__2, inputs_486__1, inputs_486__0, inputs_487__15, 
                 inputs_487__14, inputs_487__13, inputs_487__12, inputs_487__11, 
                 inputs_487__10, inputs_487__9, inputs_487__8, inputs_487__7, 
                 inputs_487__6, inputs_487__5, inputs_487__4, inputs_487__3, 
                 inputs_487__2, inputs_487__1, inputs_487__0, inputs_488__15, 
                 inputs_488__14, inputs_488__13, inputs_488__12, inputs_488__11, 
                 inputs_488__10, inputs_488__9, inputs_488__8, inputs_488__7, 
                 inputs_488__6, inputs_488__5, inputs_488__4, inputs_488__3, 
                 inputs_488__2, inputs_488__1, inputs_488__0, inputs_489__15, 
                 inputs_489__14, inputs_489__13, inputs_489__12, inputs_489__11, 
                 inputs_489__10, inputs_489__9, inputs_489__8, inputs_489__7, 
                 inputs_489__6, inputs_489__5, inputs_489__4, inputs_489__3, 
                 inputs_489__2, inputs_489__1, inputs_489__0, inputs_490__15, 
                 inputs_490__14, inputs_490__13, inputs_490__12, inputs_490__11, 
                 inputs_490__10, inputs_490__9, inputs_490__8, inputs_490__7, 
                 inputs_490__6, inputs_490__5, inputs_490__4, inputs_490__3, 
                 inputs_490__2, inputs_490__1, inputs_490__0, inputs_491__15, 
                 inputs_491__14, inputs_491__13, inputs_491__12, inputs_491__11, 
                 inputs_491__10, inputs_491__9, inputs_491__8, inputs_491__7, 
                 inputs_491__6, inputs_491__5, inputs_491__4, inputs_491__3, 
                 inputs_491__2, inputs_491__1, inputs_491__0, inputs_492__15, 
                 inputs_492__14, inputs_492__13, inputs_492__12, inputs_492__11, 
                 inputs_492__10, inputs_492__9, inputs_492__8, inputs_492__7, 
                 inputs_492__6, inputs_492__5, inputs_492__4, inputs_492__3, 
                 inputs_492__2, inputs_492__1, inputs_492__0, inputs_493__15, 
                 inputs_493__14, inputs_493__13, inputs_493__12, inputs_493__11, 
                 inputs_493__10, inputs_493__9, inputs_493__8, inputs_493__7, 
                 inputs_493__6, inputs_493__5, inputs_493__4, inputs_493__3, 
                 inputs_493__2, inputs_493__1, inputs_493__0, inputs_494__15, 
                 inputs_494__14, inputs_494__13, inputs_494__12, inputs_494__11, 
                 inputs_494__10, inputs_494__9, inputs_494__8, inputs_494__7, 
                 inputs_494__6, inputs_494__5, inputs_494__4, inputs_494__3, 
                 inputs_494__2, inputs_494__1, inputs_494__0, inputs_495__15, 
                 inputs_495__14, inputs_495__13, inputs_495__12, inputs_495__11, 
                 inputs_495__10, inputs_495__9, inputs_495__8, inputs_495__7, 
                 inputs_495__6, inputs_495__5, inputs_495__4, inputs_495__3, 
                 inputs_495__2, inputs_495__1, inputs_495__0, inputs_496__15, 
                 inputs_496__14, inputs_496__13, inputs_496__12, inputs_496__11, 
                 inputs_496__10, inputs_496__9, inputs_496__8, inputs_496__7, 
                 inputs_496__6, inputs_496__5, inputs_496__4, inputs_496__3, 
                 inputs_496__2, inputs_496__1, inputs_496__0, inputs_497__15, 
                 inputs_497__14, inputs_497__13, inputs_497__12, inputs_497__11, 
                 inputs_497__10, inputs_497__9, inputs_497__8, inputs_497__7, 
                 inputs_497__6, inputs_497__5, inputs_497__4, inputs_497__3, 
                 inputs_497__2, inputs_497__1, inputs_497__0, inputs_498__15, 
                 inputs_498__14, inputs_498__13, inputs_498__12, inputs_498__11, 
                 inputs_498__10, inputs_498__9, inputs_498__8, inputs_498__7, 
                 inputs_498__6, inputs_498__5, inputs_498__4, inputs_498__3, 
                 inputs_498__2, inputs_498__1, inputs_498__0, inputs_499__15, 
                 inputs_499__14, inputs_499__13, inputs_499__12, inputs_499__11, 
                 inputs_499__10, inputs_499__9, inputs_499__8, inputs_499__7, 
                 inputs_499__6, inputs_499__5, inputs_499__4, inputs_499__3, 
                 inputs_499__2, inputs_499__1, inputs_499__0, inputs_500__15, 
                 inputs_500__14, inputs_500__13, inputs_500__12, inputs_500__11, 
                 inputs_500__10, inputs_500__9, inputs_500__8, inputs_500__7, 
                 inputs_500__6, inputs_500__5, inputs_500__4, inputs_500__3, 
                 inputs_500__2, inputs_500__1, inputs_500__0, inputs_501__15, 
                 inputs_501__14, inputs_501__13, inputs_501__12, inputs_501__11, 
                 inputs_501__10, inputs_501__9, inputs_501__8, inputs_501__7, 
                 inputs_501__6, inputs_501__5, inputs_501__4, inputs_501__3, 
                 inputs_501__2, inputs_501__1, inputs_501__0, inputs_502__15, 
                 inputs_502__14, inputs_502__13, inputs_502__12, inputs_502__11, 
                 inputs_502__10, inputs_502__9, inputs_502__8, inputs_502__7, 
                 inputs_502__6, inputs_502__5, inputs_502__4, inputs_502__3, 
                 inputs_502__2, inputs_502__1, inputs_502__0, inputs_503__15, 
                 inputs_503__14, inputs_503__13, inputs_503__12, inputs_503__11, 
                 inputs_503__10, inputs_503__9, inputs_503__8, inputs_503__7, 
                 inputs_503__6, inputs_503__5, inputs_503__4, inputs_503__3, 
                 inputs_503__2, inputs_503__1, inputs_503__0, inputs_504__15, 
                 inputs_504__14, inputs_504__13, inputs_504__12, inputs_504__11, 
                 inputs_504__10, inputs_504__9, inputs_504__8, inputs_504__7, 
                 inputs_504__6, inputs_504__5, inputs_504__4, inputs_504__3, 
                 inputs_504__2, inputs_504__1, inputs_504__0, inputs_505__15, 
                 inputs_505__14, inputs_505__13, inputs_505__12, inputs_505__11, 
                 inputs_505__10, inputs_505__9, inputs_505__8, inputs_505__7, 
                 inputs_505__6, inputs_505__5, inputs_505__4, inputs_505__3, 
                 inputs_505__2, inputs_505__1, inputs_505__0, inputs_506__15, 
                 inputs_506__14, inputs_506__13, inputs_506__12, inputs_506__11, 
                 inputs_506__10, inputs_506__9, inputs_506__8, inputs_506__7, 
                 inputs_506__6, inputs_506__5, inputs_506__4, inputs_506__3, 
                 inputs_506__2, inputs_506__1, inputs_506__0, inputs_507__15, 
                 inputs_507__14, inputs_507__13, inputs_507__12, inputs_507__11, 
                 inputs_507__10, inputs_507__9, inputs_507__8, inputs_507__7, 
                 inputs_507__6, inputs_507__5, inputs_507__4, inputs_507__3, 
                 inputs_507__2, inputs_507__1, inputs_507__0, inputs_508__15, 
                 inputs_508__14, inputs_508__13, inputs_508__12, inputs_508__11, 
                 inputs_508__10, inputs_508__9, inputs_508__8, inputs_508__7, 
                 inputs_508__6, inputs_508__5, inputs_508__4, inputs_508__3, 
                 inputs_508__2, inputs_508__1, inputs_508__0, inputs_509__15, 
                 inputs_509__14, inputs_509__13, inputs_509__12, inputs_509__11, 
                 inputs_509__10, inputs_509__9, inputs_509__8, inputs_509__7, 
                 inputs_509__6, inputs_509__5, inputs_509__4, inputs_509__3, 
                 inputs_509__2, inputs_509__1, inputs_509__0, inputs_510__15, 
                 inputs_510__14, inputs_510__13, inputs_510__12, inputs_510__11, 
                 inputs_510__10, inputs_510__9, inputs_510__8, inputs_510__7, 
                 inputs_510__6, inputs_510__5, inputs_510__4, inputs_510__3, 
                 inputs_510__2, inputs_510__1, inputs_510__0, inputs_511__15, 
                 inputs_511__14, inputs_511__13, inputs_511__12, inputs_511__11, 
                 inputs_511__10, inputs_511__9, inputs_511__8, inputs_511__7, 
                 inputs_511__6, inputs_511__5, inputs_511__4, inputs_511__3, 
                 inputs_511__2, inputs_511__1, inputs_511__0, selectionLines, 
                 \output  ) ;

    input inputs_0__15 ;
    input inputs_0__14 ;
    input inputs_0__13 ;
    input inputs_0__12 ;
    input inputs_0__11 ;
    input inputs_0__10 ;
    input inputs_0__9 ;
    input inputs_0__8 ;
    input inputs_0__7 ;
    input inputs_0__6 ;
    input inputs_0__5 ;
    input inputs_0__4 ;
    input inputs_0__3 ;
    input inputs_0__2 ;
    input inputs_0__1 ;
    input inputs_0__0 ;
    input inputs_1__15 ;
    input inputs_1__14 ;
    input inputs_1__13 ;
    input inputs_1__12 ;
    input inputs_1__11 ;
    input inputs_1__10 ;
    input inputs_1__9 ;
    input inputs_1__8 ;
    input inputs_1__7 ;
    input inputs_1__6 ;
    input inputs_1__5 ;
    input inputs_1__4 ;
    input inputs_1__3 ;
    input inputs_1__2 ;
    input inputs_1__1 ;
    input inputs_1__0 ;
    input inputs_2__15 ;
    input inputs_2__14 ;
    input inputs_2__13 ;
    input inputs_2__12 ;
    input inputs_2__11 ;
    input inputs_2__10 ;
    input inputs_2__9 ;
    input inputs_2__8 ;
    input inputs_2__7 ;
    input inputs_2__6 ;
    input inputs_2__5 ;
    input inputs_2__4 ;
    input inputs_2__3 ;
    input inputs_2__2 ;
    input inputs_2__1 ;
    input inputs_2__0 ;
    input inputs_3__15 ;
    input inputs_3__14 ;
    input inputs_3__13 ;
    input inputs_3__12 ;
    input inputs_3__11 ;
    input inputs_3__10 ;
    input inputs_3__9 ;
    input inputs_3__8 ;
    input inputs_3__7 ;
    input inputs_3__6 ;
    input inputs_3__5 ;
    input inputs_3__4 ;
    input inputs_3__3 ;
    input inputs_3__2 ;
    input inputs_3__1 ;
    input inputs_3__0 ;
    input inputs_4__15 ;
    input inputs_4__14 ;
    input inputs_4__13 ;
    input inputs_4__12 ;
    input inputs_4__11 ;
    input inputs_4__10 ;
    input inputs_4__9 ;
    input inputs_4__8 ;
    input inputs_4__7 ;
    input inputs_4__6 ;
    input inputs_4__5 ;
    input inputs_4__4 ;
    input inputs_4__3 ;
    input inputs_4__2 ;
    input inputs_4__1 ;
    input inputs_4__0 ;
    input inputs_5__15 ;
    input inputs_5__14 ;
    input inputs_5__13 ;
    input inputs_5__12 ;
    input inputs_5__11 ;
    input inputs_5__10 ;
    input inputs_5__9 ;
    input inputs_5__8 ;
    input inputs_5__7 ;
    input inputs_5__6 ;
    input inputs_5__5 ;
    input inputs_5__4 ;
    input inputs_5__3 ;
    input inputs_5__2 ;
    input inputs_5__1 ;
    input inputs_5__0 ;
    input inputs_6__15 ;
    input inputs_6__14 ;
    input inputs_6__13 ;
    input inputs_6__12 ;
    input inputs_6__11 ;
    input inputs_6__10 ;
    input inputs_6__9 ;
    input inputs_6__8 ;
    input inputs_6__7 ;
    input inputs_6__6 ;
    input inputs_6__5 ;
    input inputs_6__4 ;
    input inputs_6__3 ;
    input inputs_6__2 ;
    input inputs_6__1 ;
    input inputs_6__0 ;
    input inputs_7__15 ;
    input inputs_7__14 ;
    input inputs_7__13 ;
    input inputs_7__12 ;
    input inputs_7__11 ;
    input inputs_7__10 ;
    input inputs_7__9 ;
    input inputs_7__8 ;
    input inputs_7__7 ;
    input inputs_7__6 ;
    input inputs_7__5 ;
    input inputs_7__4 ;
    input inputs_7__3 ;
    input inputs_7__2 ;
    input inputs_7__1 ;
    input inputs_7__0 ;
    input inputs_8__15 ;
    input inputs_8__14 ;
    input inputs_8__13 ;
    input inputs_8__12 ;
    input inputs_8__11 ;
    input inputs_8__10 ;
    input inputs_8__9 ;
    input inputs_8__8 ;
    input inputs_8__7 ;
    input inputs_8__6 ;
    input inputs_8__5 ;
    input inputs_8__4 ;
    input inputs_8__3 ;
    input inputs_8__2 ;
    input inputs_8__1 ;
    input inputs_8__0 ;
    input inputs_9__15 ;
    input inputs_9__14 ;
    input inputs_9__13 ;
    input inputs_9__12 ;
    input inputs_9__11 ;
    input inputs_9__10 ;
    input inputs_9__9 ;
    input inputs_9__8 ;
    input inputs_9__7 ;
    input inputs_9__6 ;
    input inputs_9__5 ;
    input inputs_9__4 ;
    input inputs_9__3 ;
    input inputs_9__2 ;
    input inputs_9__1 ;
    input inputs_9__0 ;
    input inputs_10__15 ;
    input inputs_10__14 ;
    input inputs_10__13 ;
    input inputs_10__12 ;
    input inputs_10__11 ;
    input inputs_10__10 ;
    input inputs_10__9 ;
    input inputs_10__8 ;
    input inputs_10__7 ;
    input inputs_10__6 ;
    input inputs_10__5 ;
    input inputs_10__4 ;
    input inputs_10__3 ;
    input inputs_10__2 ;
    input inputs_10__1 ;
    input inputs_10__0 ;
    input inputs_11__15 ;
    input inputs_11__14 ;
    input inputs_11__13 ;
    input inputs_11__12 ;
    input inputs_11__11 ;
    input inputs_11__10 ;
    input inputs_11__9 ;
    input inputs_11__8 ;
    input inputs_11__7 ;
    input inputs_11__6 ;
    input inputs_11__5 ;
    input inputs_11__4 ;
    input inputs_11__3 ;
    input inputs_11__2 ;
    input inputs_11__1 ;
    input inputs_11__0 ;
    input inputs_12__15 ;
    input inputs_12__14 ;
    input inputs_12__13 ;
    input inputs_12__12 ;
    input inputs_12__11 ;
    input inputs_12__10 ;
    input inputs_12__9 ;
    input inputs_12__8 ;
    input inputs_12__7 ;
    input inputs_12__6 ;
    input inputs_12__5 ;
    input inputs_12__4 ;
    input inputs_12__3 ;
    input inputs_12__2 ;
    input inputs_12__1 ;
    input inputs_12__0 ;
    input inputs_13__15 ;
    input inputs_13__14 ;
    input inputs_13__13 ;
    input inputs_13__12 ;
    input inputs_13__11 ;
    input inputs_13__10 ;
    input inputs_13__9 ;
    input inputs_13__8 ;
    input inputs_13__7 ;
    input inputs_13__6 ;
    input inputs_13__5 ;
    input inputs_13__4 ;
    input inputs_13__3 ;
    input inputs_13__2 ;
    input inputs_13__1 ;
    input inputs_13__0 ;
    input inputs_14__15 ;
    input inputs_14__14 ;
    input inputs_14__13 ;
    input inputs_14__12 ;
    input inputs_14__11 ;
    input inputs_14__10 ;
    input inputs_14__9 ;
    input inputs_14__8 ;
    input inputs_14__7 ;
    input inputs_14__6 ;
    input inputs_14__5 ;
    input inputs_14__4 ;
    input inputs_14__3 ;
    input inputs_14__2 ;
    input inputs_14__1 ;
    input inputs_14__0 ;
    input inputs_15__15 ;
    input inputs_15__14 ;
    input inputs_15__13 ;
    input inputs_15__12 ;
    input inputs_15__11 ;
    input inputs_15__10 ;
    input inputs_15__9 ;
    input inputs_15__8 ;
    input inputs_15__7 ;
    input inputs_15__6 ;
    input inputs_15__5 ;
    input inputs_15__4 ;
    input inputs_15__3 ;
    input inputs_15__2 ;
    input inputs_15__1 ;
    input inputs_15__0 ;
    input inputs_16__15 ;
    input inputs_16__14 ;
    input inputs_16__13 ;
    input inputs_16__12 ;
    input inputs_16__11 ;
    input inputs_16__10 ;
    input inputs_16__9 ;
    input inputs_16__8 ;
    input inputs_16__7 ;
    input inputs_16__6 ;
    input inputs_16__5 ;
    input inputs_16__4 ;
    input inputs_16__3 ;
    input inputs_16__2 ;
    input inputs_16__1 ;
    input inputs_16__0 ;
    input inputs_17__15 ;
    input inputs_17__14 ;
    input inputs_17__13 ;
    input inputs_17__12 ;
    input inputs_17__11 ;
    input inputs_17__10 ;
    input inputs_17__9 ;
    input inputs_17__8 ;
    input inputs_17__7 ;
    input inputs_17__6 ;
    input inputs_17__5 ;
    input inputs_17__4 ;
    input inputs_17__3 ;
    input inputs_17__2 ;
    input inputs_17__1 ;
    input inputs_17__0 ;
    input inputs_18__15 ;
    input inputs_18__14 ;
    input inputs_18__13 ;
    input inputs_18__12 ;
    input inputs_18__11 ;
    input inputs_18__10 ;
    input inputs_18__9 ;
    input inputs_18__8 ;
    input inputs_18__7 ;
    input inputs_18__6 ;
    input inputs_18__5 ;
    input inputs_18__4 ;
    input inputs_18__3 ;
    input inputs_18__2 ;
    input inputs_18__1 ;
    input inputs_18__0 ;
    input inputs_19__15 ;
    input inputs_19__14 ;
    input inputs_19__13 ;
    input inputs_19__12 ;
    input inputs_19__11 ;
    input inputs_19__10 ;
    input inputs_19__9 ;
    input inputs_19__8 ;
    input inputs_19__7 ;
    input inputs_19__6 ;
    input inputs_19__5 ;
    input inputs_19__4 ;
    input inputs_19__3 ;
    input inputs_19__2 ;
    input inputs_19__1 ;
    input inputs_19__0 ;
    input inputs_20__15 ;
    input inputs_20__14 ;
    input inputs_20__13 ;
    input inputs_20__12 ;
    input inputs_20__11 ;
    input inputs_20__10 ;
    input inputs_20__9 ;
    input inputs_20__8 ;
    input inputs_20__7 ;
    input inputs_20__6 ;
    input inputs_20__5 ;
    input inputs_20__4 ;
    input inputs_20__3 ;
    input inputs_20__2 ;
    input inputs_20__1 ;
    input inputs_20__0 ;
    input inputs_21__15 ;
    input inputs_21__14 ;
    input inputs_21__13 ;
    input inputs_21__12 ;
    input inputs_21__11 ;
    input inputs_21__10 ;
    input inputs_21__9 ;
    input inputs_21__8 ;
    input inputs_21__7 ;
    input inputs_21__6 ;
    input inputs_21__5 ;
    input inputs_21__4 ;
    input inputs_21__3 ;
    input inputs_21__2 ;
    input inputs_21__1 ;
    input inputs_21__0 ;
    input inputs_22__15 ;
    input inputs_22__14 ;
    input inputs_22__13 ;
    input inputs_22__12 ;
    input inputs_22__11 ;
    input inputs_22__10 ;
    input inputs_22__9 ;
    input inputs_22__8 ;
    input inputs_22__7 ;
    input inputs_22__6 ;
    input inputs_22__5 ;
    input inputs_22__4 ;
    input inputs_22__3 ;
    input inputs_22__2 ;
    input inputs_22__1 ;
    input inputs_22__0 ;
    input inputs_23__15 ;
    input inputs_23__14 ;
    input inputs_23__13 ;
    input inputs_23__12 ;
    input inputs_23__11 ;
    input inputs_23__10 ;
    input inputs_23__9 ;
    input inputs_23__8 ;
    input inputs_23__7 ;
    input inputs_23__6 ;
    input inputs_23__5 ;
    input inputs_23__4 ;
    input inputs_23__3 ;
    input inputs_23__2 ;
    input inputs_23__1 ;
    input inputs_23__0 ;
    input inputs_24__15 ;
    input inputs_24__14 ;
    input inputs_24__13 ;
    input inputs_24__12 ;
    input inputs_24__11 ;
    input inputs_24__10 ;
    input inputs_24__9 ;
    input inputs_24__8 ;
    input inputs_24__7 ;
    input inputs_24__6 ;
    input inputs_24__5 ;
    input inputs_24__4 ;
    input inputs_24__3 ;
    input inputs_24__2 ;
    input inputs_24__1 ;
    input inputs_24__0 ;
    input inputs_25__15 ;
    input inputs_25__14 ;
    input inputs_25__13 ;
    input inputs_25__12 ;
    input inputs_25__11 ;
    input inputs_25__10 ;
    input inputs_25__9 ;
    input inputs_25__8 ;
    input inputs_25__7 ;
    input inputs_25__6 ;
    input inputs_25__5 ;
    input inputs_25__4 ;
    input inputs_25__3 ;
    input inputs_25__2 ;
    input inputs_25__1 ;
    input inputs_25__0 ;
    input inputs_26__15 ;
    input inputs_26__14 ;
    input inputs_26__13 ;
    input inputs_26__12 ;
    input inputs_26__11 ;
    input inputs_26__10 ;
    input inputs_26__9 ;
    input inputs_26__8 ;
    input inputs_26__7 ;
    input inputs_26__6 ;
    input inputs_26__5 ;
    input inputs_26__4 ;
    input inputs_26__3 ;
    input inputs_26__2 ;
    input inputs_26__1 ;
    input inputs_26__0 ;
    input inputs_27__15 ;
    input inputs_27__14 ;
    input inputs_27__13 ;
    input inputs_27__12 ;
    input inputs_27__11 ;
    input inputs_27__10 ;
    input inputs_27__9 ;
    input inputs_27__8 ;
    input inputs_27__7 ;
    input inputs_27__6 ;
    input inputs_27__5 ;
    input inputs_27__4 ;
    input inputs_27__3 ;
    input inputs_27__2 ;
    input inputs_27__1 ;
    input inputs_27__0 ;
    input inputs_28__15 ;
    input inputs_28__14 ;
    input inputs_28__13 ;
    input inputs_28__12 ;
    input inputs_28__11 ;
    input inputs_28__10 ;
    input inputs_28__9 ;
    input inputs_28__8 ;
    input inputs_28__7 ;
    input inputs_28__6 ;
    input inputs_28__5 ;
    input inputs_28__4 ;
    input inputs_28__3 ;
    input inputs_28__2 ;
    input inputs_28__1 ;
    input inputs_28__0 ;
    input inputs_29__15 ;
    input inputs_29__14 ;
    input inputs_29__13 ;
    input inputs_29__12 ;
    input inputs_29__11 ;
    input inputs_29__10 ;
    input inputs_29__9 ;
    input inputs_29__8 ;
    input inputs_29__7 ;
    input inputs_29__6 ;
    input inputs_29__5 ;
    input inputs_29__4 ;
    input inputs_29__3 ;
    input inputs_29__2 ;
    input inputs_29__1 ;
    input inputs_29__0 ;
    input inputs_30__15 ;
    input inputs_30__14 ;
    input inputs_30__13 ;
    input inputs_30__12 ;
    input inputs_30__11 ;
    input inputs_30__10 ;
    input inputs_30__9 ;
    input inputs_30__8 ;
    input inputs_30__7 ;
    input inputs_30__6 ;
    input inputs_30__5 ;
    input inputs_30__4 ;
    input inputs_30__3 ;
    input inputs_30__2 ;
    input inputs_30__1 ;
    input inputs_30__0 ;
    input inputs_31__15 ;
    input inputs_31__14 ;
    input inputs_31__13 ;
    input inputs_31__12 ;
    input inputs_31__11 ;
    input inputs_31__10 ;
    input inputs_31__9 ;
    input inputs_31__8 ;
    input inputs_31__7 ;
    input inputs_31__6 ;
    input inputs_31__5 ;
    input inputs_31__4 ;
    input inputs_31__3 ;
    input inputs_31__2 ;
    input inputs_31__1 ;
    input inputs_31__0 ;
    input inputs_32__15 ;
    input inputs_32__14 ;
    input inputs_32__13 ;
    input inputs_32__12 ;
    input inputs_32__11 ;
    input inputs_32__10 ;
    input inputs_32__9 ;
    input inputs_32__8 ;
    input inputs_32__7 ;
    input inputs_32__6 ;
    input inputs_32__5 ;
    input inputs_32__4 ;
    input inputs_32__3 ;
    input inputs_32__2 ;
    input inputs_32__1 ;
    input inputs_32__0 ;
    input inputs_33__15 ;
    input inputs_33__14 ;
    input inputs_33__13 ;
    input inputs_33__12 ;
    input inputs_33__11 ;
    input inputs_33__10 ;
    input inputs_33__9 ;
    input inputs_33__8 ;
    input inputs_33__7 ;
    input inputs_33__6 ;
    input inputs_33__5 ;
    input inputs_33__4 ;
    input inputs_33__3 ;
    input inputs_33__2 ;
    input inputs_33__1 ;
    input inputs_33__0 ;
    input inputs_34__15 ;
    input inputs_34__14 ;
    input inputs_34__13 ;
    input inputs_34__12 ;
    input inputs_34__11 ;
    input inputs_34__10 ;
    input inputs_34__9 ;
    input inputs_34__8 ;
    input inputs_34__7 ;
    input inputs_34__6 ;
    input inputs_34__5 ;
    input inputs_34__4 ;
    input inputs_34__3 ;
    input inputs_34__2 ;
    input inputs_34__1 ;
    input inputs_34__0 ;
    input inputs_35__15 ;
    input inputs_35__14 ;
    input inputs_35__13 ;
    input inputs_35__12 ;
    input inputs_35__11 ;
    input inputs_35__10 ;
    input inputs_35__9 ;
    input inputs_35__8 ;
    input inputs_35__7 ;
    input inputs_35__6 ;
    input inputs_35__5 ;
    input inputs_35__4 ;
    input inputs_35__3 ;
    input inputs_35__2 ;
    input inputs_35__1 ;
    input inputs_35__0 ;
    input inputs_36__15 ;
    input inputs_36__14 ;
    input inputs_36__13 ;
    input inputs_36__12 ;
    input inputs_36__11 ;
    input inputs_36__10 ;
    input inputs_36__9 ;
    input inputs_36__8 ;
    input inputs_36__7 ;
    input inputs_36__6 ;
    input inputs_36__5 ;
    input inputs_36__4 ;
    input inputs_36__3 ;
    input inputs_36__2 ;
    input inputs_36__1 ;
    input inputs_36__0 ;
    input inputs_37__15 ;
    input inputs_37__14 ;
    input inputs_37__13 ;
    input inputs_37__12 ;
    input inputs_37__11 ;
    input inputs_37__10 ;
    input inputs_37__9 ;
    input inputs_37__8 ;
    input inputs_37__7 ;
    input inputs_37__6 ;
    input inputs_37__5 ;
    input inputs_37__4 ;
    input inputs_37__3 ;
    input inputs_37__2 ;
    input inputs_37__1 ;
    input inputs_37__0 ;
    input inputs_38__15 ;
    input inputs_38__14 ;
    input inputs_38__13 ;
    input inputs_38__12 ;
    input inputs_38__11 ;
    input inputs_38__10 ;
    input inputs_38__9 ;
    input inputs_38__8 ;
    input inputs_38__7 ;
    input inputs_38__6 ;
    input inputs_38__5 ;
    input inputs_38__4 ;
    input inputs_38__3 ;
    input inputs_38__2 ;
    input inputs_38__1 ;
    input inputs_38__0 ;
    input inputs_39__15 ;
    input inputs_39__14 ;
    input inputs_39__13 ;
    input inputs_39__12 ;
    input inputs_39__11 ;
    input inputs_39__10 ;
    input inputs_39__9 ;
    input inputs_39__8 ;
    input inputs_39__7 ;
    input inputs_39__6 ;
    input inputs_39__5 ;
    input inputs_39__4 ;
    input inputs_39__3 ;
    input inputs_39__2 ;
    input inputs_39__1 ;
    input inputs_39__0 ;
    input inputs_40__15 ;
    input inputs_40__14 ;
    input inputs_40__13 ;
    input inputs_40__12 ;
    input inputs_40__11 ;
    input inputs_40__10 ;
    input inputs_40__9 ;
    input inputs_40__8 ;
    input inputs_40__7 ;
    input inputs_40__6 ;
    input inputs_40__5 ;
    input inputs_40__4 ;
    input inputs_40__3 ;
    input inputs_40__2 ;
    input inputs_40__1 ;
    input inputs_40__0 ;
    input inputs_41__15 ;
    input inputs_41__14 ;
    input inputs_41__13 ;
    input inputs_41__12 ;
    input inputs_41__11 ;
    input inputs_41__10 ;
    input inputs_41__9 ;
    input inputs_41__8 ;
    input inputs_41__7 ;
    input inputs_41__6 ;
    input inputs_41__5 ;
    input inputs_41__4 ;
    input inputs_41__3 ;
    input inputs_41__2 ;
    input inputs_41__1 ;
    input inputs_41__0 ;
    input inputs_42__15 ;
    input inputs_42__14 ;
    input inputs_42__13 ;
    input inputs_42__12 ;
    input inputs_42__11 ;
    input inputs_42__10 ;
    input inputs_42__9 ;
    input inputs_42__8 ;
    input inputs_42__7 ;
    input inputs_42__6 ;
    input inputs_42__5 ;
    input inputs_42__4 ;
    input inputs_42__3 ;
    input inputs_42__2 ;
    input inputs_42__1 ;
    input inputs_42__0 ;
    input inputs_43__15 ;
    input inputs_43__14 ;
    input inputs_43__13 ;
    input inputs_43__12 ;
    input inputs_43__11 ;
    input inputs_43__10 ;
    input inputs_43__9 ;
    input inputs_43__8 ;
    input inputs_43__7 ;
    input inputs_43__6 ;
    input inputs_43__5 ;
    input inputs_43__4 ;
    input inputs_43__3 ;
    input inputs_43__2 ;
    input inputs_43__1 ;
    input inputs_43__0 ;
    input inputs_44__15 ;
    input inputs_44__14 ;
    input inputs_44__13 ;
    input inputs_44__12 ;
    input inputs_44__11 ;
    input inputs_44__10 ;
    input inputs_44__9 ;
    input inputs_44__8 ;
    input inputs_44__7 ;
    input inputs_44__6 ;
    input inputs_44__5 ;
    input inputs_44__4 ;
    input inputs_44__3 ;
    input inputs_44__2 ;
    input inputs_44__1 ;
    input inputs_44__0 ;
    input inputs_45__15 ;
    input inputs_45__14 ;
    input inputs_45__13 ;
    input inputs_45__12 ;
    input inputs_45__11 ;
    input inputs_45__10 ;
    input inputs_45__9 ;
    input inputs_45__8 ;
    input inputs_45__7 ;
    input inputs_45__6 ;
    input inputs_45__5 ;
    input inputs_45__4 ;
    input inputs_45__3 ;
    input inputs_45__2 ;
    input inputs_45__1 ;
    input inputs_45__0 ;
    input inputs_46__15 ;
    input inputs_46__14 ;
    input inputs_46__13 ;
    input inputs_46__12 ;
    input inputs_46__11 ;
    input inputs_46__10 ;
    input inputs_46__9 ;
    input inputs_46__8 ;
    input inputs_46__7 ;
    input inputs_46__6 ;
    input inputs_46__5 ;
    input inputs_46__4 ;
    input inputs_46__3 ;
    input inputs_46__2 ;
    input inputs_46__1 ;
    input inputs_46__0 ;
    input inputs_47__15 ;
    input inputs_47__14 ;
    input inputs_47__13 ;
    input inputs_47__12 ;
    input inputs_47__11 ;
    input inputs_47__10 ;
    input inputs_47__9 ;
    input inputs_47__8 ;
    input inputs_47__7 ;
    input inputs_47__6 ;
    input inputs_47__5 ;
    input inputs_47__4 ;
    input inputs_47__3 ;
    input inputs_47__2 ;
    input inputs_47__1 ;
    input inputs_47__0 ;
    input inputs_48__15 ;
    input inputs_48__14 ;
    input inputs_48__13 ;
    input inputs_48__12 ;
    input inputs_48__11 ;
    input inputs_48__10 ;
    input inputs_48__9 ;
    input inputs_48__8 ;
    input inputs_48__7 ;
    input inputs_48__6 ;
    input inputs_48__5 ;
    input inputs_48__4 ;
    input inputs_48__3 ;
    input inputs_48__2 ;
    input inputs_48__1 ;
    input inputs_48__0 ;
    input inputs_49__15 ;
    input inputs_49__14 ;
    input inputs_49__13 ;
    input inputs_49__12 ;
    input inputs_49__11 ;
    input inputs_49__10 ;
    input inputs_49__9 ;
    input inputs_49__8 ;
    input inputs_49__7 ;
    input inputs_49__6 ;
    input inputs_49__5 ;
    input inputs_49__4 ;
    input inputs_49__3 ;
    input inputs_49__2 ;
    input inputs_49__1 ;
    input inputs_49__0 ;
    input inputs_50__15 ;
    input inputs_50__14 ;
    input inputs_50__13 ;
    input inputs_50__12 ;
    input inputs_50__11 ;
    input inputs_50__10 ;
    input inputs_50__9 ;
    input inputs_50__8 ;
    input inputs_50__7 ;
    input inputs_50__6 ;
    input inputs_50__5 ;
    input inputs_50__4 ;
    input inputs_50__3 ;
    input inputs_50__2 ;
    input inputs_50__1 ;
    input inputs_50__0 ;
    input inputs_51__15 ;
    input inputs_51__14 ;
    input inputs_51__13 ;
    input inputs_51__12 ;
    input inputs_51__11 ;
    input inputs_51__10 ;
    input inputs_51__9 ;
    input inputs_51__8 ;
    input inputs_51__7 ;
    input inputs_51__6 ;
    input inputs_51__5 ;
    input inputs_51__4 ;
    input inputs_51__3 ;
    input inputs_51__2 ;
    input inputs_51__1 ;
    input inputs_51__0 ;
    input inputs_52__15 ;
    input inputs_52__14 ;
    input inputs_52__13 ;
    input inputs_52__12 ;
    input inputs_52__11 ;
    input inputs_52__10 ;
    input inputs_52__9 ;
    input inputs_52__8 ;
    input inputs_52__7 ;
    input inputs_52__6 ;
    input inputs_52__5 ;
    input inputs_52__4 ;
    input inputs_52__3 ;
    input inputs_52__2 ;
    input inputs_52__1 ;
    input inputs_52__0 ;
    input inputs_53__15 ;
    input inputs_53__14 ;
    input inputs_53__13 ;
    input inputs_53__12 ;
    input inputs_53__11 ;
    input inputs_53__10 ;
    input inputs_53__9 ;
    input inputs_53__8 ;
    input inputs_53__7 ;
    input inputs_53__6 ;
    input inputs_53__5 ;
    input inputs_53__4 ;
    input inputs_53__3 ;
    input inputs_53__2 ;
    input inputs_53__1 ;
    input inputs_53__0 ;
    input inputs_54__15 ;
    input inputs_54__14 ;
    input inputs_54__13 ;
    input inputs_54__12 ;
    input inputs_54__11 ;
    input inputs_54__10 ;
    input inputs_54__9 ;
    input inputs_54__8 ;
    input inputs_54__7 ;
    input inputs_54__6 ;
    input inputs_54__5 ;
    input inputs_54__4 ;
    input inputs_54__3 ;
    input inputs_54__2 ;
    input inputs_54__1 ;
    input inputs_54__0 ;
    input inputs_55__15 ;
    input inputs_55__14 ;
    input inputs_55__13 ;
    input inputs_55__12 ;
    input inputs_55__11 ;
    input inputs_55__10 ;
    input inputs_55__9 ;
    input inputs_55__8 ;
    input inputs_55__7 ;
    input inputs_55__6 ;
    input inputs_55__5 ;
    input inputs_55__4 ;
    input inputs_55__3 ;
    input inputs_55__2 ;
    input inputs_55__1 ;
    input inputs_55__0 ;
    input inputs_56__15 ;
    input inputs_56__14 ;
    input inputs_56__13 ;
    input inputs_56__12 ;
    input inputs_56__11 ;
    input inputs_56__10 ;
    input inputs_56__9 ;
    input inputs_56__8 ;
    input inputs_56__7 ;
    input inputs_56__6 ;
    input inputs_56__5 ;
    input inputs_56__4 ;
    input inputs_56__3 ;
    input inputs_56__2 ;
    input inputs_56__1 ;
    input inputs_56__0 ;
    input inputs_57__15 ;
    input inputs_57__14 ;
    input inputs_57__13 ;
    input inputs_57__12 ;
    input inputs_57__11 ;
    input inputs_57__10 ;
    input inputs_57__9 ;
    input inputs_57__8 ;
    input inputs_57__7 ;
    input inputs_57__6 ;
    input inputs_57__5 ;
    input inputs_57__4 ;
    input inputs_57__3 ;
    input inputs_57__2 ;
    input inputs_57__1 ;
    input inputs_57__0 ;
    input inputs_58__15 ;
    input inputs_58__14 ;
    input inputs_58__13 ;
    input inputs_58__12 ;
    input inputs_58__11 ;
    input inputs_58__10 ;
    input inputs_58__9 ;
    input inputs_58__8 ;
    input inputs_58__7 ;
    input inputs_58__6 ;
    input inputs_58__5 ;
    input inputs_58__4 ;
    input inputs_58__3 ;
    input inputs_58__2 ;
    input inputs_58__1 ;
    input inputs_58__0 ;
    input inputs_59__15 ;
    input inputs_59__14 ;
    input inputs_59__13 ;
    input inputs_59__12 ;
    input inputs_59__11 ;
    input inputs_59__10 ;
    input inputs_59__9 ;
    input inputs_59__8 ;
    input inputs_59__7 ;
    input inputs_59__6 ;
    input inputs_59__5 ;
    input inputs_59__4 ;
    input inputs_59__3 ;
    input inputs_59__2 ;
    input inputs_59__1 ;
    input inputs_59__0 ;
    input inputs_60__15 ;
    input inputs_60__14 ;
    input inputs_60__13 ;
    input inputs_60__12 ;
    input inputs_60__11 ;
    input inputs_60__10 ;
    input inputs_60__9 ;
    input inputs_60__8 ;
    input inputs_60__7 ;
    input inputs_60__6 ;
    input inputs_60__5 ;
    input inputs_60__4 ;
    input inputs_60__3 ;
    input inputs_60__2 ;
    input inputs_60__1 ;
    input inputs_60__0 ;
    input inputs_61__15 ;
    input inputs_61__14 ;
    input inputs_61__13 ;
    input inputs_61__12 ;
    input inputs_61__11 ;
    input inputs_61__10 ;
    input inputs_61__9 ;
    input inputs_61__8 ;
    input inputs_61__7 ;
    input inputs_61__6 ;
    input inputs_61__5 ;
    input inputs_61__4 ;
    input inputs_61__3 ;
    input inputs_61__2 ;
    input inputs_61__1 ;
    input inputs_61__0 ;
    input inputs_62__15 ;
    input inputs_62__14 ;
    input inputs_62__13 ;
    input inputs_62__12 ;
    input inputs_62__11 ;
    input inputs_62__10 ;
    input inputs_62__9 ;
    input inputs_62__8 ;
    input inputs_62__7 ;
    input inputs_62__6 ;
    input inputs_62__5 ;
    input inputs_62__4 ;
    input inputs_62__3 ;
    input inputs_62__2 ;
    input inputs_62__1 ;
    input inputs_62__0 ;
    input inputs_63__15 ;
    input inputs_63__14 ;
    input inputs_63__13 ;
    input inputs_63__12 ;
    input inputs_63__11 ;
    input inputs_63__10 ;
    input inputs_63__9 ;
    input inputs_63__8 ;
    input inputs_63__7 ;
    input inputs_63__6 ;
    input inputs_63__5 ;
    input inputs_63__4 ;
    input inputs_63__3 ;
    input inputs_63__2 ;
    input inputs_63__1 ;
    input inputs_63__0 ;
    input inputs_64__15 ;
    input inputs_64__14 ;
    input inputs_64__13 ;
    input inputs_64__12 ;
    input inputs_64__11 ;
    input inputs_64__10 ;
    input inputs_64__9 ;
    input inputs_64__8 ;
    input inputs_64__7 ;
    input inputs_64__6 ;
    input inputs_64__5 ;
    input inputs_64__4 ;
    input inputs_64__3 ;
    input inputs_64__2 ;
    input inputs_64__1 ;
    input inputs_64__0 ;
    input inputs_65__15 ;
    input inputs_65__14 ;
    input inputs_65__13 ;
    input inputs_65__12 ;
    input inputs_65__11 ;
    input inputs_65__10 ;
    input inputs_65__9 ;
    input inputs_65__8 ;
    input inputs_65__7 ;
    input inputs_65__6 ;
    input inputs_65__5 ;
    input inputs_65__4 ;
    input inputs_65__3 ;
    input inputs_65__2 ;
    input inputs_65__1 ;
    input inputs_65__0 ;
    input inputs_66__15 ;
    input inputs_66__14 ;
    input inputs_66__13 ;
    input inputs_66__12 ;
    input inputs_66__11 ;
    input inputs_66__10 ;
    input inputs_66__9 ;
    input inputs_66__8 ;
    input inputs_66__7 ;
    input inputs_66__6 ;
    input inputs_66__5 ;
    input inputs_66__4 ;
    input inputs_66__3 ;
    input inputs_66__2 ;
    input inputs_66__1 ;
    input inputs_66__0 ;
    input inputs_67__15 ;
    input inputs_67__14 ;
    input inputs_67__13 ;
    input inputs_67__12 ;
    input inputs_67__11 ;
    input inputs_67__10 ;
    input inputs_67__9 ;
    input inputs_67__8 ;
    input inputs_67__7 ;
    input inputs_67__6 ;
    input inputs_67__5 ;
    input inputs_67__4 ;
    input inputs_67__3 ;
    input inputs_67__2 ;
    input inputs_67__1 ;
    input inputs_67__0 ;
    input inputs_68__15 ;
    input inputs_68__14 ;
    input inputs_68__13 ;
    input inputs_68__12 ;
    input inputs_68__11 ;
    input inputs_68__10 ;
    input inputs_68__9 ;
    input inputs_68__8 ;
    input inputs_68__7 ;
    input inputs_68__6 ;
    input inputs_68__5 ;
    input inputs_68__4 ;
    input inputs_68__3 ;
    input inputs_68__2 ;
    input inputs_68__1 ;
    input inputs_68__0 ;
    input inputs_69__15 ;
    input inputs_69__14 ;
    input inputs_69__13 ;
    input inputs_69__12 ;
    input inputs_69__11 ;
    input inputs_69__10 ;
    input inputs_69__9 ;
    input inputs_69__8 ;
    input inputs_69__7 ;
    input inputs_69__6 ;
    input inputs_69__5 ;
    input inputs_69__4 ;
    input inputs_69__3 ;
    input inputs_69__2 ;
    input inputs_69__1 ;
    input inputs_69__0 ;
    input inputs_70__15 ;
    input inputs_70__14 ;
    input inputs_70__13 ;
    input inputs_70__12 ;
    input inputs_70__11 ;
    input inputs_70__10 ;
    input inputs_70__9 ;
    input inputs_70__8 ;
    input inputs_70__7 ;
    input inputs_70__6 ;
    input inputs_70__5 ;
    input inputs_70__4 ;
    input inputs_70__3 ;
    input inputs_70__2 ;
    input inputs_70__1 ;
    input inputs_70__0 ;
    input inputs_71__15 ;
    input inputs_71__14 ;
    input inputs_71__13 ;
    input inputs_71__12 ;
    input inputs_71__11 ;
    input inputs_71__10 ;
    input inputs_71__9 ;
    input inputs_71__8 ;
    input inputs_71__7 ;
    input inputs_71__6 ;
    input inputs_71__5 ;
    input inputs_71__4 ;
    input inputs_71__3 ;
    input inputs_71__2 ;
    input inputs_71__1 ;
    input inputs_71__0 ;
    input inputs_72__15 ;
    input inputs_72__14 ;
    input inputs_72__13 ;
    input inputs_72__12 ;
    input inputs_72__11 ;
    input inputs_72__10 ;
    input inputs_72__9 ;
    input inputs_72__8 ;
    input inputs_72__7 ;
    input inputs_72__6 ;
    input inputs_72__5 ;
    input inputs_72__4 ;
    input inputs_72__3 ;
    input inputs_72__2 ;
    input inputs_72__1 ;
    input inputs_72__0 ;
    input inputs_73__15 ;
    input inputs_73__14 ;
    input inputs_73__13 ;
    input inputs_73__12 ;
    input inputs_73__11 ;
    input inputs_73__10 ;
    input inputs_73__9 ;
    input inputs_73__8 ;
    input inputs_73__7 ;
    input inputs_73__6 ;
    input inputs_73__5 ;
    input inputs_73__4 ;
    input inputs_73__3 ;
    input inputs_73__2 ;
    input inputs_73__1 ;
    input inputs_73__0 ;
    input inputs_74__15 ;
    input inputs_74__14 ;
    input inputs_74__13 ;
    input inputs_74__12 ;
    input inputs_74__11 ;
    input inputs_74__10 ;
    input inputs_74__9 ;
    input inputs_74__8 ;
    input inputs_74__7 ;
    input inputs_74__6 ;
    input inputs_74__5 ;
    input inputs_74__4 ;
    input inputs_74__3 ;
    input inputs_74__2 ;
    input inputs_74__1 ;
    input inputs_74__0 ;
    input inputs_75__15 ;
    input inputs_75__14 ;
    input inputs_75__13 ;
    input inputs_75__12 ;
    input inputs_75__11 ;
    input inputs_75__10 ;
    input inputs_75__9 ;
    input inputs_75__8 ;
    input inputs_75__7 ;
    input inputs_75__6 ;
    input inputs_75__5 ;
    input inputs_75__4 ;
    input inputs_75__3 ;
    input inputs_75__2 ;
    input inputs_75__1 ;
    input inputs_75__0 ;
    input inputs_76__15 ;
    input inputs_76__14 ;
    input inputs_76__13 ;
    input inputs_76__12 ;
    input inputs_76__11 ;
    input inputs_76__10 ;
    input inputs_76__9 ;
    input inputs_76__8 ;
    input inputs_76__7 ;
    input inputs_76__6 ;
    input inputs_76__5 ;
    input inputs_76__4 ;
    input inputs_76__3 ;
    input inputs_76__2 ;
    input inputs_76__1 ;
    input inputs_76__0 ;
    input inputs_77__15 ;
    input inputs_77__14 ;
    input inputs_77__13 ;
    input inputs_77__12 ;
    input inputs_77__11 ;
    input inputs_77__10 ;
    input inputs_77__9 ;
    input inputs_77__8 ;
    input inputs_77__7 ;
    input inputs_77__6 ;
    input inputs_77__5 ;
    input inputs_77__4 ;
    input inputs_77__3 ;
    input inputs_77__2 ;
    input inputs_77__1 ;
    input inputs_77__0 ;
    input inputs_78__15 ;
    input inputs_78__14 ;
    input inputs_78__13 ;
    input inputs_78__12 ;
    input inputs_78__11 ;
    input inputs_78__10 ;
    input inputs_78__9 ;
    input inputs_78__8 ;
    input inputs_78__7 ;
    input inputs_78__6 ;
    input inputs_78__5 ;
    input inputs_78__4 ;
    input inputs_78__3 ;
    input inputs_78__2 ;
    input inputs_78__1 ;
    input inputs_78__0 ;
    input inputs_79__15 ;
    input inputs_79__14 ;
    input inputs_79__13 ;
    input inputs_79__12 ;
    input inputs_79__11 ;
    input inputs_79__10 ;
    input inputs_79__9 ;
    input inputs_79__8 ;
    input inputs_79__7 ;
    input inputs_79__6 ;
    input inputs_79__5 ;
    input inputs_79__4 ;
    input inputs_79__3 ;
    input inputs_79__2 ;
    input inputs_79__1 ;
    input inputs_79__0 ;
    input inputs_80__15 ;
    input inputs_80__14 ;
    input inputs_80__13 ;
    input inputs_80__12 ;
    input inputs_80__11 ;
    input inputs_80__10 ;
    input inputs_80__9 ;
    input inputs_80__8 ;
    input inputs_80__7 ;
    input inputs_80__6 ;
    input inputs_80__5 ;
    input inputs_80__4 ;
    input inputs_80__3 ;
    input inputs_80__2 ;
    input inputs_80__1 ;
    input inputs_80__0 ;
    input inputs_81__15 ;
    input inputs_81__14 ;
    input inputs_81__13 ;
    input inputs_81__12 ;
    input inputs_81__11 ;
    input inputs_81__10 ;
    input inputs_81__9 ;
    input inputs_81__8 ;
    input inputs_81__7 ;
    input inputs_81__6 ;
    input inputs_81__5 ;
    input inputs_81__4 ;
    input inputs_81__3 ;
    input inputs_81__2 ;
    input inputs_81__1 ;
    input inputs_81__0 ;
    input inputs_82__15 ;
    input inputs_82__14 ;
    input inputs_82__13 ;
    input inputs_82__12 ;
    input inputs_82__11 ;
    input inputs_82__10 ;
    input inputs_82__9 ;
    input inputs_82__8 ;
    input inputs_82__7 ;
    input inputs_82__6 ;
    input inputs_82__5 ;
    input inputs_82__4 ;
    input inputs_82__3 ;
    input inputs_82__2 ;
    input inputs_82__1 ;
    input inputs_82__0 ;
    input inputs_83__15 ;
    input inputs_83__14 ;
    input inputs_83__13 ;
    input inputs_83__12 ;
    input inputs_83__11 ;
    input inputs_83__10 ;
    input inputs_83__9 ;
    input inputs_83__8 ;
    input inputs_83__7 ;
    input inputs_83__6 ;
    input inputs_83__5 ;
    input inputs_83__4 ;
    input inputs_83__3 ;
    input inputs_83__2 ;
    input inputs_83__1 ;
    input inputs_83__0 ;
    input inputs_84__15 ;
    input inputs_84__14 ;
    input inputs_84__13 ;
    input inputs_84__12 ;
    input inputs_84__11 ;
    input inputs_84__10 ;
    input inputs_84__9 ;
    input inputs_84__8 ;
    input inputs_84__7 ;
    input inputs_84__6 ;
    input inputs_84__5 ;
    input inputs_84__4 ;
    input inputs_84__3 ;
    input inputs_84__2 ;
    input inputs_84__1 ;
    input inputs_84__0 ;
    input inputs_85__15 ;
    input inputs_85__14 ;
    input inputs_85__13 ;
    input inputs_85__12 ;
    input inputs_85__11 ;
    input inputs_85__10 ;
    input inputs_85__9 ;
    input inputs_85__8 ;
    input inputs_85__7 ;
    input inputs_85__6 ;
    input inputs_85__5 ;
    input inputs_85__4 ;
    input inputs_85__3 ;
    input inputs_85__2 ;
    input inputs_85__1 ;
    input inputs_85__0 ;
    input inputs_86__15 ;
    input inputs_86__14 ;
    input inputs_86__13 ;
    input inputs_86__12 ;
    input inputs_86__11 ;
    input inputs_86__10 ;
    input inputs_86__9 ;
    input inputs_86__8 ;
    input inputs_86__7 ;
    input inputs_86__6 ;
    input inputs_86__5 ;
    input inputs_86__4 ;
    input inputs_86__3 ;
    input inputs_86__2 ;
    input inputs_86__1 ;
    input inputs_86__0 ;
    input inputs_87__15 ;
    input inputs_87__14 ;
    input inputs_87__13 ;
    input inputs_87__12 ;
    input inputs_87__11 ;
    input inputs_87__10 ;
    input inputs_87__9 ;
    input inputs_87__8 ;
    input inputs_87__7 ;
    input inputs_87__6 ;
    input inputs_87__5 ;
    input inputs_87__4 ;
    input inputs_87__3 ;
    input inputs_87__2 ;
    input inputs_87__1 ;
    input inputs_87__0 ;
    input inputs_88__15 ;
    input inputs_88__14 ;
    input inputs_88__13 ;
    input inputs_88__12 ;
    input inputs_88__11 ;
    input inputs_88__10 ;
    input inputs_88__9 ;
    input inputs_88__8 ;
    input inputs_88__7 ;
    input inputs_88__6 ;
    input inputs_88__5 ;
    input inputs_88__4 ;
    input inputs_88__3 ;
    input inputs_88__2 ;
    input inputs_88__1 ;
    input inputs_88__0 ;
    input inputs_89__15 ;
    input inputs_89__14 ;
    input inputs_89__13 ;
    input inputs_89__12 ;
    input inputs_89__11 ;
    input inputs_89__10 ;
    input inputs_89__9 ;
    input inputs_89__8 ;
    input inputs_89__7 ;
    input inputs_89__6 ;
    input inputs_89__5 ;
    input inputs_89__4 ;
    input inputs_89__3 ;
    input inputs_89__2 ;
    input inputs_89__1 ;
    input inputs_89__0 ;
    input inputs_90__15 ;
    input inputs_90__14 ;
    input inputs_90__13 ;
    input inputs_90__12 ;
    input inputs_90__11 ;
    input inputs_90__10 ;
    input inputs_90__9 ;
    input inputs_90__8 ;
    input inputs_90__7 ;
    input inputs_90__6 ;
    input inputs_90__5 ;
    input inputs_90__4 ;
    input inputs_90__3 ;
    input inputs_90__2 ;
    input inputs_90__1 ;
    input inputs_90__0 ;
    input inputs_91__15 ;
    input inputs_91__14 ;
    input inputs_91__13 ;
    input inputs_91__12 ;
    input inputs_91__11 ;
    input inputs_91__10 ;
    input inputs_91__9 ;
    input inputs_91__8 ;
    input inputs_91__7 ;
    input inputs_91__6 ;
    input inputs_91__5 ;
    input inputs_91__4 ;
    input inputs_91__3 ;
    input inputs_91__2 ;
    input inputs_91__1 ;
    input inputs_91__0 ;
    input inputs_92__15 ;
    input inputs_92__14 ;
    input inputs_92__13 ;
    input inputs_92__12 ;
    input inputs_92__11 ;
    input inputs_92__10 ;
    input inputs_92__9 ;
    input inputs_92__8 ;
    input inputs_92__7 ;
    input inputs_92__6 ;
    input inputs_92__5 ;
    input inputs_92__4 ;
    input inputs_92__3 ;
    input inputs_92__2 ;
    input inputs_92__1 ;
    input inputs_92__0 ;
    input inputs_93__15 ;
    input inputs_93__14 ;
    input inputs_93__13 ;
    input inputs_93__12 ;
    input inputs_93__11 ;
    input inputs_93__10 ;
    input inputs_93__9 ;
    input inputs_93__8 ;
    input inputs_93__7 ;
    input inputs_93__6 ;
    input inputs_93__5 ;
    input inputs_93__4 ;
    input inputs_93__3 ;
    input inputs_93__2 ;
    input inputs_93__1 ;
    input inputs_93__0 ;
    input inputs_94__15 ;
    input inputs_94__14 ;
    input inputs_94__13 ;
    input inputs_94__12 ;
    input inputs_94__11 ;
    input inputs_94__10 ;
    input inputs_94__9 ;
    input inputs_94__8 ;
    input inputs_94__7 ;
    input inputs_94__6 ;
    input inputs_94__5 ;
    input inputs_94__4 ;
    input inputs_94__3 ;
    input inputs_94__2 ;
    input inputs_94__1 ;
    input inputs_94__0 ;
    input inputs_95__15 ;
    input inputs_95__14 ;
    input inputs_95__13 ;
    input inputs_95__12 ;
    input inputs_95__11 ;
    input inputs_95__10 ;
    input inputs_95__9 ;
    input inputs_95__8 ;
    input inputs_95__7 ;
    input inputs_95__6 ;
    input inputs_95__5 ;
    input inputs_95__4 ;
    input inputs_95__3 ;
    input inputs_95__2 ;
    input inputs_95__1 ;
    input inputs_95__0 ;
    input inputs_96__15 ;
    input inputs_96__14 ;
    input inputs_96__13 ;
    input inputs_96__12 ;
    input inputs_96__11 ;
    input inputs_96__10 ;
    input inputs_96__9 ;
    input inputs_96__8 ;
    input inputs_96__7 ;
    input inputs_96__6 ;
    input inputs_96__5 ;
    input inputs_96__4 ;
    input inputs_96__3 ;
    input inputs_96__2 ;
    input inputs_96__1 ;
    input inputs_96__0 ;
    input inputs_97__15 ;
    input inputs_97__14 ;
    input inputs_97__13 ;
    input inputs_97__12 ;
    input inputs_97__11 ;
    input inputs_97__10 ;
    input inputs_97__9 ;
    input inputs_97__8 ;
    input inputs_97__7 ;
    input inputs_97__6 ;
    input inputs_97__5 ;
    input inputs_97__4 ;
    input inputs_97__3 ;
    input inputs_97__2 ;
    input inputs_97__1 ;
    input inputs_97__0 ;
    input inputs_98__15 ;
    input inputs_98__14 ;
    input inputs_98__13 ;
    input inputs_98__12 ;
    input inputs_98__11 ;
    input inputs_98__10 ;
    input inputs_98__9 ;
    input inputs_98__8 ;
    input inputs_98__7 ;
    input inputs_98__6 ;
    input inputs_98__5 ;
    input inputs_98__4 ;
    input inputs_98__3 ;
    input inputs_98__2 ;
    input inputs_98__1 ;
    input inputs_98__0 ;
    input inputs_99__15 ;
    input inputs_99__14 ;
    input inputs_99__13 ;
    input inputs_99__12 ;
    input inputs_99__11 ;
    input inputs_99__10 ;
    input inputs_99__9 ;
    input inputs_99__8 ;
    input inputs_99__7 ;
    input inputs_99__6 ;
    input inputs_99__5 ;
    input inputs_99__4 ;
    input inputs_99__3 ;
    input inputs_99__2 ;
    input inputs_99__1 ;
    input inputs_99__0 ;
    input inputs_100__15 ;
    input inputs_100__14 ;
    input inputs_100__13 ;
    input inputs_100__12 ;
    input inputs_100__11 ;
    input inputs_100__10 ;
    input inputs_100__9 ;
    input inputs_100__8 ;
    input inputs_100__7 ;
    input inputs_100__6 ;
    input inputs_100__5 ;
    input inputs_100__4 ;
    input inputs_100__3 ;
    input inputs_100__2 ;
    input inputs_100__1 ;
    input inputs_100__0 ;
    input inputs_101__15 ;
    input inputs_101__14 ;
    input inputs_101__13 ;
    input inputs_101__12 ;
    input inputs_101__11 ;
    input inputs_101__10 ;
    input inputs_101__9 ;
    input inputs_101__8 ;
    input inputs_101__7 ;
    input inputs_101__6 ;
    input inputs_101__5 ;
    input inputs_101__4 ;
    input inputs_101__3 ;
    input inputs_101__2 ;
    input inputs_101__1 ;
    input inputs_101__0 ;
    input inputs_102__15 ;
    input inputs_102__14 ;
    input inputs_102__13 ;
    input inputs_102__12 ;
    input inputs_102__11 ;
    input inputs_102__10 ;
    input inputs_102__9 ;
    input inputs_102__8 ;
    input inputs_102__7 ;
    input inputs_102__6 ;
    input inputs_102__5 ;
    input inputs_102__4 ;
    input inputs_102__3 ;
    input inputs_102__2 ;
    input inputs_102__1 ;
    input inputs_102__0 ;
    input inputs_103__15 ;
    input inputs_103__14 ;
    input inputs_103__13 ;
    input inputs_103__12 ;
    input inputs_103__11 ;
    input inputs_103__10 ;
    input inputs_103__9 ;
    input inputs_103__8 ;
    input inputs_103__7 ;
    input inputs_103__6 ;
    input inputs_103__5 ;
    input inputs_103__4 ;
    input inputs_103__3 ;
    input inputs_103__2 ;
    input inputs_103__1 ;
    input inputs_103__0 ;
    input inputs_104__15 ;
    input inputs_104__14 ;
    input inputs_104__13 ;
    input inputs_104__12 ;
    input inputs_104__11 ;
    input inputs_104__10 ;
    input inputs_104__9 ;
    input inputs_104__8 ;
    input inputs_104__7 ;
    input inputs_104__6 ;
    input inputs_104__5 ;
    input inputs_104__4 ;
    input inputs_104__3 ;
    input inputs_104__2 ;
    input inputs_104__1 ;
    input inputs_104__0 ;
    input inputs_105__15 ;
    input inputs_105__14 ;
    input inputs_105__13 ;
    input inputs_105__12 ;
    input inputs_105__11 ;
    input inputs_105__10 ;
    input inputs_105__9 ;
    input inputs_105__8 ;
    input inputs_105__7 ;
    input inputs_105__6 ;
    input inputs_105__5 ;
    input inputs_105__4 ;
    input inputs_105__3 ;
    input inputs_105__2 ;
    input inputs_105__1 ;
    input inputs_105__0 ;
    input inputs_106__15 ;
    input inputs_106__14 ;
    input inputs_106__13 ;
    input inputs_106__12 ;
    input inputs_106__11 ;
    input inputs_106__10 ;
    input inputs_106__9 ;
    input inputs_106__8 ;
    input inputs_106__7 ;
    input inputs_106__6 ;
    input inputs_106__5 ;
    input inputs_106__4 ;
    input inputs_106__3 ;
    input inputs_106__2 ;
    input inputs_106__1 ;
    input inputs_106__0 ;
    input inputs_107__15 ;
    input inputs_107__14 ;
    input inputs_107__13 ;
    input inputs_107__12 ;
    input inputs_107__11 ;
    input inputs_107__10 ;
    input inputs_107__9 ;
    input inputs_107__8 ;
    input inputs_107__7 ;
    input inputs_107__6 ;
    input inputs_107__5 ;
    input inputs_107__4 ;
    input inputs_107__3 ;
    input inputs_107__2 ;
    input inputs_107__1 ;
    input inputs_107__0 ;
    input inputs_108__15 ;
    input inputs_108__14 ;
    input inputs_108__13 ;
    input inputs_108__12 ;
    input inputs_108__11 ;
    input inputs_108__10 ;
    input inputs_108__9 ;
    input inputs_108__8 ;
    input inputs_108__7 ;
    input inputs_108__6 ;
    input inputs_108__5 ;
    input inputs_108__4 ;
    input inputs_108__3 ;
    input inputs_108__2 ;
    input inputs_108__1 ;
    input inputs_108__0 ;
    input inputs_109__15 ;
    input inputs_109__14 ;
    input inputs_109__13 ;
    input inputs_109__12 ;
    input inputs_109__11 ;
    input inputs_109__10 ;
    input inputs_109__9 ;
    input inputs_109__8 ;
    input inputs_109__7 ;
    input inputs_109__6 ;
    input inputs_109__5 ;
    input inputs_109__4 ;
    input inputs_109__3 ;
    input inputs_109__2 ;
    input inputs_109__1 ;
    input inputs_109__0 ;
    input inputs_110__15 ;
    input inputs_110__14 ;
    input inputs_110__13 ;
    input inputs_110__12 ;
    input inputs_110__11 ;
    input inputs_110__10 ;
    input inputs_110__9 ;
    input inputs_110__8 ;
    input inputs_110__7 ;
    input inputs_110__6 ;
    input inputs_110__5 ;
    input inputs_110__4 ;
    input inputs_110__3 ;
    input inputs_110__2 ;
    input inputs_110__1 ;
    input inputs_110__0 ;
    input inputs_111__15 ;
    input inputs_111__14 ;
    input inputs_111__13 ;
    input inputs_111__12 ;
    input inputs_111__11 ;
    input inputs_111__10 ;
    input inputs_111__9 ;
    input inputs_111__8 ;
    input inputs_111__7 ;
    input inputs_111__6 ;
    input inputs_111__5 ;
    input inputs_111__4 ;
    input inputs_111__3 ;
    input inputs_111__2 ;
    input inputs_111__1 ;
    input inputs_111__0 ;
    input inputs_112__15 ;
    input inputs_112__14 ;
    input inputs_112__13 ;
    input inputs_112__12 ;
    input inputs_112__11 ;
    input inputs_112__10 ;
    input inputs_112__9 ;
    input inputs_112__8 ;
    input inputs_112__7 ;
    input inputs_112__6 ;
    input inputs_112__5 ;
    input inputs_112__4 ;
    input inputs_112__3 ;
    input inputs_112__2 ;
    input inputs_112__1 ;
    input inputs_112__0 ;
    input inputs_113__15 ;
    input inputs_113__14 ;
    input inputs_113__13 ;
    input inputs_113__12 ;
    input inputs_113__11 ;
    input inputs_113__10 ;
    input inputs_113__9 ;
    input inputs_113__8 ;
    input inputs_113__7 ;
    input inputs_113__6 ;
    input inputs_113__5 ;
    input inputs_113__4 ;
    input inputs_113__3 ;
    input inputs_113__2 ;
    input inputs_113__1 ;
    input inputs_113__0 ;
    input inputs_114__15 ;
    input inputs_114__14 ;
    input inputs_114__13 ;
    input inputs_114__12 ;
    input inputs_114__11 ;
    input inputs_114__10 ;
    input inputs_114__9 ;
    input inputs_114__8 ;
    input inputs_114__7 ;
    input inputs_114__6 ;
    input inputs_114__5 ;
    input inputs_114__4 ;
    input inputs_114__3 ;
    input inputs_114__2 ;
    input inputs_114__1 ;
    input inputs_114__0 ;
    input inputs_115__15 ;
    input inputs_115__14 ;
    input inputs_115__13 ;
    input inputs_115__12 ;
    input inputs_115__11 ;
    input inputs_115__10 ;
    input inputs_115__9 ;
    input inputs_115__8 ;
    input inputs_115__7 ;
    input inputs_115__6 ;
    input inputs_115__5 ;
    input inputs_115__4 ;
    input inputs_115__3 ;
    input inputs_115__2 ;
    input inputs_115__1 ;
    input inputs_115__0 ;
    input inputs_116__15 ;
    input inputs_116__14 ;
    input inputs_116__13 ;
    input inputs_116__12 ;
    input inputs_116__11 ;
    input inputs_116__10 ;
    input inputs_116__9 ;
    input inputs_116__8 ;
    input inputs_116__7 ;
    input inputs_116__6 ;
    input inputs_116__5 ;
    input inputs_116__4 ;
    input inputs_116__3 ;
    input inputs_116__2 ;
    input inputs_116__1 ;
    input inputs_116__0 ;
    input inputs_117__15 ;
    input inputs_117__14 ;
    input inputs_117__13 ;
    input inputs_117__12 ;
    input inputs_117__11 ;
    input inputs_117__10 ;
    input inputs_117__9 ;
    input inputs_117__8 ;
    input inputs_117__7 ;
    input inputs_117__6 ;
    input inputs_117__5 ;
    input inputs_117__4 ;
    input inputs_117__3 ;
    input inputs_117__2 ;
    input inputs_117__1 ;
    input inputs_117__0 ;
    input inputs_118__15 ;
    input inputs_118__14 ;
    input inputs_118__13 ;
    input inputs_118__12 ;
    input inputs_118__11 ;
    input inputs_118__10 ;
    input inputs_118__9 ;
    input inputs_118__8 ;
    input inputs_118__7 ;
    input inputs_118__6 ;
    input inputs_118__5 ;
    input inputs_118__4 ;
    input inputs_118__3 ;
    input inputs_118__2 ;
    input inputs_118__1 ;
    input inputs_118__0 ;
    input inputs_119__15 ;
    input inputs_119__14 ;
    input inputs_119__13 ;
    input inputs_119__12 ;
    input inputs_119__11 ;
    input inputs_119__10 ;
    input inputs_119__9 ;
    input inputs_119__8 ;
    input inputs_119__7 ;
    input inputs_119__6 ;
    input inputs_119__5 ;
    input inputs_119__4 ;
    input inputs_119__3 ;
    input inputs_119__2 ;
    input inputs_119__1 ;
    input inputs_119__0 ;
    input inputs_120__15 ;
    input inputs_120__14 ;
    input inputs_120__13 ;
    input inputs_120__12 ;
    input inputs_120__11 ;
    input inputs_120__10 ;
    input inputs_120__9 ;
    input inputs_120__8 ;
    input inputs_120__7 ;
    input inputs_120__6 ;
    input inputs_120__5 ;
    input inputs_120__4 ;
    input inputs_120__3 ;
    input inputs_120__2 ;
    input inputs_120__1 ;
    input inputs_120__0 ;
    input inputs_121__15 ;
    input inputs_121__14 ;
    input inputs_121__13 ;
    input inputs_121__12 ;
    input inputs_121__11 ;
    input inputs_121__10 ;
    input inputs_121__9 ;
    input inputs_121__8 ;
    input inputs_121__7 ;
    input inputs_121__6 ;
    input inputs_121__5 ;
    input inputs_121__4 ;
    input inputs_121__3 ;
    input inputs_121__2 ;
    input inputs_121__1 ;
    input inputs_121__0 ;
    input inputs_122__15 ;
    input inputs_122__14 ;
    input inputs_122__13 ;
    input inputs_122__12 ;
    input inputs_122__11 ;
    input inputs_122__10 ;
    input inputs_122__9 ;
    input inputs_122__8 ;
    input inputs_122__7 ;
    input inputs_122__6 ;
    input inputs_122__5 ;
    input inputs_122__4 ;
    input inputs_122__3 ;
    input inputs_122__2 ;
    input inputs_122__1 ;
    input inputs_122__0 ;
    input inputs_123__15 ;
    input inputs_123__14 ;
    input inputs_123__13 ;
    input inputs_123__12 ;
    input inputs_123__11 ;
    input inputs_123__10 ;
    input inputs_123__9 ;
    input inputs_123__8 ;
    input inputs_123__7 ;
    input inputs_123__6 ;
    input inputs_123__5 ;
    input inputs_123__4 ;
    input inputs_123__3 ;
    input inputs_123__2 ;
    input inputs_123__1 ;
    input inputs_123__0 ;
    input inputs_124__15 ;
    input inputs_124__14 ;
    input inputs_124__13 ;
    input inputs_124__12 ;
    input inputs_124__11 ;
    input inputs_124__10 ;
    input inputs_124__9 ;
    input inputs_124__8 ;
    input inputs_124__7 ;
    input inputs_124__6 ;
    input inputs_124__5 ;
    input inputs_124__4 ;
    input inputs_124__3 ;
    input inputs_124__2 ;
    input inputs_124__1 ;
    input inputs_124__0 ;
    input inputs_125__15 ;
    input inputs_125__14 ;
    input inputs_125__13 ;
    input inputs_125__12 ;
    input inputs_125__11 ;
    input inputs_125__10 ;
    input inputs_125__9 ;
    input inputs_125__8 ;
    input inputs_125__7 ;
    input inputs_125__6 ;
    input inputs_125__5 ;
    input inputs_125__4 ;
    input inputs_125__3 ;
    input inputs_125__2 ;
    input inputs_125__1 ;
    input inputs_125__0 ;
    input inputs_126__15 ;
    input inputs_126__14 ;
    input inputs_126__13 ;
    input inputs_126__12 ;
    input inputs_126__11 ;
    input inputs_126__10 ;
    input inputs_126__9 ;
    input inputs_126__8 ;
    input inputs_126__7 ;
    input inputs_126__6 ;
    input inputs_126__5 ;
    input inputs_126__4 ;
    input inputs_126__3 ;
    input inputs_126__2 ;
    input inputs_126__1 ;
    input inputs_126__0 ;
    input inputs_127__15 ;
    input inputs_127__14 ;
    input inputs_127__13 ;
    input inputs_127__12 ;
    input inputs_127__11 ;
    input inputs_127__10 ;
    input inputs_127__9 ;
    input inputs_127__8 ;
    input inputs_127__7 ;
    input inputs_127__6 ;
    input inputs_127__5 ;
    input inputs_127__4 ;
    input inputs_127__3 ;
    input inputs_127__2 ;
    input inputs_127__1 ;
    input inputs_127__0 ;
    input inputs_128__15 ;
    input inputs_128__14 ;
    input inputs_128__13 ;
    input inputs_128__12 ;
    input inputs_128__11 ;
    input inputs_128__10 ;
    input inputs_128__9 ;
    input inputs_128__8 ;
    input inputs_128__7 ;
    input inputs_128__6 ;
    input inputs_128__5 ;
    input inputs_128__4 ;
    input inputs_128__3 ;
    input inputs_128__2 ;
    input inputs_128__1 ;
    input inputs_128__0 ;
    input inputs_129__15 ;
    input inputs_129__14 ;
    input inputs_129__13 ;
    input inputs_129__12 ;
    input inputs_129__11 ;
    input inputs_129__10 ;
    input inputs_129__9 ;
    input inputs_129__8 ;
    input inputs_129__7 ;
    input inputs_129__6 ;
    input inputs_129__5 ;
    input inputs_129__4 ;
    input inputs_129__3 ;
    input inputs_129__2 ;
    input inputs_129__1 ;
    input inputs_129__0 ;
    input inputs_130__15 ;
    input inputs_130__14 ;
    input inputs_130__13 ;
    input inputs_130__12 ;
    input inputs_130__11 ;
    input inputs_130__10 ;
    input inputs_130__9 ;
    input inputs_130__8 ;
    input inputs_130__7 ;
    input inputs_130__6 ;
    input inputs_130__5 ;
    input inputs_130__4 ;
    input inputs_130__3 ;
    input inputs_130__2 ;
    input inputs_130__1 ;
    input inputs_130__0 ;
    input inputs_131__15 ;
    input inputs_131__14 ;
    input inputs_131__13 ;
    input inputs_131__12 ;
    input inputs_131__11 ;
    input inputs_131__10 ;
    input inputs_131__9 ;
    input inputs_131__8 ;
    input inputs_131__7 ;
    input inputs_131__6 ;
    input inputs_131__5 ;
    input inputs_131__4 ;
    input inputs_131__3 ;
    input inputs_131__2 ;
    input inputs_131__1 ;
    input inputs_131__0 ;
    input inputs_132__15 ;
    input inputs_132__14 ;
    input inputs_132__13 ;
    input inputs_132__12 ;
    input inputs_132__11 ;
    input inputs_132__10 ;
    input inputs_132__9 ;
    input inputs_132__8 ;
    input inputs_132__7 ;
    input inputs_132__6 ;
    input inputs_132__5 ;
    input inputs_132__4 ;
    input inputs_132__3 ;
    input inputs_132__2 ;
    input inputs_132__1 ;
    input inputs_132__0 ;
    input inputs_133__15 ;
    input inputs_133__14 ;
    input inputs_133__13 ;
    input inputs_133__12 ;
    input inputs_133__11 ;
    input inputs_133__10 ;
    input inputs_133__9 ;
    input inputs_133__8 ;
    input inputs_133__7 ;
    input inputs_133__6 ;
    input inputs_133__5 ;
    input inputs_133__4 ;
    input inputs_133__3 ;
    input inputs_133__2 ;
    input inputs_133__1 ;
    input inputs_133__0 ;
    input inputs_134__15 ;
    input inputs_134__14 ;
    input inputs_134__13 ;
    input inputs_134__12 ;
    input inputs_134__11 ;
    input inputs_134__10 ;
    input inputs_134__9 ;
    input inputs_134__8 ;
    input inputs_134__7 ;
    input inputs_134__6 ;
    input inputs_134__5 ;
    input inputs_134__4 ;
    input inputs_134__3 ;
    input inputs_134__2 ;
    input inputs_134__1 ;
    input inputs_134__0 ;
    input inputs_135__15 ;
    input inputs_135__14 ;
    input inputs_135__13 ;
    input inputs_135__12 ;
    input inputs_135__11 ;
    input inputs_135__10 ;
    input inputs_135__9 ;
    input inputs_135__8 ;
    input inputs_135__7 ;
    input inputs_135__6 ;
    input inputs_135__5 ;
    input inputs_135__4 ;
    input inputs_135__3 ;
    input inputs_135__2 ;
    input inputs_135__1 ;
    input inputs_135__0 ;
    input inputs_136__15 ;
    input inputs_136__14 ;
    input inputs_136__13 ;
    input inputs_136__12 ;
    input inputs_136__11 ;
    input inputs_136__10 ;
    input inputs_136__9 ;
    input inputs_136__8 ;
    input inputs_136__7 ;
    input inputs_136__6 ;
    input inputs_136__5 ;
    input inputs_136__4 ;
    input inputs_136__3 ;
    input inputs_136__2 ;
    input inputs_136__1 ;
    input inputs_136__0 ;
    input inputs_137__15 ;
    input inputs_137__14 ;
    input inputs_137__13 ;
    input inputs_137__12 ;
    input inputs_137__11 ;
    input inputs_137__10 ;
    input inputs_137__9 ;
    input inputs_137__8 ;
    input inputs_137__7 ;
    input inputs_137__6 ;
    input inputs_137__5 ;
    input inputs_137__4 ;
    input inputs_137__3 ;
    input inputs_137__2 ;
    input inputs_137__1 ;
    input inputs_137__0 ;
    input inputs_138__15 ;
    input inputs_138__14 ;
    input inputs_138__13 ;
    input inputs_138__12 ;
    input inputs_138__11 ;
    input inputs_138__10 ;
    input inputs_138__9 ;
    input inputs_138__8 ;
    input inputs_138__7 ;
    input inputs_138__6 ;
    input inputs_138__5 ;
    input inputs_138__4 ;
    input inputs_138__3 ;
    input inputs_138__2 ;
    input inputs_138__1 ;
    input inputs_138__0 ;
    input inputs_139__15 ;
    input inputs_139__14 ;
    input inputs_139__13 ;
    input inputs_139__12 ;
    input inputs_139__11 ;
    input inputs_139__10 ;
    input inputs_139__9 ;
    input inputs_139__8 ;
    input inputs_139__7 ;
    input inputs_139__6 ;
    input inputs_139__5 ;
    input inputs_139__4 ;
    input inputs_139__3 ;
    input inputs_139__2 ;
    input inputs_139__1 ;
    input inputs_139__0 ;
    input inputs_140__15 ;
    input inputs_140__14 ;
    input inputs_140__13 ;
    input inputs_140__12 ;
    input inputs_140__11 ;
    input inputs_140__10 ;
    input inputs_140__9 ;
    input inputs_140__8 ;
    input inputs_140__7 ;
    input inputs_140__6 ;
    input inputs_140__5 ;
    input inputs_140__4 ;
    input inputs_140__3 ;
    input inputs_140__2 ;
    input inputs_140__1 ;
    input inputs_140__0 ;
    input inputs_141__15 ;
    input inputs_141__14 ;
    input inputs_141__13 ;
    input inputs_141__12 ;
    input inputs_141__11 ;
    input inputs_141__10 ;
    input inputs_141__9 ;
    input inputs_141__8 ;
    input inputs_141__7 ;
    input inputs_141__6 ;
    input inputs_141__5 ;
    input inputs_141__4 ;
    input inputs_141__3 ;
    input inputs_141__2 ;
    input inputs_141__1 ;
    input inputs_141__0 ;
    input inputs_142__15 ;
    input inputs_142__14 ;
    input inputs_142__13 ;
    input inputs_142__12 ;
    input inputs_142__11 ;
    input inputs_142__10 ;
    input inputs_142__9 ;
    input inputs_142__8 ;
    input inputs_142__7 ;
    input inputs_142__6 ;
    input inputs_142__5 ;
    input inputs_142__4 ;
    input inputs_142__3 ;
    input inputs_142__2 ;
    input inputs_142__1 ;
    input inputs_142__0 ;
    input inputs_143__15 ;
    input inputs_143__14 ;
    input inputs_143__13 ;
    input inputs_143__12 ;
    input inputs_143__11 ;
    input inputs_143__10 ;
    input inputs_143__9 ;
    input inputs_143__8 ;
    input inputs_143__7 ;
    input inputs_143__6 ;
    input inputs_143__5 ;
    input inputs_143__4 ;
    input inputs_143__3 ;
    input inputs_143__2 ;
    input inputs_143__1 ;
    input inputs_143__0 ;
    input inputs_144__15 ;
    input inputs_144__14 ;
    input inputs_144__13 ;
    input inputs_144__12 ;
    input inputs_144__11 ;
    input inputs_144__10 ;
    input inputs_144__9 ;
    input inputs_144__8 ;
    input inputs_144__7 ;
    input inputs_144__6 ;
    input inputs_144__5 ;
    input inputs_144__4 ;
    input inputs_144__3 ;
    input inputs_144__2 ;
    input inputs_144__1 ;
    input inputs_144__0 ;
    input inputs_145__15 ;
    input inputs_145__14 ;
    input inputs_145__13 ;
    input inputs_145__12 ;
    input inputs_145__11 ;
    input inputs_145__10 ;
    input inputs_145__9 ;
    input inputs_145__8 ;
    input inputs_145__7 ;
    input inputs_145__6 ;
    input inputs_145__5 ;
    input inputs_145__4 ;
    input inputs_145__3 ;
    input inputs_145__2 ;
    input inputs_145__1 ;
    input inputs_145__0 ;
    input inputs_146__15 ;
    input inputs_146__14 ;
    input inputs_146__13 ;
    input inputs_146__12 ;
    input inputs_146__11 ;
    input inputs_146__10 ;
    input inputs_146__9 ;
    input inputs_146__8 ;
    input inputs_146__7 ;
    input inputs_146__6 ;
    input inputs_146__5 ;
    input inputs_146__4 ;
    input inputs_146__3 ;
    input inputs_146__2 ;
    input inputs_146__1 ;
    input inputs_146__0 ;
    input inputs_147__15 ;
    input inputs_147__14 ;
    input inputs_147__13 ;
    input inputs_147__12 ;
    input inputs_147__11 ;
    input inputs_147__10 ;
    input inputs_147__9 ;
    input inputs_147__8 ;
    input inputs_147__7 ;
    input inputs_147__6 ;
    input inputs_147__5 ;
    input inputs_147__4 ;
    input inputs_147__3 ;
    input inputs_147__2 ;
    input inputs_147__1 ;
    input inputs_147__0 ;
    input inputs_148__15 ;
    input inputs_148__14 ;
    input inputs_148__13 ;
    input inputs_148__12 ;
    input inputs_148__11 ;
    input inputs_148__10 ;
    input inputs_148__9 ;
    input inputs_148__8 ;
    input inputs_148__7 ;
    input inputs_148__6 ;
    input inputs_148__5 ;
    input inputs_148__4 ;
    input inputs_148__3 ;
    input inputs_148__2 ;
    input inputs_148__1 ;
    input inputs_148__0 ;
    input inputs_149__15 ;
    input inputs_149__14 ;
    input inputs_149__13 ;
    input inputs_149__12 ;
    input inputs_149__11 ;
    input inputs_149__10 ;
    input inputs_149__9 ;
    input inputs_149__8 ;
    input inputs_149__7 ;
    input inputs_149__6 ;
    input inputs_149__5 ;
    input inputs_149__4 ;
    input inputs_149__3 ;
    input inputs_149__2 ;
    input inputs_149__1 ;
    input inputs_149__0 ;
    input inputs_150__15 ;
    input inputs_150__14 ;
    input inputs_150__13 ;
    input inputs_150__12 ;
    input inputs_150__11 ;
    input inputs_150__10 ;
    input inputs_150__9 ;
    input inputs_150__8 ;
    input inputs_150__7 ;
    input inputs_150__6 ;
    input inputs_150__5 ;
    input inputs_150__4 ;
    input inputs_150__3 ;
    input inputs_150__2 ;
    input inputs_150__1 ;
    input inputs_150__0 ;
    input inputs_151__15 ;
    input inputs_151__14 ;
    input inputs_151__13 ;
    input inputs_151__12 ;
    input inputs_151__11 ;
    input inputs_151__10 ;
    input inputs_151__9 ;
    input inputs_151__8 ;
    input inputs_151__7 ;
    input inputs_151__6 ;
    input inputs_151__5 ;
    input inputs_151__4 ;
    input inputs_151__3 ;
    input inputs_151__2 ;
    input inputs_151__1 ;
    input inputs_151__0 ;
    input inputs_152__15 ;
    input inputs_152__14 ;
    input inputs_152__13 ;
    input inputs_152__12 ;
    input inputs_152__11 ;
    input inputs_152__10 ;
    input inputs_152__9 ;
    input inputs_152__8 ;
    input inputs_152__7 ;
    input inputs_152__6 ;
    input inputs_152__5 ;
    input inputs_152__4 ;
    input inputs_152__3 ;
    input inputs_152__2 ;
    input inputs_152__1 ;
    input inputs_152__0 ;
    input inputs_153__15 ;
    input inputs_153__14 ;
    input inputs_153__13 ;
    input inputs_153__12 ;
    input inputs_153__11 ;
    input inputs_153__10 ;
    input inputs_153__9 ;
    input inputs_153__8 ;
    input inputs_153__7 ;
    input inputs_153__6 ;
    input inputs_153__5 ;
    input inputs_153__4 ;
    input inputs_153__3 ;
    input inputs_153__2 ;
    input inputs_153__1 ;
    input inputs_153__0 ;
    input inputs_154__15 ;
    input inputs_154__14 ;
    input inputs_154__13 ;
    input inputs_154__12 ;
    input inputs_154__11 ;
    input inputs_154__10 ;
    input inputs_154__9 ;
    input inputs_154__8 ;
    input inputs_154__7 ;
    input inputs_154__6 ;
    input inputs_154__5 ;
    input inputs_154__4 ;
    input inputs_154__3 ;
    input inputs_154__2 ;
    input inputs_154__1 ;
    input inputs_154__0 ;
    input inputs_155__15 ;
    input inputs_155__14 ;
    input inputs_155__13 ;
    input inputs_155__12 ;
    input inputs_155__11 ;
    input inputs_155__10 ;
    input inputs_155__9 ;
    input inputs_155__8 ;
    input inputs_155__7 ;
    input inputs_155__6 ;
    input inputs_155__5 ;
    input inputs_155__4 ;
    input inputs_155__3 ;
    input inputs_155__2 ;
    input inputs_155__1 ;
    input inputs_155__0 ;
    input inputs_156__15 ;
    input inputs_156__14 ;
    input inputs_156__13 ;
    input inputs_156__12 ;
    input inputs_156__11 ;
    input inputs_156__10 ;
    input inputs_156__9 ;
    input inputs_156__8 ;
    input inputs_156__7 ;
    input inputs_156__6 ;
    input inputs_156__5 ;
    input inputs_156__4 ;
    input inputs_156__3 ;
    input inputs_156__2 ;
    input inputs_156__1 ;
    input inputs_156__0 ;
    input inputs_157__15 ;
    input inputs_157__14 ;
    input inputs_157__13 ;
    input inputs_157__12 ;
    input inputs_157__11 ;
    input inputs_157__10 ;
    input inputs_157__9 ;
    input inputs_157__8 ;
    input inputs_157__7 ;
    input inputs_157__6 ;
    input inputs_157__5 ;
    input inputs_157__4 ;
    input inputs_157__3 ;
    input inputs_157__2 ;
    input inputs_157__1 ;
    input inputs_157__0 ;
    input inputs_158__15 ;
    input inputs_158__14 ;
    input inputs_158__13 ;
    input inputs_158__12 ;
    input inputs_158__11 ;
    input inputs_158__10 ;
    input inputs_158__9 ;
    input inputs_158__8 ;
    input inputs_158__7 ;
    input inputs_158__6 ;
    input inputs_158__5 ;
    input inputs_158__4 ;
    input inputs_158__3 ;
    input inputs_158__2 ;
    input inputs_158__1 ;
    input inputs_158__0 ;
    input inputs_159__15 ;
    input inputs_159__14 ;
    input inputs_159__13 ;
    input inputs_159__12 ;
    input inputs_159__11 ;
    input inputs_159__10 ;
    input inputs_159__9 ;
    input inputs_159__8 ;
    input inputs_159__7 ;
    input inputs_159__6 ;
    input inputs_159__5 ;
    input inputs_159__4 ;
    input inputs_159__3 ;
    input inputs_159__2 ;
    input inputs_159__1 ;
    input inputs_159__0 ;
    input inputs_160__15 ;
    input inputs_160__14 ;
    input inputs_160__13 ;
    input inputs_160__12 ;
    input inputs_160__11 ;
    input inputs_160__10 ;
    input inputs_160__9 ;
    input inputs_160__8 ;
    input inputs_160__7 ;
    input inputs_160__6 ;
    input inputs_160__5 ;
    input inputs_160__4 ;
    input inputs_160__3 ;
    input inputs_160__2 ;
    input inputs_160__1 ;
    input inputs_160__0 ;
    input inputs_161__15 ;
    input inputs_161__14 ;
    input inputs_161__13 ;
    input inputs_161__12 ;
    input inputs_161__11 ;
    input inputs_161__10 ;
    input inputs_161__9 ;
    input inputs_161__8 ;
    input inputs_161__7 ;
    input inputs_161__6 ;
    input inputs_161__5 ;
    input inputs_161__4 ;
    input inputs_161__3 ;
    input inputs_161__2 ;
    input inputs_161__1 ;
    input inputs_161__0 ;
    input inputs_162__15 ;
    input inputs_162__14 ;
    input inputs_162__13 ;
    input inputs_162__12 ;
    input inputs_162__11 ;
    input inputs_162__10 ;
    input inputs_162__9 ;
    input inputs_162__8 ;
    input inputs_162__7 ;
    input inputs_162__6 ;
    input inputs_162__5 ;
    input inputs_162__4 ;
    input inputs_162__3 ;
    input inputs_162__2 ;
    input inputs_162__1 ;
    input inputs_162__0 ;
    input inputs_163__15 ;
    input inputs_163__14 ;
    input inputs_163__13 ;
    input inputs_163__12 ;
    input inputs_163__11 ;
    input inputs_163__10 ;
    input inputs_163__9 ;
    input inputs_163__8 ;
    input inputs_163__7 ;
    input inputs_163__6 ;
    input inputs_163__5 ;
    input inputs_163__4 ;
    input inputs_163__3 ;
    input inputs_163__2 ;
    input inputs_163__1 ;
    input inputs_163__0 ;
    input inputs_164__15 ;
    input inputs_164__14 ;
    input inputs_164__13 ;
    input inputs_164__12 ;
    input inputs_164__11 ;
    input inputs_164__10 ;
    input inputs_164__9 ;
    input inputs_164__8 ;
    input inputs_164__7 ;
    input inputs_164__6 ;
    input inputs_164__5 ;
    input inputs_164__4 ;
    input inputs_164__3 ;
    input inputs_164__2 ;
    input inputs_164__1 ;
    input inputs_164__0 ;
    input inputs_165__15 ;
    input inputs_165__14 ;
    input inputs_165__13 ;
    input inputs_165__12 ;
    input inputs_165__11 ;
    input inputs_165__10 ;
    input inputs_165__9 ;
    input inputs_165__8 ;
    input inputs_165__7 ;
    input inputs_165__6 ;
    input inputs_165__5 ;
    input inputs_165__4 ;
    input inputs_165__3 ;
    input inputs_165__2 ;
    input inputs_165__1 ;
    input inputs_165__0 ;
    input inputs_166__15 ;
    input inputs_166__14 ;
    input inputs_166__13 ;
    input inputs_166__12 ;
    input inputs_166__11 ;
    input inputs_166__10 ;
    input inputs_166__9 ;
    input inputs_166__8 ;
    input inputs_166__7 ;
    input inputs_166__6 ;
    input inputs_166__5 ;
    input inputs_166__4 ;
    input inputs_166__3 ;
    input inputs_166__2 ;
    input inputs_166__1 ;
    input inputs_166__0 ;
    input inputs_167__15 ;
    input inputs_167__14 ;
    input inputs_167__13 ;
    input inputs_167__12 ;
    input inputs_167__11 ;
    input inputs_167__10 ;
    input inputs_167__9 ;
    input inputs_167__8 ;
    input inputs_167__7 ;
    input inputs_167__6 ;
    input inputs_167__5 ;
    input inputs_167__4 ;
    input inputs_167__3 ;
    input inputs_167__2 ;
    input inputs_167__1 ;
    input inputs_167__0 ;
    input inputs_168__15 ;
    input inputs_168__14 ;
    input inputs_168__13 ;
    input inputs_168__12 ;
    input inputs_168__11 ;
    input inputs_168__10 ;
    input inputs_168__9 ;
    input inputs_168__8 ;
    input inputs_168__7 ;
    input inputs_168__6 ;
    input inputs_168__5 ;
    input inputs_168__4 ;
    input inputs_168__3 ;
    input inputs_168__2 ;
    input inputs_168__1 ;
    input inputs_168__0 ;
    input inputs_169__15 ;
    input inputs_169__14 ;
    input inputs_169__13 ;
    input inputs_169__12 ;
    input inputs_169__11 ;
    input inputs_169__10 ;
    input inputs_169__9 ;
    input inputs_169__8 ;
    input inputs_169__7 ;
    input inputs_169__6 ;
    input inputs_169__5 ;
    input inputs_169__4 ;
    input inputs_169__3 ;
    input inputs_169__2 ;
    input inputs_169__1 ;
    input inputs_169__0 ;
    input inputs_170__15 ;
    input inputs_170__14 ;
    input inputs_170__13 ;
    input inputs_170__12 ;
    input inputs_170__11 ;
    input inputs_170__10 ;
    input inputs_170__9 ;
    input inputs_170__8 ;
    input inputs_170__7 ;
    input inputs_170__6 ;
    input inputs_170__5 ;
    input inputs_170__4 ;
    input inputs_170__3 ;
    input inputs_170__2 ;
    input inputs_170__1 ;
    input inputs_170__0 ;
    input inputs_171__15 ;
    input inputs_171__14 ;
    input inputs_171__13 ;
    input inputs_171__12 ;
    input inputs_171__11 ;
    input inputs_171__10 ;
    input inputs_171__9 ;
    input inputs_171__8 ;
    input inputs_171__7 ;
    input inputs_171__6 ;
    input inputs_171__5 ;
    input inputs_171__4 ;
    input inputs_171__3 ;
    input inputs_171__2 ;
    input inputs_171__1 ;
    input inputs_171__0 ;
    input inputs_172__15 ;
    input inputs_172__14 ;
    input inputs_172__13 ;
    input inputs_172__12 ;
    input inputs_172__11 ;
    input inputs_172__10 ;
    input inputs_172__9 ;
    input inputs_172__8 ;
    input inputs_172__7 ;
    input inputs_172__6 ;
    input inputs_172__5 ;
    input inputs_172__4 ;
    input inputs_172__3 ;
    input inputs_172__2 ;
    input inputs_172__1 ;
    input inputs_172__0 ;
    input inputs_173__15 ;
    input inputs_173__14 ;
    input inputs_173__13 ;
    input inputs_173__12 ;
    input inputs_173__11 ;
    input inputs_173__10 ;
    input inputs_173__9 ;
    input inputs_173__8 ;
    input inputs_173__7 ;
    input inputs_173__6 ;
    input inputs_173__5 ;
    input inputs_173__4 ;
    input inputs_173__3 ;
    input inputs_173__2 ;
    input inputs_173__1 ;
    input inputs_173__0 ;
    input inputs_174__15 ;
    input inputs_174__14 ;
    input inputs_174__13 ;
    input inputs_174__12 ;
    input inputs_174__11 ;
    input inputs_174__10 ;
    input inputs_174__9 ;
    input inputs_174__8 ;
    input inputs_174__7 ;
    input inputs_174__6 ;
    input inputs_174__5 ;
    input inputs_174__4 ;
    input inputs_174__3 ;
    input inputs_174__2 ;
    input inputs_174__1 ;
    input inputs_174__0 ;
    input inputs_175__15 ;
    input inputs_175__14 ;
    input inputs_175__13 ;
    input inputs_175__12 ;
    input inputs_175__11 ;
    input inputs_175__10 ;
    input inputs_175__9 ;
    input inputs_175__8 ;
    input inputs_175__7 ;
    input inputs_175__6 ;
    input inputs_175__5 ;
    input inputs_175__4 ;
    input inputs_175__3 ;
    input inputs_175__2 ;
    input inputs_175__1 ;
    input inputs_175__0 ;
    input inputs_176__15 ;
    input inputs_176__14 ;
    input inputs_176__13 ;
    input inputs_176__12 ;
    input inputs_176__11 ;
    input inputs_176__10 ;
    input inputs_176__9 ;
    input inputs_176__8 ;
    input inputs_176__7 ;
    input inputs_176__6 ;
    input inputs_176__5 ;
    input inputs_176__4 ;
    input inputs_176__3 ;
    input inputs_176__2 ;
    input inputs_176__1 ;
    input inputs_176__0 ;
    input inputs_177__15 ;
    input inputs_177__14 ;
    input inputs_177__13 ;
    input inputs_177__12 ;
    input inputs_177__11 ;
    input inputs_177__10 ;
    input inputs_177__9 ;
    input inputs_177__8 ;
    input inputs_177__7 ;
    input inputs_177__6 ;
    input inputs_177__5 ;
    input inputs_177__4 ;
    input inputs_177__3 ;
    input inputs_177__2 ;
    input inputs_177__1 ;
    input inputs_177__0 ;
    input inputs_178__15 ;
    input inputs_178__14 ;
    input inputs_178__13 ;
    input inputs_178__12 ;
    input inputs_178__11 ;
    input inputs_178__10 ;
    input inputs_178__9 ;
    input inputs_178__8 ;
    input inputs_178__7 ;
    input inputs_178__6 ;
    input inputs_178__5 ;
    input inputs_178__4 ;
    input inputs_178__3 ;
    input inputs_178__2 ;
    input inputs_178__1 ;
    input inputs_178__0 ;
    input inputs_179__15 ;
    input inputs_179__14 ;
    input inputs_179__13 ;
    input inputs_179__12 ;
    input inputs_179__11 ;
    input inputs_179__10 ;
    input inputs_179__9 ;
    input inputs_179__8 ;
    input inputs_179__7 ;
    input inputs_179__6 ;
    input inputs_179__5 ;
    input inputs_179__4 ;
    input inputs_179__3 ;
    input inputs_179__2 ;
    input inputs_179__1 ;
    input inputs_179__0 ;
    input inputs_180__15 ;
    input inputs_180__14 ;
    input inputs_180__13 ;
    input inputs_180__12 ;
    input inputs_180__11 ;
    input inputs_180__10 ;
    input inputs_180__9 ;
    input inputs_180__8 ;
    input inputs_180__7 ;
    input inputs_180__6 ;
    input inputs_180__5 ;
    input inputs_180__4 ;
    input inputs_180__3 ;
    input inputs_180__2 ;
    input inputs_180__1 ;
    input inputs_180__0 ;
    input inputs_181__15 ;
    input inputs_181__14 ;
    input inputs_181__13 ;
    input inputs_181__12 ;
    input inputs_181__11 ;
    input inputs_181__10 ;
    input inputs_181__9 ;
    input inputs_181__8 ;
    input inputs_181__7 ;
    input inputs_181__6 ;
    input inputs_181__5 ;
    input inputs_181__4 ;
    input inputs_181__3 ;
    input inputs_181__2 ;
    input inputs_181__1 ;
    input inputs_181__0 ;
    input inputs_182__15 ;
    input inputs_182__14 ;
    input inputs_182__13 ;
    input inputs_182__12 ;
    input inputs_182__11 ;
    input inputs_182__10 ;
    input inputs_182__9 ;
    input inputs_182__8 ;
    input inputs_182__7 ;
    input inputs_182__6 ;
    input inputs_182__5 ;
    input inputs_182__4 ;
    input inputs_182__3 ;
    input inputs_182__2 ;
    input inputs_182__1 ;
    input inputs_182__0 ;
    input inputs_183__15 ;
    input inputs_183__14 ;
    input inputs_183__13 ;
    input inputs_183__12 ;
    input inputs_183__11 ;
    input inputs_183__10 ;
    input inputs_183__9 ;
    input inputs_183__8 ;
    input inputs_183__7 ;
    input inputs_183__6 ;
    input inputs_183__5 ;
    input inputs_183__4 ;
    input inputs_183__3 ;
    input inputs_183__2 ;
    input inputs_183__1 ;
    input inputs_183__0 ;
    input inputs_184__15 ;
    input inputs_184__14 ;
    input inputs_184__13 ;
    input inputs_184__12 ;
    input inputs_184__11 ;
    input inputs_184__10 ;
    input inputs_184__9 ;
    input inputs_184__8 ;
    input inputs_184__7 ;
    input inputs_184__6 ;
    input inputs_184__5 ;
    input inputs_184__4 ;
    input inputs_184__3 ;
    input inputs_184__2 ;
    input inputs_184__1 ;
    input inputs_184__0 ;
    input inputs_185__15 ;
    input inputs_185__14 ;
    input inputs_185__13 ;
    input inputs_185__12 ;
    input inputs_185__11 ;
    input inputs_185__10 ;
    input inputs_185__9 ;
    input inputs_185__8 ;
    input inputs_185__7 ;
    input inputs_185__6 ;
    input inputs_185__5 ;
    input inputs_185__4 ;
    input inputs_185__3 ;
    input inputs_185__2 ;
    input inputs_185__1 ;
    input inputs_185__0 ;
    input inputs_186__15 ;
    input inputs_186__14 ;
    input inputs_186__13 ;
    input inputs_186__12 ;
    input inputs_186__11 ;
    input inputs_186__10 ;
    input inputs_186__9 ;
    input inputs_186__8 ;
    input inputs_186__7 ;
    input inputs_186__6 ;
    input inputs_186__5 ;
    input inputs_186__4 ;
    input inputs_186__3 ;
    input inputs_186__2 ;
    input inputs_186__1 ;
    input inputs_186__0 ;
    input inputs_187__15 ;
    input inputs_187__14 ;
    input inputs_187__13 ;
    input inputs_187__12 ;
    input inputs_187__11 ;
    input inputs_187__10 ;
    input inputs_187__9 ;
    input inputs_187__8 ;
    input inputs_187__7 ;
    input inputs_187__6 ;
    input inputs_187__5 ;
    input inputs_187__4 ;
    input inputs_187__3 ;
    input inputs_187__2 ;
    input inputs_187__1 ;
    input inputs_187__0 ;
    input inputs_188__15 ;
    input inputs_188__14 ;
    input inputs_188__13 ;
    input inputs_188__12 ;
    input inputs_188__11 ;
    input inputs_188__10 ;
    input inputs_188__9 ;
    input inputs_188__8 ;
    input inputs_188__7 ;
    input inputs_188__6 ;
    input inputs_188__5 ;
    input inputs_188__4 ;
    input inputs_188__3 ;
    input inputs_188__2 ;
    input inputs_188__1 ;
    input inputs_188__0 ;
    input inputs_189__15 ;
    input inputs_189__14 ;
    input inputs_189__13 ;
    input inputs_189__12 ;
    input inputs_189__11 ;
    input inputs_189__10 ;
    input inputs_189__9 ;
    input inputs_189__8 ;
    input inputs_189__7 ;
    input inputs_189__6 ;
    input inputs_189__5 ;
    input inputs_189__4 ;
    input inputs_189__3 ;
    input inputs_189__2 ;
    input inputs_189__1 ;
    input inputs_189__0 ;
    input inputs_190__15 ;
    input inputs_190__14 ;
    input inputs_190__13 ;
    input inputs_190__12 ;
    input inputs_190__11 ;
    input inputs_190__10 ;
    input inputs_190__9 ;
    input inputs_190__8 ;
    input inputs_190__7 ;
    input inputs_190__6 ;
    input inputs_190__5 ;
    input inputs_190__4 ;
    input inputs_190__3 ;
    input inputs_190__2 ;
    input inputs_190__1 ;
    input inputs_190__0 ;
    input inputs_191__15 ;
    input inputs_191__14 ;
    input inputs_191__13 ;
    input inputs_191__12 ;
    input inputs_191__11 ;
    input inputs_191__10 ;
    input inputs_191__9 ;
    input inputs_191__8 ;
    input inputs_191__7 ;
    input inputs_191__6 ;
    input inputs_191__5 ;
    input inputs_191__4 ;
    input inputs_191__3 ;
    input inputs_191__2 ;
    input inputs_191__1 ;
    input inputs_191__0 ;
    input inputs_192__15 ;
    input inputs_192__14 ;
    input inputs_192__13 ;
    input inputs_192__12 ;
    input inputs_192__11 ;
    input inputs_192__10 ;
    input inputs_192__9 ;
    input inputs_192__8 ;
    input inputs_192__7 ;
    input inputs_192__6 ;
    input inputs_192__5 ;
    input inputs_192__4 ;
    input inputs_192__3 ;
    input inputs_192__2 ;
    input inputs_192__1 ;
    input inputs_192__0 ;
    input inputs_193__15 ;
    input inputs_193__14 ;
    input inputs_193__13 ;
    input inputs_193__12 ;
    input inputs_193__11 ;
    input inputs_193__10 ;
    input inputs_193__9 ;
    input inputs_193__8 ;
    input inputs_193__7 ;
    input inputs_193__6 ;
    input inputs_193__5 ;
    input inputs_193__4 ;
    input inputs_193__3 ;
    input inputs_193__2 ;
    input inputs_193__1 ;
    input inputs_193__0 ;
    input inputs_194__15 ;
    input inputs_194__14 ;
    input inputs_194__13 ;
    input inputs_194__12 ;
    input inputs_194__11 ;
    input inputs_194__10 ;
    input inputs_194__9 ;
    input inputs_194__8 ;
    input inputs_194__7 ;
    input inputs_194__6 ;
    input inputs_194__5 ;
    input inputs_194__4 ;
    input inputs_194__3 ;
    input inputs_194__2 ;
    input inputs_194__1 ;
    input inputs_194__0 ;
    input inputs_195__15 ;
    input inputs_195__14 ;
    input inputs_195__13 ;
    input inputs_195__12 ;
    input inputs_195__11 ;
    input inputs_195__10 ;
    input inputs_195__9 ;
    input inputs_195__8 ;
    input inputs_195__7 ;
    input inputs_195__6 ;
    input inputs_195__5 ;
    input inputs_195__4 ;
    input inputs_195__3 ;
    input inputs_195__2 ;
    input inputs_195__1 ;
    input inputs_195__0 ;
    input inputs_196__15 ;
    input inputs_196__14 ;
    input inputs_196__13 ;
    input inputs_196__12 ;
    input inputs_196__11 ;
    input inputs_196__10 ;
    input inputs_196__9 ;
    input inputs_196__8 ;
    input inputs_196__7 ;
    input inputs_196__6 ;
    input inputs_196__5 ;
    input inputs_196__4 ;
    input inputs_196__3 ;
    input inputs_196__2 ;
    input inputs_196__1 ;
    input inputs_196__0 ;
    input inputs_197__15 ;
    input inputs_197__14 ;
    input inputs_197__13 ;
    input inputs_197__12 ;
    input inputs_197__11 ;
    input inputs_197__10 ;
    input inputs_197__9 ;
    input inputs_197__8 ;
    input inputs_197__7 ;
    input inputs_197__6 ;
    input inputs_197__5 ;
    input inputs_197__4 ;
    input inputs_197__3 ;
    input inputs_197__2 ;
    input inputs_197__1 ;
    input inputs_197__0 ;
    input inputs_198__15 ;
    input inputs_198__14 ;
    input inputs_198__13 ;
    input inputs_198__12 ;
    input inputs_198__11 ;
    input inputs_198__10 ;
    input inputs_198__9 ;
    input inputs_198__8 ;
    input inputs_198__7 ;
    input inputs_198__6 ;
    input inputs_198__5 ;
    input inputs_198__4 ;
    input inputs_198__3 ;
    input inputs_198__2 ;
    input inputs_198__1 ;
    input inputs_198__0 ;
    input inputs_199__15 ;
    input inputs_199__14 ;
    input inputs_199__13 ;
    input inputs_199__12 ;
    input inputs_199__11 ;
    input inputs_199__10 ;
    input inputs_199__9 ;
    input inputs_199__8 ;
    input inputs_199__7 ;
    input inputs_199__6 ;
    input inputs_199__5 ;
    input inputs_199__4 ;
    input inputs_199__3 ;
    input inputs_199__2 ;
    input inputs_199__1 ;
    input inputs_199__0 ;
    input inputs_200__15 ;
    input inputs_200__14 ;
    input inputs_200__13 ;
    input inputs_200__12 ;
    input inputs_200__11 ;
    input inputs_200__10 ;
    input inputs_200__9 ;
    input inputs_200__8 ;
    input inputs_200__7 ;
    input inputs_200__6 ;
    input inputs_200__5 ;
    input inputs_200__4 ;
    input inputs_200__3 ;
    input inputs_200__2 ;
    input inputs_200__1 ;
    input inputs_200__0 ;
    input inputs_201__15 ;
    input inputs_201__14 ;
    input inputs_201__13 ;
    input inputs_201__12 ;
    input inputs_201__11 ;
    input inputs_201__10 ;
    input inputs_201__9 ;
    input inputs_201__8 ;
    input inputs_201__7 ;
    input inputs_201__6 ;
    input inputs_201__5 ;
    input inputs_201__4 ;
    input inputs_201__3 ;
    input inputs_201__2 ;
    input inputs_201__1 ;
    input inputs_201__0 ;
    input inputs_202__15 ;
    input inputs_202__14 ;
    input inputs_202__13 ;
    input inputs_202__12 ;
    input inputs_202__11 ;
    input inputs_202__10 ;
    input inputs_202__9 ;
    input inputs_202__8 ;
    input inputs_202__7 ;
    input inputs_202__6 ;
    input inputs_202__5 ;
    input inputs_202__4 ;
    input inputs_202__3 ;
    input inputs_202__2 ;
    input inputs_202__1 ;
    input inputs_202__0 ;
    input inputs_203__15 ;
    input inputs_203__14 ;
    input inputs_203__13 ;
    input inputs_203__12 ;
    input inputs_203__11 ;
    input inputs_203__10 ;
    input inputs_203__9 ;
    input inputs_203__8 ;
    input inputs_203__7 ;
    input inputs_203__6 ;
    input inputs_203__5 ;
    input inputs_203__4 ;
    input inputs_203__3 ;
    input inputs_203__2 ;
    input inputs_203__1 ;
    input inputs_203__0 ;
    input inputs_204__15 ;
    input inputs_204__14 ;
    input inputs_204__13 ;
    input inputs_204__12 ;
    input inputs_204__11 ;
    input inputs_204__10 ;
    input inputs_204__9 ;
    input inputs_204__8 ;
    input inputs_204__7 ;
    input inputs_204__6 ;
    input inputs_204__5 ;
    input inputs_204__4 ;
    input inputs_204__3 ;
    input inputs_204__2 ;
    input inputs_204__1 ;
    input inputs_204__0 ;
    input inputs_205__15 ;
    input inputs_205__14 ;
    input inputs_205__13 ;
    input inputs_205__12 ;
    input inputs_205__11 ;
    input inputs_205__10 ;
    input inputs_205__9 ;
    input inputs_205__8 ;
    input inputs_205__7 ;
    input inputs_205__6 ;
    input inputs_205__5 ;
    input inputs_205__4 ;
    input inputs_205__3 ;
    input inputs_205__2 ;
    input inputs_205__1 ;
    input inputs_205__0 ;
    input inputs_206__15 ;
    input inputs_206__14 ;
    input inputs_206__13 ;
    input inputs_206__12 ;
    input inputs_206__11 ;
    input inputs_206__10 ;
    input inputs_206__9 ;
    input inputs_206__8 ;
    input inputs_206__7 ;
    input inputs_206__6 ;
    input inputs_206__5 ;
    input inputs_206__4 ;
    input inputs_206__3 ;
    input inputs_206__2 ;
    input inputs_206__1 ;
    input inputs_206__0 ;
    input inputs_207__15 ;
    input inputs_207__14 ;
    input inputs_207__13 ;
    input inputs_207__12 ;
    input inputs_207__11 ;
    input inputs_207__10 ;
    input inputs_207__9 ;
    input inputs_207__8 ;
    input inputs_207__7 ;
    input inputs_207__6 ;
    input inputs_207__5 ;
    input inputs_207__4 ;
    input inputs_207__3 ;
    input inputs_207__2 ;
    input inputs_207__1 ;
    input inputs_207__0 ;
    input inputs_208__15 ;
    input inputs_208__14 ;
    input inputs_208__13 ;
    input inputs_208__12 ;
    input inputs_208__11 ;
    input inputs_208__10 ;
    input inputs_208__9 ;
    input inputs_208__8 ;
    input inputs_208__7 ;
    input inputs_208__6 ;
    input inputs_208__5 ;
    input inputs_208__4 ;
    input inputs_208__3 ;
    input inputs_208__2 ;
    input inputs_208__1 ;
    input inputs_208__0 ;
    input inputs_209__15 ;
    input inputs_209__14 ;
    input inputs_209__13 ;
    input inputs_209__12 ;
    input inputs_209__11 ;
    input inputs_209__10 ;
    input inputs_209__9 ;
    input inputs_209__8 ;
    input inputs_209__7 ;
    input inputs_209__6 ;
    input inputs_209__5 ;
    input inputs_209__4 ;
    input inputs_209__3 ;
    input inputs_209__2 ;
    input inputs_209__1 ;
    input inputs_209__0 ;
    input inputs_210__15 ;
    input inputs_210__14 ;
    input inputs_210__13 ;
    input inputs_210__12 ;
    input inputs_210__11 ;
    input inputs_210__10 ;
    input inputs_210__9 ;
    input inputs_210__8 ;
    input inputs_210__7 ;
    input inputs_210__6 ;
    input inputs_210__5 ;
    input inputs_210__4 ;
    input inputs_210__3 ;
    input inputs_210__2 ;
    input inputs_210__1 ;
    input inputs_210__0 ;
    input inputs_211__15 ;
    input inputs_211__14 ;
    input inputs_211__13 ;
    input inputs_211__12 ;
    input inputs_211__11 ;
    input inputs_211__10 ;
    input inputs_211__9 ;
    input inputs_211__8 ;
    input inputs_211__7 ;
    input inputs_211__6 ;
    input inputs_211__5 ;
    input inputs_211__4 ;
    input inputs_211__3 ;
    input inputs_211__2 ;
    input inputs_211__1 ;
    input inputs_211__0 ;
    input inputs_212__15 ;
    input inputs_212__14 ;
    input inputs_212__13 ;
    input inputs_212__12 ;
    input inputs_212__11 ;
    input inputs_212__10 ;
    input inputs_212__9 ;
    input inputs_212__8 ;
    input inputs_212__7 ;
    input inputs_212__6 ;
    input inputs_212__5 ;
    input inputs_212__4 ;
    input inputs_212__3 ;
    input inputs_212__2 ;
    input inputs_212__1 ;
    input inputs_212__0 ;
    input inputs_213__15 ;
    input inputs_213__14 ;
    input inputs_213__13 ;
    input inputs_213__12 ;
    input inputs_213__11 ;
    input inputs_213__10 ;
    input inputs_213__9 ;
    input inputs_213__8 ;
    input inputs_213__7 ;
    input inputs_213__6 ;
    input inputs_213__5 ;
    input inputs_213__4 ;
    input inputs_213__3 ;
    input inputs_213__2 ;
    input inputs_213__1 ;
    input inputs_213__0 ;
    input inputs_214__15 ;
    input inputs_214__14 ;
    input inputs_214__13 ;
    input inputs_214__12 ;
    input inputs_214__11 ;
    input inputs_214__10 ;
    input inputs_214__9 ;
    input inputs_214__8 ;
    input inputs_214__7 ;
    input inputs_214__6 ;
    input inputs_214__5 ;
    input inputs_214__4 ;
    input inputs_214__3 ;
    input inputs_214__2 ;
    input inputs_214__1 ;
    input inputs_214__0 ;
    input inputs_215__15 ;
    input inputs_215__14 ;
    input inputs_215__13 ;
    input inputs_215__12 ;
    input inputs_215__11 ;
    input inputs_215__10 ;
    input inputs_215__9 ;
    input inputs_215__8 ;
    input inputs_215__7 ;
    input inputs_215__6 ;
    input inputs_215__5 ;
    input inputs_215__4 ;
    input inputs_215__3 ;
    input inputs_215__2 ;
    input inputs_215__1 ;
    input inputs_215__0 ;
    input inputs_216__15 ;
    input inputs_216__14 ;
    input inputs_216__13 ;
    input inputs_216__12 ;
    input inputs_216__11 ;
    input inputs_216__10 ;
    input inputs_216__9 ;
    input inputs_216__8 ;
    input inputs_216__7 ;
    input inputs_216__6 ;
    input inputs_216__5 ;
    input inputs_216__4 ;
    input inputs_216__3 ;
    input inputs_216__2 ;
    input inputs_216__1 ;
    input inputs_216__0 ;
    input inputs_217__15 ;
    input inputs_217__14 ;
    input inputs_217__13 ;
    input inputs_217__12 ;
    input inputs_217__11 ;
    input inputs_217__10 ;
    input inputs_217__9 ;
    input inputs_217__8 ;
    input inputs_217__7 ;
    input inputs_217__6 ;
    input inputs_217__5 ;
    input inputs_217__4 ;
    input inputs_217__3 ;
    input inputs_217__2 ;
    input inputs_217__1 ;
    input inputs_217__0 ;
    input inputs_218__15 ;
    input inputs_218__14 ;
    input inputs_218__13 ;
    input inputs_218__12 ;
    input inputs_218__11 ;
    input inputs_218__10 ;
    input inputs_218__9 ;
    input inputs_218__8 ;
    input inputs_218__7 ;
    input inputs_218__6 ;
    input inputs_218__5 ;
    input inputs_218__4 ;
    input inputs_218__3 ;
    input inputs_218__2 ;
    input inputs_218__1 ;
    input inputs_218__0 ;
    input inputs_219__15 ;
    input inputs_219__14 ;
    input inputs_219__13 ;
    input inputs_219__12 ;
    input inputs_219__11 ;
    input inputs_219__10 ;
    input inputs_219__9 ;
    input inputs_219__8 ;
    input inputs_219__7 ;
    input inputs_219__6 ;
    input inputs_219__5 ;
    input inputs_219__4 ;
    input inputs_219__3 ;
    input inputs_219__2 ;
    input inputs_219__1 ;
    input inputs_219__0 ;
    input inputs_220__15 ;
    input inputs_220__14 ;
    input inputs_220__13 ;
    input inputs_220__12 ;
    input inputs_220__11 ;
    input inputs_220__10 ;
    input inputs_220__9 ;
    input inputs_220__8 ;
    input inputs_220__7 ;
    input inputs_220__6 ;
    input inputs_220__5 ;
    input inputs_220__4 ;
    input inputs_220__3 ;
    input inputs_220__2 ;
    input inputs_220__1 ;
    input inputs_220__0 ;
    input inputs_221__15 ;
    input inputs_221__14 ;
    input inputs_221__13 ;
    input inputs_221__12 ;
    input inputs_221__11 ;
    input inputs_221__10 ;
    input inputs_221__9 ;
    input inputs_221__8 ;
    input inputs_221__7 ;
    input inputs_221__6 ;
    input inputs_221__5 ;
    input inputs_221__4 ;
    input inputs_221__3 ;
    input inputs_221__2 ;
    input inputs_221__1 ;
    input inputs_221__0 ;
    input inputs_222__15 ;
    input inputs_222__14 ;
    input inputs_222__13 ;
    input inputs_222__12 ;
    input inputs_222__11 ;
    input inputs_222__10 ;
    input inputs_222__9 ;
    input inputs_222__8 ;
    input inputs_222__7 ;
    input inputs_222__6 ;
    input inputs_222__5 ;
    input inputs_222__4 ;
    input inputs_222__3 ;
    input inputs_222__2 ;
    input inputs_222__1 ;
    input inputs_222__0 ;
    input inputs_223__15 ;
    input inputs_223__14 ;
    input inputs_223__13 ;
    input inputs_223__12 ;
    input inputs_223__11 ;
    input inputs_223__10 ;
    input inputs_223__9 ;
    input inputs_223__8 ;
    input inputs_223__7 ;
    input inputs_223__6 ;
    input inputs_223__5 ;
    input inputs_223__4 ;
    input inputs_223__3 ;
    input inputs_223__2 ;
    input inputs_223__1 ;
    input inputs_223__0 ;
    input inputs_224__15 ;
    input inputs_224__14 ;
    input inputs_224__13 ;
    input inputs_224__12 ;
    input inputs_224__11 ;
    input inputs_224__10 ;
    input inputs_224__9 ;
    input inputs_224__8 ;
    input inputs_224__7 ;
    input inputs_224__6 ;
    input inputs_224__5 ;
    input inputs_224__4 ;
    input inputs_224__3 ;
    input inputs_224__2 ;
    input inputs_224__1 ;
    input inputs_224__0 ;
    input inputs_225__15 ;
    input inputs_225__14 ;
    input inputs_225__13 ;
    input inputs_225__12 ;
    input inputs_225__11 ;
    input inputs_225__10 ;
    input inputs_225__9 ;
    input inputs_225__8 ;
    input inputs_225__7 ;
    input inputs_225__6 ;
    input inputs_225__5 ;
    input inputs_225__4 ;
    input inputs_225__3 ;
    input inputs_225__2 ;
    input inputs_225__1 ;
    input inputs_225__0 ;
    input inputs_226__15 ;
    input inputs_226__14 ;
    input inputs_226__13 ;
    input inputs_226__12 ;
    input inputs_226__11 ;
    input inputs_226__10 ;
    input inputs_226__9 ;
    input inputs_226__8 ;
    input inputs_226__7 ;
    input inputs_226__6 ;
    input inputs_226__5 ;
    input inputs_226__4 ;
    input inputs_226__3 ;
    input inputs_226__2 ;
    input inputs_226__1 ;
    input inputs_226__0 ;
    input inputs_227__15 ;
    input inputs_227__14 ;
    input inputs_227__13 ;
    input inputs_227__12 ;
    input inputs_227__11 ;
    input inputs_227__10 ;
    input inputs_227__9 ;
    input inputs_227__8 ;
    input inputs_227__7 ;
    input inputs_227__6 ;
    input inputs_227__5 ;
    input inputs_227__4 ;
    input inputs_227__3 ;
    input inputs_227__2 ;
    input inputs_227__1 ;
    input inputs_227__0 ;
    input inputs_228__15 ;
    input inputs_228__14 ;
    input inputs_228__13 ;
    input inputs_228__12 ;
    input inputs_228__11 ;
    input inputs_228__10 ;
    input inputs_228__9 ;
    input inputs_228__8 ;
    input inputs_228__7 ;
    input inputs_228__6 ;
    input inputs_228__5 ;
    input inputs_228__4 ;
    input inputs_228__3 ;
    input inputs_228__2 ;
    input inputs_228__1 ;
    input inputs_228__0 ;
    input inputs_229__15 ;
    input inputs_229__14 ;
    input inputs_229__13 ;
    input inputs_229__12 ;
    input inputs_229__11 ;
    input inputs_229__10 ;
    input inputs_229__9 ;
    input inputs_229__8 ;
    input inputs_229__7 ;
    input inputs_229__6 ;
    input inputs_229__5 ;
    input inputs_229__4 ;
    input inputs_229__3 ;
    input inputs_229__2 ;
    input inputs_229__1 ;
    input inputs_229__0 ;
    input inputs_230__15 ;
    input inputs_230__14 ;
    input inputs_230__13 ;
    input inputs_230__12 ;
    input inputs_230__11 ;
    input inputs_230__10 ;
    input inputs_230__9 ;
    input inputs_230__8 ;
    input inputs_230__7 ;
    input inputs_230__6 ;
    input inputs_230__5 ;
    input inputs_230__4 ;
    input inputs_230__3 ;
    input inputs_230__2 ;
    input inputs_230__1 ;
    input inputs_230__0 ;
    input inputs_231__15 ;
    input inputs_231__14 ;
    input inputs_231__13 ;
    input inputs_231__12 ;
    input inputs_231__11 ;
    input inputs_231__10 ;
    input inputs_231__9 ;
    input inputs_231__8 ;
    input inputs_231__7 ;
    input inputs_231__6 ;
    input inputs_231__5 ;
    input inputs_231__4 ;
    input inputs_231__3 ;
    input inputs_231__2 ;
    input inputs_231__1 ;
    input inputs_231__0 ;
    input inputs_232__15 ;
    input inputs_232__14 ;
    input inputs_232__13 ;
    input inputs_232__12 ;
    input inputs_232__11 ;
    input inputs_232__10 ;
    input inputs_232__9 ;
    input inputs_232__8 ;
    input inputs_232__7 ;
    input inputs_232__6 ;
    input inputs_232__5 ;
    input inputs_232__4 ;
    input inputs_232__3 ;
    input inputs_232__2 ;
    input inputs_232__1 ;
    input inputs_232__0 ;
    input inputs_233__15 ;
    input inputs_233__14 ;
    input inputs_233__13 ;
    input inputs_233__12 ;
    input inputs_233__11 ;
    input inputs_233__10 ;
    input inputs_233__9 ;
    input inputs_233__8 ;
    input inputs_233__7 ;
    input inputs_233__6 ;
    input inputs_233__5 ;
    input inputs_233__4 ;
    input inputs_233__3 ;
    input inputs_233__2 ;
    input inputs_233__1 ;
    input inputs_233__0 ;
    input inputs_234__15 ;
    input inputs_234__14 ;
    input inputs_234__13 ;
    input inputs_234__12 ;
    input inputs_234__11 ;
    input inputs_234__10 ;
    input inputs_234__9 ;
    input inputs_234__8 ;
    input inputs_234__7 ;
    input inputs_234__6 ;
    input inputs_234__5 ;
    input inputs_234__4 ;
    input inputs_234__3 ;
    input inputs_234__2 ;
    input inputs_234__1 ;
    input inputs_234__0 ;
    input inputs_235__15 ;
    input inputs_235__14 ;
    input inputs_235__13 ;
    input inputs_235__12 ;
    input inputs_235__11 ;
    input inputs_235__10 ;
    input inputs_235__9 ;
    input inputs_235__8 ;
    input inputs_235__7 ;
    input inputs_235__6 ;
    input inputs_235__5 ;
    input inputs_235__4 ;
    input inputs_235__3 ;
    input inputs_235__2 ;
    input inputs_235__1 ;
    input inputs_235__0 ;
    input inputs_236__15 ;
    input inputs_236__14 ;
    input inputs_236__13 ;
    input inputs_236__12 ;
    input inputs_236__11 ;
    input inputs_236__10 ;
    input inputs_236__9 ;
    input inputs_236__8 ;
    input inputs_236__7 ;
    input inputs_236__6 ;
    input inputs_236__5 ;
    input inputs_236__4 ;
    input inputs_236__3 ;
    input inputs_236__2 ;
    input inputs_236__1 ;
    input inputs_236__0 ;
    input inputs_237__15 ;
    input inputs_237__14 ;
    input inputs_237__13 ;
    input inputs_237__12 ;
    input inputs_237__11 ;
    input inputs_237__10 ;
    input inputs_237__9 ;
    input inputs_237__8 ;
    input inputs_237__7 ;
    input inputs_237__6 ;
    input inputs_237__5 ;
    input inputs_237__4 ;
    input inputs_237__3 ;
    input inputs_237__2 ;
    input inputs_237__1 ;
    input inputs_237__0 ;
    input inputs_238__15 ;
    input inputs_238__14 ;
    input inputs_238__13 ;
    input inputs_238__12 ;
    input inputs_238__11 ;
    input inputs_238__10 ;
    input inputs_238__9 ;
    input inputs_238__8 ;
    input inputs_238__7 ;
    input inputs_238__6 ;
    input inputs_238__5 ;
    input inputs_238__4 ;
    input inputs_238__3 ;
    input inputs_238__2 ;
    input inputs_238__1 ;
    input inputs_238__0 ;
    input inputs_239__15 ;
    input inputs_239__14 ;
    input inputs_239__13 ;
    input inputs_239__12 ;
    input inputs_239__11 ;
    input inputs_239__10 ;
    input inputs_239__9 ;
    input inputs_239__8 ;
    input inputs_239__7 ;
    input inputs_239__6 ;
    input inputs_239__5 ;
    input inputs_239__4 ;
    input inputs_239__3 ;
    input inputs_239__2 ;
    input inputs_239__1 ;
    input inputs_239__0 ;
    input inputs_240__15 ;
    input inputs_240__14 ;
    input inputs_240__13 ;
    input inputs_240__12 ;
    input inputs_240__11 ;
    input inputs_240__10 ;
    input inputs_240__9 ;
    input inputs_240__8 ;
    input inputs_240__7 ;
    input inputs_240__6 ;
    input inputs_240__5 ;
    input inputs_240__4 ;
    input inputs_240__3 ;
    input inputs_240__2 ;
    input inputs_240__1 ;
    input inputs_240__0 ;
    input inputs_241__15 ;
    input inputs_241__14 ;
    input inputs_241__13 ;
    input inputs_241__12 ;
    input inputs_241__11 ;
    input inputs_241__10 ;
    input inputs_241__9 ;
    input inputs_241__8 ;
    input inputs_241__7 ;
    input inputs_241__6 ;
    input inputs_241__5 ;
    input inputs_241__4 ;
    input inputs_241__3 ;
    input inputs_241__2 ;
    input inputs_241__1 ;
    input inputs_241__0 ;
    input inputs_242__15 ;
    input inputs_242__14 ;
    input inputs_242__13 ;
    input inputs_242__12 ;
    input inputs_242__11 ;
    input inputs_242__10 ;
    input inputs_242__9 ;
    input inputs_242__8 ;
    input inputs_242__7 ;
    input inputs_242__6 ;
    input inputs_242__5 ;
    input inputs_242__4 ;
    input inputs_242__3 ;
    input inputs_242__2 ;
    input inputs_242__1 ;
    input inputs_242__0 ;
    input inputs_243__15 ;
    input inputs_243__14 ;
    input inputs_243__13 ;
    input inputs_243__12 ;
    input inputs_243__11 ;
    input inputs_243__10 ;
    input inputs_243__9 ;
    input inputs_243__8 ;
    input inputs_243__7 ;
    input inputs_243__6 ;
    input inputs_243__5 ;
    input inputs_243__4 ;
    input inputs_243__3 ;
    input inputs_243__2 ;
    input inputs_243__1 ;
    input inputs_243__0 ;
    input inputs_244__15 ;
    input inputs_244__14 ;
    input inputs_244__13 ;
    input inputs_244__12 ;
    input inputs_244__11 ;
    input inputs_244__10 ;
    input inputs_244__9 ;
    input inputs_244__8 ;
    input inputs_244__7 ;
    input inputs_244__6 ;
    input inputs_244__5 ;
    input inputs_244__4 ;
    input inputs_244__3 ;
    input inputs_244__2 ;
    input inputs_244__1 ;
    input inputs_244__0 ;
    input inputs_245__15 ;
    input inputs_245__14 ;
    input inputs_245__13 ;
    input inputs_245__12 ;
    input inputs_245__11 ;
    input inputs_245__10 ;
    input inputs_245__9 ;
    input inputs_245__8 ;
    input inputs_245__7 ;
    input inputs_245__6 ;
    input inputs_245__5 ;
    input inputs_245__4 ;
    input inputs_245__3 ;
    input inputs_245__2 ;
    input inputs_245__1 ;
    input inputs_245__0 ;
    input inputs_246__15 ;
    input inputs_246__14 ;
    input inputs_246__13 ;
    input inputs_246__12 ;
    input inputs_246__11 ;
    input inputs_246__10 ;
    input inputs_246__9 ;
    input inputs_246__8 ;
    input inputs_246__7 ;
    input inputs_246__6 ;
    input inputs_246__5 ;
    input inputs_246__4 ;
    input inputs_246__3 ;
    input inputs_246__2 ;
    input inputs_246__1 ;
    input inputs_246__0 ;
    input inputs_247__15 ;
    input inputs_247__14 ;
    input inputs_247__13 ;
    input inputs_247__12 ;
    input inputs_247__11 ;
    input inputs_247__10 ;
    input inputs_247__9 ;
    input inputs_247__8 ;
    input inputs_247__7 ;
    input inputs_247__6 ;
    input inputs_247__5 ;
    input inputs_247__4 ;
    input inputs_247__3 ;
    input inputs_247__2 ;
    input inputs_247__1 ;
    input inputs_247__0 ;
    input inputs_248__15 ;
    input inputs_248__14 ;
    input inputs_248__13 ;
    input inputs_248__12 ;
    input inputs_248__11 ;
    input inputs_248__10 ;
    input inputs_248__9 ;
    input inputs_248__8 ;
    input inputs_248__7 ;
    input inputs_248__6 ;
    input inputs_248__5 ;
    input inputs_248__4 ;
    input inputs_248__3 ;
    input inputs_248__2 ;
    input inputs_248__1 ;
    input inputs_248__0 ;
    input inputs_249__15 ;
    input inputs_249__14 ;
    input inputs_249__13 ;
    input inputs_249__12 ;
    input inputs_249__11 ;
    input inputs_249__10 ;
    input inputs_249__9 ;
    input inputs_249__8 ;
    input inputs_249__7 ;
    input inputs_249__6 ;
    input inputs_249__5 ;
    input inputs_249__4 ;
    input inputs_249__3 ;
    input inputs_249__2 ;
    input inputs_249__1 ;
    input inputs_249__0 ;
    input inputs_250__15 ;
    input inputs_250__14 ;
    input inputs_250__13 ;
    input inputs_250__12 ;
    input inputs_250__11 ;
    input inputs_250__10 ;
    input inputs_250__9 ;
    input inputs_250__8 ;
    input inputs_250__7 ;
    input inputs_250__6 ;
    input inputs_250__5 ;
    input inputs_250__4 ;
    input inputs_250__3 ;
    input inputs_250__2 ;
    input inputs_250__1 ;
    input inputs_250__0 ;
    input inputs_251__15 ;
    input inputs_251__14 ;
    input inputs_251__13 ;
    input inputs_251__12 ;
    input inputs_251__11 ;
    input inputs_251__10 ;
    input inputs_251__9 ;
    input inputs_251__8 ;
    input inputs_251__7 ;
    input inputs_251__6 ;
    input inputs_251__5 ;
    input inputs_251__4 ;
    input inputs_251__3 ;
    input inputs_251__2 ;
    input inputs_251__1 ;
    input inputs_251__0 ;
    input inputs_252__15 ;
    input inputs_252__14 ;
    input inputs_252__13 ;
    input inputs_252__12 ;
    input inputs_252__11 ;
    input inputs_252__10 ;
    input inputs_252__9 ;
    input inputs_252__8 ;
    input inputs_252__7 ;
    input inputs_252__6 ;
    input inputs_252__5 ;
    input inputs_252__4 ;
    input inputs_252__3 ;
    input inputs_252__2 ;
    input inputs_252__1 ;
    input inputs_252__0 ;
    input inputs_253__15 ;
    input inputs_253__14 ;
    input inputs_253__13 ;
    input inputs_253__12 ;
    input inputs_253__11 ;
    input inputs_253__10 ;
    input inputs_253__9 ;
    input inputs_253__8 ;
    input inputs_253__7 ;
    input inputs_253__6 ;
    input inputs_253__5 ;
    input inputs_253__4 ;
    input inputs_253__3 ;
    input inputs_253__2 ;
    input inputs_253__1 ;
    input inputs_253__0 ;
    input inputs_254__15 ;
    input inputs_254__14 ;
    input inputs_254__13 ;
    input inputs_254__12 ;
    input inputs_254__11 ;
    input inputs_254__10 ;
    input inputs_254__9 ;
    input inputs_254__8 ;
    input inputs_254__7 ;
    input inputs_254__6 ;
    input inputs_254__5 ;
    input inputs_254__4 ;
    input inputs_254__3 ;
    input inputs_254__2 ;
    input inputs_254__1 ;
    input inputs_254__0 ;
    input inputs_255__15 ;
    input inputs_255__14 ;
    input inputs_255__13 ;
    input inputs_255__12 ;
    input inputs_255__11 ;
    input inputs_255__10 ;
    input inputs_255__9 ;
    input inputs_255__8 ;
    input inputs_255__7 ;
    input inputs_255__6 ;
    input inputs_255__5 ;
    input inputs_255__4 ;
    input inputs_255__3 ;
    input inputs_255__2 ;
    input inputs_255__1 ;
    input inputs_255__0 ;
    input inputs_256__15 ;
    input inputs_256__14 ;
    input inputs_256__13 ;
    input inputs_256__12 ;
    input inputs_256__11 ;
    input inputs_256__10 ;
    input inputs_256__9 ;
    input inputs_256__8 ;
    input inputs_256__7 ;
    input inputs_256__6 ;
    input inputs_256__5 ;
    input inputs_256__4 ;
    input inputs_256__3 ;
    input inputs_256__2 ;
    input inputs_256__1 ;
    input inputs_256__0 ;
    input inputs_257__15 ;
    input inputs_257__14 ;
    input inputs_257__13 ;
    input inputs_257__12 ;
    input inputs_257__11 ;
    input inputs_257__10 ;
    input inputs_257__9 ;
    input inputs_257__8 ;
    input inputs_257__7 ;
    input inputs_257__6 ;
    input inputs_257__5 ;
    input inputs_257__4 ;
    input inputs_257__3 ;
    input inputs_257__2 ;
    input inputs_257__1 ;
    input inputs_257__0 ;
    input inputs_258__15 ;
    input inputs_258__14 ;
    input inputs_258__13 ;
    input inputs_258__12 ;
    input inputs_258__11 ;
    input inputs_258__10 ;
    input inputs_258__9 ;
    input inputs_258__8 ;
    input inputs_258__7 ;
    input inputs_258__6 ;
    input inputs_258__5 ;
    input inputs_258__4 ;
    input inputs_258__3 ;
    input inputs_258__2 ;
    input inputs_258__1 ;
    input inputs_258__0 ;
    input inputs_259__15 ;
    input inputs_259__14 ;
    input inputs_259__13 ;
    input inputs_259__12 ;
    input inputs_259__11 ;
    input inputs_259__10 ;
    input inputs_259__9 ;
    input inputs_259__8 ;
    input inputs_259__7 ;
    input inputs_259__6 ;
    input inputs_259__5 ;
    input inputs_259__4 ;
    input inputs_259__3 ;
    input inputs_259__2 ;
    input inputs_259__1 ;
    input inputs_259__0 ;
    input inputs_260__15 ;
    input inputs_260__14 ;
    input inputs_260__13 ;
    input inputs_260__12 ;
    input inputs_260__11 ;
    input inputs_260__10 ;
    input inputs_260__9 ;
    input inputs_260__8 ;
    input inputs_260__7 ;
    input inputs_260__6 ;
    input inputs_260__5 ;
    input inputs_260__4 ;
    input inputs_260__3 ;
    input inputs_260__2 ;
    input inputs_260__1 ;
    input inputs_260__0 ;
    input inputs_261__15 ;
    input inputs_261__14 ;
    input inputs_261__13 ;
    input inputs_261__12 ;
    input inputs_261__11 ;
    input inputs_261__10 ;
    input inputs_261__9 ;
    input inputs_261__8 ;
    input inputs_261__7 ;
    input inputs_261__6 ;
    input inputs_261__5 ;
    input inputs_261__4 ;
    input inputs_261__3 ;
    input inputs_261__2 ;
    input inputs_261__1 ;
    input inputs_261__0 ;
    input inputs_262__15 ;
    input inputs_262__14 ;
    input inputs_262__13 ;
    input inputs_262__12 ;
    input inputs_262__11 ;
    input inputs_262__10 ;
    input inputs_262__9 ;
    input inputs_262__8 ;
    input inputs_262__7 ;
    input inputs_262__6 ;
    input inputs_262__5 ;
    input inputs_262__4 ;
    input inputs_262__3 ;
    input inputs_262__2 ;
    input inputs_262__1 ;
    input inputs_262__0 ;
    input inputs_263__15 ;
    input inputs_263__14 ;
    input inputs_263__13 ;
    input inputs_263__12 ;
    input inputs_263__11 ;
    input inputs_263__10 ;
    input inputs_263__9 ;
    input inputs_263__8 ;
    input inputs_263__7 ;
    input inputs_263__6 ;
    input inputs_263__5 ;
    input inputs_263__4 ;
    input inputs_263__3 ;
    input inputs_263__2 ;
    input inputs_263__1 ;
    input inputs_263__0 ;
    input inputs_264__15 ;
    input inputs_264__14 ;
    input inputs_264__13 ;
    input inputs_264__12 ;
    input inputs_264__11 ;
    input inputs_264__10 ;
    input inputs_264__9 ;
    input inputs_264__8 ;
    input inputs_264__7 ;
    input inputs_264__6 ;
    input inputs_264__5 ;
    input inputs_264__4 ;
    input inputs_264__3 ;
    input inputs_264__2 ;
    input inputs_264__1 ;
    input inputs_264__0 ;
    input inputs_265__15 ;
    input inputs_265__14 ;
    input inputs_265__13 ;
    input inputs_265__12 ;
    input inputs_265__11 ;
    input inputs_265__10 ;
    input inputs_265__9 ;
    input inputs_265__8 ;
    input inputs_265__7 ;
    input inputs_265__6 ;
    input inputs_265__5 ;
    input inputs_265__4 ;
    input inputs_265__3 ;
    input inputs_265__2 ;
    input inputs_265__1 ;
    input inputs_265__0 ;
    input inputs_266__15 ;
    input inputs_266__14 ;
    input inputs_266__13 ;
    input inputs_266__12 ;
    input inputs_266__11 ;
    input inputs_266__10 ;
    input inputs_266__9 ;
    input inputs_266__8 ;
    input inputs_266__7 ;
    input inputs_266__6 ;
    input inputs_266__5 ;
    input inputs_266__4 ;
    input inputs_266__3 ;
    input inputs_266__2 ;
    input inputs_266__1 ;
    input inputs_266__0 ;
    input inputs_267__15 ;
    input inputs_267__14 ;
    input inputs_267__13 ;
    input inputs_267__12 ;
    input inputs_267__11 ;
    input inputs_267__10 ;
    input inputs_267__9 ;
    input inputs_267__8 ;
    input inputs_267__7 ;
    input inputs_267__6 ;
    input inputs_267__5 ;
    input inputs_267__4 ;
    input inputs_267__3 ;
    input inputs_267__2 ;
    input inputs_267__1 ;
    input inputs_267__0 ;
    input inputs_268__15 ;
    input inputs_268__14 ;
    input inputs_268__13 ;
    input inputs_268__12 ;
    input inputs_268__11 ;
    input inputs_268__10 ;
    input inputs_268__9 ;
    input inputs_268__8 ;
    input inputs_268__7 ;
    input inputs_268__6 ;
    input inputs_268__5 ;
    input inputs_268__4 ;
    input inputs_268__3 ;
    input inputs_268__2 ;
    input inputs_268__1 ;
    input inputs_268__0 ;
    input inputs_269__15 ;
    input inputs_269__14 ;
    input inputs_269__13 ;
    input inputs_269__12 ;
    input inputs_269__11 ;
    input inputs_269__10 ;
    input inputs_269__9 ;
    input inputs_269__8 ;
    input inputs_269__7 ;
    input inputs_269__6 ;
    input inputs_269__5 ;
    input inputs_269__4 ;
    input inputs_269__3 ;
    input inputs_269__2 ;
    input inputs_269__1 ;
    input inputs_269__0 ;
    input inputs_270__15 ;
    input inputs_270__14 ;
    input inputs_270__13 ;
    input inputs_270__12 ;
    input inputs_270__11 ;
    input inputs_270__10 ;
    input inputs_270__9 ;
    input inputs_270__8 ;
    input inputs_270__7 ;
    input inputs_270__6 ;
    input inputs_270__5 ;
    input inputs_270__4 ;
    input inputs_270__3 ;
    input inputs_270__2 ;
    input inputs_270__1 ;
    input inputs_270__0 ;
    input inputs_271__15 ;
    input inputs_271__14 ;
    input inputs_271__13 ;
    input inputs_271__12 ;
    input inputs_271__11 ;
    input inputs_271__10 ;
    input inputs_271__9 ;
    input inputs_271__8 ;
    input inputs_271__7 ;
    input inputs_271__6 ;
    input inputs_271__5 ;
    input inputs_271__4 ;
    input inputs_271__3 ;
    input inputs_271__2 ;
    input inputs_271__1 ;
    input inputs_271__0 ;
    input inputs_272__15 ;
    input inputs_272__14 ;
    input inputs_272__13 ;
    input inputs_272__12 ;
    input inputs_272__11 ;
    input inputs_272__10 ;
    input inputs_272__9 ;
    input inputs_272__8 ;
    input inputs_272__7 ;
    input inputs_272__6 ;
    input inputs_272__5 ;
    input inputs_272__4 ;
    input inputs_272__3 ;
    input inputs_272__2 ;
    input inputs_272__1 ;
    input inputs_272__0 ;
    input inputs_273__15 ;
    input inputs_273__14 ;
    input inputs_273__13 ;
    input inputs_273__12 ;
    input inputs_273__11 ;
    input inputs_273__10 ;
    input inputs_273__9 ;
    input inputs_273__8 ;
    input inputs_273__7 ;
    input inputs_273__6 ;
    input inputs_273__5 ;
    input inputs_273__4 ;
    input inputs_273__3 ;
    input inputs_273__2 ;
    input inputs_273__1 ;
    input inputs_273__0 ;
    input inputs_274__15 ;
    input inputs_274__14 ;
    input inputs_274__13 ;
    input inputs_274__12 ;
    input inputs_274__11 ;
    input inputs_274__10 ;
    input inputs_274__9 ;
    input inputs_274__8 ;
    input inputs_274__7 ;
    input inputs_274__6 ;
    input inputs_274__5 ;
    input inputs_274__4 ;
    input inputs_274__3 ;
    input inputs_274__2 ;
    input inputs_274__1 ;
    input inputs_274__0 ;
    input inputs_275__15 ;
    input inputs_275__14 ;
    input inputs_275__13 ;
    input inputs_275__12 ;
    input inputs_275__11 ;
    input inputs_275__10 ;
    input inputs_275__9 ;
    input inputs_275__8 ;
    input inputs_275__7 ;
    input inputs_275__6 ;
    input inputs_275__5 ;
    input inputs_275__4 ;
    input inputs_275__3 ;
    input inputs_275__2 ;
    input inputs_275__1 ;
    input inputs_275__0 ;
    input inputs_276__15 ;
    input inputs_276__14 ;
    input inputs_276__13 ;
    input inputs_276__12 ;
    input inputs_276__11 ;
    input inputs_276__10 ;
    input inputs_276__9 ;
    input inputs_276__8 ;
    input inputs_276__7 ;
    input inputs_276__6 ;
    input inputs_276__5 ;
    input inputs_276__4 ;
    input inputs_276__3 ;
    input inputs_276__2 ;
    input inputs_276__1 ;
    input inputs_276__0 ;
    input inputs_277__15 ;
    input inputs_277__14 ;
    input inputs_277__13 ;
    input inputs_277__12 ;
    input inputs_277__11 ;
    input inputs_277__10 ;
    input inputs_277__9 ;
    input inputs_277__8 ;
    input inputs_277__7 ;
    input inputs_277__6 ;
    input inputs_277__5 ;
    input inputs_277__4 ;
    input inputs_277__3 ;
    input inputs_277__2 ;
    input inputs_277__1 ;
    input inputs_277__0 ;
    input inputs_278__15 ;
    input inputs_278__14 ;
    input inputs_278__13 ;
    input inputs_278__12 ;
    input inputs_278__11 ;
    input inputs_278__10 ;
    input inputs_278__9 ;
    input inputs_278__8 ;
    input inputs_278__7 ;
    input inputs_278__6 ;
    input inputs_278__5 ;
    input inputs_278__4 ;
    input inputs_278__3 ;
    input inputs_278__2 ;
    input inputs_278__1 ;
    input inputs_278__0 ;
    input inputs_279__15 ;
    input inputs_279__14 ;
    input inputs_279__13 ;
    input inputs_279__12 ;
    input inputs_279__11 ;
    input inputs_279__10 ;
    input inputs_279__9 ;
    input inputs_279__8 ;
    input inputs_279__7 ;
    input inputs_279__6 ;
    input inputs_279__5 ;
    input inputs_279__4 ;
    input inputs_279__3 ;
    input inputs_279__2 ;
    input inputs_279__1 ;
    input inputs_279__0 ;
    input inputs_280__15 ;
    input inputs_280__14 ;
    input inputs_280__13 ;
    input inputs_280__12 ;
    input inputs_280__11 ;
    input inputs_280__10 ;
    input inputs_280__9 ;
    input inputs_280__8 ;
    input inputs_280__7 ;
    input inputs_280__6 ;
    input inputs_280__5 ;
    input inputs_280__4 ;
    input inputs_280__3 ;
    input inputs_280__2 ;
    input inputs_280__1 ;
    input inputs_280__0 ;
    input inputs_281__15 ;
    input inputs_281__14 ;
    input inputs_281__13 ;
    input inputs_281__12 ;
    input inputs_281__11 ;
    input inputs_281__10 ;
    input inputs_281__9 ;
    input inputs_281__8 ;
    input inputs_281__7 ;
    input inputs_281__6 ;
    input inputs_281__5 ;
    input inputs_281__4 ;
    input inputs_281__3 ;
    input inputs_281__2 ;
    input inputs_281__1 ;
    input inputs_281__0 ;
    input inputs_282__15 ;
    input inputs_282__14 ;
    input inputs_282__13 ;
    input inputs_282__12 ;
    input inputs_282__11 ;
    input inputs_282__10 ;
    input inputs_282__9 ;
    input inputs_282__8 ;
    input inputs_282__7 ;
    input inputs_282__6 ;
    input inputs_282__5 ;
    input inputs_282__4 ;
    input inputs_282__3 ;
    input inputs_282__2 ;
    input inputs_282__1 ;
    input inputs_282__0 ;
    input inputs_283__15 ;
    input inputs_283__14 ;
    input inputs_283__13 ;
    input inputs_283__12 ;
    input inputs_283__11 ;
    input inputs_283__10 ;
    input inputs_283__9 ;
    input inputs_283__8 ;
    input inputs_283__7 ;
    input inputs_283__6 ;
    input inputs_283__5 ;
    input inputs_283__4 ;
    input inputs_283__3 ;
    input inputs_283__2 ;
    input inputs_283__1 ;
    input inputs_283__0 ;
    input inputs_284__15 ;
    input inputs_284__14 ;
    input inputs_284__13 ;
    input inputs_284__12 ;
    input inputs_284__11 ;
    input inputs_284__10 ;
    input inputs_284__9 ;
    input inputs_284__8 ;
    input inputs_284__7 ;
    input inputs_284__6 ;
    input inputs_284__5 ;
    input inputs_284__4 ;
    input inputs_284__3 ;
    input inputs_284__2 ;
    input inputs_284__1 ;
    input inputs_284__0 ;
    input inputs_285__15 ;
    input inputs_285__14 ;
    input inputs_285__13 ;
    input inputs_285__12 ;
    input inputs_285__11 ;
    input inputs_285__10 ;
    input inputs_285__9 ;
    input inputs_285__8 ;
    input inputs_285__7 ;
    input inputs_285__6 ;
    input inputs_285__5 ;
    input inputs_285__4 ;
    input inputs_285__3 ;
    input inputs_285__2 ;
    input inputs_285__1 ;
    input inputs_285__0 ;
    input inputs_286__15 ;
    input inputs_286__14 ;
    input inputs_286__13 ;
    input inputs_286__12 ;
    input inputs_286__11 ;
    input inputs_286__10 ;
    input inputs_286__9 ;
    input inputs_286__8 ;
    input inputs_286__7 ;
    input inputs_286__6 ;
    input inputs_286__5 ;
    input inputs_286__4 ;
    input inputs_286__3 ;
    input inputs_286__2 ;
    input inputs_286__1 ;
    input inputs_286__0 ;
    input inputs_287__15 ;
    input inputs_287__14 ;
    input inputs_287__13 ;
    input inputs_287__12 ;
    input inputs_287__11 ;
    input inputs_287__10 ;
    input inputs_287__9 ;
    input inputs_287__8 ;
    input inputs_287__7 ;
    input inputs_287__6 ;
    input inputs_287__5 ;
    input inputs_287__4 ;
    input inputs_287__3 ;
    input inputs_287__2 ;
    input inputs_287__1 ;
    input inputs_287__0 ;
    input inputs_288__15 ;
    input inputs_288__14 ;
    input inputs_288__13 ;
    input inputs_288__12 ;
    input inputs_288__11 ;
    input inputs_288__10 ;
    input inputs_288__9 ;
    input inputs_288__8 ;
    input inputs_288__7 ;
    input inputs_288__6 ;
    input inputs_288__5 ;
    input inputs_288__4 ;
    input inputs_288__3 ;
    input inputs_288__2 ;
    input inputs_288__1 ;
    input inputs_288__0 ;
    input inputs_289__15 ;
    input inputs_289__14 ;
    input inputs_289__13 ;
    input inputs_289__12 ;
    input inputs_289__11 ;
    input inputs_289__10 ;
    input inputs_289__9 ;
    input inputs_289__8 ;
    input inputs_289__7 ;
    input inputs_289__6 ;
    input inputs_289__5 ;
    input inputs_289__4 ;
    input inputs_289__3 ;
    input inputs_289__2 ;
    input inputs_289__1 ;
    input inputs_289__0 ;
    input inputs_290__15 ;
    input inputs_290__14 ;
    input inputs_290__13 ;
    input inputs_290__12 ;
    input inputs_290__11 ;
    input inputs_290__10 ;
    input inputs_290__9 ;
    input inputs_290__8 ;
    input inputs_290__7 ;
    input inputs_290__6 ;
    input inputs_290__5 ;
    input inputs_290__4 ;
    input inputs_290__3 ;
    input inputs_290__2 ;
    input inputs_290__1 ;
    input inputs_290__0 ;
    input inputs_291__15 ;
    input inputs_291__14 ;
    input inputs_291__13 ;
    input inputs_291__12 ;
    input inputs_291__11 ;
    input inputs_291__10 ;
    input inputs_291__9 ;
    input inputs_291__8 ;
    input inputs_291__7 ;
    input inputs_291__6 ;
    input inputs_291__5 ;
    input inputs_291__4 ;
    input inputs_291__3 ;
    input inputs_291__2 ;
    input inputs_291__1 ;
    input inputs_291__0 ;
    input inputs_292__15 ;
    input inputs_292__14 ;
    input inputs_292__13 ;
    input inputs_292__12 ;
    input inputs_292__11 ;
    input inputs_292__10 ;
    input inputs_292__9 ;
    input inputs_292__8 ;
    input inputs_292__7 ;
    input inputs_292__6 ;
    input inputs_292__5 ;
    input inputs_292__4 ;
    input inputs_292__3 ;
    input inputs_292__2 ;
    input inputs_292__1 ;
    input inputs_292__0 ;
    input inputs_293__15 ;
    input inputs_293__14 ;
    input inputs_293__13 ;
    input inputs_293__12 ;
    input inputs_293__11 ;
    input inputs_293__10 ;
    input inputs_293__9 ;
    input inputs_293__8 ;
    input inputs_293__7 ;
    input inputs_293__6 ;
    input inputs_293__5 ;
    input inputs_293__4 ;
    input inputs_293__3 ;
    input inputs_293__2 ;
    input inputs_293__1 ;
    input inputs_293__0 ;
    input inputs_294__15 ;
    input inputs_294__14 ;
    input inputs_294__13 ;
    input inputs_294__12 ;
    input inputs_294__11 ;
    input inputs_294__10 ;
    input inputs_294__9 ;
    input inputs_294__8 ;
    input inputs_294__7 ;
    input inputs_294__6 ;
    input inputs_294__5 ;
    input inputs_294__4 ;
    input inputs_294__3 ;
    input inputs_294__2 ;
    input inputs_294__1 ;
    input inputs_294__0 ;
    input inputs_295__15 ;
    input inputs_295__14 ;
    input inputs_295__13 ;
    input inputs_295__12 ;
    input inputs_295__11 ;
    input inputs_295__10 ;
    input inputs_295__9 ;
    input inputs_295__8 ;
    input inputs_295__7 ;
    input inputs_295__6 ;
    input inputs_295__5 ;
    input inputs_295__4 ;
    input inputs_295__3 ;
    input inputs_295__2 ;
    input inputs_295__1 ;
    input inputs_295__0 ;
    input inputs_296__15 ;
    input inputs_296__14 ;
    input inputs_296__13 ;
    input inputs_296__12 ;
    input inputs_296__11 ;
    input inputs_296__10 ;
    input inputs_296__9 ;
    input inputs_296__8 ;
    input inputs_296__7 ;
    input inputs_296__6 ;
    input inputs_296__5 ;
    input inputs_296__4 ;
    input inputs_296__3 ;
    input inputs_296__2 ;
    input inputs_296__1 ;
    input inputs_296__0 ;
    input inputs_297__15 ;
    input inputs_297__14 ;
    input inputs_297__13 ;
    input inputs_297__12 ;
    input inputs_297__11 ;
    input inputs_297__10 ;
    input inputs_297__9 ;
    input inputs_297__8 ;
    input inputs_297__7 ;
    input inputs_297__6 ;
    input inputs_297__5 ;
    input inputs_297__4 ;
    input inputs_297__3 ;
    input inputs_297__2 ;
    input inputs_297__1 ;
    input inputs_297__0 ;
    input inputs_298__15 ;
    input inputs_298__14 ;
    input inputs_298__13 ;
    input inputs_298__12 ;
    input inputs_298__11 ;
    input inputs_298__10 ;
    input inputs_298__9 ;
    input inputs_298__8 ;
    input inputs_298__7 ;
    input inputs_298__6 ;
    input inputs_298__5 ;
    input inputs_298__4 ;
    input inputs_298__3 ;
    input inputs_298__2 ;
    input inputs_298__1 ;
    input inputs_298__0 ;
    input inputs_299__15 ;
    input inputs_299__14 ;
    input inputs_299__13 ;
    input inputs_299__12 ;
    input inputs_299__11 ;
    input inputs_299__10 ;
    input inputs_299__9 ;
    input inputs_299__8 ;
    input inputs_299__7 ;
    input inputs_299__6 ;
    input inputs_299__5 ;
    input inputs_299__4 ;
    input inputs_299__3 ;
    input inputs_299__2 ;
    input inputs_299__1 ;
    input inputs_299__0 ;
    input inputs_300__15 ;
    input inputs_300__14 ;
    input inputs_300__13 ;
    input inputs_300__12 ;
    input inputs_300__11 ;
    input inputs_300__10 ;
    input inputs_300__9 ;
    input inputs_300__8 ;
    input inputs_300__7 ;
    input inputs_300__6 ;
    input inputs_300__5 ;
    input inputs_300__4 ;
    input inputs_300__3 ;
    input inputs_300__2 ;
    input inputs_300__1 ;
    input inputs_300__0 ;
    input inputs_301__15 ;
    input inputs_301__14 ;
    input inputs_301__13 ;
    input inputs_301__12 ;
    input inputs_301__11 ;
    input inputs_301__10 ;
    input inputs_301__9 ;
    input inputs_301__8 ;
    input inputs_301__7 ;
    input inputs_301__6 ;
    input inputs_301__5 ;
    input inputs_301__4 ;
    input inputs_301__3 ;
    input inputs_301__2 ;
    input inputs_301__1 ;
    input inputs_301__0 ;
    input inputs_302__15 ;
    input inputs_302__14 ;
    input inputs_302__13 ;
    input inputs_302__12 ;
    input inputs_302__11 ;
    input inputs_302__10 ;
    input inputs_302__9 ;
    input inputs_302__8 ;
    input inputs_302__7 ;
    input inputs_302__6 ;
    input inputs_302__5 ;
    input inputs_302__4 ;
    input inputs_302__3 ;
    input inputs_302__2 ;
    input inputs_302__1 ;
    input inputs_302__0 ;
    input inputs_303__15 ;
    input inputs_303__14 ;
    input inputs_303__13 ;
    input inputs_303__12 ;
    input inputs_303__11 ;
    input inputs_303__10 ;
    input inputs_303__9 ;
    input inputs_303__8 ;
    input inputs_303__7 ;
    input inputs_303__6 ;
    input inputs_303__5 ;
    input inputs_303__4 ;
    input inputs_303__3 ;
    input inputs_303__2 ;
    input inputs_303__1 ;
    input inputs_303__0 ;
    input inputs_304__15 ;
    input inputs_304__14 ;
    input inputs_304__13 ;
    input inputs_304__12 ;
    input inputs_304__11 ;
    input inputs_304__10 ;
    input inputs_304__9 ;
    input inputs_304__8 ;
    input inputs_304__7 ;
    input inputs_304__6 ;
    input inputs_304__5 ;
    input inputs_304__4 ;
    input inputs_304__3 ;
    input inputs_304__2 ;
    input inputs_304__1 ;
    input inputs_304__0 ;
    input inputs_305__15 ;
    input inputs_305__14 ;
    input inputs_305__13 ;
    input inputs_305__12 ;
    input inputs_305__11 ;
    input inputs_305__10 ;
    input inputs_305__9 ;
    input inputs_305__8 ;
    input inputs_305__7 ;
    input inputs_305__6 ;
    input inputs_305__5 ;
    input inputs_305__4 ;
    input inputs_305__3 ;
    input inputs_305__2 ;
    input inputs_305__1 ;
    input inputs_305__0 ;
    input inputs_306__15 ;
    input inputs_306__14 ;
    input inputs_306__13 ;
    input inputs_306__12 ;
    input inputs_306__11 ;
    input inputs_306__10 ;
    input inputs_306__9 ;
    input inputs_306__8 ;
    input inputs_306__7 ;
    input inputs_306__6 ;
    input inputs_306__5 ;
    input inputs_306__4 ;
    input inputs_306__3 ;
    input inputs_306__2 ;
    input inputs_306__1 ;
    input inputs_306__0 ;
    input inputs_307__15 ;
    input inputs_307__14 ;
    input inputs_307__13 ;
    input inputs_307__12 ;
    input inputs_307__11 ;
    input inputs_307__10 ;
    input inputs_307__9 ;
    input inputs_307__8 ;
    input inputs_307__7 ;
    input inputs_307__6 ;
    input inputs_307__5 ;
    input inputs_307__4 ;
    input inputs_307__3 ;
    input inputs_307__2 ;
    input inputs_307__1 ;
    input inputs_307__0 ;
    input inputs_308__15 ;
    input inputs_308__14 ;
    input inputs_308__13 ;
    input inputs_308__12 ;
    input inputs_308__11 ;
    input inputs_308__10 ;
    input inputs_308__9 ;
    input inputs_308__8 ;
    input inputs_308__7 ;
    input inputs_308__6 ;
    input inputs_308__5 ;
    input inputs_308__4 ;
    input inputs_308__3 ;
    input inputs_308__2 ;
    input inputs_308__1 ;
    input inputs_308__0 ;
    input inputs_309__15 ;
    input inputs_309__14 ;
    input inputs_309__13 ;
    input inputs_309__12 ;
    input inputs_309__11 ;
    input inputs_309__10 ;
    input inputs_309__9 ;
    input inputs_309__8 ;
    input inputs_309__7 ;
    input inputs_309__6 ;
    input inputs_309__5 ;
    input inputs_309__4 ;
    input inputs_309__3 ;
    input inputs_309__2 ;
    input inputs_309__1 ;
    input inputs_309__0 ;
    input inputs_310__15 ;
    input inputs_310__14 ;
    input inputs_310__13 ;
    input inputs_310__12 ;
    input inputs_310__11 ;
    input inputs_310__10 ;
    input inputs_310__9 ;
    input inputs_310__8 ;
    input inputs_310__7 ;
    input inputs_310__6 ;
    input inputs_310__5 ;
    input inputs_310__4 ;
    input inputs_310__3 ;
    input inputs_310__2 ;
    input inputs_310__1 ;
    input inputs_310__0 ;
    input inputs_311__15 ;
    input inputs_311__14 ;
    input inputs_311__13 ;
    input inputs_311__12 ;
    input inputs_311__11 ;
    input inputs_311__10 ;
    input inputs_311__9 ;
    input inputs_311__8 ;
    input inputs_311__7 ;
    input inputs_311__6 ;
    input inputs_311__5 ;
    input inputs_311__4 ;
    input inputs_311__3 ;
    input inputs_311__2 ;
    input inputs_311__1 ;
    input inputs_311__0 ;
    input inputs_312__15 ;
    input inputs_312__14 ;
    input inputs_312__13 ;
    input inputs_312__12 ;
    input inputs_312__11 ;
    input inputs_312__10 ;
    input inputs_312__9 ;
    input inputs_312__8 ;
    input inputs_312__7 ;
    input inputs_312__6 ;
    input inputs_312__5 ;
    input inputs_312__4 ;
    input inputs_312__3 ;
    input inputs_312__2 ;
    input inputs_312__1 ;
    input inputs_312__0 ;
    input inputs_313__15 ;
    input inputs_313__14 ;
    input inputs_313__13 ;
    input inputs_313__12 ;
    input inputs_313__11 ;
    input inputs_313__10 ;
    input inputs_313__9 ;
    input inputs_313__8 ;
    input inputs_313__7 ;
    input inputs_313__6 ;
    input inputs_313__5 ;
    input inputs_313__4 ;
    input inputs_313__3 ;
    input inputs_313__2 ;
    input inputs_313__1 ;
    input inputs_313__0 ;
    input inputs_314__15 ;
    input inputs_314__14 ;
    input inputs_314__13 ;
    input inputs_314__12 ;
    input inputs_314__11 ;
    input inputs_314__10 ;
    input inputs_314__9 ;
    input inputs_314__8 ;
    input inputs_314__7 ;
    input inputs_314__6 ;
    input inputs_314__5 ;
    input inputs_314__4 ;
    input inputs_314__3 ;
    input inputs_314__2 ;
    input inputs_314__1 ;
    input inputs_314__0 ;
    input inputs_315__15 ;
    input inputs_315__14 ;
    input inputs_315__13 ;
    input inputs_315__12 ;
    input inputs_315__11 ;
    input inputs_315__10 ;
    input inputs_315__9 ;
    input inputs_315__8 ;
    input inputs_315__7 ;
    input inputs_315__6 ;
    input inputs_315__5 ;
    input inputs_315__4 ;
    input inputs_315__3 ;
    input inputs_315__2 ;
    input inputs_315__1 ;
    input inputs_315__0 ;
    input inputs_316__15 ;
    input inputs_316__14 ;
    input inputs_316__13 ;
    input inputs_316__12 ;
    input inputs_316__11 ;
    input inputs_316__10 ;
    input inputs_316__9 ;
    input inputs_316__8 ;
    input inputs_316__7 ;
    input inputs_316__6 ;
    input inputs_316__5 ;
    input inputs_316__4 ;
    input inputs_316__3 ;
    input inputs_316__2 ;
    input inputs_316__1 ;
    input inputs_316__0 ;
    input inputs_317__15 ;
    input inputs_317__14 ;
    input inputs_317__13 ;
    input inputs_317__12 ;
    input inputs_317__11 ;
    input inputs_317__10 ;
    input inputs_317__9 ;
    input inputs_317__8 ;
    input inputs_317__7 ;
    input inputs_317__6 ;
    input inputs_317__5 ;
    input inputs_317__4 ;
    input inputs_317__3 ;
    input inputs_317__2 ;
    input inputs_317__1 ;
    input inputs_317__0 ;
    input inputs_318__15 ;
    input inputs_318__14 ;
    input inputs_318__13 ;
    input inputs_318__12 ;
    input inputs_318__11 ;
    input inputs_318__10 ;
    input inputs_318__9 ;
    input inputs_318__8 ;
    input inputs_318__7 ;
    input inputs_318__6 ;
    input inputs_318__5 ;
    input inputs_318__4 ;
    input inputs_318__3 ;
    input inputs_318__2 ;
    input inputs_318__1 ;
    input inputs_318__0 ;
    input inputs_319__15 ;
    input inputs_319__14 ;
    input inputs_319__13 ;
    input inputs_319__12 ;
    input inputs_319__11 ;
    input inputs_319__10 ;
    input inputs_319__9 ;
    input inputs_319__8 ;
    input inputs_319__7 ;
    input inputs_319__6 ;
    input inputs_319__5 ;
    input inputs_319__4 ;
    input inputs_319__3 ;
    input inputs_319__2 ;
    input inputs_319__1 ;
    input inputs_319__0 ;
    input inputs_320__15 ;
    input inputs_320__14 ;
    input inputs_320__13 ;
    input inputs_320__12 ;
    input inputs_320__11 ;
    input inputs_320__10 ;
    input inputs_320__9 ;
    input inputs_320__8 ;
    input inputs_320__7 ;
    input inputs_320__6 ;
    input inputs_320__5 ;
    input inputs_320__4 ;
    input inputs_320__3 ;
    input inputs_320__2 ;
    input inputs_320__1 ;
    input inputs_320__0 ;
    input inputs_321__15 ;
    input inputs_321__14 ;
    input inputs_321__13 ;
    input inputs_321__12 ;
    input inputs_321__11 ;
    input inputs_321__10 ;
    input inputs_321__9 ;
    input inputs_321__8 ;
    input inputs_321__7 ;
    input inputs_321__6 ;
    input inputs_321__5 ;
    input inputs_321__4 ;
    input inputs_321__3 ;
    input inputs_321__2 ;
    input inputs_321__1 ;
    input inputs_321__0 ;
    input inputs_322__15 ;
    input inputs_322__14 ;
    input inputs_322__13 ;
    input inputs_322__12 ;
    input inputs_322__11 ;
    input inputs_322__10 ;
    input inputs_322__9 ;
    input inputs_322__8 ;
    input inputs_322__7 ;
    input inputs_322__6 ;
    input inputs_322__5 ;
    input inputs_322__4 ;
    input inputs_322__3 ;
    input inputs_322__2 ;
    input inputs_322__1 ;
    input inputs_322__0 ;
    input inputs_323__15 ;
    input inputs_323__14 ;
    input inputs_323__13 ;
    input inputs_323__12 ;
    input inputs_323__11 ;
    input inputs_323__10 ;
    input inputs_323__9 ;
    input inputs_323__8 ;
    input inputs_323__7 ;
    input inputs_323__6 ;
    input inputs_323__5 ;
    input inputs_323__4 ;
    input inputs_323__3 ;
    input inputs_323__2 ;
    input inputs_323__1 ;
    input inputs_323__0 ;
    input inputs_324__15 ;
    input inputs_324__14 ;
    input inputs_324__13 ;
    input inputs_324__12 ;
    input inputs_324__11 ;
    input inputs_324__10 ;
    input inputs_324__9 ;
    input inputs_324__8 ;
    input inputs_324__7 ;
    input inputs_324__6 ;
    input inputs_324__5 ;
    input inputs_324__4 ;
    input inputs_324__3 ;
    input inputs_324__2 ;
    input inputs_324__1 ;
    input inputs_324__0 ;
    input inputs_325__15 ;
    input inputs_325__14 ;
    input inputs_325__13 ;
    input inputs_325__12 ;
    input inputs_325__11 ;
    input inputs_325__10 ;
    input inputs_325__9 ;
    input inputs_325__8 ;
    input inputs_325__7 ;
    input inputs_325__6 ;
    input inputs_325__5 ;
    input inputs_325__4 ;
    input inputs_325__3 ;
    input inputs_325__2 ;
    input inputs_325__1 ;
    input inputs_325__0 ;
    input inputs_326__15 ;
    input inputs_326__14 ;
    input inputs_326__13 ;
    input inputs_326__12 ;
    input inputs_326__11 ;
    input inputs_326__10 ;
    input inputs_326__9 ;
    input inputs_326__8 ;
    input inputs_326__7 ;
    input inputs_326__6 ;
    input inputs_326__5 ;
    input inputs_326__4 ;
    input inputs_326__3 ;
    input inputs_326__2 ;
    input inputs_326__1 ;
    input inputs_326__0 ;
    input inputs_327__15 ;
    input inputs_327__14 ;
    input inputs_327__13 ;
    input inputs_327__12 ;
    input inputs_327__11 ;
    input inputs_327__10 ;
    input inputs_327__9 ;
    input inputs_327__8 ;
    input inputs_327__7 ;
    input inputs_327__6 ;
    input inputs_327__5 ;
    input inputs_327__4 ;
    input inputs_327__3 ;
    input inputs_327__2 ;
    input inputs_327__1 ;
    input inputs_327__0 ;
    input inputs_328__15 ;
    input inputs_328__14 ;
    input inputs_328__13 ;
    input inputs_328__12 ;
    input inputs_328__11 ;
    input inputs_328__10 ;
    input inputs_328__9 ;
    input inputs_328__8 ;
    input inputs_328__7 ;
    input inputs_328__6 ;
    input inputs_328__5 ;
    input inputs_328__4 ;
    input inputs_328__3 ;
    input inputs_328__2 ;
    input inputs_328__1 ;
    input inputs_328__0 ;
    input inputs_329__15 ;
    input inputs_329__14 ;
    input inputs_329__13 ;
    input inputs_329__12 ;
    input inputs_329__11 ;
    input inputs_329__10 ;
    input inputs_329__9 ;
    input inputs_329__8 ;
    input inputs_329__7 ;
    input inputs_329__6 ;
    input inputs_329__5 ;
    input inputs_329__4 ;
    input inputs_329__3 ;
    input inputs_329__2 ;
    input inputs_329__1 ;
    input inputs_329__0 ;
    input inputs_330__15 ;
    input inputs_330__14 ;
    input inputs_330__13 ;
    input inputs_330__12 ;
    input inputs_330__11 ;
    input inputs_330__10 ;
    input inputs_330__9 ;
    input inputs_330__8 ;
    input inputs_330__7 ;
    input inputs_330__6 ;
    input inputs_330__5 ;
    input inputs_330__4 ;
    input inputs_330__3 ;
    input inputs_330__2 ;
    input inputs_330__1 ;
    input inputs_330__0 ;
    input inputs_331__15 ;
    input inputs_331__14 ;
    input inputs_331__13 ;
    input inputs_331__12 ;
    input inputs_331__11 ;
    input inputs_331__10 ;
    input inputs_331__9 ;
    input inputs_331__8 ;
    input inputs_331__7 ;
    input inputs_331__6 ;
    input inputs_331__5 ;
    input inputs_331__4 ;
    input inputs_331__3 ;
    input inputs_331__2 ;
    input inputs_331__1 ;
    input inputs_331__0 ;
    input inputs_332__15 ;
    input inputs_332__14 ;
    input inputs_332__13 ;
    input inputs_332__12 ;
    input inputs_332__11 ;
    input inputs_332__10 ;
    input inputs_332__9 ;
    input inputs_332__8 ;
    input inputs_332__7 ;
    input inputs_332__6 ;
    input inputs_332__5 ;
    input inputs_332__4 ;
    input inputs_332__3 ;
    input inputs_332__2 ;
    input inputs_332__1 ;
    input inputs_332__0 ;
    input inputs_333__15 ;
    input inputs_333__14 ;
    input inputs_333__13 ;
    input inputs_333__12 ;
    input inputs_333__11 ;
    input inputs_333__10 ;
    input inputs_333__9 ;
    input inputs_333__8 ;
    input inputs_333__7 ;
    input inputs_333__6 ;
    input inputs_333__5 ;
    input inputs_333__4 ;
    input inputs_333__3 ;
    input inputs_333__2 ;
    input inputs_333__1 ;
    input inputs_333__0 ;
    input inputs_334__15 ;
    input inputs_334__14 ;
    input inputs_334__13 ;
    input inputs_334__12 ;
    input inputs_334__11 ;
    input inputs_334__10 ;
    input inputs_334__9 ;
    input inputs_334__8 ;
    input inputs_334__7 ;
    input inputs_334__6 ;
    input inputs_334__5 ;
    input inputs_334__4 ;
    input inputs_334__3 ;
    input inputs_334__2 ;
    input inputs_334__1 ;
    input inputs_334__0 ;
    input inputs_335__15 ;
    input inputs_335__14 ;
    input inputs_335__13 ;
    input inputs_335__12 ;
    input inputs_335__11 ;
    input inputs_335__10 ;
    input inputs_335__9 ;
    input inputs_335__8 ;
    input inputs_335__7 ;
    input inputs_335__6 ;
    input inputs_335__5 ;
    input inputs_335__4 ;
    input inputs_335__3 ;
    input inputs_335__2 ;
    input inputs_335__1 ;
    input inputs_335__0 ;
    input inputs_336__15 ;
    input inputs_336__14 ;
    input inputs_336__13 ;
    input inputs_336__12 ;
    input inputs_336__11 ;
    input inputs_336__10 ;
    input inputs_336__9 ;
    input inputs_336__8 ;
    input inputs_336__7 ;
    input inputs_336__6 ;
    input inputs_336__5 ;
    input inputs_336__4 ;
    input inputs_336__3 ;
    input inputs_336__2 ;
    input inputs_336__1 ;
    input inputs_336__0 ;
    input inputs_337__15 ;
    input inputs_337__14 ;
    input inputs_337__13 ;
    input inputs_337__12 ;
    input inputs_337__11 ;
    input inputs_337__10 ;
    input inputs_337__9 ;
    input inputs_337__8 ;
    input inputs_337__7 ;
    input inputs_337__6 ;
    input inputs_337__5 ;
    input inputs_337__4 ;
    input inputs_337__3 ;
    input inputs_337__2 ;
    input inputs_337__1 ;
    input inputs_337__0 ;
    input inputs_338__15 ;
    input inputs_338__14 ;
    input inputs_338__13 ;
    input inputs_338__12 ;
    input inputs_338__11 ;
    input inputs_338__10 ;
    input inputs_338__9 ;
    input inputs_338__8 ;
    input inputs_338__7 ;
    input inputs_338__6 ;
    input inputs_338__5 ;
    input inputs_338__4 ;
    input inputs_338__3 ;
    input inputs_338__2 ;
    input inputs_338__1 ;
    input inputs_338__0 ;
    input inputs_339__15 ;
    input inputs_339__14 ;
    input inputs_339__13 ;
    input inputs_339__12 ;
    input inputs_339__11 ;
    input inputs_339__10 ;
    input inputs_339__9 ;
    input inputs_339__8 ;
    input inputs_339__7 ;
    input inputs_339__6 ;
    input inputs_339__5 ;
    input inputs_339__4 ;
    input inputs_339__3 ;
    input inputs_339__2 ;
    input inputs_339__1 ;
    input inputs_339__0 ;
    input inputs_340__15 ;
    input inputs_340__14 ;
    input inputs_340__13 ;
    input inputs_340__12 ;
    input inputs_340__11 ;
    input inputs_340__10 ;
    input inputs_340__9 ;
    input inputs_340__8 ;
    input inputs_340__7 ;
    input inputs_340__6 ;
    input inputs_340__5 ;
    input inputs_340__4 ;
    input inputs_340__3 ;
    input inputs_340__2 ;
    input inputs_340__1 ;
    input inputs_340__0 ;
    input inputs_341__15 ;
    input inputs_341__14 ;
    input inputs_341__13 ;
    input inputs_341__12 ;
    input inputs_341__11 ;
    input inputs_341__10 ;
    input inputs_341__9 ;
    input inputs_341__8 ;
    input inputs_341__7 ;
    input inputs_341__6 ;
    input inputs_341__5 ;
    input inputs_341__4 ;
    input inputs_341__3 ;
    input inputs_341__2 ;
    input inputs_341__1 ;
    input inputs_341__0 ;
    input inputs_342__15 ;
    input inputs_342__14 ;
    input inputs_342__13 ;
    input inputs_342__12 ;
    input inputs_342__11 ;
    input inputs_342__10 ;
    input inputs_342__9 ;
    input inputs_342__8 ;
    input inputs_342__7 ;
    input inputs_342__6 ;
    input inputs_342__5 ;
    input inputs_342__4 ;
    input inputs_342__3 ;
    input inputs_342__2 ;
    input inputs_342__1 ;
    input inputs_342__0 ;
    input inputs_343__15 ;
    input inputs_343__14 ;
    input inputs_343__13 ;
    input inputs_343__12 ;
    input inputs_343__11 ;
    input inputs_343__10 ;
    input inputs_343__9 ;
    input inputs_343__8 ;
    input inputs_343__7 ;
    input inputs_343__6 ;
    input inputs_343__5 ;
    input inputs_343__4 ;
    input inputs_343__3 ;
    input inputs_343__2 ;
    input inputs_343__1 ;
    input inputs_343__0 ;
    input inputs_344__15 ;
    input inputs_344__14 ;
    input inputs_344__13 ;
    input inputs_344__12 ;
    input inputs_344__11 ;
    input inputs_344__10 ;
    input inputs_344__9 ;
    input inputs_344__8 ;
    input inputs_344__7 ;
    input inputs_344__6 ;
    input inputs_344__5 ;
    input inputs_344__4 ;
    input inputs_344__3 ;
    input inputs_344__2 ;
    input inputs_344__1 ;
    input inputs_344__0 ;
    input inputs_345__15 ;
    input inputs_345__14 ;
    input inputs_345__13 ;
    input inputs_345__12 ;
    input inputs_345__11 ;
    input inputs_345__10 ;
    input inputs_345__9 ;
    input inputs_345__8 ;
    input inputs_345__7 ;
    input inputs_345__6 ;
    input inputs_345__5 ;
    input inputs_345__4 ;
    input inputs_345__3 ;
    input inputs_345__2 ;
    input inputs_345__1 ;
    input inputs_345__0 ;
    input inputs_346__15 ;
    input inputs_346__14 ;
    input inputs_346__13 ;
    input inputs_346__12 ;
    input inputs_346__11 ;
    input inputs_346__10 ;
    input inputs_346__9 ;
    input inputs_346__8 ;
    input inputs_346__7 ;
    input inputs_346__6 ;
    input inputs_346__5 ;
    input inputs_346__4 ;
    input inputs_346__3 ;
    input inputs_346__2 ;
    input inputs_346__1 ;
    input inputs_346__0 ;
    input inputs_347__15 ;
    input inputs_347__14 ;
    input inputs_347__13 ;
    input inputs_347__12 ;
    input inputs_347__11 ;
    input inputs_347__10 ;
    input inputs_347__9 ;
    input inputs_347__8 ;
    input inputs_347__7 ;
    input inputs_347__6 ;
    input inputs_347__5 ;
    input inputs_347__4 ;
    input inputs_347__3 ;
    input inputs_347__2 ;
    input inputs_347__1 ;
    input inputs_347__0 ;
    input inputs_348__15 ;
    input inputs_348__14 ;
    input inputs_348__13 ;
    input inputs_348__12 ;
    input inputs_348__11 ;
    input inputs_348__10 ;
    input inputs_348__9 ;
    input inputs_348__8 ;
    input inputs_348__7 ;
    input inputs_348__6 ;
    input inputs_348__5 ;
    input inputs_348__4 ;
    input inputs_348__3 ;
    input inputs_348__2 ;
    input inputs_348__1 ;
    input inputs_348__0 ;
    input inputs_349__15 ;
    input inputs_349__14 ;
    input inputs_349__13 ;
    input inputs_349__12 ;
    input inputs_349__11 ;
    input inputs_349__10 ;
    input inputs_349__9 ;
    input inputs_349__8 ;
    input inputs_349__7 ;
    input inputs_349__6 ;
    input inputs_349__5 ;
    input inputs_349__4 ;
    input inputs_349__3 ;
    input inputs_349__2 ;
    input inputs_349__1 ;
    input inputs_349__0 ;
    input inputs_350__15 ;
    input inputs_350__14 ;
    input inputs_350__13 ;
    input inputs_350__12 ;
    input inputs_350__11 ;
    input inputs_350__10 ;
    input inputs_350__9 ;
    input inputs_350__8 ;
    input inputs_350__7 ;
    input inputs_350__6 ;
    input inputs_350__5 ;
    input inputs_350__4 ;
    input inputs_350__3 ;
    input inputs_350__2 ;
    input inputs_350__1 ;
    input inputs_350__0 ;
    input inputs_351__15 ;
    input inputs_351__14 ;
    input inputs_351__13 ;
    input inputs_351__12 ;
    input inputs_351__11 ;
    input inputs_351__10 ;
    input inputs_351__9 ;
    input inputs_351__8 ;
    input inputs_351__7 ;
    input inputs_351__6 ;
    input inputs_351__5 ;
    input inputs_351__4 ;
    input inputs_351__3 ;
    input inputs_351__2 ;
    input inputs_351__1 ;
    input inputs_351__0 ;
    input inputs_352__15 ;
    input inputs_352__14 ;
    input inputs_352__13 ;
    input inputs_352__12 ;
    input inputs_352__11 ;
    input inputs_352__10 ;
    input inputs_352__9 ;
    input inputs_352__8 ;
    input inputs_352__7 ;
    input inputs_352__6 ;
    input inputs_352__5 ;
    input inputs_352__4 ;
    input inputs_352__3 ;
    input inputs_352__2 ;
    input inputs_352__1 ;
    input inputs_352__0 ;
    input inputs_353__15 ;
    input inputs_353__14 ;
    input inputs_353__13 ;
    input inputs_353__12 ;
    input inputs_353__11 ;
    input inputs_353__10 ;
    input inputs_353__9 ;
    input inputs_353__8 ;
    input inputs_353__7 ;
    input inputs_353__6 ;
    input inputs_353__5 ;
    input inputs_353__4 ;
    input inputs_353__3 ;
    input inputs_353__2 ;
    input inputs_353__1 ;
    input inputs_353__0 ;
    input inputs_354__15 ;
    input inputs_354__14 ;
    input inputs_354__13 ;
    input inputs_354__12 ;
    input inputs_354__11 ;
    input inputs_354__10 ;
    input inputs_354__9 ;
    input inputs_354__8 ;
    input inputs_354__7 ;
    input inputs_354__6 ;
    input inputs_354__5 ;
    input inputs_354__4 ;
    input inputs_354__3 ;
    input inputs_354__2 ;
    input inputs_354__1 ;
    input inputs_354__0 ;
    input inputs_355__15 ;
    input inputs_355__14 ;
    input inputs_355__13 ;
    input inputs_355__12 ;
    input inputs_355__11 ;
    input inputs_355__10 ;
    input inputs_355__9 ;
    input inputs_355__8 ;
    input inputs_355__7 ;
    input inputs_355__6 ;
    input inputs_355__5 ;
    input inputs_355__4 ;
    input inputs_355__3 ;
    input inputs_355__2 ;
    input inputs_355__1 ;
    input inputs_355__0 ;
    input inputs_356__15 ;
    input inputs_356__14 ;
    input inputs_356__13 ;
    input inputs_356__12 ;
    input inputs_356__11 ;
    input inputs_356__10 ;
    input inputs_356__9 ;
    input inputs_356__8 ;
    input inputs_356__7 ;
    input inputs_356__6 ;
    input inputs_356__5 ;
    input inputs_356__4 ;
    input inputs_356__3 ;
    input inputs_356__2 ;
    input inputs_356__1 ;
    input inputs_356__0 ;
    input inputs_357__15 ;
    input inputs_357__14 ;
    input inputs_357__13 ;
    input inputs_357__12 ;
    input inputs_357__11 ;
    input inputs_357__10 ;
    input inputs_357__9 ;
    input inputs_357__8 ;
    input inputs_357__7 ;
    input inputs_357__6 ;
    input inputs_357__5 ;
    input inputs_357__4 ;
    input inputs_357__3 ;
    input inputs_357__2 ;
    input inputs_357__1 ;
    input inputs_357__0 ;
    input inputs_358__15 ;
    input inputs_358__14 ;
    input inputs_358__13 ;
    input inputs_358__12 ;
    input inputs_358__11 ;
    input inputs_358__10 ;
    input inputs_358__9 ;
    input inputs_358__8 ;
    input inputs_358__7 ;
    input inputs_358__6 ;
    input inputs_358__5 ;
    input inputs_358__4 ;
    input inputs_358__3 ;
    input inputs_358__2 ;
    input inputs_358__1 ;
    input inputs_358__0 ;
    input inputs_359__15 ;
    input inputs_359__14 ;
    input inputs_359__13 ;
    input inputs_359__12 ;
    input inputs_359__11 ;
    input inputs_359__10 ;
    input inputs_359__9 ;
    input inputs_359__8 ;
    input inputs_359__7 ;
    input inputs_359__6 ;
    input inputs_359__5 ;
    input inputs_359__4 ;
    input inputs_359__3 ;
    input inputs_359__2 ;
    input inputs_359__1 ;
    input inputs_359__0 ;
    input inputs_360__15 ;
    input inputs_360__14 ;
    input inputs_360__13 ;
    input inputs_360__12 ;
    input inputs_360__11 ;
    input inputs_360__10 ;
    input inputs_360__9 ;
    input inputs_360__8 ;
    input inputs_360__7 ;
    input inputs_360__6 ;
    input inputs_360__5 ;
    input inputs_360__4 ;
    input inputs_360__3 ;
    input inputs_360__2 ;
    input inputs_360__1 ;
    input inputs_360__0 ;
    input inputs_361__15 ;
    input inputs_361__14 ;
    input inputs_361__13 ;
    input inputs_361__12 ;
    input inputs_361__11 ;
    input inputs_361__10 ;
    input inputs_361__9 ;
    input inputs_361__8 ;
    input inputs_361__7 ;
    input inputs_361__6 ;
    input inputs_361__5 ;
    input inputs_361__4 ;
    input inputs_361__3 ;
    input inputs_361__2 ;
    input inputs_361__1 ;
    input inputs_361__0 ;
    input inputs_362__15 ;
    input inputs_362__14 ;
    input inputs_362__13 ;
    input inputs_362__12 ;
    input inputs_362__11 ;
    input inputs_362__10 ;
    input inputs_362__9 ;
    input inputs_362__8 ;
    input inputs_362__7 ;
    input inputs_362__6 ;
    input inputs_362__5 ;
    input inputs_362__4 ;
    input inputs_362__3 ;
    input inputs_362__2 ;
    input inputs_362__1 ;
    input inputs_362__0 ;
    input inputs_363__15 ;
    input inputs_363__14 ;
    input inputs_363__13 ;
    input inputs_363__12 ;
    input inputs_363__11 ;
    input inputs_363__10 ;
    input inputs_363__9 ;
    input inputs_363__8 ;
    input inputs_363__7 ;
    input inputs_363__6 ;
    input inputs_363__5 ;
    input inputs_363__4 ;
    input inputs_363__3 ;
    input inputs_363__2 ;
    input inputs_363__1 ;
    input inputs_363__0 ;
    input inputs_364__15 ;
    input inputs_364__14 ;
    input inputs_364__13 ;
    input inputs_364__12 ;
    input inputs_364__11 ;
    input inputs_364__10 ;
    input inputs_364__9 ;
    input inputs_364__8 ;
    input inputs_364__7 ;
    input inputs_364__6 ;
    input inputs_364__5 ;
    input inputs_364__4 ;
    input inputs_364__3 ;
    input inputs_364__2 ;
    input inputs_364__1 ;
    input inputs_364__0 ;
    input inputs_365__15 ;
    input inputs_365__14 ;
    input inputs_365__13 ;
    input inputs_365__12 ;
    input inputs_365__11 ;
    input inputs_365__10 ;
    input inputs_365__9 ;
    input inputs_365__8 ;
    input inputs_365__7 ;
    input inputs_365__6 ;
    input inputs_365__5 ;
    input inputs_365__4 ;
    input inputs_365__3 ;
    input inputs_365__2 ;
    input inputs_365__1 ;
    input inputs_365__0 ;
    input inputs_366__15 ;
    input inputs_366__14 ;
    input inputs_366__13 ;
    input inputs_366__12 ;
    input inputs_366__11 ;
    input inputs_366__10 ;
    input inputs_366__9 ;
    input inputs_366__8 ;
    input inputs_366__7 ;
    input inputs_366__6 ;
    input inputs_366__5 ;
    input inputs_366__4 ;
    input inputs_366__3 ;
    input inputs_366__2 ;
    input inputs_366__1 ;
    input inputs_366__0 ;
    input inputs_367__15 ;
    input inputs_367__14 ;
    input inputs_367__13 ;
    input inputs_367__12 ;
    input inputs_367__11 ;
    input inputs_367__10 ;
    input inputs_367__9 ;
    input inputs_367__8 ;
    input inputs_367__7 ;
    input inputs_367__6 ;
    input inputs_367__5 ;
    input inputs_367__4 ;
    input inputs_367__3 ;
    input inputs_367__2 ;
    input inputs_367__1 ;
    input inputs_367__0 ;
    input inputs_368__15 ;
    input inputs_368__14 ;
    input inputs_368__13 ;
    input inputs_368__12 ;
    input inputs_368__11 ;
    input inputs_368__10 ;
    input inputs_368__9 ;
    input inputs_368__8 ;
    input inputs_368__7 ;
    input inputs_368__6 ;
    input inputs_368__5 ;
    input inputs_368__4 ;
    input inputs_368__3 ;
    input inputs_368__2 ;
    input inputs_368__1 ;
    input inputs_368__0 ;
    input inputs_369__15 ;
    input inputs_369__14 ;
    input inputs_369__13 ;
    input inputs_369__12 ;
    input inputs_369__11 ;
    input inputs_369__10 ;
    input inputs_369__9 ;
    input inputs_369__8 ;
    input inputs_369__7 ;
    input inputs_369__6 ;
    input inputs_369__5 ;
    input inputs_369__4 ;
    input inputs_369__3 ;
    input inputs_369__2 ;
    input inputs_369__1 ;
    input inputs_369__0 ;
    input inputs_370__15 ;
    input inputs_370__14 ;
    input inputs_370__13 ;
    input inputs_370__12 ;
    input inputs_370__11 ;
    input inputs_370__10 ;
    input inputs_370__9 ;
    input inputs_370__8 ;
    input inputs_370__7 ;
    input inputs_370__6 ;
    input inputs_370__5 ;
    input inputs_370__4 ;
    input inputs_370__3 ;
    input inputs_370__2 ;
    input inputs_370__1 ;
    input inputs_370__0 ;
    input inputs_371__15 ;
    input inputs_371__14 ;
    input inputs_371__13 ;
    input inputs_371__12 ;
    input inputs_371__11 ;
    input inputs_371__10 ;
    input inputs_371__9 ;
    input inputs_371__8 ;
    input inputs_371__7 ;
    input inputs_371__6 ;
    input inputs_371__5 ;
    input inputs_371__4 ;
    input inputs_371__3 ;
    input inputs_371__2 ;
    input inputs_371__1 ;
    input inputs_371__0 ;
    input inputs_372__15 ;
    input inputs_372__14 ;
    input inputs_372__13 ;
    input inputs_372__12 ;
    input inputs_372__11 ;
    input inputs_372__10 ;
    input inputs_372__9 ;
    input inputs_372__8 ;
    input inputs_372__7 ;
    input inputs_372__6 ;
    input inputs_372__5 ;
    input inputs_372__4 ;
    input inputs_372__3 ;
    input inputs_372__2 ;
    input inputs_372__1 ;
    input inputs_372__0 ;
    input inputs_373__15 ;
    input inputs_373__14 ;
    input inputs_373__13 ;
    input inputs_373__12 ;
    input inputs_373__11 ;
    input inputs_373__10 ;
    input inputs_373__9 ;
    input inputs_373__8 ;
    input inputs_373__7 ;
    input inputs_373__6 ;
    input inputs_373__5 ;
    input inputs_373__4 ;
    input inputs_373__3 ;
    input inputs_373__2 ;
    input inputs_373__1 ;
    input inputs_373__0 ;
    input inputs_374__15 ;
    input inputs_374__14 ;
    input inputs_374__13 ;
    input inputs_374__12 ;
    input inputs_374__11 ;
    input inputs_374__10 ;
    input inputs_374__9 ;
    input inputs_374__8 ;
    input inputs_374__7 ;
    input inputs_374__6 ;
    input inputs_374__5 ;
    input inputs_374__4 ;
    input inputs_374__3 ;
    input inputs_374__2 ;
    input inputs_374__1 ;
    input inputs_374__0 ;
    input inputs_375__15 ;
    input inputs_375__14 ;
    input inputs_375__13 ;
    input inputs_375__12 ;
    input inputs_375__11 ;
    input inputs_375__10 ;
    input inputs_375__9 ;
    input inputs_375__8 ;
    input inputs_375__7 ;
    input inputs_375__6 ;
    input inputs_375__5 ;
    input inputs_375__4 ;
    input inputs_375__3 ;
    input inputs_375__2 ;
    input inputs_375__1 ;
    input inputs_375__0 ;
    input inputs_376__15 ;
    input inputs_376__14 ;
    input inputs_376__13 ;
    input inputs_376__12 ;
    input inputs_376__11 ;
    input inputs_376__10 ;
    input inputs_376__9 ;
    input inputs_376__8 ;
    input inputs_376__7 ;
    input inputs_376__6 ;
    input inputs_376__5 ;
    input inputs_376__4 ;
    input inputs_376__3 ;
    input inputs_376__2 ;
    input inputs_376__1 ;
    input inputs_376__0 ;
    input inputs_377__15 ;
    input inputs_377__14 ;
    input inputs_377__13 ;
    input inputs_377__12 ;
    input inputs_377__11 ;
    input inputs_377__10 ;
    input inputs_377__9 ;
    input inputs_377__8 ;
    input inputs_377__7 ;
    input inputs_377__6 ;
    input inputs_377__5 ;
    input inputs_377__4 ;
    input inputs_377__3 ;
    input inputs_377__2 ;
    input inputs_377__1 ;
    input inputs_377__0 ;
    input inputs_378__15 ;
    input inputs_378__14 ;
    input inputs_378__13 ;
    input inputs_378__12 ;
    input inputs_378__11 ;
    input inputs_378__10 ;
    input inputs_378__9 ;
    input inputs_378__8 ;
    input inputs_378__7 ;
    input inputs_378__6 ;
    input inputs_378__5 ;
    input inputs_378__4 ;
    input inputs_378__3 ;
    input inputs_378__2 ;
    input inputs_378__1 ;
    input inputs_378__0 ;
    input inputs_379__15 ;
    input inputs_379__14 ;
    input inputs_379__13 ;
    input inputs_379__12 ;
    input inputs_379__11 ;
    input inputs_379__10 ;
    input inputs_379__9 ;
    input inputs_379__8 ;
    input inputs_379__7 ;
    input inputs_379__6 ;
    input inputs_379__5 ;
    input inputs_379__4 ;
    input inputs_379__3 ;
    input inputs_379__2 ;
    input inputs_379__1 ;
    input inputs_379__0 ;
    input inputs_380__15 ;
    input inputs_380__14 ;
    input inputs_380__13 ;
    input inputs_380__12 ;
    input inputs_380__11 ;
    input inputs_380__10 ;
    input inputs_380__9 ;
    input inputs_380__8 ;
    input inputs_380__7 ;
    input inputs_380__6 ;
    input inputs_380__5 ;
    input inputs_380__4 ;
    input inputs_380__3 ;
    input inputs_380__2 ;
    input inputs_380__1 ;
    input inputs_380__0 ;
    input inputs_381__15 ;
    input inputs_381__14 ;
    input inputs_381__13 ;
    input inputs_381__12 ;
    input inputs_381__11 ;
    input inputs_381__10 ;
    input inputs_381__9 ;
    input inputs_381__8 ;
    input inputs_381__7 ;
    input inputs_381__6 ;
    input inputs_381__5 ;
    input inputs_381__4 ;
    input inputs_381__3 ;
    input inputs_381__2 ;
    input inputs_381__1 ;
    input inputs_381__0 ;
    input inputs_382__15 ;
    input inputs_382__14 ;
    input inputs_382__13 ;
    input inputs_382__12 ;
    input inputs_382__11 ;
    input inputs_382__10 ;
    input inputs_382__9 ;
    input inputs_382__8 ;
    input inputs_382__7 ;
    input inputs_382__6 ;
    input inputs_382__5 ;
    input inputs_382__4 ;
    input inputs_382__3 ;
    input inputs_382__2 ;
    input inputs_382__1 ;
    input inputs_382__0 ;
    input inputs_383__15 ;
    input inputs_383__14 ;
    input inputs_383__13 ;
    input inputs_383__12 ;
    input inputs_383__11 ;
    input inputs_383__10 ;
    input inputs_383__9 ;
    input inputs_383__8 ;
    input inputs_383__7 ;
    input inputs_383__6 ;
    input inputs_383__5 ;
    input inputs_383__4 ;
    input inputs_383__3 ;
    input inputs_383__2 ;
    input inputs_383__1 ;
    input inputs_383__0 ;
    input inputs_384__15 ;
    input inputs_384__14 ;
    input inputs_384__13 ;
    input inputs_384__12 ;
    input inputs_384__11 ;
    input inputs_384__10 ;
    input inputs_384__9 ;
    input inputs_384__8 ;
    input inputs_384__7 ;
    input inputs_384__6 ;
    input inputs_384__5 ;
    input inputs_384__4 ;
    input inputs_384__3 ;
    input inputs_384__2 ;
    input inputs_384__1 ;
    input inputs_384__0 ;
    input inputs_385__15 ;
    input inputs_385__14 ;
    input inputs_385__13 ;
    input inputs_385__12 ;
    input inputs_385__11 ;
    input inputs_385__10 ;
    input inputs_385__9 ;
    input inputs_385__8 ;
    input inputs_385__7 ;
    input inputs_385__6 ;
    input inputs_385__5 ;
    input inputs_385__4 ;
    input inputs_385__3 ;
    input inputs_385__2 ;
    input inputs_385__1 ;
    input inputs_385__0 ;
    input inputs_386__15 ;
    input inputs_386__14 ;
    input inputs_386__13 ;
    input inputs_386__12 ;
    input inputs_386__11 ;
    input inputs_386__10 ;
    input inputs_386__9 ;
    input inputs_386__8 ;
    input inputs_386__7 ;
    input inputs_386__6 ;
    input inputs_386__5 ;
    input inputs_386__4 ;
    input inputs_386__3 ;
    input inputs_386__2 ;
    input inputs_386__1 ;
    input inputs_386__0 ;
    input inputs_387__15 ;
    input inputs_387__14 ;
    input inputs_387__13 ;
    input inputs_387__12 ;
    input inputs_387__11 ;
    input inputs_387__10 ;
    input inputs_387__9 ;
    input inputs_387__8 ;
    input inputs_387__7 ;
    input inputs_387__6 ;
    input inputs_387__5 ;
    input inputs_387__4 ;
    input inputs_387__3 ;
    input inputs_387__2 ;
    input inputs_387__1 ;
    input inputs_387__0 ;
    input inputs_388__15 ;
    input inputs_388__14 ;
    input inputs_388__13 ;
    input inputs_388__12 ;
    input inputs_388__11 ;
    input inputs_388__10 ;
    input inputs_388__9 ;
    input inputs_388__8 ;
    input inputs_388__7 ;
    input inputs_388__6 ;
    input inputs_388__5 ;
    input inputs_388__4 ;
    input inputs_388__3 ;
    input inputs_388__2 ;
    input inputs_388__1 ;
    input inputs_388__0 ;
    input inputs_389__15 ;
    input inputs_389__14 ;
    input inputs_389__13 ;
    input inputs_389__12 ;
    input inputs_389__11 ;
    input inputs_389__10 ;
    input inputs_389__9 ;
    input inputs_389__8 ;
    input inputs_389__7 ;
    input inputs_389__6 ;
    input inputs_389__5 ;
    input inputs_389__4 ;
    input inputs_389__3 ;
    input inputs_389__2 ;
    input inputs_389__1 ;
    input inputs_389__0 ;
    input inputs_390__15 ;
    input inputs_390__14 ;
    input inputs_390__13 ;
    input inputs_390__12 ;
    input inputs_390__11 ;
    input inputs_390__10 ;
    input inputs_390__9 ;
    input inputs_390__8 ;
    input inputs_390__7 ;
    input inputs_390__6 ;
    input inputs_390__5 ;
    input inputs_390__4 ;
    input inputs_390__3 ;
    input inputs_390__2 ;
    input inputs_390__1 ;
    input inputs_390__0 ;
    input inputs_391__15 ;
    input inputs_391__14 ;
    input inputs_391__13 ;
    input inputs_391__12 ;
    input inputs_391__11 ;
    input inputs_391__10 ;
    input inputs_391__9 ;
    input inputs_391__8 ;
    input inputs_391__7 ;
    input inputs_391__6 ;
    input inputs_391__5 ;
    input inputs_391__4 ;
    input inputs_391__3 ;
    input inputs_391__2 ;
    input inputs_391__1 ;
    input inputs_391__0 ;
    input inputs_392__15 ;
    input inputs_392__14 ;
    input inputs_392__13 ;
    input inputs_392__12 ;
    input inputs_392__11 ;
    input inputs_392__10 ;
    input inputs_392__9 ;
    input inputs_392__8 ;
    input inputs_392__7 ;
    input inputs_392__6 ;
    input inputs_392__5 ;
    input inputs_392__4 ;
    input inputs_392__3 ;
    input inputs_392__2 ;
    input inputs_392__1 ;
    input inputs_392__0 ;
    input inputs_393__15 ;
    input inputs_393__14 ;
    input inputs_393__13 ;
    input inputs_393__12 ;
    input inputs_393__11 ;
    input inputs_393__10 ;
    input inputs_393__9 ;
    input inputs_393__8 ;
    input inputs_393__7 ;
    input inputs_393__6 ;
    input inputs_393__5 ;
    input inputs_393__4 ;
    input inputs_393__3 ;
    input inputs_393__2 ;
    input inputs_393__1 ;
    input inputs_393__0 ;
    input inputs_394__15 ;
    input inputs_394__14 ;
    input inputs_394__13 ;
    input inputs_394__12 ;
    input inputs_394__11 ;
    input inputs_394__10 ;
    input inputs_394__9 ;
    input inputs_394__8 ;
    input inputs_394__7 ;
    input inputs_394__6 ;
    input inputs_394__5 ;
    input inputs_394__4 ;
    input inputs_394__3 ;
    input inputs_394__2 ;
    input inputs_394__1 ;
    input inputs_394__0 ;
    input inputs_395__15 ;
    input inputs_395__14 ;
    input inputs_395__13 ;
    input inputs_395__12 ;
    input inputs_395__11 ;
    input inputs_395__10 ;
    input inputs_395__9 ;
    input inputs_395__8 ;
    input inputs_395__7 ;
    input inputs_395__6 ;
    input inputs_395__5 ;
    input inputs_395__4 ;
    input inputs_395__3 ;
    input inputs_395__2 ;
    input inputs_395__1 ;
    input inputs_395__0 ;
    input inputs_396__15 ;
    input inputs_396__14 ;
    input inputs_396__13 ;
    input inputs_396__12 ;
    input inputs_396__11 ;
    input inputs_396__10 ;
    input inputs_396__9 ;
    input inputs_396__8 ;
    input inputs_396__7 ;
    input inputs_396__6 ;
    input inputs_396__5 ;
    input inputs_396__4 ;
    input inputs_396__3 ;
    input inputs_396__2 ;
    input inputs_396__1 ;
    input inputs_396__0 ;
    input inputs_397__15 ;
    input inputs_397__14 ;
    input inputs_397__13 ;
    input inputs_397__12 ;
    input inputs_397__11 ;
    input inputs_397__10 ;
    input inputs_397__9 ;
    input inputs_397__8 ;
    input inputs_397__7 ;
    input inputs_397__6 ;
    input inputs_397__5 ;
    input inputs_397__4 ;
    input inputs_397__3 ;
    input inputs_397__2 ;
    input inputs_397__1 ;
    input inputs_397__0 ;
    input inputs_398__15 ;
    input inputs_398__14 ;
    input inputs_398__13 ;
    input inputs_398__12 ;
    input inputs_398__11 ;
    input inputs_398__10 ;
    input inputs_398__9 ;
    input inputs_398__8 ;
    input inputs_398__7 ;
    input inputs_398__6 ;
    input inputs_398__5 ;
    input inputs_398__4 ;
    input inputs_398__3 ;
    input inputs_398__2 ;
    input inputs_398__1 ;
    input inputs_398__0 ;
    input inputs_399__15 ;
    input inputs_399__14 ;
    input inputs_399__13 ;
    input inputs_399__12 ;
    input inputs_399__11 ;
    input inputs_399__10 ;
    input inputs_399__9 ;
    input inputs_399__8 ;
    input inputs_399__7 ;
    input inputs_399__6 ;
    input inputs_399__5 ;
    input inputs_399__4 ;
    input inputs_399__3 ;
    input inputs_399__2 ;
    input inputs_399__1 ;
    input inputs_399__0 ;
    input inputs_400__15 ;
    input inputs_400__14 ;
    input inputs_400__13 ;
    input inputs_400__12 ;
    input inputs_400__11 ;
    input inputs_400__10 ;
    input inputs_400__9 ;
    input inputs_400__8 ;
    input inputs_400__7 ;
    input inputs_400__6 ;
    input inputs_400__5 ;
    input inputs_400__4 ;
    input inputs_400__3 ;
    input inputs_400__2 ;
    input inputs_400__1 ;
    input inputs_400__0 ;
    input inputs_401__15 ;
    input inputs_401__14 ;
    input inputs_401__13 ;
    input inputs_401__12 ;
    input inputs_401__11 ;
    input inputs_401__10 ;
    input inputs_401__9 ;
    input inputs_401__8 ;
    input inputs_401__7 ;
    input inputs_401__6 ;
    input inputs_401__5 ;
    input inputs_401__4 ;
    input inputs_401__3 ;
    input inputs_401__2 ;
    input inputs_401__1 ;
    input inputs_401__0 ;
    input inputs_402__15 ;
    input inputs_402__14 ;
    input inputs_402__13 ;
    input inputs_402__12 ;
    input inputs_402__11 ;
    input inputs_402__10 ;
    input inputs_402__9 ;
    input inputs_402__8 ;
    input inputs_402__7 ;
    input inputs_402__6 ;
    input inputs_402__5 ;
    input inputs_402__4 ;
    input inputs_402__3 ;
    input inputs_402__2 ;
    input inputs_402__1 ;
    input inputs_402__0 ;
    input inputs_403__15 ;
    input inputs_403__14 ;
    input inputs_403__13 ;
    input inputs_403__12 ;
    input inputs_403__11 ;
    input inputs_403__10 ;
    input inputs_403__9 ;
    input inputs_403__8 ;
    input inputs_403__7 ;
    input inputs_403__6 ;
    input inputs_403__5 ;
    input inputs_403__4 ;
    input inputs_403__3 ;
    input inputs_403__2 ;
    input inputs_403__1 ;
    input inputs_403__0 ;
    input inputs_404__15 ;
    input inputs_404__14 ;
    input inputs_404__13 ;
    input inputs_404__12 ;
    input inputs_404__11 ;
    input inputs_404__10 ;
    input inputs_404__9 ;
    input inputs_404__8 ;
    input inputs_404__7 ;
    input inputs_404__6 ;
    input inputs_404__5 ;
    input inputs_404__4 ;
    input inputs_404__3 ;
    input inputs_404__2 ;
    input inputs_404__1 ;
    input inputs_404__0 ;
    input inputs_405__15 ;
    input inputs_405__14 ;
    input inputs_405__13 ;
    input inputs_405__12 ;
    input inputs_405__11 ;
    input inputs_405__10 ;
    input inputs_405__9 ;
    input inputs_405__8 ;
    input inputs_405__7 ;
    input inputs_405__6 ;
    input inputs_405__5 ;
    input inputs_405__4 ;
    input inputs_405__3 ;
    input inputs_405__2 ;
    input inputs_405__1 ;
    input inputs_405__0 ;
    input inputs_406__15 ;
    input inputs_406__14 ;
    input inputs_406__13 ;
    input inputs_406__12 ;
    input inputs_406__11 ;
    input inputs_406__10 ;
    input inputs_406__9 ;
    input inputs_406__8 ;
    input inputs_406__7 ;
    input inputs_406__6 ;
    input inputs_406__5 ;
    input inputs_406__4 ;
    input inputs_406__3 ;
    input inputs_406__2 ;
    input inputs_406__1 ;
    input inputs_406__0 ;
    input inputs_407__15 ;
    input inputs_407__14 ;
    input inputs_407__13 ;
    input inputs_407__12 ;
    input inputs_407__11 ;
    input inputs_407__10 ;
    input inputs_407__9 ;
    input inputs_407__8 ;
    input inputs_407__7 ;
    input inputs_407__6 ;
    input inputs_407__5 ;
    input inputs_407__4 ;
    input inputs_407__3 ;
    input inputs_407__2 ;
    input inputs_407__1 ;
    input inputs_407__0 ;
    input inputs_408__15 ;
    input inputs_408__14 ;
    input inputs_408__13 ;
    input inputs_408__12 ;
    input inputs_408__11 ;
    input inputs_408__10 ;
    input inputs_408__9 ;
    input inputs_408__8 ;
    input inputs_408__7 ;
    input inputs_408__6 ;
    input inputs_408__5 ;
    input inputs_408__4 ;
    input inputs_408__3 ;
    input inputs_408__2 ;
    input inputs_408__1 ;
    input inputs_408__0 ;
    input inputs_409__15 ;
    input inputs_409__14 ;
    input inputs_409__13 ;
    input inputs_409__12 ;
    input inputs_409__11 ;
    input inputs_409__10 ;
    input inputs_409__9 ;
    input inputs_409__8 ;
    input inputs_409__7 ;
    input inputs_409__6 ;
    input inputs_409__5 ;
    input inputs_409__4 ;
    input inputs_409__3 ;
    input inputs_409__2 ;
    input inputs_409__1 ;
    input inputs_409__0 ;
    input inputs_410__15 ;
    input inputs_410__14 ;
    input inputs_410__13 ;
    input inputs_410__12 ;
    input inputs_410__11 ;
    input inputs_410__10 ;
    input inputs_410__9 ;
    input inputs_410__8 ;
    input inputs_410__7 ;
    input inputs_410__6 ;
    input inputs_410__5 ;
    input inputs_410__4 ;
    input inputs_410__3 ;
    input inputs_410__2 ;
    input inputs_410__1 ;
    input inputs_410__0 ;
    input inputs_411__15 ;
    input inputs_411__14 ;
    input inputs_411__13 ;
    input inputs_411__12 ;
    input inputs_411__11 ;
    input inputs_411__10 ;
    input inputs_411__9 ;
    input inputs_411__8 ;
    input inputs_411__7 ;
    input inputs_411__6 ;
    input inputs_411__5 ;
    input inputs_411__4 ;
    input inputs_411__3 ;
    input inputs_411__2 ;
    input inputs_411__1 ;
    input inputs_411__0 ;
    input inputs_412__15 ;
    input inputs_412__14 ;
    input inputs_412__13 ;
    input inputs_412__12 ;
    input inputs_412__11 ;
    input inputs_412__10 ;
    input inputs_412__9 ;
    input inputs_412__8 ;
    input inputs_412__7 ;
    input inputs_412__6 ;
    input inputs_412__5 ;
    input inputs_412__4 ;
    input inputs_412__3 ;
    input inputs_412__2 ;
    input inputs_412__1 ;
    input inputs_412__0 ;
    input inputs_413__15 ;
    input inputs_413__14 ;
    input inputs_413__13 ;
    input inputs_413__12 ;
    input inputs_413__11 ;
    input inputs_413__10 ;
    input inputs_413__9 ;
    input inputs_413__8 ;
    input inputs_413__7 ;
    input inputs_413__6 ;
    input inputs_413__5 ;
    input inputs_413__4 ;
    input inputs_413__3 ;
    input inputs_413__2 ;
    input inputs_413__1 ;
    input inputs_413__0 ;
    input inputs_414__15 ;
    input inputs_414__14 ;
    input inputs_414__13 ;
    input inputs_414__12 ;
    input inputs_414__11 ;
    input inputs_414__10 ;
    input inputs_414__9 ;
    input inputs_414__8 ;
    input inputs_414__7 ;
    input inputs_414__6 ;
    input inputs_414__5 ;
    input inputs_414__4 ;
    input inputs_414__3 ;
    input inputs_414__2 ;
    input inputs_414__1 ;
    input inputs_414__0 ;
    input inputs_415__15 ;
    input inputs_415__14 ;
    input inputs_415__13 ;
    input inputs_415__12 ;
    input inputs_415__11 ;
    input inputs_415__10 ;
    input inputs_415__9 ;
    input inputs_415__8 ;
    input inputs_415__7 ;
    input inputs_415__6 ;
    input inputs_415__5 ;
    input inputs_415__4 ;
    input inputs_415__3 ;
    input inputs_415__2 ;
    input inputs_415__1 ;
    input inputs_415__0 ;
    input inputs_416__15 ;
    input inputs_416__14 ;
    input inputs_416__13 ;
    input inputs_416__12 ;
    input inputs_416__11 ;
    input inputs_416__10 ;
    input inputs_416__9 ;
    input inputs_416__8 ;
    input inputs_416__7 ;
    input inputs_416__6 ;
    input inputs_416__5 ;
    input inputs_416__4 ;
    input inputs_416__3 ;
    input inputs_416__2 ;
    input inputs_416__1 ;
    input inputs_416__0 ;
    input inputs_417__15 ;
    input inputs_417__14 ;
    input inputs_417__13 ;
    input inputs_417__12 ;
    input inputs_417__11 ;
    input inputs_417__10 ;
    input inputs_417__9 ;
    input inputs_417__8 ;
    input inputs_417__7 ;
    input inputs_417__6 ;
    input inputs_417__5 ;
    input inputs_417__4 ;
    input inputs_417__3 ;
    input inputs_417__2 ;
    input inputs_417__1 ;
    input inputs_417__0 ;
    input inputs_418__15 ;
    input inputs_418__14 ;
    input inputs_418__13 ;
    input inputs_418__12 ;
    input inputs_418__11 ;
    input inputs_418__10 ;
    input inputs_418__9 ;
    input inputs_418__8 ;
    input inputs_418__7 ;
    input inputs_418__6 ;
    input inputs_418__5 ;
    input inputs_418__4 ;
    input inputs_418__3 ;
    input inputs_418__2 ;
    input inputs_418__1 ;
    input inputs_418__0 ;
    input inputs_419__15 ;
    input inputs_419__14 ;
    input inputs_419__13 ;
    input inputs_419__12 ;
    input inputs_419__11 ;
    input inputs_419__10 ;
    input inputs_419__9 ;
    input inputs_419__8 ;
    input inputs_419__7 ;
    input inputs_419__6 ;
    input inputs_419__5 ;
    input inputs_419__4 ;
    input inputs_419__3 ;
    input inputs_419__2 ;
    input inputs_419__1 ;
    input inputs_419__0 ;
    input inputs_420__15 ;
    input inputs_420__14 ;
    input inputs_420__13 ;
    input inputs_420__12 ;
    input inputs_420__11 ;
    input inputs_420__10 ;
    input inputs_420__9 ;
    input inputs_420__8 ;
    input inputs_420__7 ;
    input inputs_420__6 ;
    input inputs_420__5 ;
    input inputs_420__4 ;
    input inputs_420__3 ;
    input inputs_420__2 ;
    input inputs_420__1 ;
    input inputs_420__0 ;
    input inputs_421__15 ;
    input inputs_421__14 ;
    input inputs_421__13 ;
    input inputs_421__12 ;
    input inputs_421__11 ;
    input inputs_421__10 ;
    input inputs_421__9 ;
    input inputs_421__8 ;
    input inputs_421__7 ;
    input inputs_421__6 ;
    input inputs_421__5 ;
    input inputs_421__4 ;
    input inputs_421__3 ;
    input inputs_421__2 ;
    input inputs_421__1 ;
    input inputs_421__0 ;
    input inputs_422__15 ;
    input inputs_422__14 ;
    input inputs_422__13 ;
    input inputs_422__12 ;
    input inputs_422__11 ;
    input inputs_422__10 ;
    input inputs_422__9 ;
    input inputs_422__8 ;
    input inputs_422__7 ;
    input inputs_422__6 ;
    input inputs_422__5 ;
    input inputs_422__4 ;
    input inputs_422__3 ;
    input inputs_422__2 ;
    input inputs_422__1 ;
    input inputs_422__0 ;
    input inputs_423__15 ;
    input inputs_423__14 ;
    input inputs_423__13 ;
    input inputs_423__12 ;
    input inputs_423__11 ;
    input inputs_423__10 ;
    input inputs_423__9 ;
    input inputs_423__8 ;
    input inputs_423__7 ;
    input inputs_423__6 ;
    input inputs_423__5 ;
    input inputs_423__4 ;
    input inputs_423__3 ;
    input inputs_423__2 ;
    input inputs_423__1 ;
    input inputs_423__0 ;
    input inputs_424__15 ;
    input inputs_424__14 ;
    input inputs_424__13 ;
    input inputs_424__12 ;
    input inputs_424__11 ;
    input inputs_424__10 ;
    input inputs_424__9 ;
    input inputs_424__8 ;
    input inputs_424__7 ;
    input inputs_424__6 ;
    input inputs_424__5 ;
    input inputs_424__4 ;
    input inputs_424__3 ;
    input inputs_424__2 ;
    input inputs_424__1 ;
    input inputs_424__0 ;
    input inputs_425__15 ;
    input inputs_425__14 ;
    input inputs_425__13 ;
    input inputs_425__12 ;
    input inputs_425__11 ;
    input inputs_425__10 ;
    input inputs_425__9 ;
    input inputs_425__8 ;
    input inputs_425__7 ;
    input inputs_425__6 ;
    input inputs_425__5 ;
    input inputs_425__4 ;
    input inputs_425__3 ;
    input inputs_425__2 ;
    input inputs_425__1 ;
    input inputs_425__0 ;
    input inputs_426__15 ;
    input inputs_426__14 ;
    input inputs_426__13 ;
    input inputs_426__12 ;
    input inputs_426__11 ;
    input inputs_426__10 ;
    input inputs_426__9 ;
    input inputs_426__8 ;
    input inputs_426__7 ;
    input inputs_426__6 ;
    input inputs_426__5 ;
    input inputs_426__4 ;
    input inputs_426__3 ;
    input inputs_426__2 ;
    input inputs_426__1 ;
    input inputs_426__0 ;
    input inputs_427__15 ;
    input inputs_427__14 ;
    input inputs_427__13 ;
    input inputs_427__12 ;
    input inputs_427__11 ;
    input inputs_427__10 ;
    input inputs_427__9 ;
    input inputs_427__8 ;
    input inputs_427__7 ;
    input inputs_427__6 ;
    input inputs_427__5 ;
    input inputs_427__4 ;
    input inputs_427__3 ;
    input inputs_427__2 ;
    input inputs_427__1 ;
    input inputs_427__0 ;
    input inputs_428__15 ;
    input inputs_428__14 ;
    input inputs_428__13 ;
    input inputs_428__12 ;
    input inputs_428__11 ;
    input inputs_428__10 ;
    input inputs_428__9 ;
    input inputs_428__8 ;
    input inputs_428__7 ;
    input inputs_428__6 ;
    input inputs_428__5 ;
    input inputs_428__4 ;
    input inputs_428__3 ;
    input inputs_428__2 ;
    input inputs_428__1 ;
    input inputs_428__0 ;
    input inputs_429__15 ;
    input inputs_429__14 ;
    input inputs_429__13 ;
    input inputs_429__12 ;
    input inputs_429__11 ;
    input inputs_429__10 ;
    input inputs_429__9 ;
    input inputs_429__8 ;
    input inputs_429__7 ;
    input inputs_429__6 ;
    input inputs_429__5 ;
    input inputs_429__4 ;
    input inputs_429__3 ;
    input inputs_429__2 ;
    input inputs_429__1 ;
    input inputs_429__0 ;
    input inputs_430__15 ;
    input inputs_430__14 ;
    input inputs_430__13 ;
    input inputs_430__12 ;
    input inputs_430__11 ;
    input inputs_430__10 ;
    input inputs_430__9 ;
    input inputs_430__8 ;
    input inputs_430__7 ;
    input inputs_430__6 ;
    input inputs_430__5 ;
    input inputs_430__4 ;
    input inputs_430__3 ;
    input inputs_430__2 ;
    input inputs_430__1 ;
    input inputs_430__0 ;
    input inputs_431__15 ;
    input inputs_431__14 ;
    input inputs_431__13 ;
    input inputs_431__12 ;
    input inputs_431__11 ;
    input inputs_431__10 ;
    input inputs_431__9 ;
    input inputs_431__8 ;
    input inputs_431__7 ;
    input inputs_431__6 ;
    input inputs_431__5 ;
    input inputs_431__4 ;
    input inputs_431__3 ;
    input inputs_431__2 ;
    input inputs_431__1 ;
    input inputs_431__0 ;
    input inputs_432__15 ;
    input inputs_432__14 ;
    input inputs_432__13 ;
    input inputs_432__12 ;
    input inputs_432__11 ;
    input inputs_432__10 ;
    input inputs_432__9 ;
    input inputs_432__8 ;
    input inputs_432__7 ;
    input inputs_432__6 ;
    input inputs_432__5 ;
    input inputs_432__4 ;
    input inputs_432__3 ;
    input inputs_432__2 ;
    input inputs_432__1 ;
    input inputs_432__0 ;
    input inputs_433__15 ;
    input inputs_433__14 ;
    input inputs_433__13 ;
    input inputs_433__12 ;
    input inputs_433__11 ;
    input inputs_433__10 ;
    input inputs_433__9 ;
    input inputs_433__8 ;
    input inputs_433__7 ;
    input inputs_433__6 ;
    input inputs_433__5 ;
    input inputs_433__4 ;
    input inputs_433__3 ;
    input inputs_433__2 ;
    input inputs_433__1 ;
    input inputs_433__0 ;
    input inputs_434__15 ;
    input inputs_434__14 ;
    input inputs_434__13 ;
    input inputs_434__12 ;
    input inputs_434__11 ;
    input inputs_434__10 ;
    input inputs_434__9 ;
    input inputs_434__8 ;
    input inputs_434__7 ;
    input inputs_434__6 ;
    input inputs_434__5 ;
    input inputs_434__4 ;
    input inputs_434__3 ;
    input inputs_434__2 ;
    input inputs_434__1 ;
    input inputs_434__0 ;
    input inputs_435__15 ;
    input inputs_435__14 ;
    input inputs_435__13 ;
    input inputs_435__12 ;
    input inputs_435__11 ;
    input inputs_435__10 ;
    input inputs_435__9 ;
    input inputs_435__8 ;
    input inputs_435__7 ;
    input inputs_435__6 ;
    input inputs_435__5 ;
    input inputs_435__4 ;
    input inputs_435__3 ;
    input inputs_435__2 ;
    input inputs_435__1 ;
    input inputs_435__0 ;
    input inputs_436__15 ;
    input inputs_436__14 ;
    input inputs_436__13 ;
    input inputs_436__12 ;
    input inputs_436__11 ;
    input inputs_436__10 ;
    input inputs_436__9 ;
    input inputs_436__8 ;
    input inputs_436__7 ;
    input inputs_436__6 ;
    input inputs_436__5 ;
    input inputs_436__4 ;
    input inputs_436__3 ;
    input inputs_436__2 ;
    input inputs_436__1 ;
    input inputs_436__0 ;
    input inputs_437__15 ;
    input inputs_437__14 ;
    input inputs_437__13 ;
    input inputs_437__12 ;
    input inputs_437__11 ;
    input inputs_437__10 ;
    input inputs_437__9 ;
    input inputs_437__8 ;
    input inputs_437__7 ;
    input inputs_437__6 ;
    input inputs_437__5 ;
    input inputs_437__4 ;
    input inputs_437__3 ;
    input inputs_437__2 ;
    input inputs_437__1 ;
    input inputs_437__0 ;
    input inputs_438__15 ;
    input inputs_438__14 ;
    input inputs_438__13 ;
    input inputs_438__12 ;
    input inputs_438__11 ;
    input inputs_438__10 ;
    input inputs_438__9 ;
    input inputs_438__8 ;
    input inputs_438__7 ;
    input inputs_438__6 ;
    input inputs_438__5 ;
    input inputs_438__4 ;
    input inputs_438__3 ;
    input inputs_438__2 ;
    input inputs_438__1 ;
    input inputs_438__0 ;
    input inputs_439__15 ;
    input inputs_439__14 ;
    input inputs_439__13 ;
    input inputs_439__12 ;
    input inputs_439__11 ;
    input inputs_439__10 ;
    input inputs_439__9 ;
    input inputs_439__8 ;
    input inputs_439__7 ;
    input inputs_439__6 ;
    input inputs_439__5 ;
    input inputs_439__4 ;
    input inputs_439__3 ;
    input inputs_439__2 ;
    input inputs_439__1 ;
    input inputs_439__0 ;
    input inputs_440__15 ;
    input inputs_440__14 ;
    input inputs_440__13 ;
    input inputs_440__12 ;
    input inputs_440__11 ;
    input inputs_440__10 ;
    input inputs_440__9 ;
    input inputs_440__8 ;
    input inputs_440__7 ;
    input inputs_440__6 ;
    input inputs_440__5 ;
    input inputs_440__4 ;
    input inputs_440__3 ;
    input inputs_440__2 ;
    input inputs_440__1 ;
    input inputs_440__0 ;
    input inputs_441__15 ;
    input inputs_441__14 ;
    input inputs_441__13 ;
    input inputs_441__12 ;
    input inputs_441__11 ;
    input inputs_441__10 ;
    input inputs_441__9 ;
    input inputs_441__8 ;
    input inputs_441__7 ;
    input inputs_441__6 ;
    input inputs_441__5 ;
    input inputs_441__4 ;
    input inputs_441__3 ;
    input inputs_441__2 ;
    input inputs_441__1 ;
    input inputs_441__0 ;
    input inputs_442__15 ;
    input inputs_442__14 ;
    input inputs_442__13 ;
    input inputs_442__12 ;
    input inputs_442__11 ;
    input inputs_442__10 ;
    input inputs_442__9 ;
    input inputs_442__8 ;
    input inputs_442__7 ;
    input inputs_442__6 ;
    input inputs_442__5 ;
    input inputs_442__4 ;
    input inputs_442__3 ;
    input inputs_442__2 ;
    input inputs_442__1 ;
    input inputs_442__0 ;
    input inputs_443__15 ;
    input inputs_443__14 ;
    input inputs_443__13 ;
    input inputs_443__12 ;
    input inputs_443__11 ;
    input inputs_443__10 ;
    input inputs_443__9 ;
    input inputs_443__8 ;
    input inputs_443__7 ;
    input inputs_443__6 ;
    input inputs_443__5 ;
    input inputs_443__4 ;
    input inputs_443__3 ;
    input inputs_443__2 ;
    input inputs_443__1 ;
    input inputs_443__0 ;
    input inputs_444__15 ;
    input inputs_444__14 ;
    input inputs_444__13 ;
    input inputs_444__12 ;
    input inputs_444__11 ;
    input inputs_444__10 ;
    input inputs_444__9 ;
    input inputs_444__8 ;
    input inputs_444__7 ;
    input inputs_444__6 ;
    input inputs_444__5 ;
    input inputs_444__4 ;
    input inputs_444__3 ;
    input inputs_444__2 ;
    input inputs_444__1 ;
    input inputs_444__0 ;
    input inputs_445__15 ;
    input inputs_445__14 ;
    input inputs_445__13 ;
    input inputs_445__12 ;
    input inputs_445__11 ;
    input inputs_445__10 ;
    input inputs_445__9 ;
    input inputs_445__8 ;
    input inputs_445__7 ;
    input inputs_445__6 ;
    input inputs_445__5 ;
    input inputs_445__4 ;
    input inputs_445__3 ;
    input inputs_445__2 ;
    input inputs_445__1 ;
    input inputs_445__0 ;
    input inputs_446__15 ;
    input inputs_446__14 ;
    input inputs_446__13 ;
    input inputs_446__12 ;
    input inputs_446__11 ;
    input inputs_446__10 ;
    input inputs_446__9 ;
    input inputs_446__8 ;
    input inputs_446__7 ;
    input inputs_446__6 ;
    input inputs_446__5 ;
    input inputs_446__4 ;
    input inputs_446__3 ;
    input inputs_446__2 ;
    input inputs_446__1 ;
    input inputs_446__0 ;
    input inputs_447__15 ;
    input inputs_447__14 ;
    input inputs_447__13 ;
    input inputs_447__12 ;
    input inputs_447__11 ;
    input inputs_447__10 ;
    input inputs_447__9 ;
    input inputs_447__8 ;
    input inputs_447__7 ;
    input inputs_447__6 ;
    input inputs_447__5 ;
    input inputs_447__4 ;
    input inputs_447__3 ;
    input inputs_447__2 ;
    input inputs_447__1 ;
    input inputs_447__0 ;
    input inputs_448__15 ;
    input inputs_448__14 ;
    input inputs_448__13 ;
    input inputs_448__12 ;
    input inputs_448__11 ;
    input inputs_448__10 ;
    input inputs_448__9 ;
    input inputs_448__8 ;
    input inputs_448__7 ;
    input inputs_448__6 ;
    input inputs_448__5 ;
    input inputs_448__4 ;
    input inputs_448__3 ;
    input inputs_448__2 ;
    input inputs_448__1 ;
    input inputs_448__0 ;
    input inputs_449__15 ;
    input inputs_449__14 ;
    input inputs_449__13 ;
    input inputs_449__12 ;
    input inputs_449__11 ;
    input inputs_449__10 ;
    input inputs_449__9 ;
    input inputs_449__8 ;
    input inputs_449__7 ;
    input inputs_449__6 ;
    input inputs_449__5 ;
    input inputs_449__4 ;
    input inputs_449__3 ;
    input inputs_449__2 ;
    input inputs_449__1 ;
    input inputs_449__0 ;
    input inputs_450__15 ;
    input inputs_450__14 ;
    input inputs_450__13 ;
    input inputs_450__12 ;
    input inputs_450__11 ;
    input inputs_450__10 ;
    input inputs_450__9 ;
    input inputs_450__8 ;
    input inputs_450__7 ;
    input inputs_450__6 ;
    input inputs_450__5 ;
    input inputs_450__4 ;
    input inputs_450__3 ;
    input inputs_450__2 ;
    input inputs_450__1 ;
    input inputs_450__0 ;
    input inputs_451__15 ;
    input inputs_451__14 ;
    input inputs_451__13 ;
    input inputs_451__12 ;
    input inputs_451__11 ;
    input inputs_451__10 ;
    input inputs_451__9 ;
    input inputs_451__8 ;
    input inputs_451__7 ;
    input inputs_451__6 ;
    input inputs_451__5 ;
    input inputs_451__4 ;
    input inputs_451__3 ;
    input inputs_451__2 ;
    input inputs_451__1 ;
    input inputs_451__0 ;
    input inputs_452__15 ;
    input inputs_452__14 ;
    input inputs_452__13 ;
    input inputs_452__12 ;
    input inputs_452__11 ;
    input inputs_452__10 ;
    input inputs_452__9 ;
    input inputs_452__8 ;
    input inputs_452__7 ;
    input inputs_452__6 ;
    input inputs_452__5 ;
    input inputs_452__4 ;
    input inputs_452__3 ;
    input inputs_452__2 ;
    input inputs_452__1 ;
    input inputs_452__0 ;
    input inputs_453__15 ;
    input inputs_453__14 ;
    input inputs_453__13 ;
    input inputs_453__12 ;
    input inputs_453__11 ;
    input inputs_453__10 ;
    input inputs_453__9 ;
    input inputs_453__8 ;
    input inputs_453__7 ;
    input inputs_453__6 ;
    input inputs_453__5 ;
    input inputs_453__4 ;
    input inputs_453__3 ;
    input inputs_453__2 ;
    input inputs_453__1 ;
    input inputs_453__0 ;
    input inputs_454__15 ;
    input inputs_454__14 ;
    input inputs_454__13 ;
    input inputs_454__12 ;
    input inputs_454__11 ;
    input inputs_454__10 ;
    input inputs_454__9 ;
    input inputs_454__8 ;
    input inputs_454__7 ;
    input inputs_454__6 ;
    input inputs_454__5 ;
    input inputs_454__4 ;
    input inputs_454__3 ;
    input inputs_454__2 ;
    input inputs_454__1 ;
    input inputs_454__0 ;
    input inputs_455__15 ;
    input inputs_455__14 ;
    input inputs_455__13 ;
    input inputs_455__12 ;
    input inputs_455__11 ;
    input inputs_455__10 ;
    input inputs_455__9 ;
    input inputs_455__8 ;
    input inputs_455__7 ;
    input inputs_455__6 ;
    input inputs_455__5 ;
    input inputs_455__4 ;
    input inputs_455__3 ;
    input inputs_455__2 ;
    input inputs_455__1 ;
    input inputs_455__0 ;
    input inputs_456__15 ;
    input inputs_456__14 ;
    input inputs_456__13 ;
    input inputs_456__12 ;
    input inputs_456__11 ;
    input inputs_456__10 ;
    input inputs_456__9 ;
    input inputs_456__8 ;
    input inputs_456__7 ;
    input inputs_456__6 ;
    input inputs_456__5 ;
    input inputs_456__4 ;
    input inputs_456__3 ;
    input inputs_456__2 ;
    input inputs_456__1 ;
    input inputs_456__0 ;
    input inputs_457__15 ;
    input inputs_457__14 ;
    input inputs_457__13 ;
    input inputs_457__12 ;
    input inputs_457__11 ;
    input inputs_457__10 ;
    input inputs_457__9 ;
    input inputs_457__8 ;
    input inputs_457__7 ;
    input inputs_457__6 ;
    input inputs_457__5 ;
    input inputs_457__4 ;
    input inputs_457__3 ;
    input inputs_457__2 ;
    input inputs_457__1 ;
    input inputs_457__0 ;
    input inputs_458__15 ;
    input inputs_458__14 ;
    input inputs_458__13 ;
    input inputs_458__12 ;
    input inputs_458__11 ;
    input inputs_458__10 ;
    input inputs_458__9 ;
    input inputs_458__8 ;
    input inputs_458__7 ;
    input inputs_458__6 ;
    input inputs_458__5 ;
    input inputs_458__4 ;
    input inputs_458__3 ;
    input inputs_458__2 ;
    input inputs_458__1 ;
    input inputs_458__0 ;
    input inputs_459__15 ;
    input inputs_459__14 ;
    input inputs_459__13 ;
    input inputs_459__12 ;
    input inputs_459__11 ;
    input inputs_459__10 ;
    input inputs_459__9 ;
    input inputs_459__8 ;
    input inputs_459__7 ;
    input inputs_459__6 ;
    input inputs_459__5 ;
    input inputs_459__4 ;
    input inputs_459__3 ;
    input inputs_459__2 ;
    input inputs_459__1 ;
    input inputs_459__0 ;
    input inputs_460__15 ;
    input inputs_460__14 ;
    input inputs_460__13 ;
    input inputs_460__12 ;
    input inputs_460__11 ;
    input inputs_460__10 ;
    input inputs_460__9 ;
    input inputs_460__8 ;
    input inputs_460__7 ;
    input inputs_460__6 ;
    input inputs_460__5 ;
    input inputs_460__4 ;
    input inputs_460__3 ;
    input inputs_460__2 ;
    input inputs_460__1 ;
    input inputs_460__0 ;
    input inputs_461__15 ;
    input inputs_461__14 ;
    input inputs_461__13 ;
    input inputs_461__12 ;
    input inputs_461__11 ;
    input inputs_461__10 ;
    input inputs_461__9 ;
    input inputs_461__8 ;
    input inputs_461__7 ;
    input inputs_461__6 ;
    input inputs_461__5 ;
    input inputs_461__4 ;
    input inputs_461__3 ;
    input inputs_461__2 ;
    input inputs_461__1 ;
    input inputs_461__0 ;
    input inputs_462__15 ;
    input inputs_462__14 ;
    input inputs_462__13 ;
    input inputs_462__12 ;
    input inputs_462__11 ;
    input inputs_462__10 ;
    input inputs_462__9 ;
    input inputs_462__8 ;
    input inputs_462__7 ;
    input inputs_462__6 ;
    input inputs_462__5 ;
    input inputs_462__4 ;
    input inputs_462__3 ;
    input inputs_462__2 ;
    input inputs_462__1 ;
    input inputs_462__0 ;
    input inputs_463__15 ;
    input inputs_463__14 ;
    input inputs_463__13 ;
    input inputs_463__12 ;
    input inputs_463__11 ;
    input inputs_463__10 ;
    input inputs_463__9 ;
    input inputs_463__8 ;
    input inputs_463__7 ;
    input inputs_463__6 ;
    input inputs_463__5 ;
    input inputs_463__4 ;
    input inputs_463__3 ;
    input inputs_463__2 ;
    input inputs_463__1 ;
    input inputs_463__0 ;
    input inputs_464__15 ;
    input inputs_464__14 ;
    input inputs_464__13 ;
    input inputs_464__12 ;
    input inputs_464__11 ;
    input inputs_464__10 ;
    input inputs_464__9 ;
    input inputs_464__8 ;
    input inputs_464__7 ;
    input inputs_464__6 ;
    input inputs_464__5 ;
    input inputs_464__4 ;
    input inputs_464__3 ;
    input inputs_464__2 ;
    input inputs_464__1 ;
    input inputs_464__0 ;
    input inputs_465__15 ;
    input inputs_465__14 ;
    input inputs_465__13 ;
    input inputs_465__12 ;
    input inputs_465__11 ;
    input inputs_465__10 ;
    input inputs_465__9 ;
    input inputs_465__8 ;
    input inputs_465__7 ;
    input inputs_465__6 ;
    input inputs_465__5 ;
    input inputs_465__4 ;
    input inputs_465__3 ;
    input inputs_465__2 ;
    input inputs_465__1 ;
    input inputs_465__0 ;
    input inputs_466__15 ;
    input inputs_466__14 ;
    input inputs_466__13 ;
    input inputs_466__12 ;
    input inputs_466__11 ;
    input inputs_466__10 ;
    input inputs_466__9 ;
    input inputs_466__8 ;
    input inputs_466__7 ;
    input inputs_466__6 ;
    input inputs_466__5 ;
    input inputs_466__4 ;
    input inputs_466__3 ;
    input inputs_466__2 ;
    input inputs_466__1 ;
    input inputs_466__0 ;
    input inputs_467__15 ;
    input inputs_467__14 ;
    input inputs_467__13 ;
    input inputs_467__12 ;
    input inputs_467__11 ;
    input inputs_467__10 ;
    input inputs_467__9 ;
    input inputs_467__8 ;
    input inputs_467__7 ;
    input inputs_467__6 ;
    input inputs_467__5 ;
    input inputs_467__4 ;
    input inputs_467__3 ;
    input inputs_467__2 ;
    input inputs_467__1 ;
    input inputs_467__0 ;
    input inputs_468__15 ;
    input inputs_468__14 ;
    input inputs_468__13 ;
    input inputs_468__12 ;
    input inputs_468__11 ;
    input inputs_468__10 ;
    input inputs_468__9 ;
    input inputs_468__8 ;
    input inputs_468__7 ;
    input inputs_468__6 ;
    input inputs_468__5 ;
    input inputs_468__4 ;
    input inputs_468__3 ;
    input inputs_468__2 ;
    input inputs_468__1 ;
    input inputs_468__0 ;
    input inputs_469__15 ;
    input inputs_469__14 ;
    input inputs_469__13 ;
    input inputs_469__12 ;
    input inputs_469__11 ;
    input inputs_469__10 ;
    input inputs_469__9 ;
    input inputs_469__8 ;
    input inputs_469__7 ;
    input inputs_469__6 ;
    input inputs_469__5 ;
    input inputs_469__4 ;
    input inputs_469__3 ;
    input inputs_469__2 ;
    input inputs_469__1 ;
    input inputs_469__0 ;
    input inputs_470__15 ;
    input inputs_470__14 ;
    input inputs_470__13 ;
    input inputs_470__12 ;
    input inputs_470__11 ;
    input inputs_470__10 ;
    input inputs_470__9 ;
    input inputs_470__8 ;
    input inputs_470__7 ;
    input inputs_470__6 ;
    input inputs_470__5 ;
    input inputs_470__4 ;
    input inputs_470__3 ;
    input inputs_470__2 ;
    input inputs_470__1 ;
    input inputs_470__0 ;
    input inputs_471__15 ;
    input inputs_471__14 ;
    input inputs_471__13 ;
    input inputs_471__12 ;
    input inputs_471__11 ;
    input inputs_471__10 ;
    input inputs_471__9 ;
    input inputs_471__8 ;
    input inputs_471__7 ;
    input inputs_471__6 ;
    input inputs_471__5 ;
    input inputs_471__4 ;
    input inputs_471__3 ;
    input inputs_471__2 ;
    input inputs_471__1 ;
    input inputs_471__0 ;
    input inputs_472__15 ;
    input inputs_472__14 ;
    input inputs_472__13 ;
    input inputs_472__12 ;
    input inputs_472__11 ;
    input inputs_472__10 ;
    input inputs_472__9 ;
    input inputs_472__8 ;
    input inputs_472__7 ;
    input inputs_472__6 ;
    input inputs_472__5 ;
    input inputs_472__4 ;
    input inputs_472__3 ;
    input inputs_472__2 ;
    input inputs_472__1 ;
    input inputs_472__0 ;
    input inputs_473__15 ;
    input inputs_473__14 ;
    input inputs_473__13 ;
    input inputs_473__12 ;
    input inputs_473__11 ;
    input inputs_473__10 ;
    input inputs_473__9 ;
    input inputs_473__8 ;
    input inputs_473__7 ;
    input inputs_473__6 ;
    input inputs_473__5 ;
    input inputs_473__4 ;
    input inputs_473__3 ;
    input inputs_473__2 ;
    input inputs_473__1 ;
    input inputs_473__0 ;
    input inputs_474__15 ;
    input inputs_474__14 ;
    input inputs_474__13 ;
    input inputs_474__12 ;
    input inputs_474__11 ;
    input inputs_474__10 ;
    input inputs_474__9 ;
    input inputs_474__8 ;
    input inputs_474__7 ;
    input inputs_474__6 ;
    input inputs_474__5 ;
    input inputs_474__4 ;
    input inputs_474__3 ;
    input inputs_474__2 ;
    input inputs_474__1 ;
    input inputs_474__0 ;
    input inputs_475__15 ;
    input inputs_475__14 ;
    input inputs_475__13 ;
    input inputs_475__12 ;
    input inputs_475__11 ;
    input inputs_475__10 ;
    input inputs_475__9 ;
    input inputs_475__8 ;
    input inputs_475__7 ;
    input inputs_475__6 ;
    input inputs_475__5 ;
    input inputs_475__4 ;
    input inputs_475__3 ;
    input inputs_475__2 ;
    input inputs_475__1 ;
    input inputs_475__0 ;
    input inputs_476__15 ;
    input inputs_476__14 ;
    input inputs_476__13 ;
    input inputs_476__12 ;
    input inputs_476__11 ;
    input inputs_476__10 ;
    input inputs_476__9 ;
    input inputs_476__8 ;
    input inputs_476__7 ;
    input inputs_476__6 ;
    input inputs_476__5 ;
    input inputs_476__4 ;
    input inputs_476__3 ;
    input inputs_476__2 ;
    input inputs_476__1 ;
    input inputs_476__0 ;
    input inputs_477__15 ;
    input inputs_477__14 ;
    input inputs_477__13 ;
    input inputs_477__12 ;
    input inputs_477__11 ;
    input inputs_477__10 ;
    input inputs_477__9 ;
    input inputs_477__8 ;
    input inputs_477__7 ;
    input inputs_477__6 ;
    input inputs_477__5 ;
    input inputs_477__4 ;
    input inputs_477__3 ;
    input inputs_477__2 ;
    input inputs_477__1 ;
    input inputs_477__0 ;
    input inputs_478__15 ;
    input inputs_478__14 ;
    input inputs_478__13 ;
    input inputs_478__12 ;
    input inputs_478__11 ;
    input inputs_478__10 ;
    input inputs_478__9 ;
    input inputs_478__8 ;
    input inputs_478__7 ;
    input inputs_478__6 ;
    input inputs_478__5 ;
    input inputs_478__4 ;
    input inputs_478__3 ;
    input inputs_478__2 ;
    input inputs_478__1 ;
    input inputs_478__0 ;
    input inputs_479__15 ;
    input inputs_479__14 ;
    input inputs_479__13 ;
    input inputs_479__12 ;
    input inputs_479__11 ;
    input inputs_479__10 ;
    input inputs_479__9 ;
    input inputs_479__8 ;
    input inputs_479__7 ;
    input inputs_479__6 ;
    input inputs_479__5 ;
    input inputs_479__4 ;
    input inputs_479__3 ;
    input inputs_479__2 ;
    input inputs_479__1 ;
    input inputs_479__0 ;
    input inputs_480__15 ;
    input inputs_480__14 ;
    input inputs_480__13 ;
    input inputs_480__12 ;
    input inputs_480__11 ;
    input inputs_480__10 ;
    input inputs_480__9 ;
    input inputs_480__8 ;
    input inputs_480__7 ;
    input inputs_480__6 ;
    input inputs_480__5 ;
    input inputs_480__4 ;
    input inputs_480__3 ;
    input inputs_480__2 ;
    input inputs_480__1 ;
    input inputs_480__0 ;
    input inputs_481__15 ;
    input inputs_481__14 ;
    input inputs_481__13 ;
    input inputs_481__12 ;
    input inputs_481__11 ;
    input inputs_481__10 ;
    input inputs_481__9 ;
    input inputs_481__8 ;
    input inputs_481__7 ;
    input inputs_481__6 ;
    input inputs_481__5 ;
    input inputs_481__4 ;
    input inputs_481__3 ;
    input inputs_481__2 ;
    input inputs_481__1 ;
    input inputs_481__0 ;
    input inputs_482__15 ;
    input inputs_482__14 ;
    input inputs_482__13 ;
    input inputs_482__12 ;
    input inputs_482__11 ;
    input inputs_482__10 ;
    input inputs_482__9 ;
    input inputs_482__8 ;
    input inputs_482__7 ;
    input inputs_482__6 ;
    input inputs_482__5 ;
    input inputs_482__4 ;
    input inputs_482__3 ;
    input inputs_482__2 ;
    input inputs_482__1 ;
    input inputs_482__0 ;
    input inputs_483__15 ;
    input inputs_483__14 ;
    input inputs_483__13 ;
    input inputs_483__12 ;
    input inputs_483__11 ;
    input inputs_483__10 ;
    input inputs_483__9 ;
    input inputs_483__8 ;
    input inputs_483__7 ;
    input inputs_483__6 ;
    input inputs_483__5 ;
    input inputs_483__4 ;
    input inputs_483__3 ;
    input inputs_483__2 ;
    input inputs_483__1 ;
    input inputs_483__0 ;
    input inputs_484__15 ;
    input inputs_484__14 ;
    input inputs_484__13 ;
    input inputs_484__12 ;
    input inputs_484__11 ;
    input inputs_484__10 ;
    input inputs_484__9 ;
    input inputs_484__8 ;
    input inputs_484__7 ;
    input inputs_484__6 ;
    input inputs_484__5 ;
    input inputs_484__4 ;
    input inputs_484__3 ;
    input inputs_484__2 ;
    input inputs_484__1 ;
    input inputs_484__0 ;
    input inputs_485__15 ;
    input inputs_485__14 ;
    input inputs_485__13 ;
    input inputs_485__12 ;
    input inputs_485__11 ;
    input inputs_485__10 ;
    input inputs_485__9 ;
    input inputs_485__8 ;
    input inputs_485__7 ;
    input inputs_485__6 ;
    input inputs_485__5 ;
    input inputs_485__4 ;
    input inputs_485__3 ;
    input inputs_485__2 ;
    input inputs_485__1 ;
    input inputs_485__0 ;
    input inputs_486__15 ;
    input inputs_486__14 ;
    input inputs_486__13 ;
    input inputs_486__12 ;
    input inputs_486__11 ;
    input inputs_486__10 ;
    input inputs_486__9 ;
    input inputs_486__8 ;
    input inputs_486__7 ;
    input inputs_486__6 ;
    input inputs_486__5 ;
    input inputs_486__4 ;
    input inputs_486__3 ;
    input inputs_486__2 ;
    input inputs_486__1 ;
    input inputs_486__0 ;
    input inputs_487__15 ;
    input inputs_487__14 ;
    input inputs_487__13 ;
    input inputs_487__12 ;
    input inputs_487__11 ;
    input inputs_487__10 ;
    input inputs_487__9 ;
    input inputs_487__8 ;
    input inputs_487__7 ;
    input inputs_487__6 ;
    input inputs_487__5 ;
    input inputs_487__4 ;
    input inputs_487__3 ;
    input inputs_487__2 ;
    input inputs_487__1 ;
    input inputs_487__0 ;
    input inputs_488__15 ;
    input inputs_488__14 ;
    input inputs_488__13 ;
    input inputs_488__12 ;
    input inputs_488__11 ;
    input inputs_488__10 ;
    input inputs_488__9 ;
    input inputs_488__8 ;
    input inputs_488__7 ;
    input inputs_488__6 ;
    input inputs_488__5 ;
    input inputs_488__4 ;
    input inputs_488__3 ;
    input inputs_488__2 ;
    input inputs_488__1 ;
    input inputs_488__0 ;
    input inputs_489__15 ;
    input inputs_489__14 ;
    input inputs_489__13 ;
    input inputs_489__12 ;
    input inputs_489__11 ;
    input inputs_489__10 ;
    input inputs_489__9 ;
    input inputs_489__8 ;
    input inputs_489__7 ;
    input inputs_489__6 ;
    input inputs_489__5 ;
    input inputs_489__4 ;
    input inputs_489__3 ;
    input inputs_489__2 ;
    input inputs_489__1 ;
    input inputs_489__0 ;
    input inputs_490__15 ;
    input inputs_490__14 ;
    input inputs_490__13 ;
    input inputs_490__12 ;
    input inputs_490__11 ;
    input inputs_490__10 ;
    input inputs_490__9 ;
    input inputs_490__8 ;
    input inputs_490__7 ;
    input inputs_490__6 ;
    input inputs_490__5 ;
    input inputs_490__4 ;
    input inputs_490__3 ;
    input inputs_490__2 ;
    input inputs_490__1 ;
    input inputs_490__0 ;
    input inputs_491__15 ;
    input inputs_491__14 ;
    input inputs_491__13 ;
    input inputs_491__12 ;
    input inputs_491__11 ;
    input inputs_491__10 ;
    input inputs_491__9 ;
    input inputs_491__8 ;
    input inputs_491__7 ;
    input inputs_491__6 ;
    input inputs_491__5 ;
    input inputs_491__4 ;
    input inputs_491__3 ;
    input inputs_491__2 ;
    input inputs_491__1 ;
    input inputs_491__0 ;
    input inputs_492__15 ;
    input inputs_492__14 ;
    input inputs_492__13 ;
    input inputs_492__12 ;
    input inputs_492__11 ;
    input inputs_492__10 ;
    input inputs_492__9 ;
    input inputs_492__8 ;
    input inputs_492__7 ;
    input inputs_492__6 ;
    input inputs_492__5 ;
    input inputs_492__4 ;
    input inputs_492__3 ;
    input inputs_492__2 ;
    input inputs_492__1 ;
    input inputs_492__0 ;
    input inputs_493__15 ;
    input inputs_493__14 ;
    input inputs_493__13 ;
    input inputs_493__12 ;
    input inputs_493__11 ;
    input inputs_493__10 ;
    input inputs_493__9 ;
    input inputs_493__8 ;
    input inputs_493__7 ;
    input inputs_493__6 ;
    input inputs_493__5 ;
    input inputs_493__4 ;
    input inputs_493__3 ;
    input inputs_493__2 ;
    input inputs_493__1 ;
    input inputs_493__0 ;
    input inputs_494__15 ;
    input inputs_494__14 ;
    input inputs_494__13 ;
    input inputs_494__12 ;
    input inputs_494__11 ;
    input inputs_494__10 ;
    input inputs_494__9 ;
    input inputs_494__8 ;
    input inputs_494__7 ;
    input inputs_494__6 ;
    input inputs_494__5 ;
    input inputs_494__4 ;
    input inputs_494__3 ;
    input inputs_494__2 ;
    input inputs_494__1 ;
    input inputs_494__0 ;
    input inputs_495__15 ;
    input inputs_495__14 ;
    input inputs_495__13 ;
    input inputs_495__12 ;
    input inputs_495__11 ;
    input inputs_495__10 ;
    input inputs_495__9 ;
    input inputs_495__8 ;
    input inputs_495__7 ;
    input inputs_495__6 ;
    input inputs_495__5 ;
    input inputs_495__4 ;
    input inputs_495__3 ;
    input inputs_495__2 ;
    input inputs_495__1 ;
    input inputs_495__0 ;
    input inputs_496__15 ;
    input inputs_496__14 ;
    input inputs_496__13 ;
    input inputs_496__12 ;
    input inputs_496__11 ;
    input inputs_496__10 ;
    input inputs_496__9 ;
    input inputs_496__8 ;
    input inputs_496__7 ;
    input inputs_496__6 ;
    input inputs_496__5 ;
    input inputs_496__4 ;
    input inputs_496__3 ;
    input inputs_496__2 ;
    input inputs_496__1 ;
    input inputs_496__0 ;
    input inputs_497__15 ;
    input inputs_497__14 ;
    input inputs_497__13 ;
    input inputs_497__12 ;
    input inputs_497__11 ;
    input inputs_497__10 ;
    input inputs_497__9 ;
    input inputs_497__8 ;
    input inputs_497__7 ;
    input inputs_497__6 ;
    input inputs_497__5 ;
    input inputs_497__4 ;
    input inputs_497__3 ;
    input inputs_497__2 ;
    input inputs_497__1 ;
    input inputs_497__0 ;
    input inputs_498__15 ;
    input inputs_498__14 ;
    input inputs_498__13 ;
    input inputs_498__12 ;
    input inputs_498__11 ;
    input inputs_498__10 ;
    input inputs_498__9 ;
    input inputs_498__8 ;
    input inputs_498__7 ;
    input inputs_498__6 ;
    input inputs_498__5 ;
    input inputs_498__4 ;
    input inputs_498__3 ;
    input inputs_498__2 ;
    input inputs_498__1 ;
    input inputs_498__0 ;
    input inputs_499__15 ;
    input inputs_499__14 ;
    input inputs_499__13 ;
    input inputs_499__12 ;
    input inputs_499__11 ;
    input inputs_499__10 ;
    input inputs_499__9 ;
    input inputs_499__8 ;
    input inputs_499__7 ;
    input inputs_499__6 ;
    input inputs_499__5 ;
    input inputs_499__4 ;
    input inputs_499__3 ;
    input inputs_499__2 ;
    input inputs_499__1 ;
    input inputs_499__0 ;
    input inputs_500__15 ;
    input inputs_500__14 ;
    input inputs_500__13 ;
    input inputs_500__12 ;
    input inputs_500__11 ;
    input inputs_500__10 ;
    input inputs_500__9 ;
    input inputs_500__8 ;
    input inputs_500__7 ;
    input inputs_500__6 ;
    input inputs_500__5 ;
    input inputs_500__4 ;
    input inputs_500__3 ;
    input inputs_500__2 ;
    input inputs_500__1 ;
    input inputs_500__0 ;
    input inputs_501__15 ;
    input inputs_501__14 ;
    input inputs_501__13 ;
    input inputs_501__12 ;
    input inputs_501__11 ;
    input inputs_501__10 ;
    input inputs_501__9 ;
    input inputs_501__8 ;
    input inputs_501__7 ;
    input inputs_501__6 ;
    input inputs_501__5 ;
    input inputs_501__4 ;
    input inputs_501__3 ;
    input inputs_501__2 ;
    input inputs_501__1 ;
    input inputs_501__0 ;
    input inputs_502__15 ;
    input inputs_502__14 ;
    input inputs_502__13 ;
    input inputs_502__12 ;
    input inputs_502__11 ;
    input inputs_502__10 ;
    input inputs_502__9 ;
    input inputs_502__8 ;
    input inputs_502__7 ;
    input inputs_502__6 ;
    input inputs_502__5 ;
    input inputs_502__4 ;
    input inputs_502__3 ;
    input inputs_502__2 ;
    input inputs_502__1 ;
    input inputs_502__0 ;
    input inputs_503__15 ;
    input inputs_503__14 ;
    input inputs_503__13 ;
    input inputs_503__12 ;
    input inputs_503__11 ;
    input inputs_503__10 ;
    input inputs_503__9 ;
    input inputs_503__8 ;
    input inputs_503__7 ;
    input inputs_503__6 ;
    input inputs_503__5 ;
    input inputs_503__4 ;
    input inputs_503__3 ;
    input inputs_503__2 ;
    input inputs_503__1 ;
    input inputs_503__0 ;
    input inputs_504__15 ;
    input inputs_504__14 ;
    input inputs_504__13 ;
    input inputs_504__12 ;
    input inputs_504__11 ;
    input inputs_504__10 ;
    input inputs_504__9 ;
    input inputs_504__8 ;
    input inputs_504__7 ;
    input inputs_504__6 ;
    input inputs_504__5 ;
    input inputs_504__4 ;
    input inputs_504__3 ;
    input inputs_504__2 ;
    input inputs_504__1 ;
    input inputs_504__0 ;
    input inputs_505__15 ;
    input inputs_505__14 ;
    input inputs_505__13 ;
    input inputs_505__12 ;
    input inputs_505__11 ;
    input inputs_505__10 ;
    input inputs_505__9 ;
    input inputs_505__8 ;
    input inputs_505__7 ;
    input inputs_505__6 ;
    input inputs_505__5 ;
    input inputs_505__4 ;
    input inputs_505__3 ;
    input inputs_505__2 ;
    input inputs_505__1 ;
    input inputs_505__0 ;
    input inputs_506__15 ;
    input inputs_506__14 ;
    input inputs_506__13 ;
    input inputs_506__12 ;
    input inputs_506__11 ;
    input inputs_506__10 ;
    input inputs_506__9 ;
    input inputs_506__8 ;
    input inputs_506__7 ;
    input inputs_506__6 ;
    input inputs_506__5 ;
    input inputs_506__4 ;
    input inputs_506__3 ;
    input inputs_506__2 ;
    input inputs_506__1 ;
    input inputs_506__0 ;
    input inputs_507__15 ;
    input inputs_507__14 ;
    input inputs_507__13 ;
    input inputs_507__12 ;
    input inputs_507__11 ;
    input inputs_507__10 ;
    input inputs_507__9 ;
    input inputs_507__8 ;
    input inputs_507__7 ;
    input inputs_507__6 ;
    input inputs_507__5 ;
    input inputs_507__4 ;
    input inputs_507__3 ;
    input inputs_507__2 ;
    input inputs_507__1 ;
    input inputs_507__0 ;
    input inputs_508__15 ;
    input inputs_508__14 ;
    input inputs_508__13 ;
    input inputs_508__12 ;
    input inputs_508__11 ;
    input inputs_508__10 ;
    input inputs_508__9 ;
    input inputs_508__8 ;
    input inputs_508__7 ;
    input inputs_508__6 ;
    input inputs_508__5 ;
    input inputs_508__4 ;
    input inputs_508__3 ;
    input inputs_508__2 ;
    input inputs_508__1 ;
    input inputs_508__0 ;
    input inputs_509__15 ;
    input inputs_509__14 ;
    input inputs_509__13 ;
    input inputs_509__12 ;
    input inputs_509__11 ;
    input inputs_509__10 ;
    input inputs_509__9 ;
    input inputs_509__8 ;
    input inputs_509__7 ;
    input inputs_509__6 ;
    input inputs_509__5 ;
    input inputs_509__4 ;
    input inputs_509__3 ;
    input inputs_509__2 ;
    input inputs_509__1 ;
    input inputs_509__0 ;
    input inputs_510__15 ;
    input inputs_510__14 ;
    input inputs_510__13 ;
    input inputs_510__12 ;
    input inputs_510__11 ;
    input inputs_510__10 ;
    input inputs_510__9 ;
    input inputs_510__8 ;
    input inputs_510__7 ;
    input inputs_510__6 ;
    input inputs_510__5 ;
    input inputs_510__4 ;
    input inputs_510__3 ;
    input inputs_510__2 ;
    input inputs_510__1 ;
    input inputs_510__0 ;
    input inputs_511__15 ;
    input inputs_511__14 ;
    input inputs_511__13 ;
    input inputs_511__12 ;
    input inputs_511__11 ;
    input inputs_511__10 ;
    input inputs_511__9 ;
    input inputs_511__8 ;
    input inputs_511__7 ;
    input inputs_511__6 ;
    input inputs_511__5 ;
    input inputs_511__4 ;
    input inputs_511__3 ;
    input inputs_511__2 ;
    input inputs_511__1 ;
    input inputs_511__0 ;
    input [8:0]selectionLines ;
    output [15:0]\output  ;

    wire nx6, nx18, nx22, nx34, nx46, nx50, nx54, nx66, nx78, nx82, nx94, nx106, 
         nx110, nx114, nx118, nx132, nx144, nx156, nx160, nx172, nx184, nx188, 
         nx196, nx202, nx214, nx226, nx230, nx242, nx254, nx258, nx262, nx274, 
         nx286, nx290, nx302, nx314, nx318, nx322, nx326, nx340, nx352, nx364, 
         nx368, nx380, nx392, nx396, nx404, nx410, nx414, nx426, nx438, nx442, 
         nx454, nx466, nx470, nx474, nx486, nx498, nx502, nx514, nx526, nx530, 
         nx534, nx538, nx552, nx564, nx576, nx580, nx592, nx604, nx608, nx616, 
         nx622, nx634, nx646, nx650, nx662, nx674, nx678, nx682, nx694, nx706, 
         nx710, nx722, nx734, nx738, nx742, nx746, nx760, nx772, nx784, nx788, 
         nx800, nx812, nx816, nx824, nx830, nx834, nx838, nx850, nx862, nx866, 
         nx878, nx890, nx894, nx898, nx910, nx922, nx926, nx938, nx950, nx954, 
         nx958, nx962, nx976, nx988, nx1000, nx1004, nx1016, nx1028, nx1032, 
         nx1040, nx1046, nx1058, nx1070, nx1074, nx1086, nx1098, nx1102, nx1106, 
         nx1118, nx1130, nx1134, nx1146, nx1158, nx1162, nx1166, nx1170, nx1184, 
         nx1196, nx1208, nx1212, nx1224, nx1236, nx1240, nx1248, nx1254, nx1258, 
         nx1270, nx1282, nx1286, nx1298, nx1310, nx1314, nx1318, nx1330, nx1342, 
         nx1346, nx1358, nx1370, nx1374, nx1378, nx1382, nx1396, nx1408, nx1420, 
         nx1424, nx1436, nx1448, nx1452, nx1460, nx1466, nx1478, nx1490, nx1494, 
         nx1506, nx1518, nx1522, nx1526, nx1538, nx1550, nx1554, nx1566, nx1578, 
         nx1582, nx1586, nx1590, nx1604, nx1616, nx1628, nx1632, nx1644, nx1656, 
         nx1660, nx1668, nx1674, nx1678, nx1682, nx1696, nx1708, nx1712, nx1724, 
         nx1736, nx1740, nx1744, nx1756, nx1768, nx1772, nx1784, nx1796, nx1800, 
         nx1804, nx1808, nx1820, nx1832, nx1836, nx1848, nx1860, nx1864, nx1868, 
         nx1880, nx1892, nx1896, nx1908, nx1920, nx1924, nx1928, nx1932, nx1936, 
         nx1950, nx1962, nx1966, nx1978, nx1990, nx1994, nx1998, nx2010, nx2022, 
         nx2026, nx2038, nx2050, nx2054, nx2058, nx2062, nx2074, nx2086, nx2090, 
         nx2102, nx2114, nx2118, nx2122, nx2134, nx2146, nx2150, nx2162, nx2174, 
         nx2178, nx2182, nx2186, nx2190, nx2202, nx2214, nx2218, nx2230, nx2242, 
         nx2246, nx2250, nx2262, nx2274, nx2278, nx2290, nx2302, nx2306, nx2310, 
         nx2314, nx2326, nx2338, nx2342, nx2354, nx2366, nx2370, nx2374, nx2386, 
         nx2398, nx2402, nx2414, nx2426, nx2430, nx2434, nx2438, nx2442, nx2452, 
         nx2468, nx2480, nx2484, nx2496, nx2508, nx2512, nx2516, nx2528, nx2540, 
         nx2544, nx2556, nx2568, nx2572, nx2576, nx2580, nx2594, nx2606, nx2618, 
         nx2622, nx2634, nx2646, nx2650, nx2658, nx2664, nx2676, nx2688, nx2692, 
         nx2704, nx2716, nx2720, nx2724, nx2736, nx2748, nx2752, nx2764, nx2776, 
         nx2780, nx2784, nx2788, nx2802, nx2814, nx2826, nx2830, nx2842, nx2854, 
         nx2858, nx2866, nx2872, nx2876, nx2888, nx2900, nx2904, nx2916, nx2928, 
         nx2932, nx2936, nx2948, nx2960, nx2964, nx2976, nx2988, nx2992, nx2996, 
         nx3000, nx3014, nx3026, nx3038, nx3042, nx3054, nx3066, nx3070, nx3078, 
         nx3084, nx3096, nx3108, nx3112, nx3124, nx3136, nx3140, nx3144, nx3156, 
         nx3168, nx3172, nx3184, nx3196, nx3200, nx3204, nx3208, nx3222, nx3234, 
         nx3246, nx3250, nx3262, nx3274, nx3278, nx3286, nx3292, nx3296, nx3300, 
         nx3312, nx3324, nx3328, nx3340, nx3352, nx3356, nx3360, nx3372, nx3384, 
         nx3388, nx3400, nx3412, nx3416, nx3420, nx3424, nx3438, nx3450, nx3462, 
         nx3466, nx3478, nx3490, nx3494, nx3502, nx3508, nx3520, nx3532, nx3536, 
         nx3548, nx3560, nx3564, nx3568, nx3580, nx3592, nx3596, nx3608, nx3620, 
         nx3624, nx3628, nx3632, nx3646, nx3658, nx3670, nx3674, nx3686, nx3698, 
         nx3702, nx3710, nx3716, nx3720, nx3732, nx3744, nx3748, nx3760, nx3772, 
         nx3776, nx3780, nx3792, nx3804, nx3808, nx3820, nx3832, nx3836, nx3840, 
         nx3844, nx3858, nx3870, nx3882, nx3886, nx3898, nx3910, nx3914, nx3922, 
         nx3928, nx3940, nx3952, nx3956, nx3968, nx3980, nx3984, nx3988, nx4000, 
         nx4012, nx4016, nx4028, nx4040, nx4044, nx4048, nx4052, nx4066, nx4078, 
         nx4090, nx4094, nx4106, nx4118, nx4122, nx4130, nx4136, nx4140, nx4144, 
         nx4148, nx4164, nx4176, nx4180, nx4192, nx4204, nx4208, nx4212, nx4224, 
         nx4236, nx4240, nx4252, nx4264, nx4268, nx4272, nx4276, nx4290, nx4302, 
         nx4314, nx4318, nx4330, nx4342, nx4346, nx4354, nx4360, nx4372, nx4384, 
         nx4388, nx4400, nx4412, nx4416, nx4420, nx4432, nx4444, nx4448, nx4460, 
         nx4472, nx4476, nx4480, nx4484, nx4498, nx4510, nx4522, nx4526, nx4538, 
         nx4550, nx4554, nx4562, nx4568, nx4572, nx4584, nx4596, nx4600, nx4612, 
         nx4624, nx4628, nx4632, nx4644, nx4656, nx4660, nx4672, nx4684, nx4688, 
         nx4692, nx4696, nx4710, nx4722, nx4734, nx4738, nx4750, nx4762, nx4766, 
         nx4774, nx4780, nx4792, nx4804, nx4808, nx4820, nx4832, nx4836, nx4840, 
         nx4852, nx4864, nx4868, nx4880, nx4892, nx4896, nx4900, nx4904, nx4918, 
         nx4930, nx4942, nx4946, nx4958, nx4970, nx4974, nx4982, nx4988, nx4992, 
         nx4996, nx5008, nx5020, nx5024, nx5036, nx5048, nx5052, nx5056, nx5068, 
         nx5080, nx5084, nx5096, nx5108, nx5112, nx5116, nx5120, nx5134, nx5146, 
         nx5158, nx5162, nx5174, nx5186, nx5190, nx5198, nx5204, nx5216, nx5228, 
         nx5232, nx5244, nx5256, nx5260, nx5264, nx5276, nx5288, nx5292, nx5304, 
         nx5316, nx5320, nx5324, nx5328, nx5342, nx5354, nx5366, nx5370, nx5382, 
         nx5394, nx5398, nx5406, nx5412, nx5416, nx5428, nx5440, nx5444, nx5456, 
         nx5468, nx5472, nx5476, nx5488, nx5500, nx5504, nx5516, nx5528, nx5532, 
         nx5536, nx5540, nx5554, nx5566, nx5578, nx5582, nx5594, nx5606, nx5610, 
         nx5618, nx5624, nx5636, nx5648, nx5652, nx5664, nx5676, nx5680, nx5684, 
         nx5696, nx5708, nx5712, nx5724, nx5736, nx5740, nx5744, nx5748, nx5762, 
         nx5774, nx5786, nx5790, nx5802, nx5814, nx5818, nx5826, nx5832, nx5836, 
         nx5840, nx5854, nx5866, nx5870, nx5882, nx5894, nx5898, nx5902, nx5914, 
         nx5926, nx5930, nx5942, nx5954, nx5958, nx5962, nx5966, nx5978, nx5990, 
         nx5994, nx6006, nx6018, nx6022, nx6026, nx6038, nx6050, nx6054, nx6066, 
         nx6078, nx6082, nx6086, nx6090, nx6094, nx6108, nx6120, nx6124, nx6136, 
         nx6148, nx6152, nx6156, nx6168, nx6180, nx6184, nx6196, nx6208, nx6212, 
         nx6216, nx6220, nx6232, nx6244, nx6248, nx6260, nx6272, nx6276, nx6280, 
         nx6292, nx6304, nx6308, nx6320, nx6332, nx6336, nx6340, nx6344, nx6348, 
         nx6360, nx6372, nx6376, nx6388, nx6400, nx6404, nx6408, nx6420, nx6432, 
         nx6436, nx6448, nx6460, nx6464, nx6468, nx6472, nx6484, nx6496, nx6500, 
         nx6512, nx6524, nx6528, nx6532, nx6544, nx6556, nx6560, nx6572, nx6584, 
         nx6588, nx6592, nx6596, nx6600, nx6610, nx6626, nx6638, nx6642, nx6654, 
         nx6666, nx6670, nx6674, nx6686, nx6698, nx6702, nx6714, nx6726, nx6730, 
         nx6734, nx6738, nx6752, nx6764, nx6776, nx6780, nx6792, nx6804, nx6808, 
         nx6816, nx6822, nx6834, nx6846, nx6850, nx6862, nx6874, nx6878, nx6882, 
         nx6894, nx6906, nx6910, nx6922, nx6934, nx6938, nx6942, nx6946, nx6960, 
         nx6972, nx6984, nx6988, nx7000, nx7012, nx7016, nx7024, nx7030, nx7034, 
         nx7046, nx7058, nx7062, nx7074, nx7086, nx7090, nx7094, nx7106, nx7118, 
         nx7122, nx7134, nx7146, nx7150, nx7154, nx7158, nx7172, nx7184, nx7196, 
         nx7200, nx7212, nx7224, nx7228, nx7236, nx7242, nx7254, nx7266, nx7270, 
         nx7282, nx7294, nx7298, nx7302, nx7314, nx7326, nx7330, nx7342, nx7354, 
         nx7358, nx7362, nx7366, nx7380, nx7392, nx7404, nx7408, nx7420, nx7432, 
         nx7436, nx7444, nx7450, nx7454, nx7458, nx7470, nx7482, nx7486, nx7498, 
         nx7510, nx7514, nx7518, nx7530, nx7542, nx7546, nx7558, nx7570, nx7574, 
         nx7578, nx7582, nx7596, nx7608, nx7620, nx7624, nx7636, nx7648, nx7652, 
         nx7660, nx7666, nx7678, nx7690, nx7694, nx7706, nx7718, nx7722, nx7726, 
         nx7738, nx7750, nx7754, nx7766, nx7778, nx7782, nx7786, nx7790, nx7804, 
         nx7816, nx7828, nx7832, nx7844, nx7856, nx7860, nx7868, nx7874, nx7878, 
         nx7890, nx7902, nx7906, nx7918, nx7930, nx7934, nx7938, nx7950, nx7962, 
         nx7966, nx7978, nx7990, nx7994, nx7998, nx8002, nx8016, nx8028, nx8040, 
         nx8044, nx8056, nx8068, nx8072, nx8080, nx8086, nx8098, nx8110, nx8114, 
         nx8126, nx8138, nx8142, nx8146, nx8158, nx8170, nx8174, nx8186, nx8198, 
         nx8202, nx8206, nx8210, nx8224, nx8236, nx8248, nx8252, nx8264, nx8276, 
         nx8280, nx8288, nx8294, nx8298, nx8302, nx8306, nx8322, nx8334, nx8338, 
         nx8350, nx8362, nx8366, nx8370, nx8382, nx8394, nx8398, nx8410, nx8422, 
         nx8426, nx8430, nx8434, nx8448, nx8460, nx8472, nx8476, nx8488, nx8500, 
         nx8504, nx8512, nx8518, nx8530, nx8542, nx8546, nx8558, nx8570, nx8574, 
         nx8578, nx8590, nx8602, nx8606, nx8618, nx8630, nx8634, nx8638, nx8642, 
         nx8656, nx8668, nx8680, nx8684, nx8696, nx8708, nx8712, nx8720, nx8726, 
         nx8730, nx8742, nx8754, nx8758, nx8770, nx8782, nx8786, nx8790, nx8802, 
         nx8814, nx8818, nx8830, nx8842, nx8846, nx8850, nx8854, nx8868, nx8880, 
         nx8892, nx8896, nx8908, nx8920, nx8924, nx8932, nx8938, nx8950, nx8962, 
         nx8966, nx8978, nx8990, nx8994, nx8998, nx9010, nx9022, nx9026, nx9038, 
         nx9050, nx9054, nx9058, nx9062, nx9076, nx9088, nx9100, nx9104, nx9116, 
         nx9128, nx9132, nx9140, nx9146, nx9150, nx9154, nx9166, nx9178, nx9182, 
         nx9194, nx9206, nx9210, nx9214, nx9226, nx9238, nx9242, nx9254, nx9266, 
         nx9270, nx9274, nx9278, nx9292, nx9304, nx9316, nx9320, nx9332, nx9344, 
         nx9348, nx9356, nx9362, nx9374, nx9386, nx9390, nx9402, nx9414, nx9418, 
         nx9422, nx9434, nx9446, nx9450, nx9462, nx9474, nx9478, nx9482, nx9486, 
         nx9500, nx9512, nx9524, nx9528, nx9540, nx9552, nx9556, nx9564, nx9570, 
         nx9574, nx9586, nx9598, nx9602, nx9614, nx9626, nx9630, nx9634, nx9646, 
         nx9658, nx9662, nx9674, nx9686, nx9690, nx9694, nx9698, nx9712, nx9724, 
         nx9736, nx9740, nx9752, nx9764, nx9768, nx9776, nx9782, nx9794, nx9806, 
         nx9810, nx9822, nx9834, nx9838, nx9842, nx9854, nx9866, nx9870, nx9882, 
         nx9894, nx9898, nx9902, nx9906, nx9920, nx9932, nx9944, nx9948, nx9960, 
         nx9972, nx9976, nx9984, nx9990, nx9994, nx9998, nx10012, nx10024, 
         nx10028, nx10040, nx10052, nx10056, nx10060, nx10072, nx10084, nx10088, 
         nx10100, nx10112, nx10116, nx10120, nx10124, nx10136, nx10148, nx10152, 
         nx10164, nx10176, nx10180, nx10184, nx10196, nx10208, nx10212, nx10224, 
         nx10236, nx10240, nx10244, nx10248, nx10252, nx10266, nx10278, nx10282, 
         nx10294, nx10306, nx10310, nx10314, nx10326, nx10338, nx10342, nx10354, 
         nx10366, nx10370, nx10374, nx10378, nx10390, nx10402, nx10406, nx10418, 
         nx10430, nx10434, nx10438, nx10450, nx10462, nx10466, nx10478, nx10490, 
         nx10494, nx10498, nx10502, nx10506, nx10518, nx10530, nx10534, nx10546, 
         nx10558, nx10562, nx10566, nx10578, nx10590, nx10594, nx10606, nx10618, 
         nx10622, nx10626, nx10630, nx10642, nx10654, nx10658, nx10670, nx10682, 
         nx10686, nx10690, nx10702, nx10714, nx10718, nx10730, nx10742, nx10746, 
         nx10750, nx10754, nx10758, nx10768, nx10784, nx10796, nx10800, nx10812, 
         nx10824, nx10828, nx10832, nx10844, nx10856, nx10860, nx10872, nx10884, 
         nx10888, nx10892, nx10896, nx10910, nx10922, nx10934, nx10938, nx10950, 
         nx10962, nx10966, nx10974, nx10980, nx10992, nx11004, nx11008, nx11020, 
         nx11032, nx11036, nx11040, nx11052, nx11064, nx11068, nx11080, nx11092, 
         nx11096, nx11100, nx11104, nx11118, nx11130, nx11142, nx11146, nx11158, 
         nx11170, nx11174, nx11182, nx11188, nx11192, nx11204, nx11216, nx11220, 
         nx11232, nx11244, nx11248, nx11252, nx11264, nx11276, nx11280, nx11292, 
         nx11304, nx11308, nx11312, nx11316, nx11330, nx11342, nx11354, nx11358, 
         nx11370, nx11382, nx11386, nx11394, nx11400, nx11412, nx11424, nx11428, 
         nx11440, nx11452, nx11456, nx11460, nx11472, nx11484, nx11488, nx11500, 
         nx11512, nx11516, nx11520, nx11524, nx11538, nx11550, nx11562, nx11566, 
         nx11578, nx11590, nx11594, nx11602, nx11608, nx11612, nx11616, nx11628, 
         nx11640, nx11644, nx11656, nx11668, nx11672, nx11676, nx11688, nx11700, 
         nx11704, nx11716, nx11728, nx11732, nx11736, nx11740, nx11754, nx11766, 
         nx11778, nx11782, nx11794, nx11806, nx11810, nx11818, nx11824, nx11836, 
         nx11848, nx11852, nx11864, nx11876, nx11880, nx11884, nx11896, nx11908, 
         nx11912, nx11924, nx11936, nx11940, nx11944, nx11948, nx11962, nx11974, 
         nx11986, nx11990, nx12002, nx12014, nx12018, nx12026, nx12032, nx12036, 
         nx12048, nx12060, nx12064, nx12076, nx12088, nx12092, nx12096, nx12108, 
         nx12120, nx12124, nx12136, nx12148, nx12152, nx12156, nx12160, nx12174, 
         nx12186, nx12198, nx12202, nx12214, nx12226, nx12230, nx12238, nx12244, 
         nx12256, nx12268, nx12272, nx12284, nx12296, nx12300, nx12304, nx12316, 
         nx12328, nx12332, nx12344, nx12356, nx12360, nx12364, nx12368, nx12382, 
         nx12394, nx12406, nx12410, nx12422, nx12434, nx12438, nx12446, nx12452, 
         nx12456, nx12460, nx12464, nx12480, nx12492, nx12496, nx12508, nx12520, 
         nx12524, nx12528, nx12540, nx12552, nx12556, nx12568, nx12580, nx12584, 
         nx12588, nx12592, nx12606, nx12618, nx12630, nx12634, nx12646, nx12658, 
         nx12662, nx12670, nx12676, nx12688, nx12700, nx12704, nx12716, nx12728, 
         nx12732, nx12736, nx12748, nx12760, nx12764, nx12776, nx12788, nx12792, 
         nx12796, nx12800, nx12814, nx12826, nx12838, nx12842, nx12854, nx12866, 
         nx12870, nx12878, nx12884, nx12888, nx12900, nx12912, nx12916, nx12928, 
         nx12940, nx12944, nx12948, nx12960, nx12972, nx12976, nx12988, nx13000, 
         nx13004, nx13008, nx13012, nx13026, nx13038, nx13050, nx13054, nx13066, 
         nx13078, nx13082, nx13090, nx13096, nx13108, nx13120, nx13124, nx13136, 
         nx13148, nx13152, nx13156, nx13168, nx13180, nx13184, nx13196, nx13208, 
         nx13212, nx13216, nx13220, nx13234, nx13246, nx13258, nx13262, nx13274, 
         nx13286, nx13290, nx13298, nx13304, nx13308, nx13312, nx13324, nx13336, 
         nx13340, nx13352, nx13364, nx13368, nx13372, nx13384, nx13396, nx13400, 
         nx13412, nx13424, nx13428, nx13432, nx13436, nx13450, nx13462, nx13474, 
         nx13478, nx13490, nx13502, nx13506, nx13514, nx13520, nx13532, nx13544, 
         nx13548, nx13560, nx13572, nx13576, nx13580, nx13592, nx13604, nx13608, 
         nx13620, nx13632, nx13636, nx13640, nx13644, nx13658, nx13670, nx13682, 
         nx13686, nx13698, nx13710, nx13714, nx13722, nx13728, nx13732, nx13744, 
         nx13756, nx13760, nx13772, nx13784, nx13788, nx13792, nx13804, nx13816, 
         nx13820, nx13832, nx13844, nx13848, nx13852, nx13856, nx13870, nx13882, 
         nx13894, nx13898, nx13910, nx13922, nx13926, nx13934, nx13940, nx13952, 
         nx13964, nx13968, nx13980, nx13992, nx13996, nx14000, nx14012, nx14024, 
         nx14028, nx14040, nx14052, nx14056, nx14060, nx14064, nx14078, nx14090, 
         nx14102, nx14106, nx14118, nx14130, nx14134, nx14142, nx14148, nx14152, 
         nx14156, nx14170, nx14182, nx14186, nx14198, nx14210, nx14214, nx14218, 
         nx14230, nx14242, nx14246, nx14258, nx14270, nx14274, nx14278, nx14282, 
         nx14294, nx14306, nx14310, nx14322, nx14334, nx14338, nx14342, nx14354, 
         nx14366, nx14370, nx14382, nx14394, nx14398, nx14402, nx14406, nx14410, 
         nx14424, nx14436, nx14440, nx14452, nx14464, nx14468, nx14472, nx14484, 
         nx14496, nx14500, nx14512, nx14524, nx14528, nx14532, nx14536, nx14548, 
         nx14560, nx14564, nx14576, nx14588, nx14592, nx14596, nx14608, nx14620, 
         nx14624, nx14636, nx14648, nx14652, nx14656, nx14660, nx14664, nx14676, 
         nx14688, nx14692, nx14704, nx14716, nx14720, nx14724, nx14736, nx14748, 
         nx14752, nx14764, nx14776, nx14780, nx14784, nx14788, nx14800, nx14812, 
         nx14816, nx14828, nx14840, nx14844, nx14848, nx14860, nx14872, nx14876, 
         nx14888, nx14900, nx14904, nx14908, nx14912, nx14916, nx14926, nx14942, 
         nx14954, nx14958, nx14970, nx14982, nx14986, nx14990, nx15002, nx15014, 
         nx15018, nx15030, nx15042, nx15046, nx15050, nx15054, nx15068, nx15080, 
         nx15092, nx15096, nx15108, nx15120, nx15124, nx15132, nx15138, nx15150, 
         nx15162, nx15166, nx15178, nx15190, nx15194, nx15198, nx15210, nx15222, 
         nx15226, nx15238, nx15250, nx15254, nx15258, nx15262, nx15276, nx15288, 
         nx15300, nx15304, nx15316, nx15328, nx15332, nx15340, nx15346, nx15350, 
         nx15362, nx15374, nx15378, nx15390, nx15402, nx15406, nx15410, nx15422, 
         nx15434, nx15438, nx15450, nx15462, nx15466, nx15470, nx15474, nx15488, 
         nx15500, nx15512, nx15516, nx15528, nx15540, nx15544, nx15552, nx15558, 
         nx15570, nx15582, nx15586, nx15598, nx15610, nx15614, nx15618, nx15630, 
         nx15642, nx15646, nx15658, nx15670, nx15674, nx15678, nx15682, nx15696, 
         nx15708, nx15720, nx15724, nx15736, nx15748, nx15752, nx15760, nx15766, 
         nx15770, nx15774, nx15786, nx15798, nx15802, nx15814, nx15826, nx15830, 
         nx15834, nx15846, nx15858, nx15862, nx15874, nx15886, nx15890, nx15894, 
         nx15898, nx15912, nx15924, nx15936, nx15940, nx15952, nx15964, nx15968, 
         nx15976, nx15982, nx15994, nx16006, nx16010, nx16022, nx16034, nx16038, 
         nx16042, nx16054, nx16066, nx16070, nx16082, nx16094, nx16098, nx16102, 
         nx16106, nx16120, nx16132, nx16144, nx16148, nx16160, nx16172, nx16176, 
         nx16184, nx16190, nx16194, nx16206, nx16218, nx16222, nx16234, nx16246, 
         nx16250, nx16254, nx16266, nx16278, nx16282, nx16294, nx16306, nx16310, 
         nx16314, nx16318, nx16332, nx16344, nx16356, nx16360, nx16372, nx16384, 
         nx16388, nx16396, nx16402, nx16414, nx16426, nx16430, nx16442, nx16454, 
         nx16458, nx16462, nx16474, nx16486, nx16490, nx16502, nx16514, nx16518, 
         nx16522, nx16526, nx16540, nx16552, nx16564, nx16568, nx16580, nx16592, 
         nx16596, nx16604, nx16610, nx16614, nx16618, nx16622, nx16638, nx16650, 
         nx16654, nx16666, nx16678, nx16682, nx16686, nx16698, nx16710, nx16714, 
         nx16726, nx16738, nx16742, nx16746, nx16750, nx16764, nx16776, nx16788, 
         nx16792, nx16804, nx16816, nx16820, nx16828, nx16834, nx16846, nx16858, 
         nx16862, nx16874, nx16886, nx16890, nx16894, nx16906, nx16918, nx16922, 
         nx16934, nx16946, nx16950, nx16954, nx16958, nx16972, nx16984, nx16996, 
         nx17000, nx17012, nx17024, nx17028, nx17036, nx17042, nx17046, nx17058, 
         nx17070, nx17074, nx17086, nx17098, nx17102, nx17106, nx17118, nx17130, 
         nx17134, nx17146, nx17158, nx17162, nx17166, nx17170, nx17184, nx17196, 
         nx17208, nx17212, nx17224, nx17236, nx17240, nx17248, nx17254, nx17266, 
         nx17278, nx17282, nx17294, nx17306, nx17310, nx17314, nx17326, nx17338, 
         nx17342, nx17354, nx17366, nx17370, nx17374, nx17378, nx17392, nx17404, 
         nx17416, nx17420, nx17432, nx17444, nx17448, nx17456, nx17462, nx17466, 
         nx17470, nx17482, nx17494, nx17498, nx17510, nx17522, nx17526, nx17530, 
         nx17542, nx17554, nx17558, nx17570, nx17582, nx17586, nx17590, nx17594, 
         nx17608, nx17620, nx17632, nx17636, nx17648, nx17660, nx17664, nx17672, 
         nx17678, nx17690, nx17702, nx17706, nx17718, nx17730, nx17734, nx17738, 
         nx17750, nx17762, nx17766, nx17778, nx17790, nx17794, nx17798, nx17802, 
         nx17816, nx17828, nx17840, nx17844, nx17856, nx17868, nx17872, nx17880, 
         nx17886, nx17890, nx17902, nx17914, nx17918, nx17930, nx17942, nx17946, 
         nx17950, nx17962, nx17974, nx17978, nx17990, nx18002, nx18006, nx18010, 
         nx18014, nx18028, nx18040, nx18052, nx18056, nx18068, nx18080, nx18084, 
         nx18092, nx18098, nx18110, nx18122, nx18126, nx18138, nx18150, nx18154, 
         nx18158, nx18170, nx18182, nx18186, nx18198, nx18210, nx18214, nx18218, 
         nx18222, nx18236, nx18248, nx18260, nx18264, nx18276, nx18288, nx18292, 
         nx18300, nx18306, nx18310, nx18314, nx18328, nx18340, nx18344, nx18356, 
         nx18368, nx18372, nx18376, nx18388, nx18400, nx18404, nx18416, nx18428, 
         nx18432, nx18436, nx18440, nx18452, nx18464, nx18468, nx18480, nx18492, 
         nx18496, nx18500, nx18512, nx18524, nx18528, nx18540, nx18552, nx18556, 
         nx18560, nx18564, nx18568, nx18582, nx18594, nx18598, nx18610, nx18622, 
         nx18626, nx18630, nx18642, nx18654, nx18658, nx18670, nx18682, nx18686, 
         nx18690, nx18694, nx18706, nx18718, nx18722, nx18734, nx18746, nx18750, 
         nx18754, nx18766, nx18778, nx18782, nx18794, nx18806, nx18810, nx18814, 
         nx18818, nx18822, nx18834, nx18846, nx18850, nx18862, nx18874, nx18878, 
         nx18882, nx18894, nx18906, nx18910, nx18922, nx18934, nx18938, nx18942, 
         nx18946, nx18958, nx18970, nx18974, nx18986, nx18998, nx19002, nx19006, 
         nx19018, nx19030, nx19034, nx19046, nx19058, nx19062, nx19066, nx19070, 
         nx19074, nx19084, nx19100, nx19112, nx19116, nx19128, nx19140, nx19144, 
         nx19148, nx19160, nx19172, nx19176, nx19188, nx19200, nx19204, nx19208, 
         nx19212, nx19226, nx19238, nx19250, nx19254, nx19266, nx19278, nx19282, 
         nx19290, nx19296, nx19308, nx19320, nx19324, nx19336, nx19348, nx19352, 
         nx19356, nx19368, nx19380, nx19384, nx19396, nx19408, nx19412, nx19416, 
         nx19420, nx19434, nx19446, nx19458, nx19462, nx19474, nx19486, nx19490, 
         nx19498, nx19504, nx19508, nx19520, nx19532, nx19536, nx19548, nx19560, 
         nx19564, nx19568, nx19580, nx19592, nx19596, nx19608, nx19620, nx19624, 
         nx19628, nx19632, nx19646, nx19658, nx19670, nx19674, nx19686, nx19698, 
         nx19702, nx19710, nx19716, nx19728, nx19740, nx19744, nx19756, nx19768, 
         nx19772, nx19776, nx19788, nx19800, nx19804, nx19816, nx19828, nx19832, 
         nx19836, nx19840, nx19854, nx19866, nx19878, nx19882, nx19894, nx19906, 
         nx19910, nx19918, nx19924, nx19928, nx19932, nx19944, nx19956, nx19960, 
         nx19972, nx19984, nx19988, nx19992, nx20004, nx20016, nx20020, nx20032, 
         nx20044, nx20048, nx20052, nx20056, nx20070, nx20082, nx20094, nx20098, 
         nx20110, nx20122, nx20126, nx20134, nx20140, nx20152, nx20164, nx20168, 
         nx20180, nx20192, nx20196, nx20200, nx20212, nx20224, nx20228, nx20240, 
         nx20252, nx20256, nx20260, nx20264, nx20278, nx20290, nx20302, nx20306, 
         nx20318, nx20330, nx20334, nx20342, nx20348, nx20352, nx20364, nx20376, 
         nx20380, nx20392, nx20404, nx20408, nx20412, nx20424, nx20436, nx20440, 
         nx20452, nx20464, nx20468, nx20472, nx20476, nx20490, nx20502, nx20514, 
         nx20518, nx20530, nx20542, nx20546, nx20554, nx20560, nx20572, nx20584, 
         nx20588, nx20600, nx20612, nx20616, nx20620, nx20632, nx20644, nx20648, 
         nx20660, nx20672, nx20676, nx20680, nx20684, nx20698, nx20710, nx20722, 
         nx20726, nx20738, nx20750, nx20754, nx20762, nx20768, nx20772, nx20776, 
         nx20780, nx20796, nx20808, nx20812, nx20824, nx20836, nx20840, nx20844, 
         nx20856, nx20868, nx20872, nx20884, nx20896, nx20900, nx20904, nx20908, 
         nx20922, nx20934, nx20946, nx20950, nx20962, nx20974, nx20978, nx20986, 
         nx20992, nx21004, nx21016, nx21020, nx21032, nx21044, nx21048, nx21052, 
         nx21064, nx21076, nx21080, nx21092, nx21104, nx21108, nx21112, nx21116, 
         nx21130, nx21142, nx21154, nx21158, nx21170, nx21182, nx21186, nx21194, 
         nx21200, nx21204, nx21216, nx21228, nx21232, nx21244, nx21256, nx21260, 
         nx21264, nx21276, nx21288, nx21292, nx21304, nx21316, nx21320, nx21324, 
         nx21328, nx21342, nx21354, nx21366, nx21370, nx21382, nx21394, nx21398, 
         nx21406, nx21412, nx21424, nx21436, nx21440, nx21452, nx21464, nx21468, 
         nx21472, nx21484, nx21496, nx21500, nx21512, nx21524, nx21528, nx21532, 
         nx21536, nx21550, nx21562, nx21574, nx21578, nx21590, nx21602, nx21606, 
         nx21614, nx21620, nx21624, nx21628, nx21640, nx21652, nx21656, nx21668, 
         nx21680, nx21684, nx21688, nx21700, nx21712, nx21716, nx21728, nx21740, 
         nx21744, nx21748, nx21752, nx21766, nx21778, nx21790, nx21794, nx21806, 
         nx21818, nx21822, nx21830, nx21836, nx21848, nx21860, nx21864, nx21876, 
         nx21888, nx21892, nx21896, nx21908, nx21920, nx21924, nx21936, nx21948, 
         nx21952, nx21956, nx21960, nx21974, nx21986, nx21998, nx22002, nx22014, 
         nx22026, nx22030, nx22038, nx22044, nx22048, nx22060, nx22072, nx22076, 
         nx22088, nx22100, nx22104, nx22108, nx22120, nx22132, nx22136, nx22148, 
         nx22160, nx22164, nx22168, nx22172, nx22186, nx22198, nx22210, nx22214, 
         nx22226, nx22238, nx22242, nx22250, nx22256, nx22268, nx22280, nx22284, 
         nx22296, nx22308, nx22312, nx22316, nx22328, nx22340, nx22344, nx22356, 
         nx22368, nx22372, nx22376, nx22380, nx22394, nx22406, nx22418, nx22422, 
         nx22434, nx22446, nx22450, nx22458, nx22464, nx22468, nx22472, nx22486, 
         nx22498, nx22502, nx22514, nx22526, nx22530, nx22534, nx22546, nx22558, 
         nx22562, nx22574, nx22586, nx22590, nx22594, nx22598, nx22610, nx22622, 
         nx22626, nx22638, nx22650, nx22654, nx22658, nx22670, nx22682, nx22686, 
         nx22698, nx22710, nx22714, nx22718, nx22722, nx22726, nx22740, nx22752, 
         nx22756, nx22768, nx22780, nx22784, nx22788, nx22800, nx22812, nx22816, 
         nx22828, nx22840, nx22844, nx22848, nx22852, nx22864, nx22876, nx22880, 
         nx22892, nx22904, nx22908, nx22912, nx22924, nx22936, nx22940, nx22952, 
         nx22964, nx22968, nx22972, nx22976, nx22980, nx22992, nx23004, nx23008, 
         nx23020, nx23032, nx23036, nx23040, nx23052, nx23064, nx23068, nx23080, 
         nx23092, nx23096, nx23100, nx23104, nx23116, nx23128, nx23132, nx23144, 
         nx23156, nx23160, nx23164, nx23176, nx23188, nx23192, nx23204, nx23216, 
         nx23220, nx23224, nx23228, nx23232, nx23242, nx23258, nx23270, nx23274, 
         nx23286, nx23298, nx23302, nx23306, nx23318, nx23330, nx23334, nx23346, 
         nx23358, nx23362, nx23366, nx23370, nx23384, nx23396, nx23408, nx23412, 
         nx23424, nx23436, nx23440, nx23448, nx23454, nx23466, nx23478, nx23482, 
         nx23494, nx23506, nx23510, nx23514, nx23526, nx23538, nx23542, nx23554, 
         nx23566, nx23570, nx23574, nx23578, nx23592, nx23604, nx23616, nx23620, 
         nx23632, nx23644, nx23648, nx23656, nx23662, nx23666, nx23678, nx23690, 
         nx23694, nx23706, nx23718, nx23722, nx23726, nx23738, nx23750, nx23754, 
         nx23766, nx23778, nx23782, nx23786, nx23790, nx23804, nx23816, nx23828, 
         nx23832, nx23844, nx23856, nx23860, nx23868, nx23874, nx23886, nx23898, 
         nx23902, nx23914, nx23926, nx23930, nx23934, nx23946, nx23958, nx23962, 
         nx23974, nx23986, nx23990, nx23994, nx23998, nx24012, nx24024, nx24036, 
         nx24040, nx24052, nx24064, nx24068, nx24076, nx24082, nx24086, nx24090, 
         nx24102, nx24114, nx24118, nx24130, nx24142, nx24146, nx24150, nx24162, 
         nx24174, nx24178, nx24190, nx24202, nx24206, nx24210, nx24214, nx24228, 
         nx24240, nx24252, nx24256, nx24268, nx24280, nx24284, nx24292, nx24298, 
         nx24310, nx24322, nx24326, nx24338, nx24350, nx24354, nx24358, nx24370, 
         nx24382, nx24386, nx24398, nx24410, nx24414, nx24418, nx24422, nx24436, 
         nx24448, nx24460, nx24464, nx24476, nx24488, nx24492, nx24500, nx24506, 
         nx24510, nx24522, nx24534, nx24538, nx24550, nx24562, nx24566, nx24570, 
         nx24582, nx24594, nx24598, nx24610, nx24622, nx24626, nx24630, nx24634, 
         nx24648, nx24660, nx24672, nx24676, nx24688, nx24700, nx24704, nx24712, 
         nx24718, nx24730, nx24742, nx24746, nx24758, nx24770, nx24774, nx24778, 
         nx24790, nx24802, nx24806, nx24818, nx24830, nx24834, nx24838, nx24842, 
         nx24856, nx24868, nx24880, nx24884, nx24896, nx24908, nx24912, nx24920, 
         nx24926, nx24930, nx24934, nx24938, nx24954, nx24966, nx24970, nx24982, 
         nx24994, nx24998, nx25002, nx25014, nx25026, nx25030, nx25042, nx25054, 
         nx25058, nx25062, nx25066, nx25080, nx25092, nx25104, nx25108, nx25120, 
         nx25132, nx25136, nx25144, nx25150, nx25162, nx25174, nx25178, nx25190, 
         nx25202, nx25206, nx25210, nx25222, nx25234, nx25238, nx25250, nx25262, 
         nx25266, nx25270, nx25274, nx25288, nx25300, nx25312, nx25316, nx25328, 
         nx25340, nx25344, nx25352, nx25358, nx25362, nx25374, nx25386, nx25390, 
         nx25402, nx25414, nx25418, nx25422, nx25434, nx25446, nx25450, nx25462, 
         nx25474, nx25478, nx25482, nx25486, nx25500, nx25512, nx25524, nx25528, 
         nx25540, nx25552, nx25556, nx25564, nx25570, nx25582, nx25594, nx25598, 
         nx25610, nx25622, nx25626, nx25630, nx25642, nx25654, nx25658, nx25670, 
         nx25682, nx25686, nx25690, nx25694, nx25708, nx25720, nx25732, nx25736, 
         nx25748, nx25760, nx25764, nx25772, nx25778, nx25782, nx25786, nx25798, 
         nx25810, nx25814, nx25826, nx25838, nx25842, nx25846, nx25858, nx25870, 
         nx25874, nx25886, nx25898, nx25902, nx25906, nx25910, nx25924, nx25936, 
         nx25948, nx25952, nx25964, nx25976, nx25980, nx25988, nx25994, nx26006, 
         nx26018, nx26022, nx26034, nx26046, nx26050, nx26054, nx26066, nx26078, 
         nx26082, nx26094, nx26106, nx26110, nx26114, nx26118, nx26132, nx26144, 
         nx26156, nx26160, nx26172, nx26184, nx26188, nx26196, nx26202, nx26206, 
         nx26218, nx26230, nx26234, nx26246, nx26258, nx26262, nx26266, nx26278, 
         nx26290, nx26294, nx26306, nx26318, nx26322, nx26326, nx26330, nx26344, 
         nx26356, nx26368, nx26372, nx26384, nx26396, nx26400, nx26408, nx26414, 
         nx26426, nx26438, nx26442, nx26454, nx26466, nx26470, nx26474, nx26486, 
         nx26498, nx26502, nx26514, nx26526, nx26530, nx26534, nx26538, nx26552, 
         nx26564, nx26576, nx26580, nx26592, nx26604, nx26608, nx26616, nx26622, 
         nx26626, nx26630, nx26644, nx26656, nx26660, nx26672, nx26684, nx26688, 
         nx26692, nx26704, nx26716, nx26720, nx26732, nx26744, nx26748, nx26752, 
         nx26756, nx26768, nx26780, nx26784, nx26796, nx26808, nx26812, nx26816, 
         nx26828, nx26840, nx26844, nx26856, nx26868, nx26872, nx26876, nx26880, 
         nx26884, nx26898, nx26910, nx26914, nx26926, nx26938, nx26942, nx26946, 
         nx26958, nx26970, nx26974, nx26986, nx26998, nx27002, nx27006, nx27010, 
         nx27022, nx27034, nx27038, nx27050, nx27062, nx27066, nx27070, nx27082, 
         nx27094, nx27098, nx27110, nx27122, nx27126, nx27130, nx27134, nx27138, 
         nx27150, nx27162, nx27166, nx27178, nx27190, nx27194, nx27198, nx27210, 
         nx27222, nx27226, nx27238, nx27250, nx27254, nx27258, nx27262, nx27274, 
         nx27286, nx27290, nx27302, nx27314, nx27318, nx27322, nx27334, nx27346, 
         nx27350, nx27362, nx27374, nx27378, nx27382, nx27386, nx27390, nx27400, 
         nx27416, nx27428, nx27432, nx27444, nx27456, nx27460, nx27464, nx27476, 
         nx27488, nx27492, nx27504, nx27516, nx27520, nx27524, nx27528, nx27542, 
         nx27554, nx27566, nx27570, nx27582, nx27594, nx27598, nx27606, nx27612, 
         nx27624, nx27636, nx27640, nx27652, nx27664, nx27668, nx27672, nx27684, 
         nx27696, nx27700, nx27712, nx27724, nx27728, nx27732, nx27736, nx27750, 
         nx27762, nx27774, nx27778, nx27790, nx27802, nx27806, nx27814, nx27820, 
         nx27824, nx27836, nx27848, nx27852, nx27864, nx27876, nx27880, nx27884, 
         nx27896, nx27908, nx27912, nx27924, nx27936, nx27940, nx27944, nx27948, 
         nx27962, nx27974, nx27986, nx27990, nx28002, nx28014, nx28018, nx28026, 
         nx28032, nx28044, nx28056, nx28060, nx28072, nx28084, nx28088, nx28092, 
         nx28104, nx28116, nx28120, nx28132, nx28144, nx28148, nx28152, nx28156, 
         nx28170, nx28182, nx28194, nx28198, nx28210, nx28222, nx28226, nx28234, 
         nx28240, nx28244, nx28248, nx28260, nx28272, nx28276, nx28288, nx28300, 
         nx28304, nx28308, nx28320, nx28332, nx28336, nx28348, nx28360, nx28364, 
         nx28368, nx28372, nx28386, nx28398, nx28410, nx28414, nx28426, nx28438, 
         nx28442, nx28450, nx28456, nx28468, nx28480, nx28484, nx28496, nx28508, 
         nx28512, nx28516, nx28528, nx28540, nx28544, nx28556, nx28568, nx28572, 
         nx28576, nx28580, nx28594, nx28606, nx28618, nx28622, nx28634, nx28646, 
         nx28650, nx28658, nx28664, nx28668, nx28680, nx28692, nx28696, nx28708, 
         nx28720, nx28724, nx28728, nx28740, nx28752, nx28756, nx28768, nx28780, 
         nx28784, nx28788, nx28792, nx28806, nx28818, nx28830, nx28834, nx28846, 
         nx28858, nx28862, nx28870, nx28876, nx28888, nx28900, nx28904, nx28916, 
         nx28928, nx28932, nx28936, nx28948, nx28960, nx28964, nx28976, nx28988, 
         nx28992, nx28996, nx29000, nx29014, nx29026, nx29038, nx29042, nx29054, 
         nx29066, nx29070, nx29078, nx29084, nx29088, nx29092, nx29096, nx29112, 
         nx29124, nx29128, nx29140, nx29152, nx29156, nx29160, nx29172, nx29184, 
         nx29188, nx29200, nx29212, nx29216, nx29220, nx29224, nx29238, nx29250, 
         nx29262, nx29266, nx29278, nx29290, nx29294, nx29302, nx29308, nx29320, 
         nx29332, nx29336, nx29348, nx29360, nx29364, nx29368, nx29380, nx29392, 
         nx29396, nx29408, nx29420, nx29424, nx29428, nx29432, nx29446, nx29458, 
         nx29470, nx29474, nx29486, nx29498, nx29502, nx29510, nx29516, nx29520, 
         nx29532, nx29544, nx29548, nx29560, nx29572, nx29576, nx29580, nx29592, 
         nx29604, nx29608, nx29620, nx29632, nx29636, nx29640, nx29644, nx29658, 
         nx29670, nx29682, nx29686, nx29698, nx29710, nx29714, nx29722, nx29728, 
         nx29740, nx29752, nx29756, nx29768, nx29780, nx29784, nx29788, nx29800, 
         nx29812, nx29816, nx29828, nx29840, nx29844, nx29848, nx29852, nx29866, 
         nx29878, nx29890, nx29894, nx29906, nx29918, nx29922, nx29930, nx29936, 
         nx29940, nx29944, nx29956, nx29968, nx29972, nx29984, nx29996, nx30000, 
         nx30004, nx30016, nx30028, nx30032, nx30044, nx30056, nx30060, nx30064, 
         nx30068, nx30082, nx30094, nx30106, nx30110, nx30122, nx30134, nx30138, 
         nx30146, nx30152, nx30164, nx30176, nx30180, nx30192, nx30204, nx30208, 
         nx30212, nx30224, nx30236, nx30240, nx30252, nx30264, nx30268, nx30272, 
         nx30276, nx30290, nx30302, nx30314, nx30318, nx30330, nx30342, nx30346, 
         nx30354, nx30360, nx30364, nx30376, nx30388, nx30392, nx30404, nx30416, 
         nx30420, nx30424, nx30436, nx30448, nx30452, nx30464, nx30476, nx30480, 
         nx30484, nx30488, nx30502, nx30514, nx30526, nx30530, nx30542, nx30554, 
         nx30558, nx30566, nx30572, nx30584, nx30596, nx30600, nx30612, nx30624, 
         nx30628, nx30632, nx30644, nx30656, nx30660, nx30672, nx30684, nx30688, 
         nx30692, nx30696, nx30710, nx30722, nx30734, nx30738, nx30750, nx30762, 
         nx30766, nx30774, nx30780, nx30784, nx30788, nx30802, nx30814, nx30818, 
         nx30830, nx30842, nx30846, nx30850, nx30862, nx30874, nx30878, nx30890, 
         nx30902, nx30906, nx30910, nx30914, nx30926, nx30938, nx30942, nx30954, 
         nx30966, nx30970, nx30974, nx30986, nx30998, nx31002, nx31014, nx31026, 
         nx31030, nx31034, nx31038, nx31042, nx31056, nx31068, nx31072, nx31084, 
         nx31096, nx31100, nx31104, nx31116, nx31128, nx31132, nx31144, nx31156, 
         nx31160, nx31164, nx31168, nx31180, nx31192, nx31196, nx31208, nx31220, 
         nx31224, nx31228, nx31240, nx31252, nx31256, nx31268, nx31280, nx31284, 
         nx31288, nx31292, nx31296, nx31308, nx31320, nx31324, nx31336, nx31348, 
         nx31352, nx31356, nx31368, nx31380, nx31384, nx31396, nx31408, nx31412, 
         nx31416, nx31420, nx31432, nx31444, nx31448, nx31460, nx31472, nx31476, 
         nx31480, nx31492, nx31504, nx31508, nx31520, nx31532, nx31536, nx31540, 
         nx31544, nx31548, nx31558, nx31574, nx31586, nx31590, nx31602, nx31614, 
         nx31618, nx31622, nx31634, nx31646, nx31650, nx31662, nx31674, nx31678, 
         nx31682, nx31686, nx31700, nx31712, nx31724, nx31728, nx31740, nx31752, 
         nx31756, nx31764, nx31770, nx31782, nx31794, nx31798, nx31810, nx31822, 
         nx31826, nx31830, nx31842, nx31854, nx31858, nx31870, nx31882, nx31886, 
         nx31890, nx31894, nx31908, nx31920, nx31932, nx31936, nx31948, nx31960, 
         nx31964, nx31972, nx31978, nx31982, nx31994, nx32006, nx32010, nx32022, 
         nx32034, nx32038, nx32042, nx32054, nx32066, nx32070, nx32082, nx32094, 
         nx32098, nx32102, nx32106, nx32120, nx32132, nx32144, nx32148, nx32160, 
         nx32172, nx32176, nx32184, nx32190, nx32202, nx32214, nx32218, nx32230, 
         nx32242, nx32246, nx32250, nx32262, nx32274, nx32278, nx32290, nx32302, 
         nx32306, nx32310, nx32314, nx32328, nx32340, nx32352, nx32356, nx32368, 
         nx32380, nx32384, nx32392, nx32398, nx32402, nx32406, nx32418, nx32430, 
         nx32434, nx32446, nx32458, nx32462, nx32466, nx32478, nx32490, nx32494, 
         nx32506, nx32518, nx32522, nx32526, nx32530, nx32544, nx32556, nx32568, 
         nx32572, nx32584, nx32596, nx32600, nx32608, nx32614, nx32626, nx32638, 
         nx32642, nx32654, nx32666, nx32670, nx32674, nx32686, nx32698, nx32702, 
         nx32714, nx32726, nx32730, nx32734, nx32738, nx32752, nx32764, nx32776, 
         nx32780, nx32792, nx32804, nx32808, nx32816, nx32822, nx32826, nx32838, 
         nx32850, nx32854, nx32866, nx32878, nx32882, nx32886, nx32898, nx32910, 
         nx32914, nx32926, nx32938, nx32942, nx32946, nx32950, nx32964, nx32976, 
         nx32988, nx32992, nx33004, nx33016, nx33020, nx33028, nx33034, nx33046, 
         nx33058, nx33062, nx33074, nx33086, nx33090, nx33094, nx33106, nx33118, 
         nx33122, nx33134, nx33146, nx33150, nx33154, nx33158, nx33172, nx33184, 
         nx33196, nx33200, nx33212, nx33224, nx33228, nx33236, nx33242, nx33246, 
         nx33250, nx33254, nx33270, nx33282, nx33286, nx33298, nx33310, nx33314, 
         nx33318, nx33330, nx33342, nx33346, nx33358, nx33370, nx33374, nx33378, 
         nx33382, nx33396, nx33408, nx33420, nx33424, nx33436, nx33448, nx33452, 
         nx33460, nx33466, nx33478, nx33490, nx33494, nx33506, nx33518, nx33522, 
         nx33526, nx33538, nx33550, nx33554, nx33566, nx33578, nx33582, nx33586, 
         nx33590, nx33604, nx33616, nx33628, nx33632, nx33644, nx33656, nx33660, 
         nx33668, nx33674, nx33678, nx33690, nx33702, nx33706, nx33718, nx33730, 
         nx33734, nx33738, nx33750, nx33762, nx33766, nx33778, nx33790, nx33794, 
         nx33798, nx33802, nx33816, nx33828, nx33840, nx33844, nx33856, nx33868, 
         nx33872, nx33880, nx33886, nx33898, nx33910, nx33914, nx33926, nx33938, 
         nx33942, nx33946, nx33958, nx33970, nx33974, nx33986, nx33998, nx34002, 
         nx34006, nx34010, nx34024, nx34036, nx34048, nx34052, nx34064, nx34076, 
         nx34080, nx34088, nx34094, nx34098, nx34102, nx34114, nx34126, nx34130, 
         nx34142, nx34154, nx34158, nx34162, nx34174, nx34186, nx34190, nx34202, 
         nx34214, nx34218, nx34222, nx34226, nx34240, nx34252, nx34264, nx34268, 
         nx34280, nx34292, nx34296, nx34304, nx34310, nx34322, nx34334, nx34338, 
         nx34350, nx34362, nx34366, nx34370, nx34382, nx34394, nx34398, nx34410, 
         nx34422, nx34426, nx34430, nx34434, nx34448, nx34460, nx34472, nx34476, 
         nx34488, nx34500, nx34504, nx34512, nx34518, nx34522, nx34534, nx34546, 
         nx34550, nx34562, nx34574, nx34578, nx34582, nx34594, nx34606, nx34610, 
         nx34622, nx34634, nx34638, nx34642, nx34646, nx34660, nx34672, nx34684, 
         nx34688, nx34700, nx34712, nx34716, nx34724, nx34730, nx34742, nx34754, 
         nx34758, nx34770, nx34782, nx34786, nx34790, nx34802, nx34814, nx34818, 
         nx34830, nx34842, nx34846, nx34850, nx34854, nx34868, nx34880, nx34892, 
         nx34896, nx34908, nx34920, nx34924, nx34932, nx34938, nx34942, nx34946, 
         nx34960, nx34972, nx34976, nx34988, nx35000, nx35004, nx35008, nx35020, 
         nx35032, nx35036, nx35048, nx35060, nx35064, nx35068, nx35072, nx35084, 
         nx35096, nx35100, nx35112, nx35124, nx35128, nx35132, nx35144, nx35156, 
         nx35160, nx35172, nx35184, nx35188, nx35192, nx35196, nx35200, nx35214, 
         nx35226, nx35230, nx35242, nx35254, nx35258, nx35262, nx35274, nx35286, 
         nx35290, nx35302, nx35314, nx35318, nx35322, nx35326, nx35338, nx35350, 
         nx35354, nx35366, nx35378, nx35382, nx35386, nx35398, nx35410, nx35414, 
         nx35426, nx35438, nx35442, nx35446, nx35450, nx35454, nx35466, nx35478, 
         nx35482, nx35494, nx35506, nx35510, nx35514, nx35526, nx35538, nx35542, 
         nx35554, nx35566, nx35570, nx35574, nx35578, nx35590, nx35602, nx35606, 
         nx35618, nx35630, nx35634, nx35638, nx35650, nx35662, nx35666, nx35678, 
         nx35690, nx35694, nx35698, nx35702, nx35706, nx35716, nx35732, nx35744, 
         nx35748, nx35760, nx35772, nx35776, nx35780, nx35792, nx35804, nx35808, 
         nx35820, nx35832, nx35836, nx35840, nx35844, nx35858, nx35870, nx35882, 
         nx35886, nx35898, nx35910, nx35914, nx35922, nx35928, nx35940, nx35952, 
         nx35956, nx35968, nx35980, nx35984, nx35988, nx36000, nx36012, nx36016, 
         nx36028, nx36040, nx36044, nx36048, nx36052, nx36066, nx36078, nx36090, 
         nx36094, nx36106, nx36118, nx36122, nx36130, nx36136, nx36140, nx36152, 
         nx36164, nx36168, nx36180, nx36192, nx36196, nx36200, nx36212, nx36224, 
         nx36228, nx36240, nx36252, nx36256, nx36260, nx36264, nx36278, nx36290, 
         nx36302, nx36306, nx36318, nx36330, nx36334, nx36342, nx36348, nx36360, 
         nx36372, nx36376, nx36388, nx36400, nx36404, nx36408, nx36420, nx36432, 
         nx36436, nx36448, nx36460, nx36464, nx36468, nx36472, nx36486, nx36498, 
         nx36510, nx36514, nx36526, nx36538, nx36542, nx36550, nx36556, nx36560, 
         nx36564, nx36576, nx36588, nx36592, nx36604, nx36616, nx36620, nx36624, 
         nx36636, nx36648, nx36652, nx36664, nx36676, nx36680, nx36684, nx36688, 
         nx36702, nx36714, nx36726, nx36730, nx36742, nx36754, nx36758, nx36766, 
         nx36772, nx36784, nx36796, nx36800, nx36812, nx36824, nx36828, nx36832, 
         nx36844, nx36856, nx36860, nx36872, nx36884, nx36888, nx36892, nx36896, 
         nx36910, nx36922, nx36934, nx36938, nx36950, nx36962, nx36966, nx36974, 
         nx36980, nx36984, nx36996, nx37008, nx37012, nx37024, nx37036, nx37040, 
         nx37044, nx37056, nx37068, nx37072, nx37084, nx37096, nx37100, nx37104, 
         nx37108, nx37122, nx37134, nx37146, nx37150, nx37162, nx37174, nx37178, 
         nx37186, nx37192, nx37204, nx37216, nx37220, nx37232, nx37244, nx37248, 
         nx37252, nx37264, nx37276, nx37280, nx37292, nx37304, nx37308, nx37312, 
         nx37316, nx37330, nx37342, nx37354, nx37358, nx37370, nx37382, nx37386, 
         nx37394, nx37400, nx37404, nx37408, nx37412, nx37428, nx37440, nx37444, 
         nx37456, nx37468, nx37472, nx37476, nx37488, nx37500, nx37504, nx37516, 
         nx37528, nx37532, nx37536, nx37540, nx37554, nx37566, nx37578, nx37582, 
         nx37594, nx37606, nx37610, nx37618, nx37624, nx37636, nx37648, nx37652, 
         nx37664, nx37676, nx37680, nx37684, nx37696, nx37708, nx37712, nx37724, 
         nx37736, nx37740, nx37744, nx37748, nx37762, nx37774, nx37786, nx37790, 
         nx37802, nx37814, nx37818, nx37826, nx37832, nx37836, nx37848, nx37860, 
         nx37864, nx37876, nx37888, nx37892, nx37896, nx37908, nx37920, nx37924, 
         nx37936, nx37948, nx37952, nx37956, nx37960, nx37974, nx37986, nx37998, 
         nx38002, nx38014, nx38026, nx38030, nx38038, nx38044, nx38056, nx38068, 
         nx38072, nx38084, nx38096, nx38100, nx38104, nx38116, nx38128, nx38132, 
         nx38144, nx38156, nx38160, nx38164, nx38168, nx38182, nx38194, nx38206, 
         nx38210, nx38222, nx38234, nx38238, nx38246, nx38252, nx38256, nx38260, 
         nx38272, nx38284, nx38288, nx38300, nx38312, nx38316, nx38320, nx38332, 
         nx38344, nx38348, nx38360, nx38372, nx38376, nx38380, nx38384, nx38398, 
         nx38410, nx38422, nx38426, nx38438, nx38450, nx38454, nx38462, nx38468, 
         nx38480, nx38492, nx38496, nx38508, nx38520, nx38524, nx38528, nx38540, 
         nx38552, nx38556, nx38568, nx38580, nx38584, nx38588, nx38592, nx38606, 
         nx38618, nx38630, nx38634, nx38646, nx38658, nx38662, nx38670, nx38676, 
         nx38680, nx38692, nx38704, nx38708, nx38720, nx38732, nx38736, nx38740, 
         nx38752, nx38764, nx38768, nx38780, nx38792, nx38796, nx38800, nx38804, 
         nx38818, nx38830, nx38842, nx38846, nx38858, nx38870, nx38874, nx38882, 
         nx38888, nx38900, nx38912, nx38916, nx38928, nx38940, nx38944, nx38948, 
         nx38960, nx38972, nx38976, nx38988, nx39000, nx39004, nx39008, nx39012, 
         nx39026, nx39038, nx39050, nx39054, nx39066, nx39078, nx39082, nx39090, 
         nx39096, nx39100, nx39104, nx39118, nx39130, nx39134, nx39146, nx39158, 
         nx39162, nx39166, nx39178, nx39190, nx39194, nx39206, nx39218, nx39222, 
         nx39226, nx39230, nx39242, nx39254, nx39258, nx39270, nx39282, nx39286, 
         nx39290, nx39302, nx39314, nx39318, nx39330, nx39342, nx39346, nx39350, 
         nx39354, nx39358, nx39372, nx39384, nx39388, nx39400, nx39412, nx39416, 
         nx39420, nx39432, nx39444, nx39448, nx39460, nx39472, nx39476, nx39480, 
         nx39484, nx39496, nx39508, nx39512, nx39524, nx39536, nx39540, nx39544, 
         nx39556, nx39568, nx39572, nx39584, nx39596, nx39600, nx39604, nx39608, 
         nx39612, nx39624, nx39636, nx39640, nx39652, nx39664, nx39668, nx39672, 
         nx39684, nx39696, nx39700, nx39712, nx39724, nx39728, nx39732, nx39736, 
         nx39748, nx39760, nx39764, nx39776, nx39788, nx39792, nx39796, nx39808, 
         nx39820, nx39824, nx39836, nx39848, nx39852, nx39856, nx39860, nx39864, 
         nx39874, nx39890, nx39902, nx39906, nx39918, nx39930, nx39934, nx39938, 
         nx39950, nx39962, nx39966, nx39978, nx39990, nx39994, nx39998, nx40002, 
         nx40016, nx40028, nx40040, nx40044, nx40056, nx40068, nx40072, nx40080, 
         nx40086, nx40098, nx40110, nx40114, nx40126, nx40138, nx40142, nx40146, 
         nx40158, nx40170, nx40174, nx40186, nx40198, nx40202, nx40206, nx40210, 
         nx40224, nx40236, nx40248, nx40252, nx40264, nx40276, nx40280, nx40288, 
         nx40294, nx40298, nx40310, nx40322, nx40326, nx40338, nx40350, nx40354, 
         nx40358, nx40370, nx40382, nx40386, nx40398, nx40410, nx40414, nx40418, 
         nx40422, nx40436, nx40448, nx40460, nx40464, nx40476, nx40488, nx40492, 
         nx40500, nx40506, nx40518, nx40530, nx40534, nx40546, nx40558, nx40562, 
         nx40566, nx40578, nx40590, nx40594, nx40606, nx40618, nx40622, nx40626, 
         nx40630, nx40644, nx40656, nx40668, nx40672, nx40684, nx40696, nx40700, 
         nx40708, nx40714, nx40718, nx40722, nx40734, nx40746, nx40750, nx40762, 
         nx40774, nx40778, nx40782, nx40794, nx40806, nx40810, nx40822, nx40834, 
         nx40838, nx40842, nx40846, nx40860, nx40872, nx40884, nx40888, nx40900, 
         nx40912, nx40916, nx40924, nx40930, nx40942, nx40954, nx40958, nx40970, 
         nx40982, nx40986, nx40990, nx41002, nx41014, nx41018, nx41030, nx41042, 
         nx41046, nx41050, nx41054, nx41068, nx41080, nx41092, nx41096, nx41108, 
         nx41120, nx41124, nx41132, nx41138, nx41142, nx41154, nx41166, nx41170, 
         nx41182, nx41194, nx41198, nx41202, nx41214, nx41226, nx41230, nx41242, 
         nx41254, nx41258, nx41262, nx41266, nx41280, nx41292, nx41304, nx41308, 
         nx41320, nx41332, nx41336, nx41344, nx41350, nx41362, nx41374, nx41378, 
         nx41390, nx41402, nx41406, nx41410, nx41422, nx41434, nx41438, nx41450, 
         nx41462, nx41466, nx41470, nx41474, nx41488, nx41500, nx41512, nx41516, 
         nx41528, nx41540, nx41544, nx41552, nx41558, nx41562, nx41566, nx41570, 
         nx41586, nx41598, nx41602, nx41614, nx41626, nx41630, nx41634, nx41646, 
         nx41658, nx41662, nx41674, nx41686, nx41690, nx41694, nx41698, nx41712, 
         nx41724, nx41736, nx41740, nx41752, nx41764, nx41768, nx41776, nx41782, 
         nx41794, nx41806, nx41810, nx41822, nx41834, nx41838, nx41842, nx41854, 
         nx41866, nx41870, nx41882, nx41894, nx41898, nx41902, nx41906, nx41920, 
         nx41932, nx41944, nx41948, nx41960, nx41972, nx41976, nx41984, nx41990, 
         nx41994, nx42006, nx42018, nx42022, nx42034, nx42046, nx42050, nx42054, 
         nx42066, nx42078, nx42082, nx42094, nx42106, nx42110, nx42114, nx42118, 
         nx42132, nx42144, nx42156, nx42160, nx42172, nx42184, nx42188, nx42196, 
         nx42202, nx42214, nx42226, nx42230, nx42242, nx42254, nx42258, nx42262, 
         nx42274, nx42286, nx42290, nx42302, nx42314, nx42318, nx42322, nx42326, 
         nx42340, nx42352, nx42364, nx42368, nx42380, nx42392, nx42396, nx42404, 
         nx42410, nx42414, nx42418, nx42430, nx42442, nx42446, nx42458, nx42470, 
         nx42474, nx42478, nx42490, nx42502, nx42506, nx42518, nx42530, nx42534, 
         nx42538, nx42542, nx42556, nx42568, nx42580, nx42584, nx42596, nx42608, 
         nx42612, nx42620, nx42626, nx42638, nx42650, nx42654, nx42666, nx42678, 
         nx42682, nx42686, nx42698, nx42710, nx42714, nx42726, nx42738, nx42742, 
         nx42746, nx42750, nx42764, nx42776, nx42788, nx42792, nx42804, nx42816, 
         nx42820, nx42828, nx42834, nx42838, nx42850, nx42862, nx42866, nx42878, 
         nx42890, nx42894, nx42898, nx42910, nx42922, nx42926, nx42938, nx42950, 
         nx42954, nx42958, nx42962, nx42976, nx42988, nx43000, nx43004, nx43016, 
         nx43028, nx43032, nx43040, nx43046, nx43058, nx43070, nx43074, nx43086, 
         nx43098, nx43102, nx43106, nx43118, nx43130, nx43134, nx43146, nx43158, 
         nx43162, nx43166, nx43170, nx43184, nx43196, nx43208, nx43212, nx43224, 
         nx43236, nx43240, nx43248, nx43254, nx43258, nx43262, nx43276, nx43288, 
         nx43292, nx43304, nx43316, nx43320, nx43324, nx43336, nx43348, nx43352, 
         nx43364, nx43376, nx43380, nx43384, nx43388, nx43400, nx43412, nx43416, 
         nx43428, nx43440, nx43444, nx43448, nx43460, nx43472, nx43476, nx43488, 
         nx43500, nx43504, nx43508, nx43512, nx43516, nx43530, nx43542, nx43546, 
         nx43558, nx43570, nx43574, nx43578, nx43590, nx43602, nx43606, nx43618, 
         nx43630, nx43634, nx43638, nx43642, nx43654, nx43666, nx43670, nx43682, 
         nx43694, nx43698, nx43702, nx43714, nx43726, nx43730, nx43742, nx43754, 
         nx43758, nx43762, nx43766, nx43770, nx43782, nx43794, nx43798, nx43810, 
         nx43822, nx43826, nx43830, nx43842, nx43854, nx43858, nx43870, nx43882, 
         nx43886, nx43890, nx43894, nx43906, nx43918, nx43922, nx43934, nx43946, 
         nx43950, nx43954, nx43966, nx43978, nx43982, nx43994, nx44006, nx44010, 
         nx44014, nx44018, nx44022, nx44032, nx44048, nx44060, nx44064, nx44076, 
         nx44088, nx44092, nx44096, nx44108, nx44120, nx44124, nx44136, nx44148, 
         nx44152, nx44156, nx44160, nx44174, nx44186, nx44198, nx44202, nx44214, 
         nx44226, nx44230, nx44238, nx44244, nx44256, nx44268, nx44272, nx44284, 
         nx44296, nx44300, nx44304, nx44316, nx44328, nx44332, nx44344, nx44356, 
         nx44360, nx44364, nx44368, nx44382, nx44394, nx44406, nx44410, nx44422, 
         nx44434, nx44438, nx44446, nx44452, nx44456, nx44468, nx44480, nx44484, 
         nx44496, nx44508, nx44512, nx44516, nx44528, nx44540, nx44544, nx44556, 
         nx44568, nx44572, nx44576, nx44580, nx44594, nx44606, nx44618, nx44622, 
         nx44634, nx44646, nx44650, nx44658, nx44664, nx44676, nx44688, nx44692, 
         nx44704, nx44716, nx44720, nx44724, nx44736, nx44748, nx44752, nx44764, 
         nx44776, nx44780, nx44784, nx44788, nx44802, nx44814, nx44826, nx44830, 
         nx44842, nx44854, nx44858, nx44866, nx44872, nx44876, nx44880, nx44892, 
         nx44904, nx44908, nx44920, nx44932, nx44936, nx44940, nx44952, nx44964, 
         nx44968, nx44980, nx44992, nx44996, nx45000, nx45004, nx45018, nx45030, 
         nx45042, nx45046, nx45058, nx45070, nx45074, nx45082, nx45088, nx45100, 
         nx45112, nx45116, nx45128, nx45140, nx45144, nx45148, nx45160, nx45172, 
         nx45176, nx45188, nx45200, nx45204, nx45208, nx45212, nx45226, nx45238, 
         nx45250, nx45254, nx45266, nx45278, nx45282, nx45290, nx45296, nx45300, 
         nx45312, nx45324, nx45328, nx45340, nx45352, nx45356, nx45360, nx45372, 
         nx45384, nx45388, nx45400, nx45412, nx45416, nx45420, nx45424, nx45438, 
         nx45450, nx45462, nx45466, nx45478, nx45490, nx45494, nx45502, nx45508, 
         nx45520, nx45532, nx45536, nx45548, nx45560, nx45564, nx45568, nx45580, 
         nx45592, nx45596, nx45608, nx45620, nx45624, nx45628, nx45632, nx45646, 
         nx45658, nx45670, nx45674, nx45686, nx45698, nx45702, nx45710, nx45716, 
         nx45720, nx45724, nx45728, nx45744, nx45756, nx45760, nx45772, nx45784, 
         nx45788, nx45792, nx45804, nx45816, nx45820, nx45832, nx45844, nx45848, 
         nx45852, nx45856, nx45870, nx45882, nx45894, nx45898, nx45910, nx45922, 
         nx45926, nx45934, nx45940, nx45952, nx45964, nx45968, nx45980, nx45992, 
         nx45996, nx46000, nx46012, nx46024, nx46028, nx46040, nx46052, nx46056, 
         nx46060, nx46064, nx46078, nx46090, nx46102, nx46106, nx46118, nx46130, 
         nx46134, nx46142, nx46148, nx46152, nx46164, nx46176, nx46180, nx46192, 
         nx46204, nx46208, nx46212, nx46224, nx46236, nx46240, nx46252, nx46264, 
         nx46268, nx46272, nx46276, nx46290, nx46302, nx46314, nx46318, nx46330, 
         nx46342, nx46346, nx46354, nx46360, nx46372, nx46384, nx46388, nx46400, 
         nx46412, nx46416, nx46420, nx46432, nx46444, nx46448, nx46460, nx46472, 
         nx46476, nx46480, nx46484, nx46498, nx46510, nx46522, nx46526, nx46538, 
         nx46550, nx46554, nx46562, nx46568, nx46572, nx46576, nx46588, nx46600, 
         nx46604, nx46616, nx46628, nx46632, nx46636, nx46648, nx46660, nx46664, 
         nx46676, nx46688, nx46692, nx46696, nx46700, nx46714, nx46726, nx46738, 
         nx46742, nx46754, nx46766, nx46770, nx46778, nx46784, nx46796, nx46808, 
         nx46812, nx46824, nx46836, nx46840, nx46844, nx46856, nx46868, nx46872, 
         nx46884, nx46896, nx46900, nx46904, nx46908, nx46922, nx46934, nx46946, 
         nx46950, nx46962, nx46974, nx46978, nx46986, nx46992, nx46996, nx47008, 
         nx47020, nx47024, nx47036, nx47048, nx47052, nx47056, nx47068, nx47080, 
         nx47084, nx47096, nx47108, nx47112, nx47116, nx47120, nx47134, nx47146, 
         nx47158, nx47162, nx47174, nx47186, nx47190, nx47198, nx47204, nx47216, 
         nx47228, nx47232, nx47244, nx47256, nx47260, nx47264, nx47276, nx47288, 
         nx47292, nx47304, nx47316, nx47320, nx47324, nx47328, nx47342, nx47354, 
         nx47366, nx47370, nx47382, nx47394, nx47398, nx47406, nx47412, nx47416, 
         nx47420, nx47434, nx47446, nx47450, nx47462, nx47474, nx47478, nx47482, 
         nx47494, nx47506, nx47510, nx47522, nx47534, nx47538, nx47542, nx47546, 
         nx47558, nx47570, nx47574, nx47586, nx47598, nx47602, nx47606, nx47618, 
         nx47630, nx47634, nx47646, nx47658, nx47662, nx47666, nx47670, nx47674, 
         nx47688, nx47700, nx47704, nx47716, nx47728, nx47732, nx47736, nx47748, 
         nx47760, nx47764, nx47776, nx47788, nx47792, nx47796, nx47800, nx47812, 
         nx47824, nx47828, nx47840, nx47852, nx47856, nx47860, nx47872, nx47884, 
         nx47888, nx47900, nx47912, nx47916, nx47920, nx47924, nx47928, nx47940, 
         nx47952, nx47956, nx47968, nx47980, nx47984, nx47988, nx48000, nx48012, 
         nx48016, nx48028, nx48040, nx48044, nx48048, nx48052, nx48064, nx48076, 
         nx48080, nx48092, nx48104, nx48108, nx48112, nx48124, nx48136, nx48140, 
         nx48152, nx48164, nx48168, nx48172, nx48176, nx48180, nx48190, nx48206, 
         nx48218, nx48222, nx48234, nx48246, nx48250, nx48254, nx48266, nx48278, 
         nx48282, nx48294, nx48306, nx48310, nx48314, nx48318, nx48332, nx48344, 
         nx48356, nx48360, nx48372, nx48384, nx48388, nx48396, nx48402, nx48414, 
         nx48426, nx48430, nx48442, nx48454, nx48458, nx48462, nx48474, nx48486, 
         nx48490, nx48502, nx48514, nx48518, nx48522, nx48526, nx48540, nx48552, 
         nx48564, nx48568, nx48580, nx48592, nx48596, nx48604, nx48610, nx48614, 
         nx48626, nx48638, nx48642, nx48654, nx48666, nx48670, nx48674, nx48686, 
         nx48698, nx48702, nx48714, nx48726, nx48730, nx48734, nx48738, nx48752, 
         nx48764, nx48776, nx48780, nx48792, nx48804, nx48808, nx48816, nx48822, 
         nx48834, nx48846, nx48850, nx48862, nx48874, nx48878, nx48882, nx48894, 
         nx48906, nx48910, nx48922, nx48934, nx48938, nx48942, nx48946, nx48960, 
         nx48972, nx48984, nx48988, nx49000, nx49012, nx49016, nx49024, nx49030, 
         nx49034, nx49038, nx49050, nx49062, nx49066, nx49078, nx49090, nx49094, 
         nx49098, nx49110, nx49122, nx49126, nx49138, nx49150, nx49154, nx49158, 
         nx49162, nx49176, nx49188, nx49200, nx49204, nx49216, nx49228, nx49232, 
         nx49240, nx49246, nx49258, nx49270, nx49274, nx49286, nx49298, nx49302, 
         nx49306, nx49318, nx49330, nx49334, nx49346, nx49358, nx49362, nx49366, 
         nx49370, nx49384, nx49396, nx49408, nx49412, nx49424, nx49436, nx49440, 
         nx49448, nx49454, nx49458, nx49470, nx49482, nx49486, nx49498, nx49510, 
         nx49514, nx49518, nx49530, nx49542, nx49546, nx49558, nx49570, nx49574, 
         nx49578, nx49582, nx49596, nx49608, nx49620, nx49624, nx49636, nx49648, 
         nx49652, nx49660, nx49666, nx49678, nx49690, nx49694, nx49706, nx49718, 
         nx49722, nx49726, nx49738, nx49750, nx49754, nx49766, nx49778, nx49782, 
         nx49786, nx49790, nx49804, nx49816, nx49828, nx49832, nx49844, nx49856, 
         nx49860, nx49868, nx49874, nx49878, nx49882, nx49886, nx49902, nx49914, 
         nx49918, nx49930, nx49942, nx49946, nx49950, nx49962, nx49974, nx49978, 
         nx49990, nx50002, nx50006, nx50010, nx50014, nx50028, nx50040, nx50052, 
         nx50056, nx50068, nx50080, nx50084, nx50092, nx50098, nx50110, nx50122, 
         nx50126, nx50138, nx50150, nx50154, nx50158, nx50170, nx50182, nx50186, 
         nx50198, nx50210, nx50214, nx50218, nx50222, nx50236, nx50248, nx50260, 
         nx50264, nx50276, nx50288, nx50292, nx50300, nx50306, nx50310, nx50322, 
         nx50334, nx50338, nx50350, nx50362, nx50366, nx50370, nx50382, nx50394, 
         nx50398, nx50410, nx50422, nx50426, nx50430, nx50434, nx50448, nx50460, 
         nx50472, nx50476, nx50488, nx50500, nx50504, nx50512, nx50518, nx50530, 
         nx50542, nx50546, nx50558, nx50570, nx50574, nx50578, nx50590, nx50602, 
         nx50606, nx50618, nx50630, nx50634, nx50638, nx50642, nx50656, nx50668, 
         nx50680, nx50684, nx50696, nx50708, nx50712, nx50720, nx50726, nx50730, 
         nx50734, nx50746, nx50758, nx50762, nx50774, nx50786, nx50790, nx50794, 
         nx50806, nx50818, nx50822, nx50834, nx50846, nx50850, nx50854, nx50858, 
         nx50872, nx50884, nx50896, nx50900, nx50912, nx50924, nx50928, nx50936, 
         nx50942, nx50954, nx50966, nx50970, nx50982, nx50994, nx50998, nx51002, 
         nx51014, nx51026, nx51030, nx51042, nx51054, nx51058, nx51062, nx51066, 
         nx51080, nx51092, nx51104, nx51108, nx51120, nx51132, nx51136, nx51144, 
         nx51150, nx51154, nx51166, nx51178, nx51182, nx51194, nx51206, nx51210, 
         nx51214, nx51226, nx51238, nx51242, nx51254, nx51266, nx51270, nx51274, 
         nx51278, nx51292, nx51304, nx51316, nx51320, nx51332, nx51344, nx51348, 
         nx51356, nx51362, nx51374, nx51386, nx51390, nx51402, nx51414, nx51418, 
         nx51422, nx51434, nx51446, nx51450, nx51462, nx51474, nx51478, nx51482, 
         nx51486, nx51500, nx51512, nx51524, nx51528, nx51540, nx51552, nx51556, 
         nx51564, nx51570, nx51574, nx51578, nx51592, nx51604, nx51608, nx51620, 
         nx51632, nx51636, nx51640, nx51652, nx51664, nx51668, nx51680, nx51692, 
         nx51696, nx51700, nx51704, nx51716, nx51728, nx51732, nx51744, nx51756, 
         nx51760, nx51764, nx51776, nx51788, nx51792, nx51804, nx51816, nx51820, 
         nx51824, nx51828, nx51832, nx51846, nx51858, nx51862, nx51874, nx51886, 
         nx51890, nx51894, nx51906, nx51918, nx51922, nx51934, nx51946, nx51950, 
         nx51954, nx51958, nx51970, nx51982, nx51986, nx51998, nx52010, nx52014, 
         nx52018, nx52030, nx52042, nx52046, nx52058, nx52070, nx52074, nx52078, 
         nx52082, nx52086, nx52098, nx52110, nx52114, nx52126, nx52138, nx52142, 
         nx52146, nx52158, nx52170, nx52174, nx52186, nx52198, nx52202, nx52206, 
         nx52210, nx52222, nx52234, nx52238, nx52250, nx52262, nx52266, nx52270, 
         nx52282, nx52294, nx52298, nx52310, nx52322, nx52326, nx52330, nx52334, 
         nx52338, nx52348, nx52364, nx52376, nx52380, nx52392, nx52404, nx52408, 
         nx52412, nx52424, nx52436, nx52440, nx52452, nx52464, nx52468, nx52472, 
         nx52476, nx52490, nx52502, nx52514, nx52518, nx52530, nx52542, nx52546, 
         nx52554, nx52560, nx52572, nx52584, nx52588, nx52600, nx52612, nx52616, 
         nx52620, nx52632, nx52644, nx52648, nx52660, nx52672, nx52676, nx52680, 
         nx52684, nx52698, nx52710, nx52722, nx52726, nx52738, nx52750, nx52754, 
         nx52762, nx52768, nx52772, nx52784, nx52796, nx52800, nx52812, nx52824, 
         nx52828, nx52832, nx52844, nx52856, nx52860, nx52872, nx52884, nx52888, 
         nx52892, nx52896, nx52910, nx52922, nx52934, nx52938, nx52950, nx52962, 
         nx52966, nx52974, nx52980, nx52992, nx53004, nx53008, nx53020, nx53032, 
         nx53036, nx53040, nx53052, nx53064, nx53068, nx53080, nx53092, nx53096, 
         nx53100, nx53104, nx53118, nx53130, nx53142, nx53146, nx53158, nx53170, 
         nx53174, nx53182, nx53188, nx53192, nx53196, nx53208, nx53220, nx53224, 
         nx53236, nx53248, nx53252, nx53256, nx53268, nx53280, nx53284, nx53296, 
         nx53308, nx53312, nx53316, nx53320, nx53334, nx53346, nx53358, nx53362, 
         nx53374, nx53386, nx53390, nx53398, nx53404, nx53416, nx53428, nx53432, 
         nx53444, nx53456, nx53460, nx53464, nx53476, nx53488, nx53492, nx53504, 
         nx53516, nx53520, nx53524, nx53528, nx53542, nx53554, nx53566, nx53570, 
         nx53582, nx53594, nx53598, nx53606, nx53612, nx53616, nx53628, nx53640, 
         nx53644, nx53656, nx53668, nx53672, nx53676, nx53688, nx53700, nx53704, 
         nx53716, nx53728, nx53732, nx53736, nx53740, nx53754, nx53766, nx53778, 
         nx53782, nx53794, nx53806, nx53810, nx53818, nx53824, nx53836, nx53848, 
         nx53852, nx53864, nx53876, nx53880, nx53884, nx53896, nx53908, nx53912, 
         nx53924, nx53936, nx53940, nx53944, nx53948, nx53962, nx53974, nx53986, 
         nx53990, nx54002, nx54014, nx54018, nx54026, nx54032, nx54036, nx54040, 
         nx54044, nx54060, nx54072, nx54076, nx54088, nx54100, nx54104, nx54108, 
         nx54120, nx54132, nx54136, nx54148, nx54160, nx54164, nx54168, nx54172, 
         nx54186, nx54198, nx54210, nx54214, nx54226, nx54238, nx54242, nx54250, 
         nx54256, nx54268, nx54280, nx54284, nx54296, nx54308, nx54312, nx54316, 
         nx54328, nx54340, nx54344, nx54356, nx54368, nx54372, nx54376, nx54380, 
         nx54394, nx54406, nx54418, nx54422, nx54434, nx54446, nx54450, nx54458, 
         nx54464, nx54468, nx54480, nx54492, nx54496, nx54508, nx54520, nx54524, 
         nx54528, nx54540, nx54552, nx54556, nx54568, nx54580, nx54584, nx54588, 
         nx54592, nx54606, nx54618, nx54630, nx54634, nx54646, nx54658, nx54662, 
         nx54670, nx54676, nx54688, nx54700, nx54704, nx54716, nx54728, nx54732, 
         nx54736, nx54748, nx54760, nx54764, nx54776, nx54788, nx54792, nx54796, 
         nx54800, nx54814, nx54826, nx54838, nx54842, nx54854, nx54866, nx54870, 
         nx54878, nx54884, nx54888, nx54892, nx54904, nx54916, nx54920, nx54932, 
         nx54944, nx54948, nx54952, nx54964, nx54976, nx54980, nx54992, nx55004, 
         nx55008, nx55012, nx55016, nx55030, nx55042, nx55054, nx55058, nx55070, 
         nx55082, nx55086, nx55094, nx55100, nx55112, nx55124, nx55128, nx55140, 
         nx55152, nx55156, nx55160, nx55172, nx55184, nx55188, nx55200, nx55212, 
         nx55216, nx55220, nx55224, nx55238, nx55250, nx55262, nx55266, nx55278, 
         nx55290, nx55294, nx55302, nx55308, nx55312, nx55324, nx55336, nx55340, 
         nx55352, nx55364, nx55368, nx55372, nx55384, nx55396, nx55400, nx55412, 
         nx55424, nx55428, nx55432, nx55436, nx55450, nx55462, nx55474, nx55478, 
         nx55490, nx55502, nx55506, nx55514, nx55520, nx55532, nx55544, nx55548, 
         nx55560, nx55572, nx55576, nx55580, nx55592, nx55604, nx55608, nx55620, 
         nx55632, nx55636, nx55640, nx55644, nx55658, nx55670, nx55682, nx55686, 
         nx55698, nx55710, nx55714, nx55722, nx55728, nx55732, nx55736, nx55750, 
         nx55762, nx55766, nx55778, nx55790, nx55794, nx55798, nx55810, nx55822, 
         nx55826, nx55838, nx55850, nx55854, nx55858, nx55862, nx55874, nx55886, 
         nx55890, nx55902, nx55914, nx55918, nx55922, nx55934, nx55946, nx55950, 
         nx55962, nx55974, nx55978, nx55982, nx55986, nx55990, nx56004, nx56016, 
         nx56020, nx56032, nx56044, nx56048, nx56052, nx56064, nx56076, nx56080, 
         nx56092, nx56104, nx56108, nx56112, nx56116, nx56128, nx56140, nx56144, 
         nx56156, nx56168, nx56172, nx56176, nx56188, nx56200, nx56204, nx56216, 
         nx56228, nx56232, nx56236, nx56240, nx56244, nx56256, nx56268, nx56272, 
         nx56284, nx56296, nx56300, nx56304, nx56316, nx56328, nx56332, nx56344, 
         nx56356, nx56360, nx56364, nx56368, nx56380, nx56392, nx56396, nx56408, 
         nx56420, nx56424, nx56428, nx56440, nx56452, nx56456, nx56468, nx56480, 
         nx56484, nx56488, nx56492, nx56496, nx56506, nx56522, nx56534, nx56538, 
         nx56550, nx56562, nx56566, nx56570, nx56582, nx56594, nx56598, nx56610, 
         nx56622, nx56626, nx56630, nx56634, nx56648, nx56660, nx56672, nx56676, 
         nx56688, nx56700, nx56704, nx56712, nx56718, nx56730, nx56742, nx56746, 
         nx56758, nx56770, nx56774, nx56778, nx56790, nx56802, nx56806, nx56818, 
         nx56830, nx56834, nx56838, nx56842, nx56856, nx56868, nx56880, nx56884, 
         nx56896, nx56908, nx56912, nx56920, nx56926, nx56930, nx56942, nx56954, 
         nx56958, nx56970, nx56982, nx56986, nx56990, nx57002, nx57014, nx57018, 
         nx57030, nx57042, nx57046, nx57050, nx57054, nx57068, nx57080, nx57092, 
         nx57096, nx57108, nx57120, nx57124, nx57132, nx57138, nx57150, nx57162, 
         nx57166, nx57178, nx57190, nx57194, nx57198, nx57210, nx57222, nx57226, 
         nx57238, nx57250, nx57254, nx57258, nx57262, nx57276, nx57288, nx57300, 
         nx57304, nx57316, nx57328, nx57332, nx57340, nx57346, nx57350, nx57354, 
         nx57366, nx57378, nx57382, nx57394, nx57406, nx57410, nx57414, nx57426, 
         nx57438, nx57442, nx57454, nx57466, nx57470, nx57474, nx57478, nx57492, 
         nx57504, nx57516, nx57520, nx57532, nx57544, nx57548, nx57556, nx57562, 
         nx57574, nx57586, nx57590, nx57602, nx57614, nx57618, nx57622, nx57634, 
         nx57646, nx57650, nx57662, nx57674, nx57678, nx57682, nx57686, nx57700, 
         nx57712, nx57724, nx57728, nx57740, nx57752, nx57756, nx57764, nx57770, 
         nx57774, nx57786, nx57798, nx57802, nx57814, nx57826, nx57830, nx57834, 
         nx57846, nx57858, nx57862, nx57874, nx57886, nx57890, nx57894, nx57898, 
         nx57912, nx57924, nx57936, nx57940, nx57952, nx57964, nx57968, nx57976, 
         nx57982, nx57994, nx58006, nx58010, nx58022, nx58034, nx58038, nx58042, 
         nx58054, nx58066, nx58070, nx58082, nx58094, nx58098, nx58102, nx58106, 
         nx58120, nx58132, nx58144, nx58148, nx58160, nx58172, nx58176, nx58184, 
         nx58190, nx58194, nx58198, nx58202, nx58218, nx58230, nx58234, nx58246, 
         nx58258, nx58262, nx58266, nx58278, nx58290, nx58294, nx58306, nx58318, 
         nx58322, nx58326, nx58330, nx58344, nx58356, nx58368, nx58372, nx58384, 
         nx58396, nx58400, nx58408, nx58414, nx58426, nx58438, nx58442, nx58454, 
         nx58466, nx58470, nx58474, nx58486, nx58498, nx58502, nx58514, nx58526, 
         nx58530, nx58534, nx58538, nx58552, nx58564, nx58576, nx58580, nx58592, 
         nx58604, nx58608, nx58616, nx58622, nx58626, nx58638, nx58650, nx58654, 
         nx58666, nx58678, nx58682, nx58686, nx58698, nx58710, nx58714, nx58726, 
         nx58738, nx58742, nx58746, nx58750, nx58764, nx58776, nx58788, nx58792, 
         nx58804, nx58816, nx58820, nx58828, nx58834, nx58846, nx58858, nx58862, 
         nx58874, nx58886, nx58890, nx58894, nx58906, nx58918, nx58922, nx58934, 
         nx58946, nx58950, nx58954, nx58958, nx58972, nx58984, nx58996, nx59000, 
         nx59012, nx59024, nx59028, nx59036, nx59042, nx59046, nx59050, nx59062, 
         nx59074, nx59078, nx59090, nx59102, nx59106, nx59110, nx59122, nx59134, 
         nx59138, nx59150, nx59162, nx59166, nx59170, nx59174, nx59188, nx59200, 
         nx59212, nx59216, nx59228, nx59240, nx59244, nx59252, nx59258, nx59270, 
         nx59282, nx59286, nx59298, nx59310, nx59314, nx59318, nx59330, nx59342, 
         nx59346, nx59358, nx59370, nx59374, nx59378, nx59382, nx59396, nx59408, 
         nx59420, nx59424, nx59436, nx59448, nx59452, nx59460, nx59466, nx59470, 
         nx59482, nx59494, nx59498, nx59510, nx59522, nx59526, nx59530, nx59542, 
         nx59554, nx59558, nx59570, nx59582, nx59586, nx59590, nx59594, nx59608, 
         nx59620, nx59632, nx59636, nx59648, nx59660, nx59664, nx59672, nx59678, 
         nx59690, nx59702, nx59706, nx59718, nx59730, nx59734, nx59738, nx59750, 
         nx59762, nx59766, nx59778, nx59790, nx59794, nx59798, nx59802, nx59816, 
         nx59828, nx59840, nx59844, nx59856, nx59868, nx59872, nx59880, nx59886, 
         nx59890, nx59894, nx59908, nx59920, nx59924, nx59936, nx59948, nx59952, 
         nx59956, nx59968, nx59980, nx59984, nx59996, nx60008, nx60012, nx60016, 
         nx60020, nx60032, nx60044, nx60048, nx60060, nx60072, nx60076, nx60080, 
         nx60092, nx60104, nx60108, nx60120, nx60132, nx60136, nx60140, nx60144, 
         nx60148, nx60162, nx60174, nx60178, nx60190, nx60202, nx60206, nx60210, 
         nx60222, nx60234, nx60238, nx60250, nx60262, nx60266, nx60270, nx60274, 
         nx60286, nx60298, nx60302, nx60314, nx60326, nx60330, nx60334, nx60346, 
         nx60358, nx60362, nx60374, nx60386, nx60390, nx60394, nx60398, nx60402, 
         nx60414, nx60426, nx60430, nx60442, nx60454, nx60458, nx60462, nx60474, 
         nx60486, nx60490, nx60502, nx60514, nx60518, nx60522, nx60526, nx60538, 
         nx60550, nx60554, nx60566, nx60578, nx60582, nx60586, nx60598, nx60610, 
         nx60614, nx60626, nx60638, nx60642, nx60646, nx60650, nx60654, nx60664, 
         nx60680, nx60692, nx60696, nx60708, nx60720, nx60724, nx60728, nx60740, 
         nx60752, nx60756, nx60768, nx60780, nx60784, nx60788, nx60792, nx60806, 
         nx60818, nx60830, nx60834, nx60846, nx60858, nx60862, nx60870, nx60876, 
         nx60888, nx60900, nx60904, nx60916, nx60928, nx60932, nx60936, nx60948, 
         nx60960, nx60964, nx60976, nx60988, nx60992, nx60996, nx61000, nx61014, 
         nx61026, nx61038, nx61042, nx61054, nx61066, nx61070, nx61078, nx61084, 
         nx61088, nx61100, nx61112, nx61116, nx61128, nx61140, nx61144, nx61148, 
         nx61160, nx61172, nx61176, nx61188, nx61200, nx61204, nx61208, nx61212, 
         nx61226, nx61238, nx61250, nx61254, nx61266, nx61278, nx61282, nx61290, 
         nx61296, nx61308, nx61320, nx61324, nx61336, nx61348, nx61352, nx61356, 
         nx61368, nx61380, nx61384, nx61396, nx61408, nx61412, nx61416, nx61420, 
         nx61434, nx61446, nx61458, nx61462, nx61474, nx61486, nx61490, nx61498, 
         nx61504, nx61508, nx61512, nx61524, nx61536, nx61540, nx61552, nx61564, 
         nx61568, nx61572, nx61584, nx61596, nx61600, nx61612, nx61624, nx61628, 
         nx61632, nx61636, nx61650, nx61662, nx61674, nx61678, nx61690, nx61702, 
         nx61706, nx61714, nx61720, nx61732, nx61744, nx61748, nx61760, nx61772, 
         nx61776, nx61780, nx61792, nx61804, nx61808, nx61820, nx61832, nx61836, 
         nx61840, nx61844, nx61858, nx61870, nx61882, nx61886, nx61898, nx61910, 
         nx61914, nx61922, nx61928, nx61932, nx61944, nx61956, nx61960, nx61972, 
         nx61984, nx61988, nx61992, nx62004, nx62016, nx62020, nx62032, nx62044, 
         nx62048, nx62052, nx62056, nx62070, nx62082, nx62094, nx62098, nx62110, 
         nx62122, nx62126, nx62134, nx62140, nx62152, nx62164, nx62168, nx62180, 
         nx62192, nx62196, nx62200, nx62212, nx62224, nx62228, nx62240, nx62252, 
         nx62256, nx62260, nx62264, nx62278, nx62290, nx62302, nx62306, nx62318, 
         nx62330, nx62334, nx62342, nx62348, nx62352, nx62356, nx62360, nx62376, 
         nx62388, nx62392, nx62404, nx62416, nx62420, nx62424, nx62436, nx62448, 
         nx62452, nx62464, nx62476, nx62480, nx62484, nx62488, nx62502, nx62514, 
         nx62526, nx62530, nx62542, nx62554, nx62558, nx62566, nx62572, nx62584, 
         nx62596, nx62600, nx62612, nx62624, nx62628, nx62632, nx62644, nx62656, 
         nx62660, nx62672, nx62684, nx62688, nx62692, nx62696, nx62710, nx62722, 
         nx62734, nx62738, nx62750, nx62762, nx62766, nx62774, nx62780, nx62784, 
         nx62796, nx62808, nx62812, nx62824, nx62836, nx62840, nx62844, nx62856, 
         nx62868, nx62872, nx62884, nx62896, nx62900, nx62904, nx62908, nx62922, 
         nx62934, nx62946, nx62950, nx62962, nx62974, nx62978, nx62986, nx62992, 
         nx63004, nx63016, nx63020, nx63032, nx63044, nx63048, nx63052, nx63064, 
         nx63076, nx63080, nx63092, nx63104, nx63108, nx63112, nx63116, nx63130, 
         nx63142, nx63154, nx63158, nx63170, nx63182, nx63186, nx63194, nx63200, 
         nx63204, nx63208, nx63220, nx63232, nx63236, nx63248, nx63260, nx63264, 
         nx63268, nx63280, nx63292, nx63296, nx63308, nx63320, nx63324, nx63328, 
         nx63332, nx63346, nx63358, nx63370, nx63374, nx63386, nx63398, nx63402, 
         nx63410, nx63416, nx63428, nx63440, nx63444, nx63456, nx63468, nx63472, 
         nx63476, nx63488, nx63500, nx63504, nx63516, nx63528, nx63532, nx63536, 
         nx63540, nx63554, nx63566, nx63578, nx63582, nx63594, nx63606, nx63610, 
         nx63618, nx63624, nx63628, nx63640, nx63652, nx63656, nx63668, nx63680, 
         nx63684, nx63688, nx63700, nx63712, nx63716, nx63728, nx63740, nx63744, 
         nx63748, nx63752, nx63766, nx63778, nx63790, nx63794, nx63806, nx63818, 
         nx63822, nx63830, nx63836, nx63848, nx63860, nx63864, nx63876, nx63888, 
         nx63892, nx63896, nx63908, nx63920, nx63924, nx63936, nx63948, nx63952, 
         nx63956, nx63960, nx63974, nx63986, nx63998, nx64002, nx64014, nx64026, 
         nx64030, nx64038, nx64044, nx64048, nx64052, nx64066, nx64078, nx64082, 
         nx64094, nx64106, nx64110, nx64114, nx64126, nx64138, nx64142, nx64154, 
         nx64166, nx64170, nx64174, nx64178, nx64190, nx64202, nx64206, nx64218, 
         nx64230, nx64234, nx64238, nx64250, nx64262, nx64266, nx64278, nx64290, 
         nx64294, nx64298, nx64302, nx64306, nx64320, nx64332, nx64336, nx64348, 
         nx64360, nx64364, nx64368, nx64380, nx64392, nx64396, nx64408, nx64420, 
         nx64424, nx64428, nx64432, nx64444, nx64456, nx64460, nx64472, nx64484, 
         nx64488, nx64492, nx64504, nx64516, nx64520, nx64532, nx64544, nx64548, 
         nx64552, nx64556, nx64560, nx64570, nx64582, nx64586, nx64598, nx64610, 
         nx64614, nx64618, nx64630, nx64642, nx64646, nx64658, nx64670, nx64674, 
         nx64678, nx64682, nx64694, nx64706, nx64710, nx64722, nx64734, nx64738, 
         nx64742, nx64754, nx64766, nx64770, nx64782, nx64794, nx64798, nx64802, 
         nx64806, nx64810, nx64822, nx64838, nx64850, nx64854, nx64866, nx64878, 
         nx64882, nx64886, nx64898, nx64910, nx64914, nx64926, nx64938, nx64942, 
         nx64946, nx64950, nx64964, nx64976, nx64988, nx64992, nx65004, nx65016, 
         nx65020, nx65028, nx65034, nx65046, nx65058, nx65062, nx65074, nx65086, 
         nx65090, nx65094, nx65106, nx65118, nx65122, nx65134, nx65146, nx65150, 
         nx65154, nx65158, nx65172, nx65184, nx65196, nx65200, nx65212, nx65224, 
         nx65228, nx65236, nx65242, nx65246, nx65258, nx65270, nx65274, nx65286, 
         nx65298, nx65302, nx65306, nx65318, nx65330, nx65334, nx65346, nx65358, 
         nx65362, nx65366, nx65370, nx65384, nx65396, nx65408, nx65412, nx65424, 
         nx65436, nx65440, nx65448, nx65454, nx65466, nx65478, nx65482, nx65494, 
         nx65506, nx65510, nx65514, nx65526, nx65538, nx65542, nx65554, nx65566, 
         nx65570, nx65574, nx65578, nx65592, nx65604, nx65616, nx65620, nx65632, 
         nx65644, nx65648, nx65656, nx65662, nx65666, nx65670, nx65682, nx65694, 
         nx65698, nx65710, nx65722, nx65726, nx65730, nx65742, nx65754, nx65758, 
         nx65770, nx65782, nx65786, nx65790, nx65794, nx65808, nx65820, nx65832, 
         nx65836, nx65848, nx65860, nx65864, nx65872, nx65878, nx65890, nx65902, 
         nx65906, nx65918, nx65930, nx65934, nx65938, nx65950, nx65962, nx65966, 
         nx65978, nx65990, nx65994, nx65998, nx66002, nx66016, nx66028, nx66040, 
         nx66044, nx66056, nx66068, nx66072, nx66080, nx66086, nx66090, nx66102, 
         nx66114, nx66118, nx66130, nx66142, nx66146, nx66150, nx66162, nx66174, 
         nx66178, nx66190, nx66202, nx66206, nx66210, nx66214, nx66228, nx66240, 
         nx66252, nx66256, nx66268, nx66280, nx66284, nx66292, nx66298, nx66310, 
         nx66322, nx66326, nx66338, nx66350, nx66354, nx66358, nx66370, nx66382, 
         nx66386, nx66398, nx66410, nx66414, nx66418, nx66422, nx66436, nx66448, 
         nx66460, nx66464, nx66476, nx66488, nx66492, nx66500, nx66506, nx66510, 
         nx66514, nx66518, nx8261, nx8271, nx8285, nx8319, nx8331, nx8363, 
         nx8375, nx8405, nx8417, nx8455, nx8467, nx8497, nx8511, nx8541, nx8553, 
         nx8585, nx8597, nx8625, nx8629, nx8735, nx8797, nx8809, nx8839, nx8853, 
         nx8885, nx8897, nx8927, nx8939, nx8971, nx8983, nx9015, nx9027, nx9059, 
         nx9071, nx9103, nx9113, nx9145, nx9155, nx9165, nx9195, nx9205, nx9237, 
         nx9249, nx9283, nx9295, nx9329, nx9341, nx9373, nx9383, nx9415, nx9427, 
         nx9457, nx9469, nx9499, nx9503, nx9605, nx9665, nx9677, nx9709, nx9721, 
         nx9753, nx9763, nx9795, nx9805, nx9839, nx9851, nx9881, nx9891, nx9927, 
         nx9939, nx9969, nx9983, nx10015, nx10023, nx10035, nx10067, nx10079, 
         nx10111, nx10125, nx10155, nx10167, nx10201, nx10213, nx10243, nx10257, 
         nx10289, nx10301, nx10333, nx10347, nx10375, nx10379, nx10477, nx10539, 
         nx10551, nx10583, nx10595, nx10627, nx10639, nx10669, nx10679, nx10713, 
         nx10725, nx10759, nx10771, nx10803, nx10815, nx10847, nx10859, nx10887, 
         nx10897, nx10907, nx10939, nx10949, nx10983, nx10995, nx11025, nx11037, 
         nx11071, nx11083, nx11115, nx11127, nx11159, nx11169, nx11201, nx11213, 
         nx11241, nx11245, nx11347, nx11407, nx11419, nx11449, nx11463, nx11495, 
         nx11507, nx11541, nx11553, nx11587, nx11601, nx11633, nx11645, nx11677, 
         nx11687, nx11717, nx11727, nx11759, nx11767, nx11777, nx11807, nx11821, 
         nx11853, nx11863, nx11893, nx11905, nx11939, nx11953, nx11983, nx11995, 
         nx12029, nx12041, nx12071, nx12083, nx12113, nx12117, nx12219, nx12279, 
         nx12291, nx12323, nx12337, nx12371, nx12381, nx12413, nx12425, nx12463, 
         nx12475, nx12505, nx12517, nx12549, nx12561, nx12593, nx12603, nx12633, 
         nx12641, nx12653, nx12685, nx12697, nx12729, nx12741, nx12771, nx12783, 
         nx12821, nx12833, nx12863, nx12877, nx12909, nx12921, nx12953, nx12965, 
         nx12993, nx12997, nx13101, nx13161, nx13173, nx13203, nx13217, nx13251, 
         nx13263, nx13293, nx13305, nx13339, nx13349, nx13381, nx13393, nx13425, 
         nx13439, nx13469, nx13483, nx13513, nx13521, nx13531, nx13561, nx13571, 
         nx13603, nx13615, nx13649, nx13661, nx13695, nx13707, nx13741, nx13753, 
         nx13785, nx13797, nx13827, nx13839, nx13869, nx13873, nx13973, nx14033, 
         nx14045, nx14077, nx14089, nx14121, nx14133, nx14167, nx14179, nx14213, 
         nx14225, nx14255, nx14267, nx14301, nx14315, nx14347, nx14359, nx14387, 
         nx14395, nx14409, nx14439, nx14449, nx14481, nx14493, nx14523, nx14537, 
         nx14569, nx14581, nx14613, nx14625, nx14657, nx14669, nx14699, nx14711, 
         nx14741, nx14745, nx14847, nx14905, nx14919, nx14947, nx14959, nx14991, 
         nx15001, nx15031, nx15041, nx15077, nx15089, nx15119, nx15133, nx15163, 
         nx15175, nx15207, nx15219, nx15247, nx15257, nx15269, nx15299, nx15311, 
         nx15345, nx15357, nx15387, nx15399, nx15433, nx15445, nx15479, nx15491, 
         nx15523, nx15535, nx15567, nx15579, nx15607, nx15611, nx15713, nx15775, 
         nx15785, nx15815, nx15825, nx15857, nx15869, nx15903, nx15915, nx15949, 
         nx15961, nx15993, nx16003, nx16035, nx16047, nx16077, nx16089, nx16121, 
         nx16129, nx16141, nx16171, nx16185, nx16215, nx16227, nx16259, nx16271, 
         nx16303, nx16317, nx16349, nx16361, nx16393, nx16405, nx16435, nx16447, 
         nx16475, nx16479, nx16581, nx16643, nx16655, nx16685, nx16695, nx16727, 
         nx16737, nx16771, nx16783, nx16817, nx16831, nx16861, nx16871, nx16903, 
         nx16915, nx16945, nx16959, nx16989, nx16997, nx17009, nx17041, nx17053, 
         nx17085, nx17095, nx17127, nx17139, nx17175, nx17187, nx17217, nx17229, 
         nx17263, nx17275, nx17305, nx17319, nx17347, nx17351, nx17455, nx17515, 
         nx17527, nx17557, nx17567, nx17601, nx17613, nx17643, nx17655, nx17691, 
         nx17701, nx17731, nx17743, nx17775, nx17787, nx17821, nx17833, nx17861, 
         nx17869, nx17883, nx17913, nx17925, nx17959, nx17971, nx18001, nx18015, 
         nx18049, nx18061, nx18093, nx18103, nx18135, nx18147, nx18179, nx18191, 
         nx18219, nx18223, nx18327, nx18385, nx18397, nx18427, nx18441, nx18473, 
         nx18485, nx18517, nx18529, nx18563, nx18575, nx18605, nx18617, nx18651, 
         nx18663, nx18695, nx18705, nx18733, nx18741, nx18755, nx18785, nx18797, 
         nx18831, nx18843, nx18873, nx18887, nx18919, nx18931, nx18963, nx18975, 
         nx19007, nx19017, nx19047, nx19057, nx19088, nx19091, nx19191, nx19253, 
         nx19263, nx19295, nx19305, nx19337, nx19347, nx19377, nx19389, nx19425, 
         nx19437, nx19467, nx19479, nx19513, nx19525, nx19555, nx19569, nx19597, 
         nx19605, nx19617, nx19651, nx19663, nx19695, nx19709, nx19737, nx19749, 
         nx19783, nx19795, nx19825, nx19839, nx19871, nx19883, nx19913, nx19925, 
         nx19953, nx19957, nx20059, nx20117, nx20131, nx20161, nx20173, nx20205, 
         nx20217, nx20247, nx20261, nx20295, nx20307, nx20337, nx20349, nx20381, 
         nx20391, nx20421, nx20433, nx20461, nx20471, nx20483, nx20513, nx20525, 
         nx20559, nx20569, nx20599, nx20609, nx20643, nx20655, nx20689, nx20701, 
         nx20733, nx20745, nx20781, nx20793, nx20821, nx20825, nx20927, nx20987, 
         nx20997, nx21027, nx21039, nx21073, nx21085, nx21117, nx21127, nx21163, 
         nx21175, nx21209, nx21221, nx21253, nx21267, nx21297, nx21309, nx21339, 
         nx21349, nx21361, nx21391, nx21405, nx21435, nx21447, nx21479, nx21491, 
         nx21525, nx21539, nx21569, nx21583, nx21617, nx21631, nx21661, nx21673, 
         nx21701, nx21705, nx21807, nx21867, nx21879, nx21911, nx21923, nx21955, 
         nx21967, nx21997, nx22009, nx22045, nx22057, nx22087, nx22097, nx22129, 
         nx22141, nx22173, nx22183, nx22217, nx22219, nx22221, nx22223, nx22225, 
         nx22227, nx22229, nx22231, nx22233, nx22235, nx22237, nx22239, nx22241, 
         nx22243, nx22245, nx22247, nx22249, nx22251, nx22253, nx22255, nx22257, 
         nx22259, nx22261, nx22263, nx22265, nx22267, nx22269, nx22271, nx22273, 
         nx22275, nx22277, nx22279, nx22281, nx22283, nx22285, nx22287, nx22289, 
         nx22291, nx22293, nx22295, nx22297, nx22299, nx22301, nx22303, nx22305, 
         nx22307, nx22309, nx22311, nx22313, nx22315, nx22317, nx22319, nx22321, 
         nx22323, nx22325, nx22327, nx22329, nx22331, nx22333, nx22335, nx22337, 
         nx22339, nx22341, nx22343, nx22345, nx22347, nx22349, nx22351, nx22353, 
         nx22355, nx22357, nx22359, nx22361, nx22363, nx22365, nx22367, nx22369, 
         nx22371, nx22373, nx22375, nx22377, nx22379, nx22381, nx22383, nx22385, 
         nx22387, nx22393, nx22395, nx22397, nx22399, nx22401, nx22403, nx22405, 
         nx22407, nx22411, nx22413, nx22415, nx22417, nx22419, nx22421, nx22423, 
         nx22425, nx22427, nx22429, nx22431, nx22433, nx22435, nx22437, nx22439, 
         nx22441, nx22443, nx22445, nx22447, nx22451, nx22453, nx22455, nx22457, 
         nx22459, nx22461, nx22463, nx22465, nx22467, nx22469, nx22471, nx22473, 
         nx22475, nx22477, nx22479, nx22481, nx22483, nx22485, nx22487, nx22489, 
         nx22491, nx22493, nx22495, nx22497, nx22499, nx22501, nx22503, nx22505, 
         nx22507, nx22509, nx22511, nx22513, nx22515, nx22517, nx22519, nx22521, 
         nx22523, nx22527, nx22529, nx22531, nx22533, nx22535, nx22537, nx22539, 
         nx22541, nx22543, nx22545, nx22547, nx22549, nx22551, nx22553, nx22555, 
         nx22557, nx22559, nx22561, nx22563, nx22565, nx22567, nx22569, nx22571, 
         nx22573, nx22575, nx22577, nx22579, nx22581, nx22583, nx22585, nx22587, 
         nx22589, nx22591, nx22593, nx22595, nx22597, nx22599, nx22601, nx22603, 
         nx22605, nx22607, nx22609, nx22611, nx22613, nx22615, nx22617, nx22619, 
         nx22621, nx22623, nx22625, nx22627, nx22629, nx22631, nx22633, nx22635, 
         nx22637, nx22639, nx22641, nx22643, nx22645, nx22647, nx22649, nx22651, 
         nx22653, nx22655, nx22657, nx22659, nx22661, nx22663, nx22665, nx22667, 
         nx22669, nx22671, nx22673, nx22677, nx22679, nx22681, nx22683, nx22685, 
         nx22687, nx22689, nx22691, nx22693, nx22695, nx22697, nx22699, nx22701, 
         nx22703, nx22705, nx22707, nx22709, nx22711, nx22713, nx22715, nx22717, 
         nx22719, nx22721, nx22723, nx22725, nx22727, nx22729, nx22731, nx22733, 
         nx22735, nx22737, nx22739, nx22741, nx22743, nx22745, nx22747, nx22749, 
         nx22751, nx22753, nx22755, nx22757, nx22759, nx22761, nx22763, nx22765, 
         nx22767, nx22769, nx22771, nx22773, nx22775, nx22777, nx22779, nx22781, 
         nx22783, nx22785, nx22787, nx22789, nx22791, nx22793, nx22795, nx22797, 
         nx22799, nx22801, nx22803, nx22805, nx22807, nx22809, nx22811, nx22813, 
         nx22815, nx22817, nx22819, nx22821, nx22823, nx22825, nx22827, nx22829, 
         nx22831, nx22833, nx22835, nx22837, nx22839, nx22841, nx22843, nx22845, 
         nx22847, nx22849, nx22851, nx22853, nx22855, nx22857, nx22859, nx22861, 
         nx22863, nx22865, nx22867, nx22869, nx22871, nx22873, nx22875, nx22877, 
         nx22879, nx22881, nx22883, nx22885, nx22887, nx22889, nx22891, nx22893, 
         nx22895, nx22897, nx22899, nx22901, nx22903, nx22905, nx22907, nx22909, 
         nx22911, nx22913, nx22915, nx22917, nx22919, nx22921, nx22923, nx22925, 
         nx22927, nx22929, nx22931, nx22933, nx22935, nx22937, nx22939, nx22941, 
         nx22943, nx22945, nx22947, nx22949, nx22951, nx22953, nx22955, nx22957, 
         nx22959, nx22961, nx22963, nx22965, nx22967, nx22969, nx22971, nx22973, 
         nx22975, nx22977, nx22979, nx22981, nx22983, nx22985, nx22987, nx22989, 
         nx22991, nx22993, nx22995, nx22997, nx22999, nx23001, nx23003, nx23005, 
         nx23007, nx23009, nx23011, nx23013, nx23015, nx23017, nx23019, nx23021, 
         nx23023, nx23025, nx23027, nx23029, nx23031, nx23033, nx23035, nx23037, 
         nx23039, nx23041, nx23043, nx23045, nx23047, nx23049, nx23051, nx23053, 
         nx23055, nx23057, nx23059, nx23061, nx23063, nx23065, nx23067, nx23069, 
         nx23071, nx23073, nx23075, nx23077, nx23079, nx23081, nx23083, nx23085, 
         nx23087, nx23089, nx23091, nx23093, nx23095, nx23097, nx23099, nx23101, 
         nx23103, nx23105, nx23107, nx23109, nx23111, nx23113, nx23115, nx23117, 
         nx23119, nx23121, nx23123, nx23125, nx23127, nx23129, nx23131, nx23133, 
         nx23135, nx23137, nx23139, nx23141, nx23143, nx23145, nx23147, nx23149, 
         nx23151, nx23153, nx23155, nx23157, nx23159, nx23161, nx23163, nx23165, 
         nx23167, nx23169, nx23171, nx23173, nx23175, nx23177, nx23179, nx23181, 
         nx23183, nx23185, nx23187, nx23189, nx23191, nx23193, nx23195, nx23197, 
         nx23199, nx23201, nx23203, nx23205, nx23207, nx23209, nx23211, nx23213, 
         nx23215, nx23217, nx23219, nx23221, nx23223, nx23225, nx23227, nx23229, 
         nx23231, nx23233, nx23235, nx23237, nx23239, nx23241, nx23243, nx23245, 
         nx23247, nx23249, nx23251, nx23253, nx23255, nx23257, nx23259, nx23261, 
         nx23263, nx23265, nx23267, nx23269, nx23271, nx23273, nx23275, nx23277, 
         nx23279, nx23281, nx23283, nx23285, nx23287, nx23289, nx23291, nx23293, 
         nx23295, nx23297, nx23299, nx23301, nx23303, nx23305, nx23307, nx23309, 
         nx23311, nx23313, nx23315, nx23317, nx23319, nx23321, nx23323, nx23325, 
         nx23327, nx23329, nx23331, nx23333, nx23335, nx23337, nx23339, nx23341, 
         nx23343, nx23345, nx23347, nx23349, nx23351, nx23353, nx23355, nx23357, 
         nx23361, nx23363, nx23365, nx23367, nx23369, nx23371, nx23373, nx23375, 
         nx23377, nx23379, nx23381, nx23383, nx23385, nx23387, nx23389, nx23391, 
         nx23393, nx23395, nx23397, nx23399, nx23401, nx23403, nx23405, nx23407, 
         nx23409, nx23411, nx23413, nx23415, nx23417, nx23419, nx23421, nx23423, 
         nx23425, nx23427, nx23429, nx23431, nx23433, nx23435, nx23437, nx23439, 
         nx23441, nx23443, nx23445, nx23447, nx23449, nx23451, nx23453, nx23455, 
         nx23457, nx23459, nx23461, nx23463, nx23465, nx23467, nx23469, nx23471, 
         nx23473, nx23475, nx23477, nx23479, nx23481, nx23483, nx23485, nx23487, 
         nx23489, nx23491, nx23493, nx23495, nx23497, nx23499, nx23501, nx23503, 
         nx23505, nx23507, nx23509, nx23511, nx23513, nx23515, nx23517, nx23519, 
         nx23521, nx23523, nx23525, nx23527, nx23529, nx23531, nx23533, nx23535, 
         nx23537, nx23539, nx23541, nx23543, nx23545, nx23547, nx23549, nx23551, 
         nx23553, nx23555, nx23557, nx23559, nx23561, nx23563, nx23565, nx23567, 
         nx23569, nx23571, nx23573, nx23575, nx23577, nx23579, nx23581, nx23583, 
         nx23585, nx23587, nx23589, nx23591, nx23593, nx23595, nx23597, nx23599, 
         nx23601, nx23603, nx23605, nx23607, nx23609, nx23611, nx23613, nx23615, 
         nx23617, nx23619, nx23621, nx23623, nx23625, nx23627, nx23629, nx23631, 
         nx23633, nx23635, nx23637, nx23639, nx23641, nx23643, nx23645, nx23647, 
         nx23649, nx23651, nx23653, nx23655, nx23657, nx23659, nx23661, nx23663, 
         nx23665, nx23667, nx23669, nx23671, nx23673, nx23675, nx23677, nx23679, 
         nx23681, nx23683, nx23685, nx23687, nx23689, nx23691, nx23693, nx23695, 
         nx23697, nx23699, nx23701, nx23703, nx23705, nx23707, nx23709, nx23711, 
         nx23713, nx23715, nx23717, nx23719, nx23721, nx23723, nx23725, nx23727, 
         nx23729, nx23731, nx23733, nx23735, nx23737, nx23739, nx23741, nx23743, 
         nx23745, nx23747, nx23749, nx23751, nx23753, nx23755, nx23757, nx23759, 
         nx23761, nx23763, nx23765, nx23767, nx23769, nx23771, nx23773, nx23775, 
         nx23777, nx23779, nx23781, nx23783, nx23785, nx23787, nx23789, nx23791, 
         nx23793, nx23795, nx23797, nx23799, nx23801, nx23803, nx23805, nx23807, 
         nx23809, nx23811, nx23813, nx23815, nx23817, nx23819, nx23821, nx23823, 
         nx23825, nx23827, nx23829, nx23831, nx23833, nx23835, nx23837, nx23839, 
         nx23841, nx23843, nx23845, nx23847, nx23849, nx23851, nx23853, nx23855, 
         nx23857, nx23859, nx23861, nx23863, nx23865, nx23867, nx23869, nx23871, 
         nx23873, nx23875, nx23877, nx23879, nx23881, nx23883, nx23885, nx23887, 
         nx23889, nx23891, nx23893, nx23895, nx23897, nx23899, nx23901, nx23903, 
         nx23905, nx23907, nx23909, nx23911, nx23913, nx23915, nx23917, nx23919, 
         nx23921, nx23923, nx23925, nx23927, nx23929, nx23931, nx23933, nx23935, 
         nx23937, nx23939, nx23941, nx23943, nx23945, nx23947, nx23949, nx23951, 
         nx23953, nx23955, nx23957, nx23959, nx23961, nx23963, nx23965, nx23967, 
         nx23969, nx23971, nx23973, nx23975, nx23977, nx23979, nx23981, nx23983, 
         nx23985, nx23987, nx23989, nx23991, nx23993, nx23995, nx23997, nx23999, 
         nx24001, nx24003, nx24005, nx24007, nx24009, nx24011, nx24013, nx24015, 
         nx24017, nx24019, nx24021, nx24023, nx24025, nx24027, nx24029, nx24031, 
         nx24033, nx24035, nx24037, nx24039, nx24041, nx24043, nx24045, nx24047, 
         nx24049, nx24051, nx24053, nx24055, nx24057, nx24059, nx24061, nx24063, 
         nx24065, nx24067, nx24069, nx24071, nx24073, nx24075, nx24077, nx24079, 
         nx24081, nx24083, nx24085, nx24087, nx24089, nx24091, nx24093, nx24095, 
         nx24097, nx24099, nx24101, nx24103, nx24105, nx24107, nx24109, nx24111, 
         nx24113, nx24115, nx24117, nx24119, nx24121, nx24123, nx24125, nx24127, 
         nx24129, nx24131, nx24133, nx24135, nx24137, nx24139, nx24141, nx24143, 
         nx24145, nx24147, nx24149, nx24151, nx24153, nx24155, nx24157, nx24159, 
         nx24161, nx24163, nx24165, nx24167, nx24169, nx24171, nx24173, nx24175, 
         nx24177, nx24179, nx24181, nx24183, nx24185, nx24187, nx24189, nx24191, 
         nx24193, nx24195, nx24197, nx24199, nx24201, nx24203, nx24205, nx24207, 
         nx24209, nx24211, nx24213, nx24215, nx24217, nx24219, nx24221, nx24223, 
         nx24225, nx24227, nx24229, nx24231, nx24233, nx24235, nx24237, nx24239, 
         nx24241, nx24243, nx24245, nx24247, nx24249, nx24251, nx24253, nx24255, 
         nx24257, nx24259, nx24261, nx24263, nx24265, nx24267, nx24269, nx24271, 
         nx24273, nx24275, nx24277, nx24279, nx24281, nx24283, nx24285, nx24287, 
         nx24289, nx24291, nx24293, nx24295, nx24297, nx24299, nx24301, nx24303, 
         nx24305, nx24307, nx24309, nx24311, nx24313, nx24315, nx24317, nx24319, 
         nx24321, nx24323, nx24325, nx24327, nx24329, nx24331, nx24333, nx24335, 
         nx24337, nx24339, nx24341, nx24343, nx24345, nx24347, nx24349, nx24351, 
         nx24353, nx24355, nx24357, nx24359, nx24361, nx24363, nx24365, nx24367, 
         nx24369, nx24371, nx24373, nx24375, nx24377, nx24379, nx24381, nx24383, 
         nx24385, nx24387, nx24389, nx24391, nx24393, nx24395, nx24397, nx24399, 
         nx24401, nx24403, nx24405, nx24407, nx24409, nx24411, nx24413, nx24415, 
         nx24417, nx24419, nx24421, nx24423, nx24425, nx24427, nx24429, nx24431, 
         nx24433, nx24435, nx24437, nx24439, nx24441, nx24443, nx24445, nx24447, 
         nx24449, nx24451, nx24453, nx24455, nx24457, nx24459, nx24461, nx24463, 
         nx24465, nx24467, nx24469, nx24471, nx24473, nx24475, nx24477, nx24479, 
         nx24481, nx24483, nx24485, nx24487, nx24489, nx24491, nx24493, nx24495, 
         nx24497, nx24499, nx24501, nx24503, nx24505, nx24507, nx24509, nx24511, 
         nx24513, nx24515, nx24517, nx24519, nx24521, nx24523, nx24525, nx24527, 
         nx24529, nx24531, nx24533, nx24535, nx24537, nx24539, nx24541, nx24543, 
         nx24545, nx24547, nx24549, nx24551, nx24553, nx24555, nx24557, nx24559, 
         nx24561, nx24563, nx24565, nx24567, nx24569, nx24571, nx24573, nx24575, 
         nx24577, nx24579, nx24581, nx24583, nx24585, nx24587, nx24589, nx24591, 
         nx24593, nx24595, nx24597, nx24599, nx24601, nx24603, nx24605, nx24607, 
         nx24609, nx24611, nx24613, nx24615, nx24617, nx24619, nx24621, nx24623, 
         nx24625, nx24627, nx24629, nx24631, nx24633, nx24635, nx24637, nx24639, 
         nx24641, nx24643, nx24645, nx24647, nx24649, nx24651, nx24653, nx24655, 
         nx24657, nx24659, nx24661, nx24663, nx24665, nx24667, nx24669, nx24671, 
         nx24673, nx24675, nx24677, nx24679, nx24681, nx24683, nx24685, nx24687, 
         nx24689, nx24691, nx24693, nx24695, nx24697, nx24699, nx24701, nx24703, 
         nx24705, nx24707, nx24709, nx24711, nx24713, nx24715, nx24717, nx24719, 
         nx24721, nx24723, nx24725, nx24727, nx24729, nx24731, nx24733, nx24735, 
         nx24737, nx24739, nx24741, nx24743, nx24745, nx24747, nx24749, nx24751, 
         nx24753, nx24755, nx24757, nx24759, nx24761, nx24763, nx24765, nx24767, 
         nx24769, nx24771, nx24773, nx24775, nx24777, nx24779, nx24781, nx24783, 
         nx24785, nx24787, nx24789, nx24791, nx24793, nx24795, nx24797, nx24799, 
         nx24801, nx24803, nx24805, nx24807, nx24809, nx24811, nx24813, nx24815, 
         nx24817, nx24819, nx24821, nx24823, nx24825, nx24827, nx24829, nx24831, 
         nx24833, nx24835, nx24837, nx24839, nx24841, nx24843, nx24845, nx24847, 
         nx24849, nx24851, nx24853, nx24855, nx24857, nx24859, nx24861, nx24863, 
         nx24865, nx24867, nx24869, nx24871, nx24873, nx24875, nx24877, nx24879, 
         nx24881, nx24883, nx24885, nx24887, nx24889, nx24891, nx24893, nx24895, 
         nx24897, nx24899, nx24901, nx24903, nx24905, nx24907, nx24909, nx24911, 
         nx24913, nx24915, nx24917, nx24919, nx24921, nx24923, nx24925, nx24927, 
         nx24929, nx24931, nx24933, nx24935, nx24937, nx24939, nx24941, nx24943, 
         nx24945, nx24947, nx24949, nx24951, nx24953, nx24955, nx24957, nx24959, 
         nx24961, nx24963, nx24965, nx24967, nx24969, nx24971, nx24973, nx24975, 
         nx24977, nx24979, nx24981, nx24983, nx24985, nx24987, nx24989, nx24991, 
         nx24993, nx24995, nx24997, nx24999, nx25001, nx25003, nx25005, nx25007, 
         nx25009, nx25011, nx25013, nx25015, nx25017, nx25019, nx25021, nx25023, 
         nx25025, nx25027, nx25029, nx25031, nx25033, nx25035, nx25037, nx25039, 
         nx25041, nx25043, nx25045, nx25047, nx25049, nx25051, nx25053, nx25055, 
         nx25057, nx25059, nx25061, nx25063, nx25065, nx25067, nx25069, nx25071, 
         nx25073, nx25075, nx25077, nx25079, nx25081, nx25083, nx25085, nx25087, 
         nx25089, nx25091, nx25093, nx25095, nx25097, nx25099, nx25101, nx25103, 
         nx25105, nx25107, nx25109, nx25111, nx25113, nx25115, nx25117, nx25119, 
         nx25121, nx25123, nx25125, nx25127, nx25129, nx25131, nx25133, nx25135, 
         nx25137, nx25139, nx25141, nx25143, nx25145, nx25147, nx25149, nx25151, 
         nx25153, nx25155, nx25157, nx25159, nx25161, nx25163, nx25165, nx25167, 
         nx25169, nx25171, nx25173, nx25175, nx25177, nx25179, nx25181, nx25183, 
         nx25185, nx25187, nx25189, nx25191, nx25193, nx25195, nx25201, nx25203, 
         nx25205, nx25207, nx25209, nx25211, nx25213, nx25215, nx25217, nx25219, 
         nx25221, nx25223, nx25225, nx25227, nx25229, nx25231, nx25233, nx25235, 
         nx25237, nx25239, nx25241, nx25243, nx25245, nx25247, nx25249;



    oai21 ix4157 (.Y (\output [0]), .A0 (nx24851), .A1 (nx8261), .B0 (nx8625)) ;
    mux21 ix8262 (.Y (nx8261), .A0 (nx838), .A1 (nx1682), .S0 (nx22411)) ;
    mux21_ni ix839 (.Y (nx838), .A0 (nx414), .A1 (nx834), .S0 (nx22451)) ;
    mux21_ni ix415 (.Y (nx414), .A0 (nx202), .A1 (nx410), .S0 (nx22527)) ;
    mux21_ni ix203 (.Y (nx202), .A0 (nx196), .A1 (nx118), .S0 (nx23117)) ;
    oai21 ix197 (.Y (nx196), .A0 (nx24855), .A1 (nx8271), .B0 (nx8285)) ;
    mux21 ix8272 (.Y (nx8271), .A0 (nx160), .A1 (nx188), .S0 (nx22677)) ;
    mux21_ni ix161 (.Y (nx160), .A0 (nx144), .A1 (nx156), .S0 (nx23361)) ;
    mux21_ni ix145 (.Y (nx144), .A0 (inputs_260__0), .A1 (inputs_261__0), .S0 (
             nx23883)) ;
    mux21_ni ix157 (.Y (nx156), .A0 (inputs_262__0), .A1 (inputs_263__0), .S0 (
             nx23883)) ;
    mux21_ni ix189 (.Y (nx188), .A0 (nx172), .A1 (nx184), .S0 (nx23361)) ;
    mux21_ni ix173 (.Y (nx172), .A0 (inputs_276__0), .A1 (inputs_277__0), .S0 (
             nx23883)) ;
    mux21_ni ix185 (.Y (nx184), .A0 (inputs_278__0), .A1 (inputs_279__0), .S0 (
             nx23883)) ;
    nand04 ix8286 (.Y (nx8285), .A0 (nx24855), .A1 (nx23361), .A2 (nx23883), .A3 (
           nx132)) ;
    mux21_ni ix133 (.Y (nx132), .A0 (inputs_259__0), .A1 (inputs_275__0), .S0 (
             nx22677)) ;
    mux21_ni ix119 (.Y (nx118), .A0 (nx54), .A1 (nx114), .S0 (nx22677)) ;
    mux21_ni ix55 (.Y (nx54), .A0 (nx22), .A1 (nx50), .S0 (nx23191)) ;
    mux21_ni ix23 (.Y (nx22), .A0 (nx6), .A1 (nx18), .S0 (nx23361)) ;
    mux21_ni ix7 (.Y (nx6), .A0 (inputs_264__0), .A1 (inputs_265__0), .S0 (
             nx23883)) ;
    mux21_ni ix19 (.Y (nx18), .A0 (inputs_266__0), .A1 (inputs_267__0), .S0 (
             nx23883)) ;
    mux21_ni ix51 (.Y (nx50), .A0 (nx34), .A1 (nx46), .S0 (nx23361)) ;
    mux21_ni ix35 (.Y (nx34), .A0 (inputs_268__0), .A1 (inputs_269__0), .S0 (
             nx23885)) ;
    mux21_ni ix47 (.Y (nx46), .A0 (inputs_270__0), .A1 (inputs_271__0), .S0 (
             nx23885)) ;
    mux21_ni ix115 (.Y (nx114), .A0 (nx82), .A1 (nx110), .S0 (nx23191)) ;
    mux21_ni ix83 (.Y (nx82), .A0 (nx66), .A1 (nx78), .S0 (nx23361)) ;
    mux21_ni ix67 (.Y (nx66), .A0 (inputs_280__0), .A1 (inputs_281__0), .S0 (
             nx23885)) ;
    mux21_ni ix79 (.Y (nx78), .A0 (inputs_282__0), .A1 (inputs_283__0), .S0 (
             nx23885)) ;
    mux21_ni ix111 (.Y (nx110), .A0 (nx94), .A1 (nx106), .S0 (nx23361)) ;
    mux21_ni ix95 (.Y (nx94), .A0 (inputs_284__0), .A1 (inputs_285__0), .S0 (
             nx23885)) ;
    mux21_ni ix107 (.Y (nx106), .A0 (inputs_286__0), .A1 (inputs_287__0), .S0 (
             nx23885)) ;
    mux21_ni ix411 (.Y (nx410), .A0 (nx404), .A1 (nx326), .S0 (nx23117)) ;
    oai21 ix405 (.Y (nx404), .A0 (nx24855), .A1 (nx8319), .B0 (nx8331)) ;
    mux21 ix8320 (.Y (nx8319), .A0 (nx368), .A1 (nx396), .S0 (nx22677)) ;
    mux21_ni ix369 (.Y (nx368), .A0 (nx352), .A1 (nx364), .S0 (nx23363)) ;
    mux21_ni ix353 (.Y (nx352), .A0 (inputs_292__0), .A1 (inputs_293__0), .S0 (
             nx23885)) ;
    mux21_ni ix365 (.Y (nx364), .A0 (inputs_294__0), .A1 (inputs_295__0), .S0 (
             nx23887)) ;
    mux21_ni ix397 (.Y (nx396), .A0 (nx380), .A1 (nx392), .S0 (nx23363)) ;
    mux21_ni ix381 (.Y (nx380), .A0 (inputs_308__0), .A1 (inputs_309__0), .S0 (
             nx23887)) ;
    mux21_ni ix393 (.Y (nx392), .A0 (inputs_310__0), .A1 (inputs_311__0), .S0 (
             nx23887)) ;
    nand04 ix8332 (.Y (nx8331), .A0 (nx24855), .A1 (nx23363), .A2 (nx23887), .A3 (
           nx340)) ;
    mux21_ni ix341 (.Y (nx340), .A0 (inputs_291__0), .A1 (inputs_307__0), .S0 (
             nx22677)) ;
    mux21_ni ix327 (.Y (nx326), .A0 (nx262), .A1 (nx322), .S0 (nx22677)) ;
    mux21_ni ix263 (.Y (nx262), .A0 (nx230), .A1 (nx258), .S0 (nx23191)) ;
    mux21_ni ix231 (.Y (nx230), .A0 (nx214), .A1 (nx226), .S0 (nx23363)) ;
    mux21_ni ix215 (.Y (nx214), .A0 (inputs_296__0), .A1 (inputs_297__0), .S0 (
             nx23887)) ;
    mux21_ni ix227 (.Y (nx226), .A0 (inputs_298__0), .A1 (inputs_299__0), .S0 (
             nx23887)) ;
    mux21_ni ix259 (.Y (nx258), .A0 (nx242), .A1 (nx254), .S0 (nx23363)) ;
    mux21_ni ix243 (.Y (nx242), .A0 (inputs_300__0), .A1 (inputs_301__0), .S0 (
             nx23887)) ;
    mux21_ni ix255 (.Y (nx254), .A0 (inputs_302__0), .A1 (inputs_303__0), .S0 (
             nx23889)) ;
    mux21_ni ix323 (.Y (nx322), .A0 (nx290), .A1 (nx318), .S0 (nx23191)) ;
    mux21_ni ix291 (.Y (nx290), .A0 (nx274), .A1 (nx286), .S0 (nx23363)) ;
    mux21_ni ix275 (.Y (nx274), .A0 (inputs_312__0), .A1 (inputs_313__0), .S0 (
             nx23889)) ;
    mux21_ni ix287 (.Y (nx286), .A0 (inputs_314__0), .A1 (inputs_315__0), .S0 (
             nx23889)) ;
    mux21_ni ix319 (.Y (nx318), .A0 (nx302), .A1 (nx314), .S0 (nx23363)) ;
    mux21_ni ix303 (.Y (nx302), .A0 (inputs_316__0), .A1 (inputs_317__0), .S0 (
             nx23889)) ;
    mux21_ni ix315 (.Y (nx314), .A0 (inputs_318__0), .A1 (inputs_319__0), .S0 (
             nx23889)) ;
    mux21_ni ix835 (.Y (nx834), .A0 (nx622), .A1 (nx830), .S0 (nx22527)) ;
    mux21_ni ix623 (.Y (nx622), .A0 (nx616), .A1 (nx538), .S0 (nx23117)) ;
    oai21 ix617 (.Y (nx616), .A0 (nx24855), .A1 (nx8363), .B0 (nx8375)) ;
    mux21 ix8364 (.Y (nx8363), .A0 (nx580), .A1 (nx608), .S0 (nx22677)) ;
    mux21_ni ix581 (.Y (nx580), .A0 (nx564), .A1 (nx576), .S0 (nx23365)) ;
    mux21_ni ix565 (.Y (nx564), .A0 (inputs_324__0), .A1 (inputs_325__0), .S0 (
             nx23889)) ;
    mux21_ni ix577 (.Y (nx576), .A0 (inputs_326__0), .A1 (inputs_327__0), .S0 (
             nx23889)) ;
    mux21_ni ix609 (.Y (nx608), .A0 (nx592), .A1 (nx604), .S0 (nx23365)) ;
    mux21_ni ix593 (.Y (nx592), .A0 (inputs_340__0), .A1 (inputs_341__0), .S0 (
             nx23891)) ;
    mux21_ni ix605 (.Y (nx604), .A0 (inputs_342__0), .A1 (inputs_343__0), .S0 (
             nx23891)) ;
    nand04 ix8376 (.Y (nx8375), .A0 (nx24855), .A1 (nx23365), .A2 (nx23891), .A3 (
           nx552)) ;
    mux21_ni ix553 (.Y (nx552), .A0 (inputs_323__0), .A1 (inputs_339__0), .S0 (
             nx22679)) ;
    mux21_ni ix539 (.Y (nx538), .A0 (nx474), .A1 (nx534), .S0 (nx22679)) ;
    mux21_ni ix475 (.Y (nx474), .A0 (nx442), .A1 (nx470), .S0 (nx23191)) ;
    mux21_ni ix443 (.Y (nx442), .A0 (nx426), .A1 (nx438), .S0 (nx23365)) ;
    mux21_ni ix427 (.Y (nx426), .A0 (inputs_328__0), .A1 (inputs_329__0), .S0 (
             nx23891)) ;
    mux21_ni ix439 (.Y (nx438), .A0 (inputs_330__0), .A1 (inputs_331__0), .S0 (
             nx23891)) ;
    mux21_ni ix471 (.Y (nx470), .A0 (nx454), .A1 (nx466), .S0 (nx23365)) ;
    mux21_ni ix455 (.Y (nx454), .A0 (inputs_332__0), .A1 (inputs_333__0), .S0 (
             nx23891)) ;
    mux21_ni ix467 (.Y (nx466), .A0 (inputs_334__0), .A1 (inputs_335__0), .S0 (
             nx23891)) ;
    mux21_ni ix535 (.Y (nx534), .A0 (nx502), .A1 (nx530), .S0 (nx23191)) ;
    mux21_ni ix503 (.Y (nx502), .A0 (nx486), .A1 (nx498), .S0 (nx23365)) ;
    mux21_ni ix487 (.Y (nx486), .A0 (inputs_344__0), .A1 (inputs_345__0), .S0 (
             nx23893)) ;
    mux21_ni ix499 (.Y (nx498), .A0 (inputs_346__0), .A1 (inputs_347__0), .S0 (
             nx23893)) ;
    mux21_ni ix531 (.Y (nx530), .A0 (nx514), .A1 (nx526), .S0 (nx23365)) ;
    mux21_ni ix515 (.Y (nx514), .A0 (inputs_348__0), .A1 (inputs_349__0), .S0 (
             nx23893)) ;
    mux21_ni ix527 (.Y (nx526), .A0 (inputs_350__0), .A1 (inputs_351__0), .S0 (
             nx23893)) ;
    mux21_ni ix831 (.Y (nx830), .A0 (nx824), .A1 (nx746), .S0 (nx23117)) ;
    oai21 ix825 (.Y (nx824), .A0 (nx24855), .A1 (nx8405), .B0 (nx8417)) ;
    mux21 ix8406 (.Y (nx8405), .A0 (nx788), .A1 (nx816), .S0 (nx22679)) ;
    mux21_ni ix789 (.Y (nx788), .A0 (nx772), .A1 (nx784), .S0 (nx23367)) ;
    mux21_ni ix773 (.Y (nx772), .A0 (inputs_356__0), .A1 (inputs_357__0), .S0 (
             nx23893)) ;
    mux21_ni ix785 (.Y (nx784), .A0 (inputs_358__0), .A1 (inputs_359__0), .S0 (
             nx23893)) ;
    mux21_ni ix817 (.Y (nx816), .A0 (nx800), .A1 (nx812), .S0 (nx23367)) ;
    mux21_ni ix801 (.Y (nx800), .A0 (inputs_372__0), .A1 (inputs_373__0), .S0 (
             nx23893)) ;
    mux21_ni ix813 (.Y (nx812), .A0 (inputs_374__0), .A1 (inputs_375__0), .S0 (
             nx23895)) ;
    nand04 ix8418 (.Y (nx8417), .A0 (nx22229), .A1 (nx23367), .A2 (nx23895), .A3 (
           nx760)) ;
    mux21_ni ix761 (.Y (nx760), .A0 (inputs_355__0), .A1 (inputs_371__0), .S0 (
             nx22679)) ;
    mux21_ni ix747 (.Y (nx746), .A0 (nx682), .A1 (nx742), .S0 (nx22679)) ;
    mux21_ni ix683 (.Y (nx682), .A0 (nx650), .A1 (nx678), .S0 (nx23191)) ;
    mux21_ni ix651 (.Y (nx650), .A0 (nx634), .A1 (nx646), .S0 (nx23367)) ;
    mux21_ni ix635 (.Y (nx634), .A0 (inputs_360__0), .A1 (inputs_361__0), .S0 (
             nx23895)) ;
    mux21_ni ix647 (.Y (nx646), .A0 (inputs_362__0), .A1 (inputs_363__0), .S0 (
             nx23895)) ;
    mux21_ni ix679 (.Y (nx678), .A0 (nx662), .A1 (nx674), .S0 (nx23367)) ;
    mux21_ni ix663 (.Y (nx662), .A0 (inputs_364__0), .A1 (inputs_365__0), .S0 (
             nx23895)) ;
    mux21_ni ix675 (.Y (nx674), .A0 (inputs_366__0), .A1 (inputs_367__0), .S0 (
             nx23895)) ;
    mux21_ni ix743 (.Y (nx742), .A0 (nx710), .A1 (nx738), .S0 (nx23193)) ;
    mux21_ni ix711 (.Y (nx710), .A0 (nx694), .A1 (nx706), .S0 (nx23367)) ;
    mux21_ni ix695 (.Y (nx694), .A0 (inputs_376__0), .A1 (inputs_377__0), .S0 (
             nx23895)) ;
    mux21_ni ix707 (.Y (nx706), .A0 (inputs_378__0), .A1 (inputs_379__0), .S0 (
             nx23897)) ;
    mux21_ni ix739 (.Y (nx738), .A0 (nx722), .A1 (nx734), .S0 (nx23367)) ;
    mux21_ni ix723 (.Y (nx722), .A0 (inputs_380__0), .A1 (inputs_381__0), .S0 (
             nx23897)) ;
    mux21_ni ix735 (.Y (nx734), .A0 (inputs_382__0), .A1 (inputs_383__0), .S0 (
             nx23897)) ;
    mux21_ni ix1683 (.Y (nx1682), .A0 (nx1258), .A1 (nx1678), .S0 (nx22451)) ;
    mux21_ni ix1259 (.Y (nx1258), .A0 (nx1046), .A1 (nx1254), .S0 (nx22527)) ;
    mux21_ni ix1047 (.Y (nx1046), .A0 (nx1040), .A1 (nx962), .S0 (nx23117)) ;
    oai21 ix1041 (.Y (nx1040), .A0 (nx22229), .A1 (nx8455), .B0 (nx8467)) ;
    mux21 ix8456 (.Y (nx8455), .A0 (nx1004), .A1 (nx1032), .S0 (nx22679)) ;
    mux21_ni ix1005 (.Y (nx1004), .A0 (nx988), .A1 (nx1000), .S0 (nx23369)) ;
    mux21_ni ix989 (.Y (nx988), .A0 (inputs_388__0), .A1 (inputs_389__0), .S0 (
             nx23897)) ;
    mux21_ni ix1001 (.Y (nx1000), .A0 (inputs_390__0), .A1 (inputs_391__0), .S0 (
             nx23897)) ;
    mux21_ni ix1033 (.Y (nx1032), .A0 (nx1016), .A1 (nx1028), .S0 (nx23369)) ;
    mux21_ni ix1017 (.Y (nx1016), .A0 (inputs_404__0), .A1 (inputs_405__0), .S0 (
             nx23897)) ;
    mux21_ni ix1029 (.Y (nx1028), .A0 (inputs_406__0), .A1 (inputs_407__0), .S0 (
             nx23897)) ;
    nand04 ix8468 (.Y (nx8467), .A0 (nx22229), .A1 (nx23369), .A2 (nx23899), .A3 (
           nx976)) ;
    mux21_ni ix977 (.Y (nx976), .A0 (inputs_387__0), .A1 (inputs_403__0), .S0 (
             nx22679)) ;
    mux21_ni ix963 (.Y (nx962), .A0 (nx898), .A1 (nx958), .S0 (nx22681)) ;
    mux21_ni ix899 (.Y (nx898), .A0 (nx866), .A1 (nx894), .S0 (nx23193)) ;
    mux21_ni ix867 (.Y (nx866), .A0 (nx850), .A1 (nx862), .S0 (nx23369)) ;
    mux21_ni ix851 (.Y (nx850), .A0 (inputs_392__0), .A1 (inputs_393__0), .S0 (
             nx23899)) ;
    mux21_ni ix863 (.Y (nx862), .A0 (inputs_394__0), .A1 (inputs_395__0), .S0 (
             nx23899)) ;
    mux21_ni ix895 (.Y (nx894), .A0 (nx878), .A1 (nx890), .S0 (nx23369)) ;
    mux21_ni ix879 (.Y (nx878), .A0 (inputs_396__0), .A1 (inputs_397__0), .S0 (
             nx23899)) ;
    mux21_ni ix891 (.Y (nx890), .A0 (inputs_398__0), .A1 (inputs_399__0), .S0 (
             nx23899)) ;
    mux21_ni ix959 (.Y (nx958), .A0 (nx926), .A1 (nx954), .S0 (nx23193)) ;
    mux21_ni ix927 (.Y (nx926), .A0 (nx910), .A1 (nx922), .S0 (nx23369)) ;
    mux21_ni ix911 (.Y (nx910), .A0 (inputs_408__0), .A1 (inputs_409__0), .S0 (
             nx23899)) ;
    mux21_ni ix923 (.Y (nx922), .A0 (inputs_410__0), .A1 (inputs_411__0), .S0 (
             nx23899)) ;
    mux21_ni ix955 (.Y (nx954), .A0 (nx938), .A1 (nx950), .S0 (nx23369)) ;
    mux21_ni ix939 (.Y (nx938), .A0 (inputs_412__0), .A1 (inputs_413__0), .S0 (
             nx23901)) ;
    mux21_ni ix951 (.Y (nx950), .A0 (inputs_414__0), .A1 (inputs_415__0), .S0 (
             nx23901)) ;
    mux21_ni ix1255 (.Y (nx1254), .A0 (nx1248), .A1 (nx1170), .S0 (nx23117)) ;
    oai21 ix1249 (.Y (nx1248), .A0 (nx22229), .A1 (nx8497), .B0 (nx8511)) ;
    mux21 ix8498 (.Y (nx8497), .A0 (nx1212), .A1 (nx1240), .S0 (nx22681)) ;
    mux21_ni ix1213 (.Y (nx1212), .A0 (nx1196), .A1 (nx1208), .S0 (nx23371)) ;
    mux21_ni ix1197 (.Y (nx1196), .A0 (inputs_420__0), .A1 (inputs_421__0), .S0 (
             nx23901)) ;
    mux21_ni ix1209 (.Y (nx1208), .A0 (inputs_422__0), .A1 (inputs_423__0), .S0 (
             nx23901)) ;
    mux21_ni ix1241 (.Y (nx1240), .A0 (nx1224), .A1 (nx1236), .S0 (nx23371)) ;
    mux21_ni ix1225 (.Y (nx1224), .A0 (inputs_436__0), .A1 (inputs_437__0), .S0 (
             nx23901)) ;
    mux21_ni ix1237 (.Y (nx1236), .A0 (inputs_438__0), .A1 (inputs_439__0), .S0 (
             nx23901)) ;
    nand04 ix8512 (.Y (nx8511), .A0 (nx22229), .A1 (nx23371), .A2 (nx23901), .A3 (
           nx1184)) ;
    mux21_ni ix1185 (.Y (nx1184), .A0 (inputs_419__0), .A1 (inputs_435__0), .S0 (
             nx22681)) ;
    mux21_ni ix1171 (.Y (nx1170), .A0 (nx1106), .A1 (nx1166), .S0 (nx22681)) ;
    mux21_ni ix1107 (.Y (nx1106), .A0 (nx1074), .A1 (nx1102), .S0 (nx23193)) ;
    mux21_ni ix1075 (.Y (nx1074), .A0 (nx1058), .A1 (nx1070), .S0 (nx23371)) ;
    mux21_ni ix1059 (.Y (nx1058), .A0 (inputs_424__0), .A1 (inputs_425__0), .S0 (
             nx23903)) ;
    mux21_ni ix1071 (.Y (nx1070), .A0 (inputs_426__0), .A1 (inputs_427__0), .S0 (
             nx23903)) ;
    mux21_ni ix1103 (.Y (nx1102), .A0 (nx1086), .A1 (nx1098), .S0 (nx23371)) ;
    mux21_ni ix1087 (.Y (nx1086), .A0 (inputs_428__0), .A1 (inputs_429__0), .S0 (
             nx23903)) ;
    mux21_ni ix1099 (.Y (nx1098), .A0 (inputs_430__0), .A1 (inputs_431__0), .S0 (
             nx23903)) ;
    mux21_ni ix1167 (.Y (nx1166), .A0 (nx1134), .A1 (nx1162), .S0 (nx23193)) ;
    mux21_ni ix1135 (.Y (nx1134), .A0 (nx1118), .A1 (nx1130), .S0 (nx23371)) ;
    mux21_ni ix1119 (.Y (nx1118), .A0 (inputs_440__0), .A1 (inputs_441__0), .S0 (
             nx23903)) ;
    mux21_ni ix1131 (.Y (nx1130), .A0 (inputs_442__0), .A1 (inputs_443__0), .S0 (
             nx23903)) ;
    mux21_ni ix1163 (.Y (nx1162), .A0 (nx1146), .A1 (nx1158), .S0 (nx23371)) ;
    mux21_ni ix1147 (.Y (nx1146), .A0 (inputs_444__0), .A1 (inputs_445__0), .S0 (
             nx23903)) ;
    mux21_ni ix1159 (.Y (nx1158), .A0 (inputs_446__0), .A1 (inputs_447__0), .S0 (
             nx23905)) ;
    mux21_ni ix1679 (.Y (nx1678), .A0 (nx1466), .A1 (nx1674), .S0 (nx22527)) ;
    mux21_ni ix1467 (.Y (nx1466), .A0 (nx1460), .A1 (nx1382), .S0 (nx23117)) ;
    oai21 ix1461 (.Y (nx1460), .A0 (nx22229), .A1 (nx8541), .B0 (nx8553)) ;
    mux21 ix8542 (.Y (nx8541), .A0 (nx1424), .A1 (nx1452), .S0 (nx22681)) ;
    mux21_ni ix1425 (.Y (nx1424), .A0 (nx1408), .A1 (nx1420), .S0 (nx23373)) ;
    mux21_ni ix1409 (.Y (nx1408), .A0 (inputs_452__0), .A1 (inputs_453__0), .S0 (
             nx23905)) ;
    mux21_ni ix1421 (.Y (nx1420), .A0 (inputs_454__0), .A1 (inputs_455__0), .S0 (
             nx23905)) ;
    mux21_ni ix1453 (.Y (nx1452), .A0 (nx1436), .A1 (nx1448), .S0 (nx23373)) ;
    mux21_ni ix1437 (.Y (nx1436), .A0 (inputs_468__0), .A1 (inputs_469__0), .S0 (
             nx23905)) ;
    mux21_ni ix1449 (.Y (nx1448), .A0 (inputs_470__0), .A1 (inputs_471__0), .S0 (
             nx23905)) ;
    nand04 ix8554 (.Y (nx8553), .A0 (nx22229), .A1 (nx23373), .A2 (nx23905), .A3 (
           nx1396)) ;
    mux21_ni ix1397 (.Y (nx1396), .A0 (inputs_451__0), .A1 (inputs_467__0), .S0 (
             nx22681)) ;
    mux21_ni ix1383 (.Y (nx1382), .A0 (nx1318), .A1 (nx1378), .S0 (nx22681)) ;
    mux21_ni ix1319 (.Y (nx1318), .A0 (nx1286), .A1 (nx1314), .S0 (nx23193)) ;
    mux21_ni ix1287 (.Y (nx1286), .A0 (nx1270), .A1 (nx1282), .S0 (nx23373)) ;
    mux21_ni ix1271 (.Y (nx1270), .A0 (inputs_456__0), .A1 (inputs_457__0), .S0 (
             nx23905)) ;
    mux21_ni ix1283 (.Y (nx1282), .A0 (inputs_458__0), .A1 (inputs_459__0), .S0 (
             nx23907)) ;
    mux21_ni ix1315 (.Y (nx1314), .A0 (nx1298), .A1 (nx1310), .S0 (nx23373)) ;
    mux21_ni ix1299 (.Y (nx1298), .A0 (inputs_460__0), .A1 (inputs_461__0), .S0 (
             nx23907)) ;
    mux21_ni ix1311 (.Y (nx1310), .A0 (inputs_462__0), .A1 (inputs_463__0), .S0 (
             nx23907)) ;
    mux21_ni ix1379 (.Y (nx1378), .A0 (nx1346), .A1 (nx1374), .S0 (nx23193)) ;
    mux21_ni ix1347 (.Y (nx1346), .A0 (nx1330), .A1 (nx1342), .S0 (nx23373)) ;
    mux21_ni ix1331 (.Y (nx1330), .A0 (inputs_472__0), .A1 (inputs_473__0), .S0 (
             nx23907)) ;
    mux21_ni ix1343 (.Y (nx1342), .A0 (inputs_474__0), .A1 (inputs_475__0), .S0 (
             nx23907)) ;
    mux21_ni ix1375 (.Y (nx1374), .A0 (nx1358), .A1 (nx1370), .S0 (nx23373)) ;
    mux21_ni ix1359 (.Y (nx1358), .A0 (inputs_476__0), .A1 (inputs_477__0), .S0 (
             nx23907)) ;
    mux21_ni ix1371 (.Y (nx1370), .A0 (inputs_478__0), .A1 (inputs_479__0), .S0 (
             nx23907)) ;
    mux21_ni ix1675 (.Y (nx1674), .A0 (nx1668), .A1 (nx1590), .S0 (nx23119)) ;
    oai21 ix1669 (.Y (nx1668), .A0 (nx22231), .A1 (nx8585), .B0 (nx8597)) ;
    mux21 ix8586 (.Y (nx8585), .A0 (nx1632), .A1 (nx1660), .S0 (nx22683)) ;
    mux21_ni ix1633 (.Y (nx1632), .A0 (nx1616), .A1 (nx1628), .S0 (nx23375)) ;
    mux21_ni ix1617 (.Y (nx1616), .A0 (inputs_484__0), .A1 (inputs_485__0), .S0 (
             nx23909)) ;
    mux21_ni ix1629 (.Y (nx1628), .A0 (inputs_486__0), .A1 (inputs_487__0), .S0 (
             nx23909)) ;
    mux21_ni ix1661 (.Y (nx1660), .A0 (nx1644), .A1 (nx1656), .S0 (nx23375)) ;
    mux21_ni ix1645 (.Y (nx1644), .A0 (inputs_500__0), .A1 (inputs_501__0), .S0 (
             nx23909)) ;
    mux21_ni ix1657 (.Y (nx1656), .A0 (inputs_502__0), .A1 (inputs_503__0), .S0 (
             nx23909)) ;
    nand04 ix8598 (.Y (nx8597), .A0 (nx22231), .A1 (nx23375), .A2 (nx23909), .A3 (
           nx1604)) ;
    mux21_ni ix1605 (.Y (nx1604), .A0 (inputs_483__0), .A1 (inputs_499__0), .S0 (
             nx22683)) ;
    mux21_ni ix1591 (.Y (nx1590), .A0 (nx1526), .A1 (nx1586), .S0 (nx22683)) ;
    mux21_ni ix1527 (.Y (nx1526), .A0 (nx1494), .A1 (nx1522), .S0 (nx23195)) ;
    mux21_ni ix1495 (.Y (nx1494), .A0 (nx1478), .A1 (nx1490), .S0 (nx23375)) ;
    mux21_ni ix1479 (.Y (nx1478), .A0 (inputs_488__0), .A1 (inputs_489__0), .S0 (
             nx23909)) ;
    mux21_ni ix1491 (.Y (nx1490), .A0 (inputs_490__0), .A1 (inputs_491__0), .S0 (
             nx23909)) ;
    mux21_ni ix1523 (.Y (nx1522), .A0 (nx1506), .A1 (nx1518), .S0 (nx23375)) ;
    mux21_ni ix1507 (.Y (nx1506), .A0 (inputs_492__0), .A1 (inputs_493__0), .S0 (
             nx23911)) ;
    mux21_ni ix1519 (.Y (nx1518), .A0 (inputs_494__0), .A1 (inputs_495__0), .S0 (
             nx23911)) ;
    mux21_ni ix1587 (.Y (nx1586), .A0 (nx1554), .A1 (nx1582), .S0 (nx23195)) ;
    mux21_ni ix1555 (.Y (nx1554), .A0 (nx1538), .A1 (nx1550), .S0 (nx23375)) ;
    mux21_ni ix1539 (.Y (nx1538), .A0 (inputs_504__0), .A1 (inputs_505__0), .S0 (
             nx23911)) ;
    mux21_ni ix1551 (.Y (nx1550), .A0 (inputs_506__0), .A1 (inputs_507__0), .S0 (
             nx23911)) ;
    mux21_ni ix1583 (.Y (nx1582), .A0 (nx1566), .A1 (nx1578), .S0 (nx23375)) ;
    mux21_ni ix1567 (.Y (nx1566), .A0 (inputs_508__0), .A1 (inputs_509__0), .S0 (
             nx23911)) ;
    mux21_ni ix1579 (.Y (nx1578), .A0 (inputs_510__0), .A1 (inputs_511__0), .S0 (
             nx23911)) ;
    aoi32 ix8626 (.Y (nx8625), .A0 (nx2452), .A1 (nx22385), .A2 (nx22231), .B0 (
          nx24851), .B1 (nx4148)) ;
    oai21 ix2453 (.Y (nx2452), .A0 (nx23377), .A1 (nx8629), .B0 (nx8735)) ;
    mux21 ix8630 (.Y (nx8629), .A0 (nx2190), .A1 (nx2442), .S0 (nx23911)) ;
    mux21_ni ix2191 (.Y (nx2190), .A0 (nx2062), .A1 (nx2186), .S0 (nx22393)) ;
    mux21_ni ix2063 (.Y (nx2062), .A0 (nx1998), .A1 (nx2058), .S0 (nx22411)) ;
    mux21_ni ix1999 (.Y (nx1998), .A0 (nx1966), .A1 (nx1994), .S0 (nx22451)) ;
    mux21_ni ix1967 (.Y (nx1966), .A0 (nx1950), .A1 (nx1962), .S0 (nx22527)) ;
    mux21_ni ix1951 (.Y (nx1950), .A0 (inputs_0__0), .A1 (inputs_16__0), .S0 (
             nx22683)) ;
    mux21_ni ix1963 (.Y (nx1962), .A0 (inputs_32__0), .A1 (inputs_48__0), .S0 (
             nx22683)) ;
    mux21_ni ix1995 (.Y (nx1994), .A0 (nx1978), .A1 (nx1990), .S0 (nx22527)) ;
    mux21_ni ix1979 (.Y (nx1978), .A0 (inputs_64__0), .A1 (inputs_80__0), .S0 (
             nx22683)) ;
    mux21_ni ix1991 (.Y (nx1990), .A0 (inputs_96__0), .A1 (inputs_112__0), .S0 (
             nx22683)) ;
    mux21_ni ix2059 (.Y (nx2058), .A0 (nx2026), .A1 (nx2054), .S0 (nx22451)) ;
    mux21_ni ix2027 (.Y (nx2026), .A0 (nx2010), .A1 (nx2022), .S0 (nx22527)) ;
    mux21_ni ix2011 (.Y (nx2010), .A0 (inputs_128__0), .A1 (inputs_144__0), .S0 (
             nx22685)) ;
    mux21_ni ix2023 (.Y (nx2022), .A0 (inputs_160__0), .A1 (inputs_176__0), .S0 (
             nx22685)) ;
    mux21_ni ix2055 (.Y (nx2054), .A0 (nx2038), .A1 (nx2050), .S0 (nx22529)) ;
    mux21_ni ix2039 (.Y (nx2038), .A0 (inputs_192__0), .A1 (inputs_208__0), .S0 (
             nx22685)) ;
    mux21_ni ix2051 (.Y (nx2050), .A0 (inputs_224__0), .A1 (inputs_240__0), .S0 (
             nx22685)) ;
    mux21_ni ix2187 (.Y (nx2186), .A0 (nx2122), .A1 (nx2182), .S0 (nx22411)) ;
    mux21_ni ix2123 (.Y (nx2122), .A0 (nx2090), .A1 (nx2118), .S0 (nx22451)) ;
    mux21_ni ix2091 (.Y (nx2090), .A0 (nx2074), .A1 (nx2086), .S0 (nx22529)) ;
    mux21_ni ix2075 (.Y (nx2074), .A0 (inputs_256__0), .A1 (inputs_272__0), .S0 (
             nx22685)) ;
    mux21_ni ix2087 (.Y (nx2086), .A0 (inputs_288__0), .A1 (inputs_304__0), .S0 (
             nx22685)) ;
    mux21_ni ix2119 (.Y (nx2118), .A0 (nx2102), .A1 (nx2114), .S0 (nx22529)) ;
    mux21_ni ix2103 (.Y (nx2102), .A0 (inputs_320__0), .A1 (inputs_336__0), .S0 (
             nx22685)) ;
    mux21_ni ix2115 (.Y (nx2114), .A0 (inputs_352__0), .A1 (inputs_368__0), .S0 (
             nx22687)) ;
    mux21_ni ix2183 (.Y (nx2182), .A0 (nx2150), .A1 (nx2178), .S0 (nx22451)) ;
    mux21_ni ix2151 (.Y (nx2150), .A0 (nx2134), .A1 (nx2146), .S0 (nx22529)) ;
    mux21_ni ix2135 (.Y (nx2134), .A0 (inputs_384__0), .A1 (inputs_400__0), .S0 (
             nx22687)) ;
    mux21_ni ix2147 (.Y (nx2146), .A0 (inputs_416__0), .A1 (inputs_432__0), .S0 (
             nx22687)) ;
    mux21_ni ix2179 (.Y (nx2178), .A0 (nx2162), .A1 (nx2174), .S0 (nx22529)) ;
    mux21_ni ix2163 (.Y (nx2162), .A0 (inputs_448__0), .A1 (inputs_464__0), .S0 (
             nx22687)) ;
    mux21_ni ix2175 (.Y (nx2174), .A0 (inputs_480__0), .A1 (inputs_496__0), .S0 (
             nx22687)) ;
    mux21_ni ix2443 (.Y (nx2442), .A0 (nx2314), .A1 (nx2438), .S0 (nx22393)) ;
    mux21_ni ix2315 (.Y (nx2314), .A0 (nx2250), .A1 (nx2310), .S0 (nx22411)) ;
    mux21_ni ix2251 (.Y (nx2250), .A0 (nx2218), .A1 (nx2246), .S0 (nx22451)) ;
    mux21_ni ix2219 (.Y (nx2218), .A0 (nx2202), .A1 (nx2214), .S0 (nx22529)) ;
    mux21_ni ix2203 (.Y (nx2202), .A0 (inputs_1__0), .A1 (inputs_17__0), .S0 (
             nx22687)) ;
    mux21_ni ix2215 (.Y (nx2214), .A0 (inputs_33__0), .A1 (inputs_49__0), .S0 (
             nx22687)) ;
    mux21_ni ix2247 (.Y (nx2246), .A0 (nx2230), .A1 (nx2242), .S0 (nx22529)) ;
    mux21_ni ix2231 (.Y (nx2230), .A0 (inputs_65__0), .A1 (inputs_81__0), .S0 (
             nx22689)) ;
    mux21_ni ix2243 (.Y (nx2242), .A0 (inputs_97__0), .A1 (inputs_113__0), .S0 (
             nx22689)) ;
    mux21_ni ix2311 (.Y (nx2310), .A0 (nx2278), .A1 (nx2306), .S0 (nx22453)) ;
    mux21_ni ix2279 (.Y (nx2278), .A0 (nx2262), .A1 (nx2274), .S0 (nx22531)) ;
    mux21_ni ix2263 (.Y (nx2262), .A0 (inputs_129__0), .A1 (inputs_145__0), .S0 (
             nx22689)) ;
    mux21_ni ix2275 (.Y (nx2274), .A0 (inputs_161__0), .A1 (inputs_177__0), .S0 (
             nx22689)) ;
    mux21_ni ix2307 (.Y (nx2306), .A0 (nx2290), .A1 (nx2302), .S0 (nx22531)) ;
    mux21_ni ix2291 (.Y (nx2290), .A0 (inputs_193__0), .A1 (inputs_209__0), .S0 (
             nx22689)) ;
    mux21_ni ix2303 (.Y (nx2302), .A0 (inputs_225__0), .A1 (inputs_241__0), .S0 (
             nx22689)) ;
    mux21_ni ix2439 (.Y (nx2438), .A0 (nx2374), .A1 (nx2434), .S0 (nx22411)) ;
    mux21_ni ix2375 (.Y (nx2374), .A0 (nx2342), .A1 (nx2370), .S0 (nx22453)) ;
    mux21_ni ix2343 (.Y (nx2342), .A0 (nx2326), .A1 (nx2338), .S0 (nx22531)) ;
    mux21_ni ix2327 (.Y (nx2326), .A0 (inputs_257__0), .A1 (inputs_273__0), .S0 (
             nx22689)) ;
    mux21_ni ix2339 (.Y (nx2338), .A0 (inputs_289__0), .A1 (inputs_305__0), .S0 (
             nx22691)) ;
    mux21_ni ix2371 (.Y (nx2370), .A0 (nx2354), .A1 (nx2366), .S0 (nx22531)) ;
    mux21_ni ix2355 (.Y (nx2354), .A0 (inputs_321__0), .A1 (inputs_337__0), .S0 (
             nx22691)) ;
    mux21_ni ix2367 (.Y (nx2366), .A0 (inputs_353__0), .A1 (inputs_369__0), .S0 (
             nx22691)) ;
    mux21_ni ix2435 (.Y (nx2434), .A0 (nx2402), .A1 (nx2430), .S0 (nx22453)) ;
    mux21_ni ix2403 (.Y (nx2402), .A0 (nx2386), .A1 (nx2398), .S0 (nx22531)) ;
    mux21_ni ix2387 (.Y (nx2386), .A0 (inputs_385__0), .A1 (inputs_401__0), .S0 (
             nx22691)) ;
    mux21_ni ix2399 (.Y (nx2398), .A0 (inputs_417__0), .A1 (inputs_433__0), .S0 (
             nx22691)) ;
    mux21_ni ix2431 (.Y (nx2430), .A0 (nx2414), .A1 (nx2426), .S0 (nx22531)) ;
    mux21_ni ix2415 (.Y (nx2414), .A0 (inputs_449__0), .A1 (inputs_465__0), .S0 (
             nx22691)) ;
    mux21_ni ix2427 (.Y (nx2426), .A0 (inputs_481__0), .A1 (inputs_497__0), .S0 (
             nx22691)) ;
    nand03 ix8736 (.Y (nx8735), .A0 (nx1936), .A1 (nx23377), .A2 (nx24879)) ;
    mux21_ni ix1937 (.Y (nx1936), .A0 (nx1808), .A1 (nx1932), .S0 (nx22393)) ;
    mux21_ni ix1809 (.Y (nx1808), .A0 (nx1744), .A1 (nx1804), .S0 (nx22411)) ;
    mux21_ni ix1745 (.Y (nx1744), .A0 (nx1712), .A1 (nx1740), .S0 (nx22453)) ;
    mux21_ni ix1713 (.Y (nx1712), .A0 (nx1696), .A1 (nx1708), .S0 (nx22531)) ;
    mux21_ni ix1697 (.Y (nx1696), .A0 (inputs_2__0), .A1 (inputs_18__0), .S0 (
             nx22693)) ;
    mux21_ni ix1709 (.Y (nx1708), .A0 (inputs_34__0), .A1 (inputs_50__0), .S0 (
             nx22693)) ;
    mux21_ni ix1741 (.Y (nx1740), .A0 (nx1724), .A1 (nx1736), .S0 (nx22533)) ;
    mux21_ni ix1725 (.Y (nx1724), .A0 (inputs_66__0), .A1 (inputs_82__0), .S0 (
             nx22693)) ;
    mux21_ni ix1737 (.Y (nx1736), .A0 (inputs_98__0), .A1 (inputs_114__0), .S0 (
             nx22693)) ;
    mux21_ni ix1805 (.Y (nx1804), .A0 (nx1772), .A1 (nx1800), .S0 (nx22453)) ;
    mux21_ni ix1773 (.Y (nx1772), .A0 (nx1756), .A1 (nx1768), .S0 (nx22533)) ;
    mux21_ni ix1757 (.Y (nx1756), .A0 (inputs_130__0), .A1 (inputs_146__0), .S0 (
             nx22693)) ;
    mux21_ni ix1769 (.Y (nx1768), .A0 (inputs_162__0), .A1 (inputs_178__0), .S0 (
             nx22693)) ;
    mux21_ni ix1801 (.Y (nx1800), .A0 (nx1784), .A1 (nx1796), .S0 (nx22533)) ;
    mux21_ni ix1785 (.Y (nx1784), .A0 (inputs_194__0), .A1 (inputs_210__0), .S0 (
             nx22693)) ;
    mux21_ni ix1797 (.Y (nx1796), .A0 (inputs_226__0), .A1 (inputs_242__0), .S0 (
             nx22695)) ;
    mux21_ni ix1933 (.Y (nx1932), .A0 (nx1868), .A1 (nx1928), .S0 (nx22411)) ;
    mux21_ni ix1869 (.Y (nx1868), .A0 (nx1836), .A1 (nx1864), .S0 (nx22453)) ;
    mux21_ni ix1837 (.Y (nx1836), .A0 (nx1820), .A1 (nx1832), .S0 (nx22533)) ;
    mux21_ni ix1821 (.Y (nx1820), .A0 (inputs_258__0), .A1 (inputs_274__0), .S0 (
             nx22695)) ;
    mux21_ni ix1833 (.Y (nx1832), .A0 (inputs_290__0), .A1 (inputs_306__0), .S0 (
             nx22695)) ;
    mux21_ni ix1865 (.Y (nx1864), .A0 (nx1848), .A1 (nx1860), .S0 (nx22533)) ;
    mux21_ni ix1849 (.Y (nx1848), .A0 (inputs_322__0), .A1 (inputs_338__0), .S0 (
             nx22695)) ;
    mux21_ni ix1861 (.Y (nx1860), .A0 (inputs_354__0), .A1 (inputs_370__0), .S0 (
             nx22695)) ;
    mux21_ni ix1929 (.Y (nx1928), .A0 (nx1896), .A1 (nx1924), .S0 (nx22453)) ;
    mux21_ni ix1897 (.Y (nx1896), .A0 (nx1880), .A1 (nx1892), .S0 (nx22533)) ;
    mux21_ni ix1881 (.Y (nx1880), .A0 (inputs_386__0), .A1 (inputs_402__0), .S0 (
             nx22695)) ;
    mux21_ni ix1893 (.Y (nx1892), .A0 (inputs_418__0), .A1 (inputs_434__0), .S0 (
             nx22695)) ;
    mux21_ni ix1925 (.Y (nx1924), .A0 (nx1908), .A1 (nx1920), .S0 (nx22533)) ;
    mux21_ni ix1909 (.Y (nx1908), .A0 (inputs_450__0), .A1 (inputs_466__0), .S0 (
             nx22697)) ;
    mux21_ni ix1921 (.Y (nx1920), .A0 (inputs_482__0), .A1 (inputs_498__0), .S0 (
             nx22697)) ;
    mux21_ni ix4149 (.Y (nx4148), .A0 (nx3300), .A1 (nx4144), .S0 (nx22413)) ;
    mux21_ni ix3301 (.Y (nx3300), .A0 (nx2876), .A1 (nx3296), .S0 (nx22455)) ;
    mux21_ni ix2877 (.Y (nx2876), .A0 (nx2664), .A1 (nx2872), .S0 (nx22535)) ;
    mux21_ni ix2665 (.Y (nx2664), .A0 (nx2658), .A1 (nx2580), .S0 (nx23119)) ;
    oai21 ix2659 (.Y (nx2658), .A0 (nx22231), .A1 (nx8797), .B0 (nx8809)) ;
    mux21 ix8798 (.Y (nx8797), .A0 (nx2622), .A1 (nx2650), .S0 (nx22697)) ;
    mux21_ni ix2623 (.Y (nx2622), .A0 (nx2606), .A1 (nx2618), .S0 (nx23377)) ;
    mux21_ni ix2607 (.Y (nx2606), .A0 (inputs_4__0), .A1 (inputs_5__0), .S0 (
             nx23913)) ;
    mux21_ni ix2619 (.Y (nx2618), .A0 (inputs_6__0), .A1 (inputs_7__0), .S0 (
             nx23913)) ;
    mux21_ni ix2651 (.Y (nx2650), .A0 (nx2634), .A1 (nx2646), .S0 (nx23377)) ;
    mux21_ni ix2635 (.Y (nx2634), .A0 (inputs_20__0), .A1 (inputs_21__0), .S0 (
             nx23913)) ;
    mux21_ni ix2647 (.Y (nx2646), .A0 (inputs_22__0), .A1 (inputs_23__0), .S0 (
             nx23913)) ;
    nand04 ix8810 (.Y (nx8809), .A0 (nx22231), .A1 (nx23377), .A2 (nx23913), .A3 (
           nx2594)) ;
    mux21_ni ix2595 (.Y (nx2594), .A0 (inputs_3__0), .A1 (inputs_19__0), .S0 (
             nx22697)) ;
    mux21_ni ix2581 (.Y (nx2580), .A0 (nx2516), .A1 (nx2576), .S0 (nx22697)) ;
    mux21_ni ix2517 (.Y (nx2516), .A0 (nx2484), .A1 (nx2512), .S0 (nx23195)) ;
    mux21_ni ix2485 (.Y (nx2484), .A0 (nx2468), .A1 (nx2480), .S0 (nx23377)) ;
    mux21_ni ix2469 (.Y (nx2468), .A0 (inputs_8__0), .A1 (inputs_9__0), .S0 (
             nx23913)) ;
    mux21_ni ix2481 (.Y (nx2480), .A0 (inputs_10__0), .A1 (inputs_11__0), .S0 (
             nx23913)) ;
    mux21_ni ix2513 (.Y (nx2512), .A0 (nx2496), .A1 (nx2508), .S0 (nx23377)) ;
    mux21_ni ix2497 (.Y (nx2496), .A0 (inputs_12__0), .A1 (inputs_13__0), .S0 (
             nx23915)) ;
    mux21_ni ix2509 (.Y (nx2508), .A0 (inputs_14__0), .A1 (inputs_15__0), .S0 (
             nx23915)) ;
    mux21_ni ix2577 (.Y (nx2576), .A0 (nx2544), .A1 (nx2572), .S0 (nx23195)) ;
    mux21_ni ix2545 (.Y (nx2544), .A0 (nx2528), .A1 (nx2540), .S0 (nx23379)) ;
    mux21_ni ix2529 (.Y (nx2528), .A0 (inputs_24__0), .A1 (inputs_25__0), .S0 (
             nx23915)) ;
    mux21_ni ix2541 (.Y (nx2540), .A0 (inputs_26__0), .A1 (inputs_27__0), .S0 (
             nx23915)) ;
    mux21_ni ix2573 (.Y (nx2572), .A0 (nx2556), .A1 (nx2568), .S0 (nx23379)) ;
    mux21_ni ix2557 (.Y (nx2556), .A0 (inputs_28__0), .A1 (inputs_29__0), .S0 (
             nx23915)) ;
    mux21_ni ix2569 (.Y (nx2568), .A0 (inputs_30__0), .A1 (inputs_31__0), .S0 (
             nx23915)) ;
    mux21_ni ix2873 (.Y (nx2872), .A0 (nx2866), .A1 (nx2788), .S0 (nx23119)) ;
    oai21 ix2867 (.Y (nx2866), .A0 (nx22231), .A1 (nx8839), .B0 (nx8853)) ;
    mux21 ix8840 (.Y (nx8839), .A0 (nx2830), .A1 (nx2858), .S0 (nx22697)) ;
    mux21_ni ix2831 (.Y (nx2830), .A0 (nx2814), .A1 (nx2826), .S0 (nx23379)) ;
    mux21_ni ix2815 (.Y (nx2814), .A0 (inputs_36__0), .A1 (inputs_37__0), .S0 (
             nx23915)) ;
    mux21_ni ix2827 (.Y (nx2826), .A0 (inputs_38__0), .A1 (inputs_39__0), .S0 (
             nx23917)) ;
    mux21_ni ix2859 (.Y (nx2858), .A0 (nx2842), .A1 (nx2854), .S0 (nx23379)) ;
    mux21_ni ix2843 (.Y (nx2842), .A0 (inputs_52__0), .A1 (inputs_53__0), .S0 (
             nx23917)) ;
    mux21_ni ix2855 (.Y (nx2854), .A0 (inputs_54__0), .A1 (inputs_55__0), .S0 (
             nx23917)) ;
    nand04 ix8854 (.Y (nx8853), .A0 (nx22231), .A1 (nx23379), .A2 (nx23917), .A3 (
           nx2802)) ;
    mux21_ni ix2803 (.Y (nx2802), .A0 (inputs_35__0), .A1 (inputs_51__0), .S0 (
             nx22697)) ;
    mux21_ni ix2789 (.Y (nx2788), .A0 (nx2724), .A1 (nx2784), .S0 (nx22699)) ;
    mux21_ni ix2725 (.Y (nx2724), .A0 (nx2692), .A1 (nx2720), .S0 (nx23195)) ;
    mux21_ni ix2693 (.Y (nx2692), .A0 (nx2676), .A1 (nx2688), .S0 (nx23379)) ;
    mux21_ni ix2677 (.Y (nx2676), .A0 (inputs_40__0), .A1 (inputs_41__0), .S0 (
             nx23917)) ;
    mux21_ni ix2689 (.Y (nx2688), .A0 (inputs_42__0), .A1 (inputs_43__0), .S0 (
             nx23917)) ;
    mux21_ni ix2721 (.Y (nx2720), .A0 (nx2704), .A1 (nx2716), .S0 (nx23379)) ;
    mux21_ni ix2705 (.Y (nx2704), .A0 (inputs_44__0), .A1 (inputs_45__0), .S0 (
             nx23917)) ;
    mux21_ni ix2717 (.Y (nx2716), .A0 (inputs_46__0), .A1 (inputs_47__0), .S0 (
             nx23919)) ;
    mux21_ni ix2785 (.Y (nx2784), .A0 (nx2752), .A1 (nx2780), .S0 (nx23195)) ;
    mux21_ni ix2753 (.Y (nx2752), .A0 (nx2736), .A1 (nx2748), .S0 (nx23381)) ;
    mux21_ni ix2737 (.Y (nx2736), .A0 (inputs_56__0), .A1 (inputs_57__0), .S0 (
             nx23919)) ;
    mux21_ni ix2749 (.Y (nx2748), .A0 (inputs_58__0), .A1 (inputs_59__0), .S0 (
             nx23919)) ;
    mux21_ni ix2781 (.Y (nx2780), .A0 (nx2764), .A1 (nx2776), .S0 (nx23381)) ;
    mux21_ni ix2765 (.Y (nx2764), .A0 (inputs_60__0), .A1 (inputs_61__0), .S0 (
             nx23919)) ;
    mux21_ni ix2777 (.Y (nx2776), .A0 (inputs_62__0), .A1 (inputs_63__0), .S0 (
             nx23919)) ;
    mux21_ni ix3297 (.Y (nx3296), .A0 (nx3084), .A1 (nx3292), .S0 (nx22535)) ;
    mux21_ni ix3085 (.Y (nx3084), .A0 (nx3078), .A1 (nx3000), .S0 (nx23119)) ;
    oai21 ix3079 (.Y (nx3078), .A0 (nx22233), .A1 (nx8885), .B0 (nx8897)) ;
    mux21 ix8886 (.Y (nx8885), .A0 (nx3042), .A1 (nx3070), .S0 (nx22699)) ;
    mux21_ni ix3043 (.Y (nx3042), .A0 (nx3026), .A1 (nx3038), .S0 (nx23381)) ;
    mux21_ni ix3027 (.Y (nx3026), .A0 (inputs_68__0), .A1 (inputs_69__0), .S0 (
             nx23919)) ;
    mux21_ni ix3039 (.Y (nx3038), .A0 (inputs_70__0), .A1 (inputs_71__0), .S0 (
             nx23919)) ;
    mux21_ni ix3071 (.Y (nx3070), .A0 (nx3054), .A1 (nx3066), .S0 (nx23381)) ;
    mux21_ni ix3055 (.Y (nx3054), .A0 (inputs_84__0), .A1 (inputs_85__0), .S0 (
             nx23921)) ;
    mux21_ni ix3067 (.Y (nx3066), .A0 (inputs_86__0), .A1 (inputs_87__0), .S0 (
             nx23921)) ;
    nand04 ix8898 (.Y (nx8897), .A0 (nx22233), .A1 (nx23381), .A2 (nx23921), .A3 (
           nx3014)) ;
    mux21_ni ix3015 (.Y (nx3014), .A0 (inputs_67__0), .A1 (inputs_83__0), .S0 (
             nx22699)) ;
    mux21_ni ix3001 (.Y (nx3000), .A0 (nx2936), .A1 (nx2996), .S0 (nx22699)) ;
    mux21_ni ix2937 (.Y (nx2936), .A0 (nx2904), .A1 (nx2932), .S0 (nx23195)) ;
    mux21_ni ix2905 (.Y (nx2904), .A0 (nx2888), .A1 (nx2900), .S0 (nx23381)) ;
    mux21_ni ix2889 (.Y (nx2888), .A0 (inputs_72__0), .A1 (inputs_73__0), .S0 (
             nx23921)) ;
    mux21_ni ix2901 (.Y (nx2900), .A0 (inputs_74__0), .A1 (inputs_75__0), .S0 (
             nx23921)) ;
    mux21_ni ix2933 (.Y (nx2932), .A0 (nx2916), .A1 (nx2928), .S0 (nx23381)) ;
    mux21_ni ix2917 (.Y (nx2916), .A0 (inputs_76__0), .A1 (inputs_77__0), .S0 (
             nx23921)) ;
    mux21_ni ix2929 (.Y (nx2928), .A0 (inputs_78__0), .A1 (inputs_79__0), .S0 (
             nx23921)) ;
    mux21_ni ix2997 (.Y (nx2996), .A0 (nx2964), .A1 (nx2992), .S0 (nx23197)) ;
    mux21_ni ix2965 (.Y (nx2964), .A0 (nx2948), .A1 (nx2960), .S0 (nx23383)) ;
    mux21_ni ix2949 (.Y (nx2948), .A0 (inputs_88__0), .A1 (inputs_89__0), .S0 (
             nx23923)) ;
    mux21_ni ix2961 (.Y (nx2960), .A0 (inputs_90__0), .A1 (inputs_91__0), .S0 (
             nx23923)) ;
    mux21_ni ix2993 (.Y (nx2992), .A0 (nx2976), .A1 (nx2988), .S0 (nx23383)) ;
    mux21_ni ix2977 (.Y (nx2976), .A0 (inputs_92__0), .A1 (inputs_93__0), .S0 (
             nx23923)) ;
    mux21_ni ix2989 (.Y (nx2988), .A0 (inputs_94__0), .A1 (inputs_95__0), .S0 (
             nx23923)) ;
    mux21_ni ix3293 (.Y (nx3292), .A0 (nx3286), .A1 (nx3208), .S0 (nx23119)) ;
    oai21 ix3287 (.Y (nx3286), .A0 (nx22233), .A1 (nx8927), .B0 (nx8939)) ;
    mux21 ix8928 (.Y (nx8927), .A0 (nx3250), .A1 (nx3278), .S0 (nx22699)) ;
    mux21_ni ix3251 (.Y (nx3250), .A0 (nx3234), .A1 (nx3246), .S0 (nx23383)) ;
    mux21_ni ix3235 (.Y (nx3234), .A0 (inputs_100__0), .A1 (inputs_101__0), .S0 (
             nx23923)) ;
    mux21_ni ix3247 (.Y (nx3246), .A0 (inputs_102__0), .A1 (inputs_103__0), .S0 (
             nx23923)) ;
    mux21_ni ix3279 (.Y (nx3278), .A0 (nx3262), .A1 (nx3274), .S0 (nx23383)) ;
    mux21_ni ix3263 (.Y (nx3262), .A0 (inputs_116__0), .A1 (inputs_117__0), .S0 (
             nx23923)) ;
    mux21_ni ix3275 (.Y (nx3274), .A0 (inputs_118__0), .A1 (inputs_119__0), .S0 (
             nx23925)) ;
    nand04 ix8940 (.Y (nx8939), .A0 (nx22233), .A1 (nx23383), .A2 (nx23925), .A3 (
           nx3222)) ;
    mux21_ni ix3223 (.Y (nx3222), .A0 (inputs_99__0), .A1 (inputs_115__0), .S0 (
             nx22699)) ;
    mux21_ni ix3209 (.Y (nx3208), .A0 (nx3144), .A1 (nx3204), .S0 (nx22699)) ;
    mux21_ni ix3145 (.Y (nx3144), .A0 (nx3112), .A1 (nx3140), .S0 (nx23197)) ;
    mux21_ni ix3113 (.Y (nx3112), .A0 (nx3096), .A1 (nx3108), .S0 (nx23383)) ;
    mux21_ni ix3097 (.Y (nx3096), .A0 (inputs_104__0), .A1 (inputs_105__0), .S0 (
             nx23925)) ;
    mux21_ni ix3109 (.Y (nx3108), .A0 (inputs_106__0), .A1 (inputs_107__0), .S0 (
             nx23925)) ;
    mux21_ni ix3141 (.Y (nx3140), .A0 (nx3124), .A1 (nx3136), .S0 (nx23383)) ;
    mux21_ni ix3125 (.Y (nx3124), .A0 (inputs_108__0), .A1 (inputs_109__0), .S0 (
             nx23925)) ;
    mux21_ni ix3137 (.Y (nx3136), .A0 (inputs_110__0), .A1 (inputs_111__0), .S0 (
             nx23925)) ;
    mux21_ni ix3205 (.Y (nx3204), .A0 (nx3172), .A1 (nx3200), .S0 (nx23197)) ;
    mux21_ni ix3173 (.Y (nx3172), .A0 (nx3156), .A1 (nx3168), .S0 (nx23385)) ;
    mux21_ni ix3157 (.Y (nx3156), .A0 (inputs_120__0), .A1 (inputs_121__0), .S0 (
             nx23925)) ;
    mux21_ni ix3169 (.Y (nx3168), .A0 (inputs_122__0), .A1 (inputs_123__0), .S0 (
             nx23927)) ;
    mux21_ni ix3201 (.Y (nx3200), .A0 (nx3184), .A1 (nx3196), .S0 (nx23385)) ;
    mux21_ni ix3185 (.Y (nx3184), .A0 (inputs_124__0), .A1 (inputs_125__0), .S0 (
             nx23927)) ;
    mux21_ni ix3197 (.Y (nx3196), .A0 (inputs_126__0), .A1 (inputs_127__0), .S0 (
             nx23927)) ;
    mux21_ni ix4145 (.Y (nx4144), .A0 (nx3720), .A1 (nx4140), .S0 (nx22455)) ;
    mux21_ni ix3721 (.Y (nx3720), .A0 (nx3508), .A1 (nx3716), .S0 (nx22535)) ;
    mux21_ni ix3509 (.Y (nx3508), .A0 (nx3502), .A1 (nx3424), .S0 (nx23119)) ;
    oai21 ix3503 (.Y (nx3502), .A0 (nx22233), .A1 (nx8971), .B0 (nx8983)) ;
    mux21 ix8972 (.Y (nx8971), .A0 (nx3466), .A1 (nx3494), .S0 (nx22701)) ;
    mux21_ni ix3467 (.Y (nx3466), .A0 (nx3450), .A1 (nx3462), .S0 (nx23385)) ;
    mux21_ni ix3451 (.Y (nx3450), .A0 (inputs_132__0), .A1 (inputs_133__0), .S0 (
             nx23927)) ;
    mux21_ni ix3463 (.Y (nx3462), .A0 (inputs_134__0), .A1 (inputs_135__0), .S0 (
             nx23927)) ;
    mux21_ni ix3495 (.Y (nx3494), .A0 (nx3478), .A1 (nx3490), .S0 (nx23385)) ;
    mux21_ni ix3479 (.Y (nx3478), .A0 (inputs_148__0), .A1 (inputs_149__0), .S0 (
             nx23927)) ;
    mux21_ni ix3491 (.Y (nx3490), .A0 (inputs_150__0), .A1 (inputs_151__0), .S0 (
             nx23927)) ;
    nand04 ix8984 (.Y (nx8983), .A0 (nx22233), .A1 (nx23385), .A2 (nx23929), .A3 (
           nx3438)) ;
    mux21_ni ix3439 (.Y (nx3438), .A0 (inputs_131__0), .A1 (inputs_147__0), .S0 (
             nx22701)) ;
    mux21_ni ix3425 (.Y (nx3424), .A0 (nx3360), .A1 (nx3420), .S0 (nx22701)) ;
    mux21_ni ix3361 (.Y (nx3360), .A0 (nx3328), .A1 (nx3356), .S0 (nx23197)) ;
    mux21_ni ix3329 (.Y (nx3328), .A0 (nx3312), .A1 (nx3324), .S0 (nx23385)) ;
    mux21_ni ix3313 (.Y (nx3312), .A0 (inputs_136__0), .A1 (inputs_137__0), .S0 (
             nx23929)) ;
    mux21_ni ix3325 (.Y (nx3324), .A0 (inputs_138__0), .A1 (inputs_139__0), .S0 (
             nx23929)) ;
    mux21_ni ix3357 (.Y (nx3356), .A0 (nx3340), .A1 (nx3352), .S0 (nx23385)) ;
    mux21_ni ix3341 (.Y (nx3340), .A0 (inputs_140__0), .A1 (inputs_141__0), .S0 (
             nx23929)) ;
    mux21_ni ix3353 (.Y (nx3352), .A0 (inputs_142__0), .A1 (inputs_143__0), .S0 (
             nx23929)) ;
    mux21_ni ix3421 (.Y (nx3420), .A0 (nx3388), .A1 (nx3416), .S0 (nx23197)) ;
    mux21_ni ix3389 (.Y (nx3388), .A0 (nx3372), .A1 (nx3384), .S0 (nx23387)) ;
    mux21_ni ix3373 (.Y (nx3372), .A0 (inputs_152__0), .A1 (inputs_153__0), .S0 (
             nx23929)) ;
    mux21_ni ix3385 (.Y (nx3384), .A0 (inputs_154__0), .A1 (inputs_155__0), .S0 (
             nx23929)) ;
    mux21_ni ix3417 (.Y (nx3416), .A0 (nx3400), .A1 (nx3412), .S0 (nx23387)) ;
    mux21_ni ix3401 (.Y (nx3400), .A0 (inputs_156__0), .A1 (inputs_157__0), .S0 (
             nx23931)) ;
    mux21_ni ix3413 (.Y (nx3412), .A0 (inputs_158__0), .A1 (inputs_159__0), .S0 (
             nx23931)) ;
    mux21_ni ix3717 (.Y (nx3716), .A0 (nx3710), .A1 (nx3632), .S0 (nx23119)) ;
    oai21 ix3711 (.Y (nx3710), .A0 (nx22233), .A1 (nx9015), .B0 (nx9027)) ;
    mux21 ix9016 (.Y (nx9015), .A0 (nx3674), .A1 (nx3702), .S0 (nx22701)) ;
    mux21_ni ix3675 (.Y (nx3674), .A0 (nx3658), .A1 (nx3670), .S0 (nx23387)) ;
    mux21_ni ix3659 (.Y (nx3658), .A0 (inputs_164__0), .A1 (inputs_165__0), .S0 (
             nx23931)) ;
    mux21_ni ix3671 (.Y (nx3670), .A0 (inputs_166__0), .A1 (inputs_167__0), .S0 (
             nx23931)) ;
    mux21_ni ix3703 (.Y (nx3702), .A0 (nx3686), .A1 (nx3698), .S0 (nx23387)) ;
    mux21_ni ix3687 (.Y (nx3686), .A0 (inputs_180__0), .A1 (inputs_181__0), .S0 (
             nx23931)) ;
    mux21_ni ix3699 (.Y (nx3698), .A0 (inputs_182__0), .A1 (inputs_183__0), .S0 (
             nx23931)) ;
    nand04 ix9028 (.Y (nx9027), .A0 (nx22235), .A1 (nx23387), .A2 (nx23931), .A3 (
           nx3646)) ;
    mux21_ni ix3647 (.Y (nx3646), .A0 (inputs_163__0), .A1 (inputs_179__0), .S0 (
             nx22701)) ;
    mux21_ni ix3633 (.Y (nx3632), .A0 (nx3568), .A1 (nx3628), .S0 (nx22701)) ;
    mux21_ni ix3569 (.Y (nx3568), .A0 (nx3536), .A1 (nx3564), .S0 (nx23197)) ;
    mux21_ni ix3537 (.Y (nx3536), .A0 (nx3520), .A1 (nx3532), .S0 (nx23387)) ;
    mux21_ni ix3521 (.Y (nx3520), .A0 (inputs_168__0), .A1 (inputs_169__0), .S0 (
             nx23933)) ;
    mux21_ni ix3533 (.Y (nx3532), .A0 (inputs_170__0), .A1 (inputs_171__0), .S0 (
             nx23933)) ;
    mux21_ni ix3565 (.Y (nx3564), .A0 (nx3548), .A1 (nx3560), .S0 (nx23387)) ;
    mux21_ni ix3549 (.Y (nx3548), .A0 (inputs_172__0), .A1 (inputs_173__0), .S0 (
             nx23933)) ;
    mux21_ni ix3561 (.Y (nx3560), .A0 (inputs_174__0), .A1 (inputs_175__0), .S0 (
             nx23933)) ;
    mux21_ni ix3629 (.Y (nx3628), .A0 (nx3596), .A1 (nx3624), .S0 (nx23197)) ;
    mux21_ni ix3597 (.Y (nx3596), .A0 (nx3580), .A1 (nx3592), .S0 (nx23389)) ;
    mux21_ni ix3581 (.Y (nx3580), .A0 (inputs_184__0), .A1 (inputs_185__0), .S0 (
             nx23933)) ;
    mux21_ni ix3593 (.Y (nx3592), .A0 (inputs_186__0), .A1 (inputs_187__0), .S0 (
             nx23933)) ;
    mux21_ni ix3625 (.Y (nx3624), .A0 (nx3608), .A1 (nx3620), .S0 (nx23389)) ;
    mux21_ni ix3609 (.Y (nx3608), .A0 (inputs_188__0), .A1 (inputs_189__0), .S0 (
             nx23933)) ;
    mux21_ni ix3621 (.Y (nx3620), .A0 (inputs_190__0), .A1 (inputs_191__0), .S0 (
             nx23935)) ;
    mux21_ni ix4141 (.Y (nx4140), .A0 (nx3928), .A1 (nx4136), .S0 (nx22535)) ;
    mux21_ni ix3929 (.Y (nx3928), .A0 (nx3922), .A1 (nx3844), .S0 (nx23121)) ;
    oai21 ix3923 (.Y (nx3922), .A0 (nx22235), .A1 (nx9059), .B0 (nx9071)) ;
    mux21 ix9060 (.Y (nx9059), .A0 (nx3886), .A1 (nx3914), .S0 (nx22701)) ;
    mux21_ni ix3887 (.Y (nx3886), .A0 (nx3870), .A1 (nx3882), .S0 (nx23389)) ;
    mux21_ni ix3871 (.Y (nx3870), .A0 (inputs_196__0), .A1 (inputs_197__0), .S0 (
             nx23935)) ;
    mux21_ni ix3883 (.Y (nx3882), .A0 (inputs_198__0), .A1 (inputs_199__0), .S0 (
             nx23935)) ;
    mux21_ni ix3915 (.Y (nx3914), .A0 (nx3898), .A1 (nx3910), .S0 (nx23389)) ;
    mux21_ni ix3899 (.Y (nx3898), .A0 (inputs_212__0), .A1 (inputs_213__0), .S0 (
             nx23935)) ;
    mux21_ni ix3911 (.Y (nx3910), .A0 (inputs_214__0), .A1 (inputs_215__0), .S0 (
             nx23935)) ;
    nand04 ix9072 (.Y (nx9071), .A0 (nx22235), .A1 (nx23389), .A2 (nx23935), .A3 (
           nx3858)) ;
    mux21_ni ix3859 (.Y (nx3858), .A0 (inputs_195__0), .A1 (inputs_211__0), .S0 (
             nx22703)) ;
    mux21_ni ix3845 (.Y (nx3844), .A0 (nx3780), .A1 (nx3840), .S0 (nx22703)) ;
    mux21_ni ix3781 (.Y (nx3780), .A0 (nx3748), .A1 (nx3776), .S0 (nx23199)) ;
    mux21_ni ix3749 (.Y (nx3748), .A0 (nx3732), .A1 (nx3744), .S0 (nx23389)) ;
    mux21_ni ix3733 (.Y (nx3732), .A0 (inputs_200__0), .A1 (inputs_201__0), .S0 (
             nx23935)) ;
    mux21_ni ix3745 (.Y (nx3744), .A0 (inputs_202__0), .A1 (inputs_203__0), .S0 (
             nx23937)) ;
    mux21_ni ix3777 (.Y (nx3776), .A0 (nx3760), .A1 (nx3772), .S0 (nx23389)) ;
    mux21_ni ix3761 (.Y (nx3760), .A0 (inputs_204__0), .A1 (inputs_205__0), .S0 (
             nx23937)) ;
    mux21_ni ix3773 (.Y (nx3772), .A0 (inputs_206__0), .A1 (inputs_207__0), .S0 (
             nx23937)) ;
    mux21_ni ix3841 (.Y (nx3840), .A0 (nx3808), .A1 (nx3836), .S0 (nx23199)) ;
    mux21_ni ix3809 (.Y (nx3808), .A0 (nx3792), .A1 (nx3804), .S0 (nx23391)) ;
    mux21_ni ix3793 (.Y (nx3792), .A0 (inputs_216__0), .A1 (inputs_217__0), .S0 (
             nx23937)) ;
    mux21_ni ix3805 (.Y (nx3804), .A0 (inputs_218__0), .A1 (inputs_219__0), .S0 (
             nx23937)) ;
    mux21_ni ix3837 (.Y (nx3836), .A0 (nx3820), .A1 (nx3832), .S0 (nx23391)) ;
    mux21_ni ix3821 (.Y (nx3820), .A0 (inputs_220__0), .A1 (inputs_221__0), .S0 (
             nx23937)) ;
    mux21_ni ix3833 (.Y (nx3832), .A0 (inputs_222__0), .A1 (inputs_223__0), .S0 (
             nx23937)) ;
    mux21_ni ix4137 (.Y (nx4136), .A0 (nx4130), .A1 (nx4052), .S0 (nx23121)) ;
    oai21 ix4131 (.Y (nx4130), .A0 (nx22235), .A1 (nx9103), .B0 (nx9113)) ;
    mux21 ix9104 (.Y (nx9103), .A0 (nx4094), .A1 (nx4122), .S0 (nx22703)) ;
    mux21_ni ix4095 (.Y (nx4094), .A0 (nx4078), .A1 (nx4090), .S0 (nx23391)) ;
    mux21_ni ix4079 (.Y (nx4078), .A0 (inputs_228__0), .A1 (inputs_229__0), .S0 (
             nx23939)) ;
    mux21_ni ix4091 (.Y (nx4090), .A0 (inputs_230__0), .A1 (inputs_231__0), .S0 (
             nx23939)) ;
    mux21_ni ix4123 (.Y (nx4122), .A0 (nx4106), .A1 (nx4118), .S0 (nx23391)) ;
    mux21_ni ix4107 (.Y (nx4106), .A0 (inputs_244__0), .A1 (inputs_245__0), .S0 (
             nx23939)) ;
    mux21_ni ix4119 (.Y (nx4118), .A0 (inputs_246__0), .A1 (inputs_247__0), .S0 (
             nx23939)) ;
    nand04 ix9114 (.Y (nx9113), .A0 (nx22235), .A1 (nx23391), .A2 (nx23939), .A3 (
           nx4066)) ;
    mux21_ni ix4067 (.Y (nx4066), .A0 (inputs_227__0), .A1 (inputs_243__0), .S0 (
             nx22703)) ;
    mux21_ni ix4053 (.Y (nx4052), .A0 (nx3988), .A1 (nx4048), .S0 (nx22703)) ;
    mux21_ni ix3989 (.Y (nx3988), .A0 (nx3956), .A1 (nx3984), .S0 (nx23199)) ;
    mux21_ni ix3957 (.Y (nx3956), .A0 (nx3940), .A1 (nx3952), .S0 (nx23391)) ;
    mux21_ni ix3941 (.Y (nx3940), .A0 (inputs_232__0), .A1 (inputs_233__0), .S0 (
             nx23939)) ;
    mux21_ni ix3953 (.Y (nx3952), .A0 (inputs_234__0), .A1 (inputs_235__0), .S0 (
             nx23939)) ;
    mux21_ni ix3985 (.Y (nx3984), .A0 (nx3968), .A1 (nx3980), .S0 (nx23391)) ;
    mux21_ni ix3969 (.Y (nx3968), .A0 (inputs_236__0), .A1 (inputs_237__0), .S0 (
             nx23941)) ;
    mux21_ni ix3981 (.Y (nx3980), .A0 (inputs_238__0), .A1 (inputs_239__0), .S0 (
             nx23941)) ;
    mux21_ni ix4049 (.Y (nx4048), .A0 (nx4016), .A1 (nx4044), .S0 (nx23199)) ;
    mux21_ni ix4017 (.Y (nx4016), .A0 (nx4000), .A1 (nx4012), .S0 (nx23393)) ;
    mux21_ni ix4001 (.Y (nx4000), .A0 (inputs_248__0), .A1 (inputs_249__0), .S0 (
             nx23941)) ;
    mux21_ni ix4013 (.Y (nx4012), .A0 (inputs_250__0), .A1 (inputs_251__0), .S0 (
             nx23941)) ;
    mux21_ni ix4045 (.Y (nx4044), .A0 (nx4028), .A1 (nx4040), .S0 (nx23393)) ;
    mux21_ni ix4029 (.Y (nx4028), .A0 (inputs_252__0), .A1 (inputs_253__0), .S0 (
             nx23941)) ;
    mux21_ni ix4041 (.Y (nx4040), .A0 (inputs_254__0), .A1 (inputs_255__0), .S0 (
             nx23941)) ;
    oai21 ix8315 (.Y (\output [1]), .A0 (nx24851), .A1 (nx9145), .B0 (nx9499)) ;
    mux21 ix9146 (.Y (nx9145), .A0 (nx4996), .A1 (nx5840), .S0 (nx22413)) ;
    mux21_ni ix4997 (.Y (nx4996), .A0 (nx4572), .A1 (nx4992), .S0 (nx22455)) ;
    mux21_ni ix4573 (.Y (nx4572), .A0 (nx4360), .A1 (nx4568), .S0 (nx22535)) ;
    mux21_ni ix4361 (.Y (nx4360), .A0 (nx4354), .A1 (nx4276), .S0 (nx23121)) ;
    oai21 ix4355 (.Y (nx4354), .A0 (nx22235), .A1 (nx9155), .B0 (nx9165)) ;
    mux21 ix9156 (.Y (nx9155), .A0 (nx4318), .A1 (nx4346), .S0 (nx22703)) ;
    mux21_ni ix4319 (.Y (nx4318), .A0 (nx4302), .A1 (nx4314), .S0 (nx23393)) ;
    mux21_ni ix4303 (.Y (nx4302), .A0 (inputs_260__1), .A1 (inputs_261__1), .S0 (
             nx23941)) ;
    mux21_ni ix4315 (.Y (nx4314), .A0 (inputs_262__1), .A1 (inputs_263__1), .S0 (
             nx23943)) ;
    mux21_ni ix4347 (.Y (nx4346), .A0 (nx4330), .A1 (nx4342), .S0 (nx23393)) ;
    mux21_ni ix4331 (.Y (nx4330), .A0 (inputs_276__1), .A1 (inputs_277__1), .S0 (
             nx23943)) ;
    mux21_ni ix4343 (.Y (nx4342), .A0 (inputs_278__1), .A1 (inputs_279__1), .S0 (
             nx23943)) ;
    nand04 ix9166 (.Y (nx9165), .A0 (nx22235), .A1 (nx23393), .A2 (nx23943), .A3 (
           nx4290)) ;
    mux21_ni ix4291 (.Y (nx4290), .A0 (inputs_259__1), .A1 (inputs_275__1), .S0 (
             nx22703)) ;
    mux21_ni ix4277 (.Y (nx4276), .A0 (nx4212), .A1 (nx4272), .S0 (nx22705)) ;
    mux21_ni ix4213 (.Y (nx4212), .A0 (nx4180), .A1 (nx4208), .S0 (nx23199)) ;
    mux21_ni ix4181 (.Y (nx4180), .A0 (nx4164), .A1 (nx4176), .S0 (nx23393)) ;
    mux21_ni ix4165 (.Y (nx4164), .A0 (inputs_264__1), .A1 (inputs_265__1), .S0 (
             nx23943)) ;
    mux21_ni ix4177 (.Y (nx4176), .A0 (inputs_266__1), .A1 (inputs_267__1), .S0 (
             nx23943)) ;
    mux21_ni ix4209 (.Y (nx4208), .A0 (nx4192), .A1 (nx4204), .S0 (nx23393)) ;
    mux21_ni ix4193 (.Y (nx4192), .A0 (inputs_268__1), .A1 (inputs_269__1), .S0 (
             nx23943)) ;
    mux21_ni ix4205 (.Y (nx4204), .A0 (inputs_270__1), .A1 (inputs_271__1), .S0 (
             nx23945)) ;
    mux21_ni ix4273 (.Y (nx4272), .A0 (nx4240), .A1 (nx4268), .S0 (nx23199)) ;
    mux21_ni ix4241 (.Y (nx4240), .A0 (nx4224), .A1 (nx4236), .S0 (nx23395)) ;
    mux21_ni ix4225 (.Y (nx4224), .A0 (inputs_280__1), .A1 (inputs_281__1), .S0 (
             nx23945)) ;
    mux21_ni ix4237 (.Y (nx4236), .A0 (inputs_282__1), .A1 (inputs_283__1), .S0 (
             nx23945)) ;
    mux21_ni ix4269 (.Y (nx4268), .A0 (nx4252), .A1 (nx4264), .S0 (nx23395)) ;
    mux21_ni ix4253 (.Y (nx4252), .A0 (inputs_284__1), .A1 (inputs_285__1), .S0 (
             nx23945)) ;
    mux21_ni ix4265 (.Y (nx4264), .A0 (inputs_286__1), .A1 (inputs_287__1), .S0 (
             nx23945)) ;
    mux21_ni ix4569 (.Y (nx4568), .A0 (nx4562), .A1 (nx4484), .S0 (nx23121)) ;
    oai21 ix4563 (.Y (nx4562), .A0 (nx22237), .A1 (nx9195), .B0 (nx9205)) ;
    mux21 ix9196 (.Y (nx9195), .A0 (nx4526), .A1 (nx4554), .S0 (nx22705)) ;
    mux21_ni ix4527 (.Y (nx4526), .A0 (nx4510), .A1 (nx4522), .S0 (nx23395)) ;
    mux21_ni ix4511 (.Y (nx4510), .A0 (inputs_292__1), .A1 (inputs_293__1), .S0 (
             nx23945)) ;
    mux21_ni ix4523 (.Y (nx4522), .A0 (inputs_294__1), .A1 (inputs_295__1), .S0 (
             nx23945)) ;
    mux21_ni ix4555 (.Y (nx4554), .A0 (nx4538), .A1 (nx4550), .S0 (nx23395)) ;
    mux21_ni ix4539 (.Y (nx4538), .A0 (inputs_308__1), .A1 (inputs_309__1), .S0 (
             nx23947)) ;
    mux21_ni ix4551 (.Y (nx4550), .A0 (inputs_310__1), .A1 (inputs_311__1), .S0 (
             nx23947)) ;
    nand04 ix9206 (.Y (nx9205), .A0 (nx22237), .A1 (nx23395), .A2 (nx23947), .A3 (
           nx4498)) ;
    mux21_ni ix4499 (.Y (nx4498), .A0 (inputs_291__1), .A1 (inputs_307__1), .S0 (
             nx22705)) ;
    mux21_ni ix4485 (.Y (nx4484), .A0 (nx4420), .A1 (nx4480), .S0 (nx22705)) ;
    mux21_ni ix4421 (.Y (nx4420), .A0 (nx4388), .A1 (nx4416), .S0 (nx23199)) ;
    mux21_ni ix4389 (.Y (nx4388), .A0 (nx4372), .A1 (nx4384), .S0 (nx23395)) ;
    mux21_ni ix4373 (.Y (nx4372), .A0 (inputs_296__1), .A1 (inputs_297__1), .S0 (
             nx23947)) ;
    mux21_ni ix4385 (.Y (nx4384), .A0 (inputs_298__1), .A1 (inputs_299__1), .S0 (
             nx23947)) ;
    mux21_ni ix4417 (.Y (nx4416), .A0 (nx4400), .A1 (nx4412), .S0 (nx23395)) ;
    mux21_ni ix4401 (.Y (nx4400), .A0 (inputs_300__1), .A1 (inputs_301__1), .S0 (
             nx23947)) ;
    mux21_ni ix4413 (.Y (nx4412), .A0 (inputs_302__1), .A1 (inputs_303__1), .S0 (
             nx23947)) ;
    mux21_ni ix4481 (.Y (nx4480), .A0 (nx4448), .A1 (nx4476), .S0 (nx23201)) ;
    mux21_ni ix4449 (.Y (nx4448), .A0 (nx4432), .A1 (nx4444), .S0 (nx23397)) ;
    mux21_ni ix4433 (.Y (nx4432), .A0 (inputs_312__1), .A1 (inputs_313__1), .S0 (
             nx23949)) ;
    mux21_ni ix4445 (.Y (nx4444), .A0 (inputs_314__1), .A1 (inputs_315__1), .S0 (
             nx23949)) ;
    mux21_ni ix4477 (.Y (nx4476), .A0 (nx4460), .A1 (nx4472), .S0 (nx23397)) ;
    mux21_ni ix4461 (.Y (nx4460), .A0 (inputs_316__1), .A1 (inputs_317__1), .S0 (
             nx23949)) ;
    mux21_ni ix4473 (.Y (nx4472), .A0 (inputs_318__1), .A1 (inputs_319__1), .S0 (
             nx23949)) ;
    mux21_ni ix4993 (.Y (nx4992), .A0 (nx4780), .A1 (nx4988), .S0 (nx22535)) ;
    mux21_ni ix4781 (.Y (nx4780), .A0 (nx4774), .A1 (nx4696), .S0 (nx23121)) ;
    oai21 ix4775 (.Y (nx4774), .A0 (nx22237), .A1 (nx9237), .B0 (nx9249)) ;
    mux21 ix9238 (.Y (nx9237), .A0 (nx4738), .A1 (nx4766), .S0 (nx22705)) ;
    mux21_ni ix4739 (.Y (nx4738), .A0 (nx4722), .A1 (nx4734), .S0 (nx23397)) ;
    mux21_ni ix4723 (.Y (nx4722), .A0 (inputs_324__1), .A1 (inputs_325__1), .S0 (
             nx23949)) ;
    mux21_ni ix4735 (.Y (nx4734), .A0 (inputs_326__1), .A1 (inputs_327__1), .S0 (
             nx23949)) ;
    mux21_ni ix4767 (.Y (nx4766), .A0 (nx4750), .A1 (nx4762), .S0 (nx23397)) ;
    mux21_ni ix4751 (.Y (nx4750), .A0 (inputs_340__1), .A1 (inputs_341__1), .S0 (
             nx23949)) ;
    mux21_ni ix4763 (.Y (nx4762), .A0 (inputs_342__1), .A1 (inputs_343__1), .S0 (
             nx23951)) ;
    nand04 ix9250 (.Y (nx9249), .A0 (nx22237), .A1 (nx23397), .A2 (nx23951), .A3 (
           nx4710)) ;
    mux21_ni ix4711 (.Y (nx4710), .A0 (inputs_323__1), .A1 (inputs_339__1), .S0 (
             nx22705)) ;
    mux21_ni ix4697 (.Y (nx4696), .A0 (nx4632), .A1 (nx4692), .S0 (nx22705)) ;
    mux21_ni ix4633 (.Y (nx4632), .A0 (nx4600), .A1 (nx4628), .S0 (nx23201)) ;
    mux21_ni ix4601 (.Y (nx4600), .A0 (nx4584), .A1 (nx4596), .S0 (nx23397)) ;
    mux21_ni ix4585 (.Y (nx4584), .A0 (inputs_328__1), .A1 (inputs_329__1), .S0 (
             nx23951)) ;
    mux21_ni ix4597 (.Y (nx4596), .A0 (inputs_330__1), .A1 (inputs_331__1), .S0 (
             nx23951)) ;
    mux21_ni ix4629 (.Y (nx4628), .A0 (nx4612), .A1 (nx4624), .S0 (nx23397)) ;
    mux21_ni ix4613 (.Y (nx4612), .A0 (inputs_332__1), .A1 (inputs_333__1), .S0 (
             nx23951)) ;
    mux21_ni ix4625 (.Y (nx4624), .A0 (inputs_334__1), .A1 (inputs_335__1), .S0 (
             nx23951)) ;
    mux21_ni ix4693 (.Y (nx4692), .A0 (nx4660), .A1 (nx4688), .S0 (nx23201)) ;
    mux21_ni ix4661 (.Y (nx4660), .A0 (nx4644), .A1 (nx4656), .S0 (nx23399)) ;
    mux21_ni ix4645 (.Y (nx4644), .A0 (inputs_344__1), .A1 (inputs_345__1), .S0 (
             nx23951)) ;
    mux21_ni ix4657 (.Y (nx4656), .A0 (inputs_346__1), .A1 (inputs_347__1), .S0 (
             nx23953)) ;
    mux21_ni ix4689 (.Y (nx4688), .A0 (nx4672), .A1 (nx4684), .S0 (nx23399)) ;
    mux21_ni ix4673 (.Y (nx4672), .A0 (inputs_348__1), .A1 (inputs_349__1), .S0 (
             nx23953)) ;
    mux21_ni ix4685 (.Y (nx4684), .A0 (inputs_350__1), .A1 (inputs_351__1), .S0 (
             nx23953)) ;
    mux21_ni ix4989 (.Y (nx4988), .A0 (nx4982), .A1 (nx4904), .S0 (nx23121)) ;
    oai21 ix4983 (.Y (nx4982), .A0 (nx22237), .A1 (nx9283), .B0 (nx9295)) ;
    mux21 ix9284 (.Y (nx9283), .A0 (nx4946), .A1 (nx4974), .S0 (nx22707)) ;
    mux21_ni ix4947 (.Y (nx4946), .A0 (nx4930), .A1 (nx4942), .S0 (nx23399)) ;
    mux21_ni ix4931 (.Y (nx4930), .A0 (inputs_356__1), .A1 (inputs_357__1), .S0 (
             nx23953)) ;
    mux21_ni ix4943 (.Y (nx4942), .A0 (inputs_358__1), .A1 (inputs_359__1), .S0 (
             nx23953)) ;
    mux21_ni ix4975 (.Y (nx4974), .A0 (nx4958), .A1 (nx4970), .S0 (nx23399)) ;
    mux21_ni ix4959 (.Y (nx4958), .A0 (inputs_372__1), .A1 (inputs_373__1), .S0 (
             nx23953)) ;
    mux21_ni ix4971 (.Y (nx4970), .A0 (inputs_374__1), .A1 (inputs_375__1), .S0 (
             nx23953)) ;
    nand04 ix9296 (.Y (nx9295), .A0 (nx22237), .A1 (nx23399), .A2 (nx23955), .A3 (
           nx4918)) ;
    mux21_ni ix4919 (.Y (nx4918), .A0 (inputs_355__1), .A1 (inputs_371__1), .S0 (
             nx22707)) ;
    mux21_ni ix4905 (.Y (nx4904), .A0 (nx4840), .A1 (nx4900), .S0 (nx22707)) ;
    mux21_ni ix4841 (.Y (nx4840), .A0 (nx4808), .A1 (nx4836), .S0 (nx23201)) ;
    mux21_ni ix4809 (.Y (nx4808), .A0 (nx4792), .A1 (nx4804), .S0 (nx23399)) ;
    mux21_ni ix4793 (.Y (nx4792), .A0 (inputs_360__1), .A1 (inputs_361__1), .S0 (
             nx23955)) ;
    mux21_ni ix4805 (.Y (nx4804), .A0 (inputs_362__1), .A1 (inputs_363__1), .S0 (
             nx23955)) ;
    mux21_ni ix4837 (.Y (nx4836), .A0 (nx4820), .A1 (nx4832), .S0 (nx23399)) ;
    mux21_ni ix4821 (.Y (nx4820), .A0 (inputs_364__1), .A1 (inputs_365__1), .S0 (
             nx23955)) ;
    mux21_ni ix4833 (.Y (nx4832), .A0 (inputs_366__1), .A1 (inputs_367__1), .S0 (
             nx23955)) ;
    mux21_ni ix4901 (.Y (nx4900), .A0 (nx4868), .A1 (nx4896), .S0 (nx23201)) ;
    mux21_ni ix4869 (.Y (nx4868), .A0 (nx4852), .A1 (nx4864), .S0 (nx23401)) ;
    mux21_ni ix4853 (.Y (nx4852), .A0 (inputs_376__1), .A1 (inputs_377__1), .S0 (
             nx23955)) ;
    mux21_ni ix4865 (.Y (nx4864), .A0 (inputs_378__1), .A1 (inputs_379__1), .S0 (
             nx23955)) ;
    mux21_ni ix4897 (.Y (nx4896), .A0 (nx4880), .A1 (nx4892), .S0 (nx23401)) ;
    mux21_ni ix4881 (.Y (nx4880), .A0 (inputs_380__1), .A1 (inputs_381__1), .S0 (
             nx23957)) ;
    mux21_ni ix4893 (.Y (nx4892), .A0 (inputs_382__1), .A1 (inputs_383__1), .S0 (
             nx23957)) ;
    mux21_ni ix5841 (.Y (nx5840), .A0 (nx5416), .A1 (nx5836), .S0 (nx22455)) ;
    mux21_ni ix5417 (.Y (nx5416), .A0 (nx5204), .A1 (nx5412), .S0 (nx22535)) ;
    mux21_ni ix5205 (.Y (nx5204), .A0 (nx5198), .A1 (nx5120), .S0 (nx23121)) ;
    oai21 ix5199 (.Y (nx5198), .A0 (nx22237), .A1 (nx9329), .B0 (nx9341)) ;
    mux21 ix9330 (.Y (nx9329), .A0 (nx5162), .A1 (nx5190), .S0 (nx22707)) ;
    mux21_ni ix5163 (.Y (nx5162), .A0 (nx5146), .A1 (nx5158), .S0 (nx23401)) ;
    mux21_ni ix5147 (.Y (nx5146), .A0 (inputs_388__1), .A1 (inputs_389__1), .S0 (
             nx23957)) ;
    mux21_ni ix5159 (.Y (nx5158), .A0 (inputs_390__1), .A1 (inputs_391__1), .S0 (
             nx23957)) ;
    mux21_ni ix5191 (.Y (nx5190), .A0 (nx5174), .A1 (nx5186), .S0 (nx23401)) ;
    mux21_ni ix5175 (.Y (nx5174), .A0 (inputs_404__1), .A1 (inputs_405__1), .S0 (
             nx23957)) ;
    mux21_ni ix5187 (.Y (nx5186), .A0 (inputs_406__1), .A1 (inputs_407__1), .S0 (
             nx23957)) ;
    nand04 ix9342 (.Y (nx9341), .A0 (nx22239), .A1 (nx23401), .A2 (nx23957), .A3 (
           nx5134)) ;
    mux21_ni ix5135 (.Y (nx5134), .A0 (inputs_387__1), .A1 (inputs_403__1), .S0 (
             nx22707)) ;
    mux21_ni ix5121 (.Y (nx5120), .A0 (nx5056), .A1 (nx5116), .S0 (nx22707)) ;
    mux21_ni ix5057 (.Y (nx5056), .A0 (nx5024), .A1 (nx5052), .S0 (nx23201)) ;
    mux21_ni ix5025 (.Y (nx5024), .A0 (nx5008), .A1 (nx5020), .S0 (nx23401)) ;
    mux21_ni ix5009 (.Y (nx5008), .A0 (inputs_392__1), .A1 (inputs_393__1), .S0 (
             nx23959)) ;
    mux21_ni ix5021 (.Y (nx5020), .A0 (inputs_394__1), .A1 (inputs_395__1), .S0 (
             nx23959)) ;
    mux21_ni ix5053 (.Y (nx5052), .A0 (nx5036), .A1 (nx5048), .S0 (nx23401)) ;
    mux21_ni ix5037 (.Y (nx5036), .A0 (inputs_396__1), .A1 (inputs_397__1), .S0 (
             nx23959)) ;
    mux21_ni ix5049 (.Y (nx5048), .A0 (inputs_398__1), .A1 (inputs_399__1), .S0 (
             nx23959)) ;
    mux21_ni ix5117 (.Y (nx5116), .A0 (nx5084), .A1 (nx5112), .S0 (nx23201)) ;
    mux21_ni ix5085 (.Y (nx5084), .A0 (nx5068), .A1 (nx5080), .S0 (nx23403)) ;
    mux21_ni ix5069 (.Y (nx5068), .A0 (inputs_408__1), .A1 (inputs_409__1), .S0 (
             nx23959)) ;
    mux21_ni ix5081 (.Y (nx5080), .A0 (inputs_410__1), .A1 (inputs_411__1), .S0 (
             nx23959)) ;
    mux21_ni ix5113 (.Y (nx5112), .A0 (nx5096), .A1 (nx5108), .S0 (nx23403)) ;
    mux21_ni ix5097 (.Y (nx5096), .A0 (inputs_412__1), .A1 (inputs_413__1), .S0 (
             nx23959)) ;
    mux21_ni ix5109 (.Y (nx5108), .A0 (inputs_414__1), .A1 (inputs_415__1), .S0 (
             nx23961)) ;
    mux21_ni ix5413 (.Y (nx5412), .A0 (nx5406), .A1 (nx5328), .S0 (nx23123)) ;
    oai21 ix5407 (.Y (nx5406), .A0 (nx22239), .A1 (nx9373), .B0 (nx9383)) ;
    mux21 ix9374 (.Y (nx9373), .A0 (nx5370), .A1 (nx5398), .S0 (nx22707)) ;
    mux21_ni ix5371 (.Y (nx5370), .A0 (nx5354), .A1 (nx5366), .S0 (nx23403)) ;
    mux21_ni ix5355 (.Y (nx5354), .A0 (inputs_420__1), .A1 (inputs_421__1), .S0 (
             nx23961)) ;
    mux21_ni ix5367 (.Y (nx5366), .A0 (inputs_422__1), .A1 (inputs_423__1), .S0 (
             nx23961)) ;
    mux21_ni ix5399 (.Y (nx5398), .A0 (nx5382), .A1 (nx5394), .S0 (nx23403)) ;
    mux21_ni ix5383 (.Y (nx5382), .A0 (inputs_436__1), .A1 (inputs_437__1), .S0 (
             nx23961)) ;
    mux21_ni ix5395 (.Y (nx5394), .A0 (inputs_438__1), .A1 (inputs_439__1), .S0 (
             nx23961)) ;
    nand04 ix9384 (.Y (nx9383), .A0 (nx22239), .A1 (nx23403), .A2 (nx23961), .A3 (
           nx5342)) ;
    mux21_ni ix5343 (.Y (nx5342), .A0 (inputs_419__1), .A1 (inputs_435__1), .S0 (
             nx22709)) ;
    mux21_ni ix5329 (.Y (nx5328), .A0 (nx5264), .A1 (nx5324), .S0 (nx22709)) ;
    mux21_ni ix5265 (.Y (nx5264), .A0 (nx5232), .A1 (nx5260), .S0 (nx23203)) ;
    mux21_ni ix5233 (.Y (nx5232), .A0 (nx5216), .A1 (nx5228), .S0 (nx23403)) ;
    mux21_ni ix5217 (.Y (nx5216), .A0 (inputs_424__1), .A1 (inputs_425__1), .S0 (
             nx23961)) ;
    mux21_ni ix5229 (.Y (nx5228), .A0 (inputs_426__1), .A1 (inputs_427__1), .S0 (
             nx23963)) ;
    mux21_ni ix5261 (.Y (nx5260), .A0 (nx5244), .A1 (nx5256), .S0 (nx23403)) ;
    mux21_ni ix5245 (.Y (nx5244), .A0 (inputs_428__1), .A1 (inputs_429__1), .S0 (
             nx23963)) ;
    mux21_ni ix5257 (.Y (nx5256), .A0 (inputs_430__1), .A1 (inputs_431__1), .S0 (
             nx23963)) ;
    mux21_ni ix5325 (.Y (nx5324), .A0 (nx5292), .A1 (nx5320), .S0 (nx23203)) ;
    mux21_ni ix5293 (.Y (nx5292), .A0 (nx5276), .A1 (nx5288), .S0 (nx23405)) ;
    mux21_ni ix5277 (.Y (nx5276), .A0 (inputs_440__1), .A1 (inputs_441__1), .S0 (
             nx23963)) ;
    mux21_ni ix5289 (.Y (nx5288), .A0 (inputs_442__1), .A1 (inputs_443__1), .S0 (
             nx23963)) ;
    mux21_ni ix5321 (.Y (nx5320), .A0 (nx5304), .A1 (nx5316), .S0 (nx23405)) ;
    mux21_ni ix5305 (.Y (nx5304), .A0 (inputs_444__1), .A1 (inputs_445__1), .S0 (
             nx23963)) ;
    mux21_ni ix5317 (.Y (nx5316), .A0 (inputs_446__1), .A1 (inputs_447__1), .S0 (
             nx23963)) ;
    mux21_ni ix5837 (.Y (nx5836), .A0 (nx5624), .A1 (nx5832), .S0 (nx22537)) ;
    mux21_ni ix5625 (.Y (nx5624), .A0 (nx5618), .A1 (nx5540), .S0 (nx23123)) ;
    oai21 ix5619 (.Y (nx5618), .A0 (nx22239), .A1 (nx9415), .B0 (nx9427)) ;
    mux21 ix9416 (.Y (nx9415), .A0 (nx5582), .A1 (nx5610), .S0 (nx22709)) ;
    mux21_ni ix5583 (.Y (nx5582), .A0 (nx5566), .A1 (nx5578), .S0 (nx23405)) ;
    mux21_ni ix5567 (.Y (nx5566), .A0 (inputs_452__1), .A1 (inputs_453__1), .S0 (
             nx23965)) ;
    mux21_ni ix5579 (.Y (nx5578), .A0 (inputs_454__1), .A1 (inputs_455__1), .S0 (
             nx23965)) ;
    mux21_ni ix5611 (.Y (nx5610), .A0 (nx5594), .A1 (nx5606), .S0 (nx23405)) ;
    mux21_ni ix5595 (.Y (nx5594), .A0 (inputs_468__1), .A1 (inputs_469__1), .S0 (
             nx23965)) ;
    mux21_ni ix5607 (.Y (nx5606), .A0 (inputs_470__1), .A1 (inputs_471__1), .S0 (
             nx23965)) ;
    nand04 ix9428 (.Y (nx9427), .A0 (nx22239), .A1 (nx23405), .A2 (nx23965), .A3 (
           nx5554)) ;
    mux21_ni ix5555 (.Y (nx5554), .A0 (inputs_451__1), .A1 (inputs_467__1), .S0 (
             nx22709)) ;
    mux21_ni ix5541 (.Y (nx5540), .A0 (nx5476), .A1 (nx5536), .S0 (nx22709)) ;
    mux21_ni ix5477 (.Y (nx5476), .A0 (nx5444), .A1 (nx5472), .S0 (nx23203)) ;
    mux21_ni ix5445 (.Y (nx5444), .A0 (nx5428), .A1 (nx5440), .S0 (nx23405)) ;
    mux21_ni ix5429 (.Y (nx5428), .A0 (inputs_456__1), .A1 (inputs_457__1), .S0 (
             nx23965)) ;
    mux21_ni ix5441 (.Y (nx5440), .A0 (inputs_458__1), .A1 (inputs_459__1), .S0 (
             nx23965)) ;
    mux21_ni ix5473 (.Y (nx5472), .A0 (nx5456), .A1 (nx5468), .S0 (nx23405)) ;
    mux21_ni ix5457 (.Y (nx5456), .A0 (inputs_460__1), .A1 (inputs_461__1), .S0 (
             nx23967)) ;
    mux21_ni ix5469 (.Y (nx5468), .A0 (inputs_462__1), .A1 (inputs_463__1), .S0 (
             nx23967)) ;
    mux21_ni ix5537 (.Y (nx5536), .A0 (nx5504), .A1 (nx5532), .S0 (nx23203)) ;
    mux21_ni ix5505 (.Y (nx5504), .A0 (nx5488), .A1 (nx5500), .S0 (nx23407)) ;
    mux21_ni ix5489 (.Y (nx5488), .A0 (inputs_472__1), .A1 (inputs_473__1), .S0 (
             nx23967)) ;
    mux21_ni ix5501 (.Y (nx5500), .A0 (inputs_474__1), .A1 (inputs_475__1), .S0 (
             nx23967)) ;
    mux21_ni ix5533 (.Y (nx5532), .A0 (nx5516), .A1 (nx5528), .S0 (nx23407)) ;
    mux21_ni ix5517 (.Y (nx5516), .A0 (inputs_476__1), .A1 (inputs_477__1), .S0 (
             nx23967)) ;
    mux21_ni ix5529 (.Y (nx5528), .A0 (inputs_478__1), .A1 (inputs_479__1), .S0 (
             nx23967)) ;
    mux21_ni ix5833 (.Y (nx5832), .A0 (nx5826), .A1 (nx5748), .S0 (nx23123)) ;
    oai21 ix5827 (.Y (nx5826), .A0 (nx22239), .A1 (nx9457), .B0 (nx9469)) ;
    mux21 ix9458 (.Y (nx9457), .A0 (nx5790), .A1 (nx5818), .S0 (nx22709)) ;
    mux21_ni ix5791 (.Y (nx5790), .A0 (nx5774), .A1 (nx5786), .S0 (nx23407)) ;
    mux21_ni ix5775 (.Y (nx5774), .A0 (inputs_484__1), .A1 (inputs_485__1), .S0 (
             nx23967)) ;
    mux21_ni ix5787 (.Y (nx5786), .A0 (inputs_486__1), .A1 (inputs_487__1), .S0 (
             nx23969)) ;
    mux21_ni ix5819 (.Y (nx5818), .A0 (nx5802), .A1 (nx5814), .S0 (nx23407)) ;
    mux21_ni ix5803 (.Y (nx5802), .A0 (inputs_500__1), .A1 (inputs_501__1), .S0 (
             nx23969)) ;
    mux21_ni ix5815 (.Y (nx5814), .A0 (inputs_502__1), .A1 (inputs_503__1), .S0 (
             nx23969)) ;
    nand04 ix9470 (.Y (nx9469), .A0 (nx22239), .A1 (nx23407), .A2 (nx23969), .A3 (
           nx5762)) ;
    mux21_ni ix5763 (.Y (nx5762), .A0 (inputs_483__1), .A1 (inputs_499__1), .S0 (
             nx22709)) ;
    mux21_ni ix5749 (.Y (nx5748), .A0 (nx5684), .A1 (nx5744), .S0 (nx22711)) ;
    mux21_ni ix5685 (.Y (nx5684), .A0 (nx5652), .A1 (nx5680), .S0 (nx23203)) ;
    mux21_ni ix5653 (.Y (nx5652), .A0 (nx5636), .A1 (nx5648), .S0 (nx23407)) ;
    mux21_ni ix5637 (.Y (nx5636), .A0 (inputs_488__1), .A1 (inputs_489__1), .S0 (
             nx23969)) ;
    mux21_ni ix5649 (.Y (nx5648), .A0 (inputs_490__1), .A1 (inputs_491__1), .S0 (
             nx23969)) ;
    mux21_ni ix5681 (.Y (nx5680), .A0 (nx5664), .A1 (nx5676), .S0 (nx23407)) ;
    mux21_ni ix5665 (.Y (nx5664), .A0 (inputs_492__1), .A1 (inputs_493__1), .S0 (
             nx23969)) ;
    mux21_ni ix5677 (.Y (nx5676), .A0 (inputs_494__1), .A1 (inputs_495__1), .S0 (
             nx23971)) ;
    mux21_ni ix5745 (.Y (nx5744), .A0 (nx5712), .A1 (nx5740), .S0 (nx23203)) ;
    mux21_ni ix5713 (.Y (nx5712), .A0 (nx5696), .A1 (nx5708), .S0 (nx23409)) ;
    mux21_ni ix5697 (.Y (nx5696), .A0 (inputs_504__1), .A1 (inputs_505__1), .S0 (
             nx23971)) ;
    mux21_ni ix5709 (.Y (nx5708), .A0 (inputs_506__1), .A1 (inputs_507__1), .S0 (
             nx23971)) ;
    mux21_ni ix5741 (.Y (nx5740), .A0 (nx5724), .A1 (nx5736), .S0 (nx23409)) ;
    mux21_ni ix5725 (.Y (nx5724), .A0 (inputs_508__1), .A1 (inputs_509__1), .S0 (
             nx23971)) ;
    mux21_ni ix5737 (.Y (nx5736), .A0 (inputs_510__1), .A1 (inputs_511__1), .S0 (
             nx23971)) ;
    aoi32 ix9500 (.Y (nx9499), .A0 (nx6610), .A1 (nx22385), .A2 (nx22241), .B0 (
          nx24851), .B1 (nx8306)) ;
    oai21 ix6611 (.Y (nx6610), .A0 (nx23409), .A1 (nx9503), .B0 (nx9605)) ;
    mux21 ix9504 (.Y (nx9503), .A0 (nx6348), .A1 (nx6600), .S0 (nx23971)) ;
    mux21_ni ix6349 (.Y (nx6348), .A0 (nx6220), .A1 (nx6344), .S0 (nx22393)) ;
    mux21_ni ix6221 (.Y (nx6220), .A0 (nx6156), .A1 (nx6216), .S0 (nx22413)) ;
    mux21_ni ix6157 (.Y (nx6156), .A0 (nx6124), .A1 (nx6152), .S0 (nx22455)) ;
    mux21_ni ix6125 (.Y (nx6124), .A0 (nx6108), .A1 (nx6120), .S0 (nx22537)) ;
    mux21_ni ix6109 (.Y (nx6108), .A0 (inputs_0__1), .A1 (inputs_16__1), .S0 (
             nx22711)) ;
    mux21_ni ix6121 (.Y (nx6120), .A0 (inputs_32__1), .A1 (inputs_48__1), .S0 (
             nx22711)) ;
    mux21_ni ix6153 (.Y (nx6152), .A0 (nx6136), .A1 (nx6148), .S0 (nx22537)) ;
    mux21_ni ix6137 (.Y (nx6136), .A0 (inputs_64__1), .A1 (inputs_80__1), .S0 (
             nx22711)) ;
    mux21_ni ix6149 (.Y (nx6148), .A0 (inputs_96__1), .A1 (inputs_112__1), .S0 (
             nx22711)) ;
    mux21_ni ix6217 (.Y (nx6216), .A0 (nx6184), .A1 (nx6212), .S0 (nx22455)) ;
    mux21_ni ix6185 (.Y (nx6184), .A0 (nx6168), .A1 (nx6180), .S0 (nx22537)) ;
    mux21_ni ix6169 (.Y (nx6168), .A0 (inputs_128__1), .A1 (inputs_144__1), .S0 (
             nx22711)) ;
    mux21_ni ix6181 (.Y (nx6180), .A0 (inputs_160__1), .A1 (inputs_176__1), .S0 (
             nx22711)) ;
    mux21_ni ix6213 (.Y (nx6212), .A0 (nx6196), .A1 (nx6208), .S0 (nx22537)) ;
    mux21_ni ix6197 (.Y (nx6196), .A0 (inputs_192__1), .A1 (inputs_208__1), .S0 (
             nx22713)) ;
    mux21_ni ix6209 (.Y (nx6208), .A0 (inputs_224__1), .A1 (inputs_240__1), .S0 (
             nx22713)) ;
    mux21_ni ix6345 (.Y (nx6344), .A0 (nx6280), .A1 (nx6340), .S0 (nx22413)) ;
    mux21_ni ix6281 (.Y (nx6280), .A0 (nx6248), .A1 (nx6276), .S0 (nx22455)) ;
    mux21_ni ix6249 (.Y (nx6248), .A0 (nx6232), .A1 (nx6244), .S0 (nx22537)) ;
    mux21_ni ix6233 (.Y (nx6232), .A0 (inputs_256__1), .A1 (inputs_272__1), .S0 (
             nx22713)) ;
    mux21_ni ix6245 (.Y (nx6244), .A0 (inputs_288__1), .A1 (inputs_304__1), .S0 (
             nx22713)) ;
    mux21_ni ix6277 (.Y (nx6276), .A0 (nx6260), .A1 (nx6272), .S0 (nx22537)) ;
    mux21_ni ix6261 (.Y (nx6260), .A0 (inputs_320__1), .A1 (inputs_336__1), .S0 (
             nx22713)) ;
    mux21_ni ix6273 (.Y (nx6272), .A0 (inputs_352__1), .A1 (inputs_368__1), .S0 (
             nx22713)) ;
    mux21_ni ix6341 (.Y (nx6340), .A0 (nx6308), .A1 (nx6336), .S0 (nx22457)) ;
    mux21_ni ix6309 (.Y (nx6308), .A0 (nx6292), .A1 (nx6304), .S0 (nx22539)) ;
    mux21_ni ix6293 (.Y (nx6292), .A0 (inputs_384__1), .A1 (inputs_400__1), .S0 (
             nx22713)) ;
    mux21_ni ix6305 (.Y (nx6304), .A0 (inputs_416__1), .A1 (inputs_432__1), .S0 (
             nx22715)) ;
    mux21_ni ix6337 (.Y (nx6336), .A0 (nx6320), .A1 (nx6332), .S0 (nx22539)) ;
    mux21_ni ix6321 (.Y (nx6320), .A0 (inputs_448__1), .A1 (inputs_464__1), .S0 (
             nx22715)) ;
    mux21_ni ix6333 (.Y (nx6332), .A0 (inputs_480__1), .A1 (inputs_496__1), .S0 (
             nx22715)) ;
    mux21_ni ix6601 (.Y (nx6600), .A0 (nx6472), .A1 (nx6596), .S0 (nx22393)) ;
    mux21_ni ix6473 (.Y (nx6472), .A0 (nx6408), .A1 (nx6468), .S0 (nx22413)) ;
    mux21_ni ix6409 (.Y (nx6408), .A0 (nx6376), .A1 (nx6404), .S0 (nx22457)) ;
    mux21_ni ix6377 (.Y (nx6376), .A0 (nx6360), .A1 (nx6372), .S0 (nx22539)) ;
    mux21_ni ix6361 (.Y (nx6360), .A0 (inputs_1__1), .A1 (inputs_17__1), .S0 (
             nx22715)) ;
    mux21_ni ix6373 (.Y (nx6372), .A0 (inputs_33__1), .A1 (inputs_49__1), .S0 (
             nx22715)) ;
    mux21_ni ix6405 (.Y (nx6404), .A0 (nx6388), .A1 (nx6400), .S0 (nx22539)) ;
    mux21_ni ix6389 (.Y (nx6388), .A0 (inputs_65__1), .A1 (inputs_81__1), .S0 (
             nx22715)) ;
    mux21_ni ix6401 (.Y (nx6400), .A0 (inputs_97__1), .A1 (inputs_113__1), .S0 (
             nx22715)) ;
    mux21_ni ix6469 (.Y (nx6468), .A0 (nx6436), .A1 (nx6464), .S0 (nx22457)) ;
    mux21_ni ix6437 (.Y (nx6436), .A0 (nx6420), .A1 (nx6432), .S0 (nx22539)) ;
    mux21_ni ix6421 (.Y (nx6420), .A0 (inputs_129__1), .A1 (inputs_145__1), .S0 (
             nx22717)) ;
    mux21_ni ix6433 (.Y (nx6432), .A0 (inputs_161__1), .A1 (inputs_177__1), .S0 (
             nx22717)) ;
    mux21_ni ix6465 (.Y (nx6464), .A0 (nx6448), .A1 (nx6460), .S0 (nx22539)) ;
    mux21_ni ix6449 (.Y (nx6448), .A0 (inputs_193__1), .A1 (inputs_209__1), .S0 (
             nx22717)) ;
    mux21_ni ix6461 (.Y (nx6460), .A0 (inputs_225__1), .A1 (inputs_241__1), .S0 (
             nx22717)) ;
    mux21_ni ix6597 (.Y (nx6596), .A0 (nx6532), .A1 (nx6592), .S0 (nx22413)) ;
    mux21_ni ix6533 (.Y (nx6532), .A0 (nx6500), .A1 (nx6528), .S0 (nx22457)) ;
    mux21_ni ix6501 (.Y (nx6500), .A0 (nx6484), .A1 (nx6496), .S0 (nx22539)) ;
    mux21_ni ix6485 (.Y (nx6484), .A0 (inputs_257__1), .A1 (inputs_273__1), .S0 (
             nx22717)) ;
    mux21_ni ix6497 (.Y (nx6496), .A0 (inputs_289__1), .A1 (inputs_305__1), .S0 (
             nx22717)) ;
    mux21_ni ix6529 (.Y (nx6528), .A0 (nx6512), .A1 (nx6524), .S0 (nx22541)) ;
    mux21_ni ix6513 (.Y (nx6512), .A0 (inputs_321__1), .A1 (inputs_337__1), .S0 (
             nx22717)) ;
    mux21_ni ix6525 (.Y (nx6524), .A0 (inputs_353__1), .A1 (inputs_369__1), .S0 (
             nx22719)) ;
    mux21_ni ix6593 (.Y (nx6592), .A0 (nx6560), .A1 (nx6588), .S0 (nx22457)) ;
    mux21_ni ix6561 (.Y (nx6560), .A0 (nx6544), .A1 (nx6556), .S0 (nx22541)) ;
    mux21_ni ix6545 (.Y (nx6544), .A0 (inputs_385__1), .A1 (inputs_401__1), .S0 (
             nx22719)) ;
    mux21_ni ix6557 (.Y (nx6556), .A0 (inputs_417__1), .A1 (inputs_433__1), .S0 (
             nx22719)) ;
    mux21_ni ix6589 (.Y (nx6588), .A0 (nx6572), .A1 (nx6584), .S0 (nx22541)) ;
    mux21_ni ix6573 (.Y (nx6572), .A0 (inputs_449__1), .A1 (inputs_465__1), .S0 (
             nx22719)) ;
    mux21_ni ix6585 (.Y (nx6584), .A0 (inputs_481__1), .A1 (inputs_497__1), .S0 (
             nx22719)) ;
    nand03 ix9606 (.Y (nx9605), .A0 (nx6094), .A1 (nx23409), .A2 (nx24879)) ;
    mux21_ni ix6095 (.Y (nx6094), .A0 (nx5966), .A1 (nx6090), .S0 (nx22393)) ;
    mux21_ni ix5967 (.Y (nx5966), .A0 (nx5902), .A1 (nx5962), .S0 (nx22413)) ;
    mux21_ni ix5903 (.Y (nx5902), .A0 (nx5870), .A1 (nx5898), .S0 (nx22457)) ;
    mux21_ni ix5871 (.Y (nx5870), .A0 (nx5854), .A1 (nx5866), .S0 (nx22541)) ;
    mux21_ni ix5855 (.Y (nx5854), .A0 (inputs_2__1), .A1 (inputs_18__1), .S0 (
             nx22719)) ;
    mux21_ni ix5867 (.Y (nx5866), .A0 (inputs_34__1), .A1 (inputs_50__1), .S0 (
             nx22719)) ;
    mux21_ni ix5899 (.Y (nx5898), .A0 (nx5882), .A1 (nx5894), .S0 (nx22541)) ;
    mux21_ni ix5883 (.Y (nx5882), .A0 (inputs_66__1), .A1 (inputs_82__1), .S0 (
             nx22721)) ;
    mux21_ni ix5895 (.Y (nx5894), .A0 (inputs_98__1), .A1 (inputs_114__1), .S0 (
             nx22721)) ;
    mux21_ni ix5963 (.Y (nx5962), .A0 (nx5930), .A1 (nx5958), .S0 (nx22457)) ;
    mux21_ni ix5931 (.Y (nx5930), .A0 (nx5914), .A1 (nx5926), .S0 (nx22541)) ;
    mux21_ni ix5915 (.Y (nx5914), .A0 (inputs_130__1), .A1 (inputs_146__1), .S0 (
             nx22721)) ;
    mux21_ni ix5927 (.Y (nx5926), .A0 (inputs_162__1), .A1 (inputs_178__1), .S0 (
             nx22721)) ;
    mux21_ni ix5959 (.Y (nx5958), .A0 (nx5942), .A1 (nx5954), .S0 (nx22541)) ;
    mux21_ni ix5943 (.Y (nx5942), .A0 (inputs_194__1), .A1 (inputs_210__1), .S0 (
             nx22721)) ;
    mux21_ni ix5955 (.Y (nx5954), .A0 (inputs_226__1), .A1 (inputs_242__1), .S0 (
             nx22721)) ;
    mux21_ni ix6091 (.Y (nx6090), .A0 (nx6026), .A1 (nx6086), .S0 (nx22415)) ;
    mux21_ni ix6027 (.Y (nx6026), .A0 (nx5994), .A1 (nx6022), .S0 (nx22459)) ;
    mux21_ni ix5995 (.Y (nx5994), .A0 (nx5978), .A1 (nx5990), .S0 (nx22543)) ;
    mux21_ni ix5979 (.Y (nx5978), .A0 (inputs_258__1), .A1 (inputs_274__1), .S0 (
             nx22721)) ;
    mux21_ni ix5991 (.Y (nx5990), .A0 (inputs_290__1), .A1 (inputs_306__1), .S0 (
             nx22723)) ;
    mux21_ni ix6023 (.Y (nx6022), .A0 (nx6006), .A1 (nx6018), .S0 (nx22543)) ;
    mux21_ni ix6007 (.Y (nx6006), .A0 (inputs_322__1), .A1 (inputs_338__1), .S0 (
             nx22723)) ;
    mux21_ni ix6019 (.Y (nx6018), .A0 (inputs_354__1), .A1 (inputs_370__1), .S0 (
             nx22723)) ;
    mux21_ni ix6087 (.Y (nx6086), .A0 (nx6054), .A1 (nx6082), .S0 (nx22459)) ;
    mux21_ni ix6055 (.Y (nx6054), .A0 (nx6038), .A1 (nx6050), .S0 (nx22543)) ;
    mux21_ni ix6039 (.Y (nx6038), .A0 (inputs_386__1), .A1 (inputs_402__1), .S0 (
             nx22723)) ;
    mux21_ni ix6051 (.Y (nx6050), .A0 (inputs_418__1), .A1 (inputs_434__1), .S0 (
             nx22723)) ;
    mux21_ni ix6083 (.Y (nx6082), .A0 (nx6066), .A1 (nx6078), .S0 (nx22543)) ;
    mux21_ni ix6067 (.Y (nx6066), .A0 (inputs_450__1), .A1 (inputs_466__1), .S0 (
             nx22723)) ;
    mux21_ni ix6079 (.Y (nx6078), .A0 (inputs_482__1), .A1 (inputs_498__1), .S0 (
             nx22723)) ;
    mux21_ni ix8307 (.Y (nx8306), .A0 (nx7458), .A1 (nx8302), .S0 (nx22415)) ;
    mux21_ni ix7459 (.Y (nx7458), .A0 (nx7034), .A1 (nx7454), .S0 (nx22459)) ;
    mux21_ni ix7035 (.Y (nx7034), .A0 (nx6822), .A1 (nx7030), .S0 (nx22543)) ;
    mux21_ni ix6823 (.Y (nx6822), .A0 (nx6816), .A1 (nx6738), .S0 (nx23123)) ;
    oai21 ix6817 (.Y (nx6816), .A0 (nx22241), .A1 (nx9665), .B0 (nx9677)) ;
    mux21 ix9666 (.Y (nx9665), .A0 (nx6780), .A1 (nx6808), .S0 (nx22725)) ;
    mux21_ni ix6781 (.Y (nx6780), .A0 (nx6764), .A1 (nx6776), .S0 (nx23409)) ;
    mux21_ni ix6765 (.Y (nx6764), .A0 (inputs_4__1), .A1 (inputs_5__1), .S0 (
             nx23971)) ;
    mux21_ni ix6777 (.Y (nx6776), .A0 (inputs_6__1), .A1 (inputs_7__1), .S0 (
             nx23973)) ;
    mux21_ni ix6809 (.Y (nx6808), .A0 (nx6792), .A1 (nx6804), .S0 (nx23409)) ;
    mux21_ni ix6793 (.Y (nx6792), .A0 (inputs_20__1), .A1 (inputs_21__1), .S0 (
             nx23973)) ;
    mux21_ni ix6805 (.Y (nx6804), .A0 (inputs_22__1), .A1 (inputs_23__1), .S0 (
             nx23973)) ;
    nand04 ix9678 (.Y (nx9677), .A0 (nx22241), .A1 (nx23409), .A2 (nx23973), .A3 (
           nx6752)) ;
    mux21_ni ix6753 (.Y (nx6752), .A0 (inputs_3__1), .A1 (inputs_19__1), .S0 (
             nx22725)) ;
    mux21_ni ix6739 (.Y (nx6738), .A0 (nx6674), .A1 (nx6734), .S0 (nx22725)) ;
    mux21_ni ix6675 (.Y (nx6674), .A0 (nx6642), .A1 (nx6670), .S0 (nx23203)) ;
    mux21_ni ix6643 (.Y (nx6642), .A0 (nx6626), .A1 (nx6638), .S0 (nx23411)) ;
    mux21_ni ix6627 (.Y (nx6626), .A0 (inputs_8__1), .A1 (inputs_9__1), .S0 (
             nx23973)) ;
    mux21_ni ix6639 (.Y (nx6638), .A0 (inputs_10__1), .A1 (inputs_11__1), .S0 (
             nx23973)) ;
    mux21_ni ix6671 (.Y (nx6670), .A0 (nx6654), .A1 (nx6666), .S0 (nx23411)) ;
    mux21_ni ix6655 (.Y (nx6654), .A0 (inputs_12__1), .A1 (inputs_13__1), .S0 (
             nx23973)) ;
    mux21_ni ix6667 (.Y (nx6666), .A0 (inputs_14__1), .A1 (inputs_15__1), .S0 (
             nx23975)) ;
    mux21_ni ix6735 (.Y (nx6734), .A0 (nx6702), .A1 (nx6730), .S0 (nx23205)) ;
    mux21_ni ix6703 (.Y (nx6702), .A0 (nx6686), .A1 (nx6698), .S0 (nx23411)) ;
    mux21_ni ix6687 (.Y (nx6686), .A0 (inputs_24__1), .A1 (inputs_25__1), .S0 (
             nx23975)) ;
    mux21_ni ix6699 (.Y (nx6698), .A0 (inputs_26__1), .A1 (inputs_27__1), .S0 (
             nx23975)) ;
    mux21_ni ix6731 (.Y (nx6730), .A0 (nx6714), .A1 (nx6726), .S0 (nx23411)) ;
    mux21_ni ix6715 (.Y (nx6714), .A0 (inputs_28__1), .A1 (inputs_29__1), .S0 (
             nx23975)) ;
    mux21_ni ix6727 (.Y (nx6726), .A0 (inputs_30__1), .A1 (inputs_31__1), .S0 (
             nx23975)) ;
    mux21_ni ix7031 (.Y (nx7030), .A0 (nx7024), .A1 (nx6946), .S0 (nx23123)) ;
    oai21 ix7025 (.Y (nx7024), .A0 (nx22241), .A1 (nx9709), .B0 (nx9721)) ;
    mux21 ix9710 (.Y (nx9709), .A0 (nx6988), .A1 (nx7016), .S0 (nx22725)) ;
    mux21_ni ix6989 (.Y (nx6988), .A0 (nx6972), .A1 (nx6984), .S0 (nx23411)) ;
    mux21_ni ix6973 (.Y (nx6972), .A0 (inputs_36__1), .A1 (inputs_37__1), .S0 (
             nx23975)) ;
    mux21_ni ix6985 (.Y (nx6984), .A0 (inputs_38__1), .A1 (inputs_39__1), .S0 (
             nx23975)) ;
    mux21_ni ix7017 (.Y (nx7016), .A0 (nx7000), .A1 (nx7012), .S0 (nx23411)) ;
    mux21_ni ix7001 (.Y (nx7000), .A0 (inputs_52__1), .A1 (inputs_53__1), .S0 (
             nx23977)) ;
    mux21_ni ix7013 (.Y (nx7012), .A0 (inputs_54__1), .A1 (inputs_55__1), .S0 (
             nx23977)) ;
    nand04 ix9722 (.Y (nx9721), .A0 (nx22241), .A1 (nx23411), .A2 (nx23977), .A3 (
           nx6960)) ;
    mux21_ni ix6961 (.Y (nx6960), .A0 (inputs_35__1), .A1 (inputs_51__1), .S0 (
             nx22725)) ;
    mux21_ni ix6947 (.Y (nx6946), .A0 (nx6882), .A1 (nx6942), .S0 (nx22725)) ;
    mux21_ni ix6883 (.Y (nx6882), .A0 (nx6850), .A1 (nx6878), .S0 (nx23205)) ;
    mux21_ni ix6851 (.Y (nx6850), .A0 (nx6834), .A1 (nx6846), .S0 (nx23413)) ;
    mux21_ni ix6835 (.Y (nx6834), .A0 (inputs_40__1), .A1 (inputs_41__1), .S0 (
             nx23977)) ;
    mux21_ni ix6847 (.Y (nx6846), .A0 (inputs_42__1), .A1 (inputs_43__1), .S0 (
             nx23977)) ;
    mux21_ni ix6879 (.Y (nx6878), .A0 (nx6862), .A1 (nx6874), .S0 (nx23413)) ;
    mux21_ni ix6863 (.Y (nx6862), .A0 (inputs_44__1), .A1 (inputs_45__1), .S0 (
             nx23977)) ;
    mux21_ni ix6875 (.Y (nx6874), .A0 (inputs_46__1), .A1 (inputs_47__1), .S0 (
             nx23977)) ;
    mux21_ni ix6943 (.Y (nx6942), .A0 (nx6910), .A1 (nx6938), .S0 (nx23205)) ;
    mux21_ni ix6911 (.Y (nx6910), .A0 (nx6894), .A1 (nx6906), .S0 (nx23413)) ;
    mux21_ni ix6895 (.Y (nx6894), .A0 (inputs_56__1), .A1 (inputs_57__1), .S0 (
             nx23979)) ;
    mux21_ni ix6907 (.Y (nx6906), .A0 (inputs_58__1), .A1 (inputs_59__1), .S0 (
             nx23979)) ;
    mux21_ni ix6939 (.Y (nx6938), .A0 (nx6922), .A1 (nx6934), .S0 (nx23413)) ;
    mux21_ni ix6923 (.Y (nx6922), .A0 (inputs_60__1), .A1 (inputs_61__1), .S0 (
             nx23979)) ;
    mux21_ni ix6935 (.Y (nx6934), .A0 (inputs_62__1), .A1 (inputs_63__1), .S0 (
             nx23979)) ;
    mux21_ni ix7455 (.Y (nx7454), .A0 (nx7242), .A1 (nx7450), .S0 (nx22543)) ;
    mux21_ni ix7243 (.Y (nx7242), .A0 (nx7236), .A1 (nx7158), .S0 (nx23123)) ;
    oai21 ix7237 (.Y (nx7236), .A0 (nx22241), .A1 (nx9753), .B0 (nx9763)) ;
    mux21 ix9754 (.Y (nx9753), .A0 (nx7200), .A1 (nx7228), .S0 (nx22725)) ;
    mux21_ni ix7201 (.Y (nx7200), .A0 (nx7184), .A1 (nx7196), .S0 (nx23413)) ;
    mux21_ni ix7185 (.Y (nx7184), .A0 (inputs_68__1), .A1 (inputs_69__1), .S0 (
             nx23979)) ;
    mux21_ni ix7197 (.Y (nx7196), .A0 (inputs_70__1), .A1 (inputs_71__1), .S0 (
             nx23979)) ;
    mux21_ni ix7229 (.Y (nx7228), .A0 (nx7212), .A1 (nx7224), .S0 (nx23413)) ;
    mux21_ni ix7213 (.Y (nx7212), .A0 (inputs_84__1), .A1 (inputs_85__1), .S0 (
             nx23979)) ;
    mux21_ni ix7225 (.Y (nx7224), .A0 (inputs_86__1), .A1 (inputs_87__1), .S0 (
             nx23981)) ;
    nand04 ix9764 (.Y (nx9763), .A0 (nx22241), .A1 (nx23413), .A2 (nx23981), .A3 (
           nx7172)) ;
    mux21_ni ix7173 (.Y (nx7172), .A0 (inputs_67__1), .A1 (inputs_83__1), .S0 (
             nx22727)) ;
    mux21_ni ix7159 (.Y (nx7158), .A0 (nx7094), .A1 (nx7154), .S0 (nx22727)) ;
    mux21_ni ix7095 (.Y (nx7094), .A0 (nx7062), .A1 (nx7090), .S0 (nx23205)) ;
    mux21_ni ix7063 (.Y (nx7062), .A0 (nx7046), .A1 (nx7058), .S0 (nx23415)) ;
    mux21_ni ix7047 (.Y (nx7046), .A0 (inputs_72__1), .A1 (inputs_73__1), .S0 (
             nx23981)) ;
    mux21_ni ix7059 (.Y (nx7058), .A0 (inputs_74__1), .A1 (inputs_75__1), .S0 (
             nx23981)) ;
    mux21_ni ix7091 (.Y (nx7090), .A0 (nx7074), .A1 (nx7086), .S0 (nx23415)) ;
    mux21_ni ix7075 (.Y (nx7074), .A0 (inputs_76__1), .A1 (inputs_77__1), .S0 (
             nx23981)) ;
    mux21_ni ix7087 (.Y (nx7086), .A0 (inputs_78__1), .A1 (inputs_79__1), .S0 (
             nx23981)) ;
    mux21_ni ix7155 (.Y (nx7154), .A0 (nx7122), .A1 (nx7150), .S0 (nx23205)) ;
    mux21_ni ix7123 (.Y (nx7122), .A0 (nx7106), .A1 (nx7118), .S0 (nx23415)) ;
    mux21_ni ix7107 (.Y (nx7106), .A0 (inputs_88__1), .A1 (inputs_89__1), .S0 (
             nx23981)) ;
    mux21_ni ix7119 (.Y (nx7118), .A0 (inputs_90__1), .A1 (inputs_91__1), .S0 (
             nx23983)) ;
    mux21_ni ix7151 (.Y (nx7150), .A0 (nx7134), .A1 (nx7146), .S0 (nx23415)) ;
    mux21_ni ix7135 (.Y (nx7134), .A0 (inputs_92__1), .A1 (inputs_93__1), .S0 (
             nx23983)) ;
    mux21_ni ix7147 (.Y (nx7146), .A0 (inputs_94__1), .A1 (inputs_95__1), .S0 (
             nx23983)) ;
    mux21_ni ix7451 (.Y (nx7450), .A0 (nx7444), .A1 (nx7366), .S0 (nx23123)) ;
    oai21 ix7445 (.Y (nx7444), .A0 (nx22243), .A1 (nx9795), .B0 (nx9805)) ;
    mux21 ix9796 (.Y (nx9795), .A0 (nx7408), .A1 (nx7436), .S0 (nx22727)) ;
    mux21_ni ix7409 (.Y (nx7408), .A0 (nx7392), .A1 (nx7404), .S0 (nx23415)) ;
    mux21_ni ix7393 (.Y (nx7392), .A0 (inputs_100__1), .A1 (inputs_101__1), .S0 (
             nx23983)) ;
    mux21_ni ix7405 (.Y (nx7404), .A0 (inputs_102__1), .A1 (inputs_103__1), .S0 (
             nx23983)) ;
    mux21_ni ix7437 (.Y (nx7436), .A0 (nx7420), .A1 (nx7432), .S0 (nx23415)) ;
    mux21_ni ix7421 (.Y (nx7420), .A0 (inputs_116__1), .A1 (inputs_117__1), .S0 (
             nx23983)) ;
    mux21_ni ix7433 (.Y (nx7432), .A0 (inputs_118__1), .A1 (inputs_119__1), .S0 (
             nx23983)) ;
    nand04 ix9806 (.Y (nx9805), .A0 (nx22243), .A1 (nx23415), .A2 (nx23985), .A3 (
           nx7380)) ;
    mux21_ni ix7381 (.Y (nx7380), .A0 (inputs_99__1), .A1 (inputs_115__1), .S0 (
             nx22727)) ;
    mux21_ni ix7367 (.Y (nx7366), .A0 (nx7302), .A1 (nx7362), .S0 (nx22727)) ;
    mux21_ni ix7303 (.Y (nx7302), .A0 (nx7270), .A1 (nx7298), .S0 (nx23205)) ;
    mux21_ni ix7271 (.Y (nx7270), .A0 (nx7254), .A1 (nx7266), .S0 (nx23417)) ;
    mux21_ni ix7255 (.Y (nx7254), .A0 (inputs_104__1), .A1 (inputs_105__1), .S0 (
             nx23985)) ;
    mux21_ni ix7267 (.Y (nx7266), .A0 (inputs_106__1), .A1 (inputs_107__1), .S0 (
             nx23985)) ;
    mux21_ni ix7299 (.Y (nx7298), .A0 (nx7282), .A1 (nx7294), .S0 (nx23417)) ;
    mux21_ni ix7283 (.Y (nx7282), .A0 (inputs_108__1), .A1 (inputs_109__1), .S0 (
             nx23985)) ;
    mux21_ni ix7295 (.Y (nx7294), .A0 (inputs_110__1), .A1 (inputs_111__1), .S0 (
             nx23985)) ;
    mux21_ni ix7363 (.Y (nx7362), .A0 (nx7330), .A1 (nx7358), .S0 (nx23205)) ;
    mux21_ni ix7331 (.Y (nx7330), .A0 (nx7314), .A1 (nx7326), .S0 (nx23417)) ;
    mux21_ni ix7315 (.Y (nx7314), .A0 (inputs_120__1), .A1 (inputs_121__1), .S0 (
             nx23985)) ;
    mux21_ni ix7327 (.Y (nx7326), .A0 (inputs_122__1), .A1 (inputs_123__1), .S0 (
             nx23985)) ;
    mux21_ni ix7359 (.Y (nx7358), .A0 (nx7342), .A1 (nx7354), .S0 (nx23417)) ;
    mux21_ni ix7343 (.Y (nx7342), .A0 (inputs_124__1), .A1 (inputs_125__1), .S0 (
             nx23987)) ;
    mux21_ni ix7355 (.Y (nx7354), .A0 (inputs_126__1), .A1 (inputs_127__1), .S0 (
             nx23987)) ;
    mux21_ni ix8303 (.Y (nx8302), .A0 (nx7878), .A1 (nx8298), .S0 (nx22459)) ;
    mux21_ni ix7879 (.Y (nx7878), .A0 (nx7666), .A1 (nx7874), .S0 (nx22543)) ;
    mux21_ni ix7667 (.Y (nx7666), .A0 (nx7660), .A1 (nx7582), .S0 (nx23125)) ;
    oai21 ix7661 (.Y (nx7660), .A0 (nx22243), .A1 (nx9839), .B0 (nx9851)) ;
    mux21 ix9840 (.Y (nx9839), .A0 (nx7624), .A1 (nx7652), .S0 (nx22727)) ;
    mux21_ni ix7625 (.Y (nx7624), .A0 (nx7608), .A1 (nx7620), .S0 (nx23417)) ;
    mux21_ni ix7609 (.Y (nx7608), .A0 (inputs_132__1), .A1 (inputs_133__1), .S0 (
             nx23987)) ;
    mux21_ni ix7621 (.Y (nx7620), .A0 (inputs_134__1), .A1 (inputs_135__1), .S0 (
             nx23987)) ;
    mux21_ni ix7653 (.Y (nx7652), .A0 (nx7636), .A1 (nx7648), .S0 (nx23417)) ;
    mux21_ni ix7637 (.Y (nx7636), .A0 (inputs_148__1), .A1 (inputs_149__1), .S0 (
             nx23987)) ;
    mux21_ni ix7649 (.Y (nx7648), .A0 (inputs_150__1), .A1 (inputs_151__1), .S0 (
             nx23987)) ;
    nand04 ix9852 (.Y (nx9851), .A0 (nx22243), .A1 (nx23417), .A2 (nx23987), .A3 (
           nx7596)) ;
    mux21_ni ix7597 (.Y (nx7596), .A0 (inputs_131__1), .A1 (inputs_147__1), .S0 (
             nx22727)) ;
    mux21_ni ix7583 (.Y (nx7582), .A0 (nx7518), .A1 (nx7578), .S0 (nx22729)) ;
    mux21_ni ix7519 (.Y (nx7518), .A0 (nx7486), .A1 (nx7514), .S0 (nx23207)) ;
    mux21_ni ix7487 (.Y (nx7486), .A0 (nx7470), .A1 (nx7482), .S0 (nx23419)) ;
    mux21_ni ix7471 (.Y (nx7470), .A0 (inputs_136__1), .A1 (inputs_137__1), .S0 (
             nx23989)) ;
    mux21_ni ix7483 (.Y (nx7482), .A0 (inputs_138__1), .A1 (inputs_139__1), .S0 (
             nx23989)) ;
    mux21_ni ix7515 (.Y (nx7514), .A0 (nx7498), .A1 (nx7510), .S0 (nx23419)) ;
    mux21_ni ix7499 (.Y (nx7498), .A0 (inputs_140__1), .A1 (inputs_141__1), .S0 (
             nx23989)) ;
    mux21_ni ix7511 (.Y (nx7510), .A0 (inputs_142__1), .A1 (inputs_143__1), .S0 (
             nx23989)) ;
    mux21_ni ix7579 (.Y (nx7578), .A0 (nx7546), .A1 (nx7574), .S0 (nx23207)) ;
    mux21_ni ix7547 (.Y (nx7546), .A0 (nx7530), .A1 (nx7542), .S0 (nx23419)) ;
    mux21_ni ix7531 (.Y (nx7530), .A0 (inputs_152__1), .A1 (inputs_153__1), .S0 (
             nx23989)) ;
    mux21_ni ix7543 (.Y (nx7542), .A0 (inputs_154__1), .A1 (inputs_155__1), .S0 (
             nx23989)) ;
    mux21_ni ix7575 (.Y (nx7574), .A0 (nx7558), .A1 (nx7570), .S0 (nx23419)) ;
    mux21_ni ix7559 (.Y (nx7558), .A0 (inputs_156__1), .A1 (inputs_157__1), .S0 (
             nx23989)) ;
    mux21_ni ix7571 (.Y (nx7570), .A0 (inputs_158__1), .A1 (inputs_159__1), .S0 (
             nx23991)) ;
    mux21_ni ix7875 (.Y (nx7874), .A0 (nx7868), .A1 (nx7790), .S0 (nx23125)) ;
    oai21 ix7869 (.Y (nx7868), .A0 (nx22243), .A1 (nx9881), .B0 (nx9891)) ;
    mux21 ix9882 (.Y (nx9881), .A0 (nx7832), .A1 (nx7860), .S0 (nx22729)) ;
    mux21_ni ix7833 (.Y (nx7832), .A0 (nx7816), .A1 (nx7828), .S0 (nx23419)) ;
    mux21_ni ix7817 (.Y (nx7816), .A0 (inputs_164__1), .A1 (inputs_165__1), .S0 (
             nx23991)) ;
    mux21_ni ix7829 (.Y (nx7828), .A0 (inputs_166__1), .A1 (inputs_167__1), .S0 (
             nx23991)) ;
    mux21_ni ix7861 (.Y (nx7860), .A0 (nx7844), .A1 (nx7856), .S0 (nx23419)) ;
    mux21_ni ix7845 (.Y (nx7844), .A0 (inputs_180__1), .A1 (inputs_181__1), .S0 (
             nx23991)) ;
    mux21_ni ix7857 (.Y (nx7856), .A0 (inputs_182__1), .A1 (inputs_183__1), .S0 (
             nx23991)) ;
    nand04 ix9892 (.Y (nx9891), .A0 (nx22243), .A1 (nx23419), .A2 (nx23991), .A3 (
           nx7804)) ;
    mux21_ni ix7805 (.Y (nx7804), .A0 (inputs_163__1), .A1 (inputs_179__1), .S0 (
             nx22729)) ;
    mux21_ni ix7791 (.Y (nx7790), .A0 (nx7726), .A1 (nx7786), .S0 (nx22729)) ;
    mux21_ni ix7727 (.Y (nx7726), .A0 (nx7694), .A1 (nx7722), .S0 (nx23207)) ;
    mux21_ni ix7695 (.Y (nx7694), .A0 (nx7678), .A1 (nx7690), .S0 (nx23421)) ;
    mux21_ni ix7679 (.Y (nx7678), .A0 (inputs_168__1), .A1 (inputs_169__1), .S0 (
             nx23991)) ;
    mux21_ni ix7691 (.Y (nx7690), .A0 (inputs_170__1), .A1 (inputs_171__1), .S0 (
             nx23993)) ;
    mux21_ni ix7723 (.Y (nx7722), .A0 (nx7706), .A1 (nx7718), .S0 (nx23421)) ;
    mux21_ni ix7707 (.Y (nx7706), .A0 (inputs_172__1), .A1 (inputs_173__1), .S0 (
             nx23993)) ;
    mux21_ni ix7719 (.Y (nx7718), .A0 (inputs_174__1), .A1 (inputs_175__1), .S0 (
             nx23993)) ;
    mux21_ni ix7787 (.Y (nx7786), .A0 (nx7754), .A1 (nx7782), .S0 (nx23207)) ;
    mux21_ni ix7755 (.Y (nx7754), .A0 (nx7738), .A1 (nx7750), .S0 (nx23421)) ;
    mux21_ni ix7739 (.Y (nx7738), .A0 (inputs_184__1), .A1 (inputs_185__1), .S0 (
             nx23993)) ;
    mux21_ni ix7751 (.Y (nx7750), .A0 (inputs_186__1), .A1 (inputs_187__1), .S0 (
             nx23993)) ;
    mux21_ni ix7783 (.Y (nx7782), .A0 (nx7766), .A1 (nx7778), .S0 (nx23421)) ;
    mux21_ni ix7767 (.Y (nx7766), .A0 (inputs_188__1), .A1 (inputs_189__1), .S0 (
             nx23993)) ;
    mux21_ni ix7779 (.Y (nx7778), .A0 (inputs_190__1), .A1 (inputs_191__1), .S0 (
             nx23993)) ;
    mux21_ni ix8299 (.Y (nx8298), .A0 (nx8086), .A1 (nx8294), .S0 (nx22545)) ;
    mux21_ni ix8087 (.Y (nx8086), .A0 (nx8080), .A1 (nx8002), .S0 (nx23125)) ;
    oai21 ix8081 (.Y (nx8080), .A0 (nx22243), .A1 (nx9927), .B0 (nx9939)) ;
    mux21 ix9928 (.Y (nx9927), .A0 (nx8044), .A1 (nx8072), .S0 (nx22729)) ;
    mux21_ni ix8045 (.Y (nx8044), .A0 (nx8028), .A1 (nx8040), .S0 (nx23421)) ;
    mux21_ni ix8029 (.Y (nx8028), .A0 (inputs_196__1), .A1 (inputs_197__1), .S0 (
             nx23995)) ;
    mux21_ni ix8041 (.Y (nx8040), .A0 (inputs_198__1), .A1 (inputs_199__1), .S0 (
             nx23995)) ;
    mux21_ni ix8073 (.Y (nx8072), .A0 (nx8056), .A1 (nx8068), .S0 (nx23421)) ;
    mux21_ni ix8057 (.Y (nx8056), .A0 (inputs_212__1), .A1 (inputs_213__1), .S0 (
             nx23995)) ;
    mux21_ni ix8069 (.Y (nx8068), .A0 (inputs_214__1), .A1 (inputs_215__1), .S0 (
             nx23995)) ;
    nand04 ix9940 (.Y (nx9939), .A0 (nx22245), .A1 (nx23421), .A2 (nx23995), .A3 (
           nx8016)) ;
    mux21_ni ix8017 (.Y (nx8016), .A0 (inputs_195__1), .A1 (inputs_211__1), .S0 (
             nx22729)) ;
    mux21_ni ix8003 (.Y (nx8002), .A0 (nx7938), .A1 (nx7998), .S0 (nx22729)) ;
    mux21_ni ix7939 (.Y (nx7938), .A0 (nx7906), .A1 (nx7934), .S0 (nx23207)) ;
    mux21_ni ix7907 (.Y (nx7906), .A0 (nx7890), .A1 (nx7902), .S0 (nx23423)) ;
    mux21_ni ix7891 (.Y (nx7890), .A0 (inputs_200__1), .A1 (inputs_201__1), .S0 (
             nx23995)) ;
    mux21_ni ix7903 (.Y (nx7902), .A0 (inputs_202__1), .A1 (inputs_203__1), .S0 (
             nx23995)) ;
    mux21_ni ix7935 (.Y (nx7934), .A0 (nx7918), .A1 (nx7930), .S0 (nx23423)) ;
    mux21_ni ix7919 (.Y (nx7918), .A0 (inputs_204__1), .A1 (inputs_205__1), .S0 (
             nx23997)) ;
    mux21_ni ix7931 (.Y (nx7930), .A0 (inputs_206__1), .A1 (inputs_207__1), .S0 (
             nx23997)) ;
    mux21_ni ix7999 (.Y (nx7998), .A0 (nx7966), .A1 (nx7994), .S0 (nx23207)) ;
    mux21_ni ix7967 (.Y (nx7966), .A0 (nx7950), .A1 (nx7962), .S0 (nx23423)) ;
    mux21_ni ix7951 (.Y (nx7950), .A0 (inputs_216__1), .A1 (inputs_217__1), .S0 (
             nx23997)) ;
    mux21_ni ix7963 (.Y (nx7962), .A0 (inputs_218__1), .A1 (inputs_219__1), .S0 (
             nx23997)) ;
    mux21_ni ix7995 (.Y (nx7994), .A0 (nx7978), .A1 (nx7990), .S0 (nx23423)) ;
    mux21_ni ix7979 (.Y (nx7978), .A0 (inputs_220__1), .A1 (inputs_221__1), .S0 (
             nx23997)) ;
    mux21_ni ix7991 (.Y (nx7990), .A0 (inputs_222__1), .A1 (inputs_223__1), .S0 (
             nx23997)) ;
    mux21_ni ix8295 (.Y (nx8294), .A0 (nx8288), .A1 (nx8210), .S0 (nx23125)) ;
    oai21 ix8289 (.Y (nx8288), .A0 (nx22245), .A1 (nx9969), .B0 (nx9983)) ;
    mux21 ix9970 (.Y (nx9969), .A0 (nx8252), .A1 (nx8280), .S0 (nx22731)) ;
    mux21_ni ix8253 (.Y (nx8252), .A0 (nx8236), .A1 (nx8248), .S0 (nx23423)) ;
    mux21_ni ix8237 (.Y (nx8236), .A0 (inputs_228__1), .A1 (inputs_229__1), .S0 (
             nx23997)) ;
    mux21_ni ix8249 (.Y (nx8248), .A0 (inputs_230__1), .A1 (inputs_231__1), .S0 (
             nx23999)) ;
    mux21_ni ix8281 (.Y (nx8280), .A0 (nx8264), .A1 (nx8276), .S0 (nx23423)) ;
    mux21_ni ix8265 (.Y (nx8264), .A0 (inputs_244__1), .A1 (inputs_245__1), .S0 (
             nx23999)) ;
    mux21_ni ix8277 (.Y (nx8276), .A0 (inputs_246__1), .A1 (inputs_247__1), .S0 (
             nx23999)) ;
    nand04 ix9984 (.Y (nx9983), .A0 (nx22245), .A1 (nx23423), .A2 (nx23999), .A3 (
           nx8224)) ;
    mux21_ni ix8225 (.Y (nx8224), .A0 (inputs_227__1), .A1 (inputs_243__1), .S0 (
             nx22731)) ;
    mux21_ni ix8211 (.Y (nx8210), .A0 (nx8146), .A1 (nx8206), .S0 (nx22731)) ;
    mux21_ni ix8147 (.Y (nx8146), .A0 (nx8114), .A1 (nx8142), .S0 (nx23207)) ;
    mux21_ni ix8115 (.Y (nx8114), .A0 (nx8098), .A1 (nx8110), .S0 (nx23425)) ;
    mux21_ni ix8099 (.Y (nx8098), .A0 (inputs_232__1), .A1 (inputs_233__1), .S0 (
             nx23999)) ;
    mux21_ni ix8111 (.Y (nx8110), .A0 (inputs_234__1), .A1 (inputs_235__1), .S0 (
             nx23999)) ;
    mux21_ni ix8143 (.Y (nx8142), .A0 (nx8126), .A1 (nx8138), .S0 (nx23425)) ;
    mux21_ni ix8127 (.Y (nx8126), .A0 (inputs_236__1), .A1 (inputs_237__1), .S0 (
             nx23999)) ;
    mux21_ni ix8139 (.Y (nx8138), .A0 (inputs_238__1), .A1 (inputs_239__1), .S0 (
             nx24001)) ;
    mux21_ni ix8207 (.Y (nx8206), .A0 (nx8174), .A1 (nx8202), .S0 (nx23209)) ;
    mux21_ni ix8175 (.Y (nx8174), .A0 (nx8158), .A1 (nx8170), .S0 (nx23425)) ;
    mux21_ni ix8159 (.Y (nx8158), .A0 (inputs_248__1), .A1 (inputs_249__1), .S0 (
             nx24001)) ;
    mux21_ni ix8171 (.Y (nx8170), .A0 (inputs_250__1), .A1 (inputs_251__1), .S0 (
             nx24001)) ;
    mux21_ni ix8203 (.Y (nx8202), .A0 (nx8186), .A1 (nx8198), .S0 (nx23425)) ;
    mux21_ni ix8187 (.Y (nx8186), .A0 (inputs_252__1), .A1 (inputs_253__1), .S0 (
             nx24001)) ;
    mux21_ni ix8199 (.Y (nx8198), .A0 (inputs_254__1), .A1 (inputs_255__1), .S0 (
             nx24001)) ;
    oai21 ix12473 (.Y (\output [2]), .A0 (nx24851), .A1 (nx10015), .B0 (nx10375)
          ) ;
    mux21 ix10016 (.Y (nx10015), .A0 (nx9154), .A1 (nx9998), .S0 (nx22415)) ;
    mux21_ni ix9155 (.Y (nx9154), .A0 (nx8730), .A1 (nx9150), .S0 (nx22459)) ;
    mux21_ni ix8731 (.Y (nx8730), .A0 (nx8518), .A1 (nx8726), .S0 (nx22545)) ;
    mux21_ni ix8519 (.Y (nx8518), .A0 (nx8512), .A1 (nx8434), .S0 (nx23125)) ;
    oai21 ix8513 (.Y (nx8512), .A0 (nx22245), .A1 (nx10023), .B0 (nx10035)) ;
    mux21 ix10024 (.Y (nx10023), .A0 (nx8476), .A1 (nx8504), .S0 (nx22731)) ;
    mux21_ni ix8477 (.Y (nx8476), .A0 (nx8460), .A1 (nx8472), .S0 (nx23425)) ;
    mux21_ni ix8461 (.Y (nx8460), .A0 (inputs_260__2), .A1 (inputs_261__2), .S0 (
             nx24001)) ;
    mux21_ni ix8473 (.Y (nx8472), .A0 (inputs_262__2), .A1 (inputs_263__2), .S0 (
             nx24001)) ;
    mux21_ni ix8505 (.Y (nx8504), .A0 (nx8488), .A1 (nx8500), .S0 (nx23425)) ;
    mux21_ni ix8489 (.Y (nx8488), .A0 (inputs_276__2), .A1 (inputs_277__2), .S0 (
             nx24003)) ;
    mux21_ni ix8501 (.Y (nx8500), .A0 (inputs_278__2), .A1 (inputs_279__2), .S0 (
             nx24003)) ;
    nand04 ix10036 (.Y (nx10035), .A0 (nx22245), .A1 (nx23425), .A2 (nx24003), .A3 (
           nx8448)) ;
    mux21_ni ix8449 (.Y (nx8448), .A0 (inputs_259__2), .A1 (inputs_275__2), .S0 (
             nx22731)) ;
    mux21_ni ix8435 (.Y (nx8434), .A0 (nx8370), .A1 (nx8430), .S0 (nx22731)) ;
    mux21_ni ix8371 (.Y (nx8370), .A0 (nx8338), .A1 (nx8366), .S0 (nx23209)) ;
    mux21_ni ix8339 (.Y (nx8338), .A0 (nx8322), .A1 (nx8334), .S0 (nx23427)) ;
    mux21_ni ix8323 (.Y (nx8322), .A0 (inputs_264__2), .A1 (inputs_265__2), .S0 (
             nx24003)) ;
    mux21_ni ix8335 (.Y (nx8334), .A0 (inputs_266__2), .A1 (inputs_267__2), .S0 (
             nx24003)) ;
    mux21_ni ix8367 (.Y (nx8366), .A0 (nx8350), .A1 (nx8362), .S0 (nx23427)) ;
    mux21_ni ix8351 (.Y (nx8350), .A0 (inputs_268__2), .A1 (inputs_269__2), .S0 (
             nx24003)) ;
    mux21_ni ix8363 (.Y (nx8362), .A0 (inputs_270__2), .A1 (inputs_271__2), .S0 (
             nx24003)) ;
    mux21_ni ix8431 (.Y (nx8430), .A0 (nx8398), .A1 (nx8426), .S0 (nx23209)) ;
    mux21_ni ix8399 (.Y (nx8398), .A0 (nx8382), .A1 (nx8394), .S0 (nx23427)) ;
    mux21_ni ix8383 (.Y (nx8382), .A0 (inputs_280__2), .A1 (inputs_281__2), .S0 (
             nx24005)) ;
    mux21_ni ix8395 (.Y (nx8394), .A0 (inputs_282__2), .A1 (inputs_283__2), .S0 (
             nx24005)) ;
    mux21_ni ix8427 (.Y (nx8426), .A0 (nx8410), .A1 (nx8422), .S0 (nx23427)) ;
    mux21_ni ix8411 (.Y (nx8410), .A0 (inputs_284__2), .A1 (inputs_285__2), .S0 (
             nx24005)) ;
    mux21_ni ix8423 (.Y (nx8422), .A0 (inputs_286__2), .A1 (inputs_287__2), .S0 (
             nx24005)) ;
    mux21_ni ix8727 (.Y (nx8726), .A0 (nx8720), .A1 (nx8642), .S0 (nx23125)) ;
    oai21 ix8721 (.Y (nx8720), .A0 (nx22245), .A1 (nx10067), .B0 (nx10079)) ;
    mux21 ix10068 (.Y (nx10067), .A0 (nx8684), .A1 (nx8712), .S0 (nx22731)) ;
    mux21_ni ix8685 (.Y (nx8684), .A0 (nx8668), .A1 (nx8680), .S0 (nx23427)) ;
    mux21_ni ix8669 (.Y (nx8668), .A0 (inputs_292__2), .A1 (inputs_293__2), .S0 (
             nx24005)) ;
    mux21_ni ix8681 (.Y (nx8680), .A0 (inputs_294__2), .A1 (inputs_295__2), .S0 (
             nx24005)) ;
    mux21_ni ix8713 (.Y (nx8712), .A0 (nx8696), .A1 (nx8708), .S0 (nx23427)) ;
    mux21_ni ix8697 (.Y (nx8696), .A0 (inputs_308__2), .A1 (inputs_309__2), .S0 (
             nx24005)) ;
    mux21_ni ix8709 (.Y (nx8708), .A0 (inputs_310__2), .A1 (inputs_311__2), .S0 (
             nx24007)) ;
    nand04 ix10080 (.Y (nx10079), .A0 (nx22245), .A1 (nx23427), .A2 (nx24007), .A3 (
           nx8656)) ;
    mux21_ni ix8657 (.Y (nx8656), .A0 (inputs_291__2), .A1 (inputs_307__2), .S0 (
             nx22733)) ;
    mux21_ni ix8643 (.Y (nx8642), .A0 (nx8578), .A1 (nx8638), .S0 (nx22733)) ;
    mux21_ni ix8579 (.Y (nx8578), .A0 (nx8546), .A1 (nx8574), .S0 (nx23209)) ;
    mux21_ni ix8547 (.Y (nx8546), .A0 (nx8530), .A1 (nx8542), .S0 (nx23429)) ;
    mux21_ni ix8531 (.Y (nx8530), .A0 (inputs_296__2), .A1 (inputs_297__2), .S0 (
             nx24007)) ;
    mux21_ni ix8543 (.Y (nx8542), .A0 (inputs_298__2), .A1 (inputs_299__2), .S0 (
             nx24007)) ;
    mux21_ni ix8575 (.Y (nx8574), .A0 (nx8558), .A1 (nx8570), .S0 (nx23429)) ;
    mux21_ni ix8559 (.Y (nx8558), .A0 (inputs_300__2), .A1 (inputs_301__2), .S0 (
             nx24007)) ;
    mux21_ni ix8571 (.Y (nx8570), .A0 (inputs_302__2), .A1 (inputs_303__2), .S0 (
             nx24007)) ;
    mux21_ni ix8639 (.Y (nx8638), .A0 (nx8606), .A1 (nx8634), .S0 (nx23209)) ;
    mux21_ni ix8607 (.Y (nx8606), .A0 (nx8590), .A1 (nx8602), .S0 (nx23429)) ;
    mux21_ni ix8591 (.Y (nx8590), .A0 (inputs_312__2), .A1 (inputs_313__2), .S0 (
             nx24007)) ;
    mux21_ni ix8603 (.Y (nx8602), .A0 (inputs_314__2), .A1 (inputs_315__2), .S0 (
             nx24009)) ;
    mux21_ni ix8635 (.Y (nx8634), .A0 (nx8618), .A1 (nx8630), .S0 (nx23429)) ;
    mux21_ni ix8619 (.Y (nx8618), .A0 (inputs_316__2), .A1 (inputs_317__2), .S0 (
             nx24009)) ;
    mux21_ni ix8631 (.Y (nx8630), .A0 (inputs_318__2), .A1 (inputs_319__2), .S0 (
             nx24009)) ;
    mux21_ni ix9151 (.Y (nx9150), .A0 (nx8938), .A1 (nx9146), .S0 (nx22545)) ;
    mux21_ni ix8939 (.Y (nx8938), .A0 (nx8932), .A1 (nx8854), .S0 (nx23125)) ;
    oai21 ix8933 (.Y (nx8932), .A0 (nx22247), .A1 (nx10111), .B0 (nx10125)) ;
    mux21 ix10112 (.Y (nx10111), .A0 (nx8896), .A1 (nx8924), .S0 (nx22733)) ;
    mux21_ni ix8897 (.Y (nx8896), .A0 (nx8880), .A1 (nx8892), .S0 (nx23429)) ;
    mux21_ni ix8881 (.Y (nx8880), .A0 (inputs_324__2), .A1 (inputs_325__2), .S0 (
             nx24009)) ;
    mux21_ni ix8893 (.Y (nx8892), .A0 (inputs_326__2), .A1 (inputs_327__2), .S0 (
             nx24009)) ;
    mux21_ni ix8925 (.Y (nx8924), .A0 (nx8908), .A1 (nx8920), .S0 (nx23429)) ;
    mux21_ni ix8909 (.Y (nx8908), .A0 (inputs_340__2), .A1 (inputs_341__2), .S0 (
             nx24009)) ;
    mux21_ni ix8921 (.Y (nx8920), .A0 (inputs_342__2), .A1 (inputs_343__2), .S0 (
             nx24009)) ;
    nand04 ix10126 (.Y (nx10125), .A0 (nx22247), .A1 (nx23429), .A2 (nx24011), .A3 (
           nx8868)) ;
    mux21_ni ix8869 (.Y (nx8868), .A0 (inputs_323__2), .A1 (inputs_339__2), .S0 (
             nx22733)) ;
    mux21_ni ix8855 (.Y (nx8854), .A0 (nx8790), .A1 (nx8850), .S0 (nx22733)) ;
    mux21_ni ix8791 (.Y (nx8790), .A0 (nx8758), .A1 (nx8786), .S0 (nx23209)) ;
    mux21_ni ix8759 (.Y (nx8758), .A0 (nx8742), .A1 (nx8754), .S0 (nx23431)) ;
    mux21_ni ix8743 (.Y (nx8742), .A0 (inputs_328__2), .A1 (inputs_329__2), .S0 (
             nx24011)) ;
    mux21_ni ix8755 (.Y (nx8754), .A0 (inputs_330__2), .A1 (inputs_331__2), .S0 (
             nx24011)) ;
    mux21_ni ix8787 (.Y (nx8786), .A0 (nx8770), .A1 (nx8782), .S0 (nx23431)) ;
    mux21_ni ix8771 (.Y (nx8770), .A0 (inputs_332__2), .A1 (inputs_333__2), .S0 (
             nx24011)) ;
    mux21_ni ix8783 (.Y (nx8782), .A0 (inputs_334__2), .A1 (inputs_335__2), .S0 (
             nx24011)) ;
    mux21_ni ix8851 (.Y (nx8850), .A0 (nx8818), .A1 (nx8846), .S0 (nx23209)) ;
    mux21_ni ix8819 (.Y (nx8818), .A0 (nx8802), .A1 (nx8814), .S0 (nx23431)) ;
    mux21_ni ix8803 (.Y (nx8802), .A0 (inputs_344__2), .A1 (inputs_345__2), .S0 (
             nx24011)) ;
    mux21_ni ix8815 (.Y (nx8814), .A0 (inputs_346__2), .A1 (inputs_347__2), .S0 (
             nx24011)) ;
    mux21_ni ix8847 (.Y (nx8846), .A0 (nx8830), .A1 (nx8842), .S0 (nx23431)) ;
    mux21_ni ix8831 (.Y (nx8830), .A0 (inputs_348__2), .A1 (inputs_349__2), .S0 (
             nx24013)) ;
    mux21_ni ix8843 (.Y (nx8842), .A0 (inputs_350__2), .A1 (inputs_351__2), .S0 (
             nx24013)) ;
    mux21_ni ix9147 (.Y (nx9146), .A0 (nx9140), .A1 (nx9062), .S0 (nx23127)) ;
    oai21 ix9141 (.Y (nx9140), .A0 (nx22247), .A1 (nx10155), .B0 (nx10167)) ;
    mux21 ix10156 (.Y (nx10155), .A0 (nx9104), .A1 (nx9132), .S0 (nx22733)) ;
    mux21_ni ix9105 (.Y (nx9104), .A0 (nx9088), .A1 (nx9100), .S0 (nx23431)) ;
    mux21_ni ix9089 (.Y (nx9088), .A0 (inputs_356__2), .A1 (inputs_357__2), .S0 (
             nx24013)) ;
    mux21_ni ix9101 (.Y (nx9100), .A0 (inputs_358__2), .A1 (inputs_359__2), .S0 (
             nx24013)) ;
    mux21_ni ix9133 (.Y (nx9132), .A0 (nx9116), .A1 (nx9128), .S0 (nx23431)) ;
    mux21_ni ix9117 (.Y (nx9116), .A0 (inputs_372__2), .A1 (inputs_373__2), .S0 (
             nx24013)) ;
    mux21_ni ix9129 (.Y (nx9128), .A0 (inputs_374__2), .A1 (inputs_375__2), .S0 (
             nx24013)) ;
    nand04 ix10168 (.Y (nx10167), .A0 (nx22247), .A1 (nx23431), .A2 (nx24013), .A3 (
           nx9076)) ;
    mux21_ni ix9077 (.Y (nx9076), .A0 (inputs_355__2), .A1 (inputs_371__2), .S0 (
             nx22733)) ;
    mux21_ni ix9063 (.Y (nx9062), .A0 (nx8998), .A1 (nx9058), .S0 (nx22735)) ;
    mux21_ni ix8999 (.Y (nx8998), .A0 (nx8966), .A1 (nx8994), .S0 (nx23211)) ;
    mux21_ni ix8967 (.Y (nx8966), .A0 (nx8950), .A1 (nx8962), .S0 (nx23433)) ;
    mux21_ni ix8951 (.Y (nx8950), .A0 (inputs_360__2), .A1 (inputs_361__2), .S0 (
             nx24015)) ;
    mux21_ni ix8963 (.Y (nx8962), .A0 (inputs_362__2), .A1 (inputs_363__2), .S0 (
             nx24015)) ;
    mux21_ni ix8995 (.Y (nx8994), .A0 (nx8978), .A1 (nx8990), .S0 (nx23433)) ;
    mux21_ni ix8979 (.Y (nx8978), .A0 (inputs_364__2), .A1 (inputs_365__2), .S0 (
             nx24015)) ;
    mux21_ni ix8991 (.Y (nx8990), .A0 (inputs_366__2), .A1 (inputs_367__2), .S0 (
             nx24015)) ;
    mux21_ni ix9059 (.Y (nx9058), .A0 (nx9026), .A1 (nx9054), .S0 (nx23211)) ;
    mux21_ni ix9027 (.Y (nx9026), .A0 (nx9010), .A1 (nx9022), .S0 (nx23433)) ;
    mux21_ni ix9011 (.Y (nx9010), .A0 (inputs_376__2), .A1 (inputs_377__2), .S0 (
             nx24015)) ;
    mux21_ni ix9023 (.Y (nx9022), .A0 (inputs_378__2), .A1 (inputs_379__2), .S0 (
             nx24015)) ;
    mux21_ni ix9055 (.Y (nx9054), .A0 (nx9038), .A1 (nx9050), .S0 (nx23433)) ;
    mux21_ni ix9039 (.Y (nx9038), .A0 (inputs_380__2), .A1 (inputs_381__2), .S0 (
             nx24015)) ;
    mux21_ni ix9051 (.Y (nx9050), .A0 (inputs_382__2), .A1 (inputs_383__2), .S0 (
             nx24017)) ;
    mux21_ni ix9999 (.Y (nx9998), .A0 (nx9574), .A1 (nx9994), .S0 (nx22459)) ;
    mux21_ni ix9575 (.Y (nx9574), .A0 (nx9362), .A1 (nx9570), .S0 (nx22545)) ;
    mux21_ni ix9363 (.Y (nx9362), .A0 (nx9356), .A1 (nx9278), .S0 (nx23127)) ;
    oai21 ix9357 (.Y (nx9356), .A0 (nx22247), .A1 (nx10201), .B0 (nx10213)) ;
    mux21 ix10202 (.Y (nx10201), .A0 (nx9320), .A1 (nx9348), .S0 (nx22735)) ;
    mux21_ni ix9321 (.Y (nx9320), .A0 (nx9304), .A1 (nx9316), .S0 (nx23433)) ;
    mux21_ni ix9305 (.Y (nx9304), .A0 (inputs_388__2), .A1 (inputs_389__2), .S0 (
             nx24017)) ;
    mux21_ni ix9317 (.Y (nx9316), .A0 (inputs_390__2), .A1 (inputs_391__2), .S0 (
             nx24017)) ;
    mux21_ni ix9349 (.Y (nx9348), .A0 (nx9332), .A1 (nx9344), .S0 (nx23433)) ;
    mux21_ni ix9333 (.Y (nx9332), .A0 (inputs_404__2), .A1 (inputs_405__2), .S0 (
             nx24017)) ;
    mux21_ni ix9345 (.Y (nx9344), .A0 (inputs_406__2), .A1 (inputs_407__2), .S0 (
             nx24017)) ;
    nand04 ix10214 (.Y (nx10213), .A0 (nx22247), .A1 (nx23433), .A2 (nx24017), .A3 (
           nx9292)) ;
    mux21_ni ix9293 (.Y (nx9292), .A0 (inputs_387__2), .A1 (inputs_403__2), .S0 (
             nx22735)) ;
    mux21_ni ix9279 (.Y (nx9278), .A0 (nx9214), .A1 (nx9274), .S0 (nx22735)) ;
    mux21_ni ix9215 (.Y (nx9214), .A0 (nx9182), .A1 (nx9210), .S0 (nx23211)) ;
    mux21_ni ix9183 (.Y (nx9182), .A0 (nx9166), .A1 (nx9178), .S0 (nx23435)) ;
    mux21_ni ix9167 (.Y (nx9166), .A0 (inputs_392__2), .A1 (inputs_393__2), .S0 (
             nx24017)) ;
    mux21_ni ix9179 (.Y (nx9178), .A0 (inputs_394__2), .A1 (inputs_395__2), .S0 (
             nx24019)) ;
    mux21_ni ix9211 (.Y (nx9210), .A0 (nx9194), .A1 (nx9206), .S0 (nx23435)) ;
    mux21_ni ix9195 (.Y (nx9194), .A0 (inputs_396__2), .A1 (inputs_397__2), .S0 (
             nx24019)) ;
    mux21_ni ix9207 (.Y (nx9206), .A0 (inputs_398__2), .A1 (inputs_399__2), .S0 (
             nx24019)) ;
    mux21_ni ix9275 (.Y (nx9274), .A0 (nx9242), .A1 (nx9270), .S0 (nx23211)) ;
    mux21_ni ix9243 (.Y (nx9242), .A0 (nx9226), .A1 (nx9238), .S0 (nx23435)) ;
    mux21_ni ix9227 (.Y (nx9226), .A0 (inputs_408__2), .A1 (inputs_409__2), .S0 (
             nx24019)) ;
    mux21_ni ix9239 (.Y (nx9238), .A0 (inputs_410__2), .A1 (inputs_411__2), .S0 (
             nx24019)) ;
    mux21_ni ix9271 (.Y (nx9270), .A0 (nx9254), .A1 (nx9266), .S0 (nx23435)) ;
    mux21_ni ix9255 (.Y (nx9254), .A0 (inputs_412__2), .A1 (inputs_413__2), .S0 (
             nx24019)) ;
    mux21_ni ix9267 (.Y (nx9266), .A0 (inputs_414__2), .A1 (inputs_415__2), .S0 (
             nx24019)) ;
    mux21_ni ix9571 (.Y (nx9570), .A0 (nx9564), .A1 (nx9486), .S0 (nx23127)) ;
    oai21 ix9565 (.Y (nx9564), .A0 (nx22247), .A1 (nx10243), .B0 (nx10257)) ;
    mux21 ix10244 (.Y (nx10243), .A0 (nx9528), .A1 (nx9556), .S0 (nx22735)) ;
    mux21_ni ix9529 (.Y (nx9528), .A0 (nx9512), .A1 (nx9524), .S0 (nx23435)) ;
    mux21_ni ix9513 (.Y (nx9512), .A0 (inputs_420__2), .A1 (inputs_421__2), .S0 (
             nx24021)) ;
    mux21_ni ix9525 (.Y (nx9524), .A0 (inputs_422__2), .A1 (inputs_423__2), .S0 (
             nx24021)) ;
    mux21_ni ix9557 (.Y (nx9556), .A0 (nx9540), .A1 (nx9552), .S0 (nx23435)) ;
    mux21_ni ix9541 (.Y (nx9540), .A0 (inputs_436__2), .A1 (inputs_437__2), .S0 (
             nx24021)) ;
    mux21_ni ix9553 (.Y (nx9552), .A0 (inputs_438__2), .A1 (inputs_439__2), .S0 (
             nx24021)) ;
    nand04 ix10258 (.Y (nx10257), .A0 (nx22249), .A1 (nx23435), .A2 (nx24021), .A3 (
           nx9500)) ;
    mux21_ni ix9501 (.Y (nx9500), .A0 (inputs_419__2), .A1 (inputs_435__2), .S0 (
             nx22735)) ;
    mux21_ni ix9487 (.Y (nx9486), .A0 (nx9422), .A1 (nx9482), .S0 (nx22735)) ;
    mux21_ni ix9423 (.Y (nx9422), .A0 (nx9390), .A1 (nx9418), .S0 (nx23211)) ;
    mux21_ni ix9391 (.Y (nx9390), .A0 (nx9374), .A1 (nx9386), .S0 (nx23437)) ;
    mux21_ni ix9375 (.Y (nx9374), .A0 (inputs_424__2), .A1 (inputs_425__2), .S0 (
             nx24021)) ;
    mux21_ni ix9387 (.Y (nx9386), .A0 (inputs_426__2), .A1 (inputs_427__2), .S0 (
             nx24021)) ;
    mux21_ni ix9419 (.Y (nx9418), .A0 (nx9402), .A1 (nx9414), .S0 (nx23437)) ;
    mux21_ni ix9403 (.Y (nx9402), .A0 (inputs_428__2), .A1 (inputs_429__2), .S0 (
             nx24023)) ;
    mux21_ni ix9415 (.Y (nx9414), .A0 (inputs_430__2), .A1 (inputs_431__2), .S0 (
             nx24023)) ;
    mux21_ni ix9483 (.Y (nx9482), .A0 (nx9450), .A1 (nx9478), .S0 (nx23211)) ;
    mux21_ni ix9451 (.Y (nx9450), .A0 (nx9434), .A1 (nx9446), .S0 (nx23437)) ;
    mux21_ni ix9435 (.Y (nx9434), .A0 (inputs_440__2), .A1 (inputs_441__2), .S0 (
             nx24023)) ;
    mux21_ni ix9447 (.Y (nx9446), .A0 (inputs_442__2), .A1 (inputs_443__2), .S0 (
             nx24023)) ;
    mux21_ni ix9479 (.Y (nx9478), .A0 (nx9462), .A1 (nx9474), .S0 (nx23437)) ;
    mux21_ni ix9463 (.Y (nx9462), .A0 (inputs_444__2), .A1 (inputs_445__2), .S0 (
             nx24023)) ;
    mux21_ni ix9475 (.Y (nx9474), .A0 (inputs_446__2), .A1 (inputs_447__2), .S0 (
             nx24023)) ;
    mux21_ni ix9995 (.Y (nx9994), .A0 (nx9782), .A1 (nx9990), .S0 (nx22545)) ;
    mux21_ni ix9783 (.Y (nx9782), .A0 (nx9776), .A1 (nx9698), .S0 (nx23127)) ;
    oai21 ix9777 (.Y (nx9776), .A0 (nx22249), .A1 (nx10289), .B0 (nx10301)) ;
    mux21 ix10290 (.Y (nx10289), .A0 (nx9740), .A1 (nx9768), .S0 (nx22737)) ;
    mux21_ni ix9741 (.Y (nx9740), .A0 (nx9724), .A1 (nx9736), .S0 (nx23437)) ;
    mux21_ni ix9725 (.Y (nx9724), .A0 (inputs_452__2), .A1 (inputs_453__2), .S0 (
             nx24023)) ;
    mux21_ni ix9737 (.Y (nx9736), .A0 (inputs_454__2), .A1 (inputs_455__2), .S0 (
             nx24025)) ;
    mux21_ni ix9769 (.Y (nx9768), .A0 (nx9752), .A1 (nx9764), .S0 (nx23437)) ;
    mux21_ni ix9753 (.Y (nx9752), .A0 (inputs_468__2), .A1 (inputs_469__2), .S0 (
             nx24025)) ;
    mux21_ni ix9765 (.Y (nx9764), .A0 (inputs_470__2), .A1 (inputs_471__2), .S0 (
             nx24025)) ;
    nand04 ix10302 (.Y (nx10301), .A0 (nx22249), .A1 (nx23437), .A2 (nx24025), .A3 (
           nx9712)) ;
    mux21_ni ix9713 (.Y (nx9712), .A0 (inputs_451__2), .A1 (inputs_467__2), .S0 (
             nx22737)) ;
    mux21_ni ix9699 (.Y (nx9698), .A0 (nx9634), .A1 (nx9694), .S0 (nx22737)) ;
    mux21_ni ix9635 (.Y (nx9634), .A0 (nx9602), .A1 (nx9630), .S0 (nx23211)) ;
    mux21_ni ix9603 (.Y (nx9602), .A0 (nx9586), .A1 (nx9598), .S0 (nx23439)) ;
    mux21_ni ix9587 (.Y (nx9586), .A0 (inputs_456__2), .A1 (inputs_457__2), .S0 (
             nx24025)) ;
    mux21_ni ix9599 (.Y (nx9598), .A0 (inputs_458__2), .A1 (inputs_459__2), .S0 (
             nx24025)) ;
    mux21_ni ix9631 (.Y (nx9630), .A0 (nx9614), .A1 (nx9626), .S0 (nx23439)) ;
    mux21_ni ix9615 (.Y (nx9614), .A0 (inputs_460__2), .A1 (inputs_461__2), .S0 (
             nx24025)) ;
    mux21_ni ix9627 (.Y (nx9626), .A0 (inputs_462__2), .A1 (inputs_463__2), .S0 (
             nx24027)) ;
    mux21_ni ix9695 (.Y (nx9694), .A0 (nx9662), .A1 (nx9690), .S0 (nx23213)) ;
    mux21_ni ix9663 (.Y (nx9662), .A0 (nx9646), .A1 (nx9658), .S0 (nx23439)) ;
    mux21_ni ix9647 (.Y (nx9646), .A0 (inputs_472__2), .A1 (inputs_473__2), .S0 (
             nx24027)) ;
    mux21_ni ix9659 (.Y (nx9658), .A0 (inputs_474__2), .A1 (inputs_475__2), .S0 (
             nx24027)) ;
    mux21_ni ix9691 (.Y (nx9690), .A0 (nx9674), .A1 (nx9686), .S0 (nx23439)) ;
    mux21_ni ix9675 (.Y (nx9674), .A0 (inputs_476__2), .A1 (inputs_477__2), .S0 (
             nx24027)) ;
    mux21_ni ix9687 (.Y (nx9686), .A0 (inputs_478__2), .A1 (inputs_479__2), .S0 (
             nx24027)) ;
    mux21_ni ix9991 (.Y (nx9990), .A0 (nx9984), .A1 (nx9906), .S0 (nx23127)) ;
    oai21 ix9985 (.Y (nx9984), .A0 (nx22249), .A1 (nx10333), .B0 (nx10347)) ;
    mux21 ix10334 (.Y (nx10333), .A0 (nx9948), .A1 (nx9976), .S0 (nx22737)) ;
    mux21_ni ix9949 (.Y (nx9948), .A0 (nx9932), .A1 (nx9944), .S0 (nx23439)) ;
    mux21_ni ix9933 (.Y (nx9932), .A0 (inputs_484__2), .A1 (inputs_485__2), .S0 (
             nx24027)) ;
    mux21_ni ix9945 (.Y (nx9944), .A0 (inputs_486__2), .A1 (inputs_487__2), .S0 (
             nx24027)) ;
    mux21_ni ix9977 (.Y (nx9976), .A0 (nx9960), .A1 (nx9972), .S0 (nx23439)) ;
    mux21_ni ix9961 (.Y (nx9960), .A0 (inputs_500__2), .A1 (inputs_501__2), .S0 (
             nx24029)) ;
    mux21_ni ix9973 (.Y (nx9972), .A0 (inputs_502__2), .A1 (inputs_503__2), .S0 (
             nx24029)) ;
    nand04 ix10348 (.Y (nx10347), .A0 (nx22249), .A1 (nx23439), .A2 (nx24029), .A3 (
           nx9920)) ;
    mux21_ni ix9921 (.Y (nx9920), .A0 (inputs_483__2), .A1 (inputs_499__2), .S0 (
             nx22737)) ;
    mux21_ni ix9907 (.Y (nx9906), .A0 (nx9842), .A1 (nx9902), .S0 (nx22737)) ;
    mux21_ni ix9843 (.Y (nx9842), .A0 (nx9810), .A1 (nx9838), .S0 (nx23213)) ;
    mux21_ni ix9811 (.Y (nx9810), .A0 (nx9794), .A1 (nx9806), .S0 (nx23441)) ;
    mux21_ni ix9795 (.Y (nx9794), .A0 (inputs_488__2), .A1 (inputs_489__2), .S0 (
             nx24029)) ;
    mux21_ni ix9807 (.Y (nx9806), .A0 (inputs_490__2), .A1 (inputs_491__2), .S0 (
             nx24029)) ;
    mux21_ni ix9839 (.Y (nx9838), .A0 (nx9822), .A1 (nx9834), .S0 (nx23441)) ;
    mux21_ni ix9823 (.Y (nx9822), .A0 (inputs_492__2), .A1 (inputs_493__2), .S0 (
             nx24029)) ;
    mux21_ni ix9835 (.Y (nx9834), .A0 (inputs_494__2), .A1 (inputs_495__2), .S0 (
             nx24029)) ;
    mux21_ni ix9903 (.Y (nx9902), .A0 (nx9870), .A1 (nx9898), .S0 (nx23213)) ;
    mux21_ni ix9871 (.Y (nx9870), .A0 (nx9854), .A1 (nx9866), .S0 (nx23441)) ;
    mux21_ni ix9855 (.Y (nx9854), .A0 (inputs_504__2), .A1 (inputs_505__2), .S0 (
             nx24031)) ;
    mux21_ni ix9867 (.Y (nx9866), .A0 (inputs_506__2), .A1 (inputs_507__2), .S0 (
             nx24031)) ;
    mux21_ni ix9899 (.Y (nx9898), .A0 (nx9882), .A1 (nx9894), .S0 (nx23441)) ;
    mux21_ni ix9883 (.Y (nx9882), .A0 (inputs_508__2), .A1 (inputs_509__2), .S0 (
             nx24031)) ;
    mux21_ni ix9895 (.Y (nx9894), .A0 (inputs_510__2), .A1 (inputs_511__2), .S0 (
             nx24031)) ;
    aoi32 ix10376 (.Y (nx10375), .A0 (nx10768), .A1 (nx22385), .A2 (nx22249), .B0 (
          nx24851), .B1 (nx12464)) ;
    oai21 ix10769 (.Y (nx10768), .A0 (nx23441), .A1 (nx10379), .B0 (nx10477)) ;
    mux21 ix10380 (.Y (nx10379), .A0 (nx10506), .A1 (nx10758), .S0 (nx24031)) ;
    mux21_ni ix10507 (.Y (nx10506), .A0 (nx10378), .A1 (nx10502), .S0 (nx22393)
             ) ;
    mux21_ni ix10379 (.Y (nx10378), .A0 (nx10314), .A1 (nx10374), .S0 (nx22415)
             ) ;
    mux21_ni ix10315 (.Y (nx10314), .A0 (nx10282), .A1 (nx10310), .S0 (nx22459)
             ) ;
    mux21_ni ix10283 (.Y (nx10282), .A0 (nx10266), .A1 (nx10278), .S0 (nx22545)
             ) ;
    mux21_ni ix10267 (.Y (nx10266), .A0 (inputs_0__2), .A1 (inputs_16__2), .S0 (
             nx22737)) ;
    mux21_ni ix10279 (.Y (nx10278), .A0 (inputs_32__2), .A1 (inputs_48__2), .S0 (
             nx22739)) ;
    mux21_ni ix10311 (.Y (nx10310), .A0 (nx10294), .A1 (nx10306), .S0 (nx22545)
             ) ;
    mux21_ni ix10295 (.Y (nx10294), .A0 (inputs_64__2), .A1 (inputs_80__2), .S0 (
             nx22739)) ;
    mux21_ni ix10307 (.Y (nx10306), .A0 (inputs_96__2), .A1 (inputs_112__2), .S0 (
             nx22739)) ;
    mux21_ni ix10375 (.Y (nx10374), .A0 (nx10342), .A1 (nx10370), .S0 (nx22461)
             ) ;
    mux21_ni ix10343 (.Y (nx10342), .A0 (nx10326), .A1 (nx10338), .S0 (nx22547)
             ) ;
    mux21_ni ix10327 (.Y (nx10326), .A0 (inputs_128__2), .A1 (inputs_144__2), .S0 (
             nx22739)) ;
    mux21_ni ix10339 (.Y (nx10338), .A0 (inputs_160__2), .A1 (inputs_176__2), .S0 (
             nx22739)) ;
    mux21_ni ix10371 (.Y (nx10370), .A0 (nx10354), .A1 (nx10366), .S0 (nx22547)
             ) ;
    mux21_ni ix10355 (.Y (nx10354), .A0 (inputs_192__2), .A1 (inputs_208__2), .S0 (
             nx22739)) ;
    mux21_ni ix10367 (.Y (nx10366), .A0 (inputs_224__2), .A1 (inputs_240__2), .S0 (
             nx22739)) ;
    mux21_ni ix10503 (.Y (nx10502), .A0 (nx10438), .A1 (nx10498), .S0 (nx22415)
             ) ;
    mux21_ni ix10439 (.Y (nx10438), .A0 (nx10406), .A1 (nx10434), .S0 (nx22461)
             ) ;
    mux21_ni ix10407 (.Y (nx10406), .A0 (nx10390), .A1 (nx10402), .S0 (nx22547)
             ) ;
    mux21_ni ix10391 (.Y (nx10390), .A0 (inputs_256__2), .A1 (inputs_272__2), .S0 (
             nx22741)) ;
    mux21_ni ix10403 (.Y (nx10402), .A0 (inputs_288__2), .A1 (inputs_304__2), .S0 (
             nx22741)) ;
    mux21_ni ix10435 (.Y (nx10434), .A0 (nx10418), .A1 (nx10430), .S0 (nx22547)
             ) ;
    mux21_ni ix10419 (.Y (nx10418), .A0 (inputs_320__2), .A1 (inputs_336__2), .S0 (
             nx22741)) ;
    mux21_ni ix10431 (.Y (nx10430), .A0 (inputs_352__2), .A1 (inputs_368__2), .S0 (
             nx22741)) ;
    mux21_ni ix10499 (.Y (nx10498), .A0 (nx10466), .A1 (nx10494), .S0 (nx22461)
             ) ;
    mux21_ni ix10467 (.Y (nx10466), .A0 (nx10450), .A1 (nx10462), .S0 (nx22547)
             ) ;
    mux21_ni ix10451 (.Y (nx10450), .A0 (inputs_384__2), .A1 (inputs_400__2), .S0 (
             nx22741)) ;
    mux21_ni ix10463 (.Y (nx10462), .A0 (inputs_416__2), .A1 (inputs_432__2), .S0 (
             nx22741)) ;
    mux21_ni ix10495 (.Y (nx10494), .A0 (nx10478), .A1 (nx10490), .S0 (nx22547)
             ) ;
    mux21_ni ix10479 (.Y (nx10478), .A0 (inputs_448__2), .A1 (inputs_464__2), .S0 (
             nx22741)) ;
    mux21_ni ix10491 (.Y (nx10490), .A0 (inputs_480__2), .A1 (inputs_496__2), .S0 (
             nx22743)) ;
    mux21_ni ix10759 (.Y (nx10758), .A0 (nx10630), .A1 (nx10754), .S0 (nx22395)
             ) ;
    mux21_ni ix10631 (.Y (nx10630), .A0 (nx10566), .A1 (nx10626), .S0 (nx22415)
             ) ;
    mux21_ni ix10567 (.Y (nx10566), .A0 (nx10534), .A1 (nx10562), .S0 (nx22461)
             ) ;
    mux21_ni ix10535 (.Y (nx10534), .A0 (nx10518), .A1 (nx10530), .S0 (nx22547)
             ) ;
    mux21_ni ix10519 (.Y (nx10518), .A0 (inputs_1__2), .A1 (inputs_17__2), .S0 (
             nx22743)) ;
    mux21_ni ix10531 (.Y (nx10530), .A0 (inputs_33__2), .A1 (inputs_49__2), .S0 (
             nx22743)) ;
    mux21_ni ix10563 (.Y (nx10562), .A0 (nx10546), .A1 (nx10558), .S0 (nx22549)
             ) ;
    mux21_ni ix10547 (.Y (nx10546), .A0 (inputs_65__2), .A1 (inputs_81__2), .S0 (
             nx22743)) ;
    mux21_ni ix10559 (.Y (nx10558), .A0 (inputs_97__2), .A1 (inputs_113__2), .S0 (
             nx22743)) ;
    mux21_ni ix10627 (.Y (nx10626), .A0 (nx10594), .A1 (nx10622), .S0 (nx22461)
             ) ;
    mux21_ni ix10595 (.Y (nx10594), .A0 (nx10578), .A1 (nx10590), .S0 (nx22549)
             ) ;
    mux21_ni ix10579 (.Y (nx10578), .A0 (inputs_129__2), .A1 (inputs_145__2), .S0 (
             nx22743)) ;
    mux21_ni ix10591 (.Y (nx10590), .A0 (inputs_161__2), .A1 (inputs_177__2), .S0 (
             nx22743)) ;
    mux21_ni ix10623 (.Y (nx10622), .A0 (nx10606), .A1 (nx10618), .S0 (nx22549)
             ) ;
    mux21_ni ix10607 (.Y (nx10606), .A0 (inputs_193__2), .A1 (inputs_209__2), .S0 (
             nx22745)) ;
    mux21_ni ix10619 (.Y (nx10618), .A0 (inputs_225__2), .A1 (inputs_241__2), .S0 (
             nx22745)) ;
    mux21_ni ix10755 (.Y (nx10754), .A0 (nx10690), .A1 (nx10750), .S0 (nx22415)
             ) ;
    mux21_ni ix10691 (.Y (nx10690), .A0 (nx10658), .A1 (nx10686), .S0 (nx22461)
             ) ;
    mux21_ni ix10659 (.Y (nx10658), .A0 (nx10642), .A1 (nx10654), .S0 (nx22549)
             ) ;
    mux21_ni ix10643 (.Y (nx10642), .A0 (inputs_257__2), .A1 (inputs_273__2), .S0 (
             nx22745)) ;
    mux21_ni ix10655 (.Y (nx10654), .A0 (inputs_289__2), .A1 (inputs_305__2), .S0 (
             nx22745)) ;
    mux21_ni ix10687 (.Y (nx10686), .A0 (nx10670), .A1 (nx10682), .S0 (nx22549)
             ) ;
    mux21_ni ix10671 (.Y (nx10670), .A0 (inputs_321__2), .A1 (inputs_337__2), .S0 (
             nx22745)) ;
    mux21_ni ix10683 (.Y (nx10682), .A0 (inputs_353__2), .A1 (inputs_369__2), .S0 (
             nx22745)) ;
    mux21_ni ix10751 (.Y (nx10750), .A0 (nx10718), .A1 (nx10746), .S0 (nx22461)
             ) ;
    mux21_ni ix10719 (.Y (nx10718), .A0 (nx10702), .A1 (nx10714), .S0 (nx22549)
             ) ;
    mux21_ni ix10703 (.Y (nx10702), .A0 (inputs_385__2), .A1 (inputs_401__2), .S0 (
             nx22745)) ;
    mux21_ni ix10715 (.Y (nx10714), .A0 (inputs_417__2), .A1 (inputs_433__2), .S0 (
             nx22747)) ;
    mux21_ni ix10747 (.Y (nx10746), .A0 (nx10730), .A1 (nx10742), .S0 (nx22549)
             ) ;
    mux21_ni ix10731 (.Y (nx10730), .A0 (inputs_449__2), .A1 (inputs_465__2), .S0 (
             nx22747)) ;
    mux21_ni ix10743 (.Y (nx10742), .A0 (inputs_481__2), .A1 (inputs_497__2), .S0 (
             nx22747)) ;
    nand03 ix10478 (.Y (nx10477), .A0 (nx10252), .A1 (nx23441), .A2 (nx24879)) ;
    mux21_ni ix10253 (.Y (nx10252), .A0 (nx10124), .A1 (nx10248), .S0 (nx22395)
             ) ;
    mux21_ni ix10125 (.Y (nx10124), .A0 (nx10060), .A1 (nx10120), .S0 (nx22417)
             ) ;
    mux21_ni ix10061 (.Y (nx10060), .A0 (nx10028), .A1 (nx10056), .S0 (nx22463)
             ) ;
    mux21_ni ix10029 (.Y (nx10028), .A0 (nx10012), .A1 (nx10024), .S0 (nx22551)
             ) ;
    mux21_ni ix10013 (.Y (nx10012), .A0 (inputs_2__2), .A1 (inputs_18__2), .S0 (
             nx22747)) ;
    mux21_ni ix10025 (.Y (nx10024), .A0 (inputs_34__2), .A1 (inputs_50__2), .S0 (
             nx22747)) ;
    mux21_ni ix10057 (.Y (nx10056), .A0 (nx10040), .A1 (nx10052), .S0 (nx22551)
             ) ;
    mux21_ni ix10041 (.Y (nx10040), .A0 (inputs_66__2), .A1 (inputs_82__2), .S0 (
             nx22747)) ;
    mux21_ni ix10053 (.Y (nx10052), .A0 (inputs_98__2), .A1 (inputs_114__2), .S0 (
             nx22747)) ;
    mux21_ni ix10121 (.Y (nx10120), .A0 (nx10088), .A1 (nx10116), .S0 (nx22463)
             ) ;
    mux21_ni ix10089 (.Y (nx10088), .A0 (nx10072), .A1 (nx10084), .S0 (nx22551)
             ) ;
    mux21_ni ix10073 (.Y (nx10072), .A0 (inputs_130__2), .A1 (inputs_146__2), .S0 (
             nx22749)) ;
    mux21_ni ix10085 (.Y (nx10084), .A0 (inputs_162__2), .A1 (inputs_178__2), .S0 (
             nx22749)) ;
    mux21_ni ix10117 (.Y (nx10116), .A0 (nx10100), .A1 (nx10112), .S0 (nx22551)
             ) ;
    mux21_ni ix10101 (.Y (nx10100), .A0 (inputs_194__2), .A1 (inputs_210__2), .S0 (
             nx22749)) ;
    mux21_ni ix10113 (.Y (nx10112), .A0 (inputs_226__2), .A1 (inputs_242__2), .S0 (
             nx22749)) ;
    mux21_ni ix10249 (.Y (nx10248), .A0 (nx10184), .A1 (nx10244), .S0 (nx22417)
             ) ;
    mux21_ni ix10185 (.Y (nx10184), .A0 (nx10152), .A1 (nx10180), .S0 (nx22463)
             ) ;
    mux21_ni ix10153 (.Y (nx10152), .A0 (nx10136), .A1 (nx10148), .S0 (nx22551)
             ) ;
    mux21_ni ix10137 (.Y (nx10136), .A0 (inputs_258__2), .A1 (inputs_274__2), .S0 (
             nx22749)) ;
    mux21_ni ix10149 (.Y (nx10148), .A0 (inputs_290__2), .A1 (inputs_306__2), .S0 (
             nx22749)) ;
    mux21_ni ix10181 (.Y (nx10180), .A0 (nx10164), .A1 (nx10176), .S0 (nx22551)
             ) ;
    mux21_ni ix10165 (.Y (nx10164), .A0 (inputs_322__2), .A1 (inputs_338__2), .S0 (
             nx22749)) ;
    mux21_ni ix10177 (.Y (nx10176), .A0 (inputs_354__2), .A1 (inputs_370__2), .S0 (
             nx22751)) ;
    mux21_ni ix10245 (.Y (nx10244), .A0 (nx10212), .A1 (nx10240), .S0 (nx22463)
             ) ;
    mux21_ni ix10213 (.Y (nx10212), .A0 (nx10196), .A1 (nx10208), .S0 (nx22551)
             ) ;
    mux21_ni ix10197 (.Y (nx10196), .A0 (inputs_386__2), .A1 (inputs_402__2), .S0 (
             nx22751)) ;
    mux21_ni ix10209 (.Y (nx10208), .A0 (inputs_418__2), .A1 (inputs_434__2), .S0 (
             nx22751)) ;
    mux21_ni ix10241 (.Y (nx10240), .A0 (nx10224), .A1 (nx10236), .S0 (nx22553)
             ) ;
    mux21_ni ix10225 (.Y (nx10224), .A0 (inputs_450__2), .A1 (inputs_466__2), .S0 (
             nx22751)) ;
    mux21_ni ix10237 (.Y (nx10236), .A0 (inputs_482__2), .A1 (inputs_498__2), .S0 (
             nx22751)) ;
    mux21_ni ix12465 (.Y (nx12464), .A0 (nx11616), .A1 (nx12460), .S0 (nx22417)
             ) ;
    mux21_ni ix11617 (.Y (nx11616), .A0 (nx11192), .A1 (nx11612), .S0 (nx22463)
             ) ;
    mux21_ni ix11193 (.Y (nx11192), .A0 (nx10980), .A1 (nx11188), .S0 (nx22553)
             ) ;
    mux21_ni ix10981 (.Y (nx10980), .A0 (nx10974), .A1 (nx10896), .S0 (nx23127)
             ) ;
    oai21 ix10975 (.Y (nx10974), .A0 (nx22249), .A1 (nx10539), .B0 (nx10551)) ;
    mux21 ix10540 (.Y (nx10539), .A0 (nx10938), .A1 (nx10966), .S0 (nx22751)) ;
    mux21_ni ix10939 (.Y (nx10938), .A0 (nx10922), .A1 (nx10934), .S0 (nx23441)
             ) ;
    mux21_ni ix10923 (.Y (nx10922), .A0 (inputs_4__2), .A1 (inputs_5__2), .S0 (
             nx24031)) ;
    mux21_ni ix10935 (.Y (nx10934), .A0 (inputs_6__2), .A1 (inputs_7__2), .S0 (
             nx24031)) ;
    mux21_ni ix10967 (.Y (nx10966), .A0 (nx10950), .A1 (nx10962), .S0 (nx23443)
             ) ;
    mux21_ni ix10951 (.Y (nx10950), .A0 (inputs_20__2), .A1 (inputs_21__2), .S0 (
             nx24033)) ;
    mux21_ni ix10963 (.Y (nx10962), .A0 (inputs_22__2), .A1 (inputs_23__2), .S0 (
             nx24033)) ;
    nand04 ix10552 (.Y (nx10551), .A0 (nx22251), .A1 (nx23443), .A2 (nx24033), .A3 (
           nx10910)) ;
    mux21_ni ix10911 (.Y (nx10910), .A0 (inputs_3__2), .A1 (inputs_19__2), .S0 (
             nx22751)) ;
    mux21_ni ix10897 (.Y (nx10896), .A0 (nx10832), .A1 (nx10892), .S0 (nx22753)
             ) ;
    mux21_ni ix10833 (.Y (nx10832), .A0 (nx10800), .A1 (nx10828), .S0 (nx23213)
             ) ;
    mux21_ni ix10801 (.Y (nx10800), .A0 (nx10784), .A1 (nx10796), .S0 (nx23443)
             ) ;
    mux21_ni ix10785 (.Y (nx10784), .A0 (inputs_8__2), .A1 (inputs_9__2), .S0 (
             nx24033)) ;
    mux21_ni ix10797 (.Y (nx10796), .A0 (inputs_10__2), .A1 (inputs_11__2), .S0 (
             nx24033)) ;
    mux21_ni ix10829 (.Y (nx10828), .A0 (nx10812), .A1 (nx10824), .S0 (nx23443)
             ) ;
    mux21_ni ix10813 (.Y (nx10812), .A0 (inputs_12__2), .A1 (inputs_13__2), .S0 (
             nx24033)) ;
    mux21_ni ix10825 (.Y (nx10824), .A0 (inputs_14__2), .A1 (inputs_15__2), .S0 (
             nx24033)) ;
    mux21_ni ix10893 (.Y (nx10892), .A0 (nx10860), .A1 (nx10888), .S0 (nx23213)
             ) ;
    mux21_ni ix10861 (.Y (nx10860), .A0 (nx10844), .A1 (nx10856), .S0 (nx23443)
             ) ;
    mux21_ni ix10845 (.Y (nx10844), .A0 (inputs_24__2), .A1 (inputs_25__2), .S0 (
             nx24035)) ;
    mux21_ni ix10857 (.Y (nx10856), .A0 (inputs_26__2), .A1 (inputs_27__2), .S0 (
             nx24035)) ;
    mux21_ni ix10889 (.Y (nx10888), .A0 (nx10872), .A1 (nx10884), .S0 (nx23443)
             ) ;
    mux21_ni ix10873 (.Y (nx10872), .A0 (inputs_28__2), .A1 (inputs_29__2), .S0 (
             nx24035)) ;
    mux21_ni ix10885 (.Y (nx10884), .A0 (inputs_30__2), .A1 (inputs_31__2), .S0 (
             nx24035)) ;
    mux21_ni ix11189 (.Y (nx11188), .A0 (nx11182), .A1 (nx11104), .S0 (nx23127)
             ) ;
    oai21 ix11183 (.Y (nx11182), .A0 (nx22251), .A1 (nx10583), .B0 (nx10595)) ;
    mux21 ix10584 (.Y (nx10583), .A0 (nx11146), .A1 (nx11174), .S0 (nx22753)) ;
    mux21_ni ix11147 (.Y (nx11146), .A0 (nx11130), .A1 (nx11142), .S0 (nx23443)
             ) ;
    mux21_ni ix11131 (.Y (nx11130), .A0 (inputs_36__2), .A1 (inputs_37__2), .S0 (
             nx24035)) ;
    mux21_ni ix11143 (.Y (nx11142), .A0 (inputs_38__2), .A1 (inputs_39__2), .S0 (
             nx24035)) ;
    mux21_ni ix11175 (.Y (nx11174), .A0 (nx11158), .A1 (nx11170), .S0 (nx23445)
             ) ;
    mux21_ni ix11159 (.Y (nx11158), .A0 (inputs_52__2), .A1 (inputs_53__2), .S0 (
             nx24035)) ;
    mux21_ni ix11171 (.Y (nx11170), .A0 (inputs_54__2), .A1 (inputs_55__2), .S0 (
             nx24037)) ;
    nand04 ix10596 (.Y (nx10595), .A0 (nx22251), .A1 (nx23445), .A2 (nx24037), .A3 (
           nx11118)) ;
    mux21_ni ix11119 (.Y (nx11118), .A0 (inputs_35__2), .A1 (inputs_51__2), .S0 (
             nx22753)) ;
    mux21_ni ix11105 (.Y (nx11104), .A0 (nx11040), .A1 (nx11100), .S0 (nx22753)
             ) ;
    mux21_ni ix11041 (.Y (nx11040), .A0 (nx11008), .A1 (nx11036), .S0 (nx23213)
             ) ;
    mux21_ni ix11009 (.Y (nx11008), .A0 (nx10992), .A1 (nx11004), .S0 (nx23445)
             ) ;
    mux21_ni ix10993 (.Y (nx10992), .A0 (inputs_40__2), .A1 (inputs_41__2), .S0 (
             nx24037)) ;
    mux21_ni ix11005 (.Y (nx11004), .A0 (inputs_42__2), .A1 (inputs_43__2), .S0 (
             nx24037)) ;
    mux21_ni ix11037 (.Y (nx11036), .A0 (nx11020), .A1 (nx11032), .S0 (nx23445)
             ) ;
    mux21_ni ix11021 (.Y (nx11020), .A0 (inputs_44__2), .A1 (inputs_45__2), .S0 (
             nx24037)) ;
    mux21_ni ix11033 (.Y (nx11032), .A0 (inputs_46__2), .A1 (inputs_47__2), .S0 (
             nx24037)) ;
    mux21_ni ix11101 (.Y (nx11100), .A0 (nx11068), .A1 (nx11096), .S0 (nx23213)
             ) ;
    mux21_ni ix11069 (.Y (nx11068), .A0 (nx11052), .A1 (nx11064), .S0 (nx23445)
             ) ;
    mux21_ni ix11053 (.Y (nx11052), .A0 (inputs_56__2), .A1 (inputs_57__2), .S0 (
             nx24037)) ;
    mux21_ni ix11065 (.Y (nx11064), .A0 (inputs_58__2), .A1 (inputs_59__2), .S0 (
             nx24039)) ;
    mux21_ni ix11097 (.Y (nx11096), .A0 (nx11080), .A1 (nx11092), .S0 (nx23445)
             ) ;
    mux21_ni ix11081 (.Y (nx11080), .A0 (inputs_60__2), .A1 (inputs_61__2), .S0 (
             nx24039)) ;
    mux21_ni ix11093 (.Y (nx11092), .A0 (inputs_62__2), .A1 (inputs_63__2), .S0 (
             nx24039)) ;
    mux21_ni ix11613 (.Y (nx11612), .A0 (nx11400), .A1 (nx11608), .S0 (nx22553)
             ) ;
    mux21_ni ix11401 (.Y (nx11400), .A0 (nx11394), .A1 (nx11316), .S0 (nx23129)
             ) ;
    oai21 ix11395 (.Y (nx11394), .A0 (nx22251), .A1 (nx10627), .B0 (nx10639)) ;
    mux21 ix10628 (.Y (nx10627), .A0 (nx11358), .A1 (nx11386), .S0 (nx22753)) ;
    mux21_ni ix11359 (.Y (nx11358), .A0 (nx11342), .A1 (nx11354), .S0 (nx23445)
             ) ;
    mux21_ni ix11343 (.Y (nx11342), .A0 (inputs_68__2), .A1 (inputs_69__2), .S0 (
             nx24039)) ;
    mux21_ni ix11355 (.Y (nx11354), .A0 (inputs_70__2), .A1 (inputs_71__2), .S0 (
             nx24039)) ;
    mux21_ni ix11387 (.Y (nx11386), .A0 (nx11370), .A1 (nx11382), .S0 (nx23447)
             ) ;
    mux21_ni ix11371 (.Y (nx11370), .A0 (inputs_84__2), .A1 (inputs_85__2), .S0 (
             nx24039)) ;
    mux21_ni ix11383 (.Y (nx11382), .A0 (inputs_86__2), .A1 (inputs_87__2), .S0 (
             nx24039)) ;
    nand04 ix10640 (.Y (nx10639), .A0 (nx22251), .A1 (nx23447), .A2 (nx24041), .A3 (
           nx11330)) ;
    mux21_ni ix11331 (.Y (nx11330), .A0 (inputs_67__2), .A1 (inputs_83__2), .S0 (
             nx22753)) ;
    mux21_ni ix11317 (.Y (nx11316), .A0 (nx11252), .A1 (nx11312), .S0 (nx22753)
             ) ;
    mux21_ni ix11253 (.Y (nx11252), .A0 (nx11220), .A1 (nx11248), .S0 (nx23215)
             ) ;
    mux21_ni ix11221 (.Y (nx11220), .A0 (nx11204), .A1 (nx11216), .S0 (nx23447)
             ) ;
    mux21_ni ix11205 (.Y (nx11204), .A0 (inputs_72__2), .A1 (inputs_73__2), .S0 (
             nx24041)) ;
    mux21_ni ix11217 (.Y (nx11216), .A0 (inputs_74__2), .A1 (inputs_75__2), .S0 (
             nx24041)) ;
    mux21_ni ix11249 (.Y (nx11248), .A0 (nx11232), .A1 (nx11244), .S0 (nx23447)
             ) ;
    mux21_ni ix11233 (.Y (nx11232), .A0 (inputs_76__2), .A1 (inputs_77__2), .S0 (
             nx24041)) ;
    mux21_ni ix11245 (.Y (nx11244), .A0 (inputs_78__2), .A1 (inputs_79__2), .S0 (
             nx24041)) ;
    mux21_ni ix11313 (.Y (nx11312), .A0 (nx11280), .A1 (nx11308), .S0 (nx23215)
             ) ;
    mux21_ni ix11281 (.Y (nx11280), .A0 (nx11264), .A1 (nx11276), .S0 (nx23447)
             ) ;
    mux21_ni ix11265 (.Y (nx11264), .A0 (inputs_88__2), .A1 (inputs_89__2), .S0 (
             nx24041)) ;
    mux21_ni ix11277 (.Y (nx11276), .A0 (inputs_90__2), .A1 (inputs_91__2), .S0 (
             nx24041)) ;
    mux21_ni ix11309 (.Y (nx11308), .A0 (nx11292), .A1 (nx11304), .S0 (nx23447)
             ) ;
    mux21_ni ix11293 (.Y (nx11292), .A0 (inputs_92__2), .A1 (inputs_93__2), .S0 (
             nx24043)) ;
    mux21_ni ix11305 (.Y (nx11304), .A0 (inputs_94__2), .A1 (inputs_95__2), .S0 (
             nx24043)) ;
    mux21_ni ix11609 (.Y (nx11608), .A0 (nx11602), .A1 (nx11524), .S0 (nx23129)
             ) ;
    oai21 ix11603 (.Y (nx11602), .A0 (nx22251), .A1 (nx10669), .B0 (nx10679)) ;
    mux21 ix10670 (.Y (nx10669), .A0 (nx11566), .A1 (nx11594), .S0 (nx22755)) ;
    mux21_ni ix11567 (.Y (nx11566), .A0 (nx11550), .A1 (nx11562), .S0 (nx23447)
             ) ;
    mux21_ni ix11551 (.Y (nx11550), .A0 (inputs_100__2), .A1 (inputs_101__2), .S0 (
             nx24043)) ;
    mux21_ni ix11563 (.Y (nx11562), .A0 (inputs_102__2), .A1 (inputs_103__2), .S0 (
             nx24043)) ;
    mux21_ni ix11595 (.Y (nx11594), .A0 (nx11578), .A1 (nx11590), .S0 (nx23449)
             ) ;
    mux21_ni ix11579 (.Y (nx11578), .A0 (inputs_116__2), .A1 (inputs_117__2), .S0 (
             nx24043)) ;
    mux21_ni ix11591 (.Y (nx11590), .A0 (inputs_118__2), .A1 (inputs_119__2), .S0 (
             nx24043)) ;
    nand04 ix10680 (.Y (nx10679), .A0 (nx22251), .A1 (nx23449), .A2 (nx24043), .A3 (
           nx11538)) ;
    mux21_ni ix11539 (.Y (nx11538), .A0 (inputs_99__2), .A1 (inputs_115__2), .S0 (
             nx22755)) ;
    mux21_ni ix11525 (.Y (nx11524), .A0 (nx11460), .A1 (nx11520), .S0 (nx22755)
             ) ;
    mux21_ni ix11461 (.Y (nx11460), .A0 (nx11428), .A1 (nx11456), .S0 (nx23215)
             ) ;
    mux21_ni ix11429 (.Y (nx11428), .A0 (nx11412), .A1 (nx11424), .S0 (nx23449)
             ) ;
    mux21_ni ix11413 (.Y (nx11412), .A0 (inputs_104__2), .A1 (inputs_105__2), .S0 (
             nx24045)) ;
    mux21_ni ix11425 (.Y (nx11424), .A0 (inputs_106__2), .A1 (inputs_107__2), .S0 (
             nx24045)) ;
    mux21_ni ix11457 (.Y (nx11456), .A0 (nx11440), .A1 (nx11452), .S0 (nx23449)
             ) ;
    mux21_ni ix11441 (.Y (nx11440), .A0 (inputs_108__2), .A1 (inputs_109__2), .S0 (
             nx24045)) ;
    mux21_ni ix11453 (.Y (nx11452), .A0 (inputs_110__2), .A1 (inputs_111__2), .S0 (
             nx24045)) ;
    mux21_ni ix11521 (.Y (nx11520), .A0 (nx11488), .A1 (nx11516), .S0 (nx23215)
             ) ;
    mux21_ni ix11489 (.Y (nx11488), .A0 (nx11472), .A1 (nx11484), .S0 (nx23449)
             ) ;
    mux21_ni ix11473 (.Y (nx11472), .A0 (inputs_120__2), .A1 (inputs_121__2), .S0 (
             nx24045)) ;
    mux21_ni ix11485 (.Y (nx11484), .A0 (inputs_122__2), .A1 (inputs_123__2), .S0 (
             nx24045)) ;
    mux21_ni ix11517 (.Y (nx11516), .A0 (nx11500), .A1 (nx11512), .S0 (nx23449)
             ) ;
    mux21_ni ix11501 (.Y (nx11500), .A0 (inputs_124__2), .A1 (inputs_125__2), .S0 (
             nx24045)) ;
    mux21_ni ix11513 (.Y (nx11512), .A0 (inputs_126__2), .A1 (inputs_127__2), .S0 (
             nx24047)) ;
    mux21_ni ix12461 (.Y (nx12460), .A0 (nx12036), .A1 (nx12456), .S0 (nx22463)
             ) ;
    mux21_ni ix12037 (.Y (nx12036), .A0 (nx11824), .A1 (nx12032), .S0 (nx22553)
             ) ;
    mux21_ni ix11825 (.Y (nx11824), .A0 (nx11818), .A1 (nx11740), .S0 (nx23129)
             ) ;
    oai21 ix11819 (.Y (nx11818), .A0 (nx22253), .A1 (nx10713), .B0 (nx10725)) ;
    mux21 ix10714 (.Y (nx10713), .A0 (nx11782), .A1 (nx11810), .S0 (nx22755)) ;
    mux21_ni ix11783 (.Y (nx11782), .A0 (nx11766), .A1 (nx11778), .S0 (nx23449)
             ) ;
    mux21_ni ix11767 (.Y (nx11766), .A0 (inputs_132__2), .A1 (inputs_133__2), .S0 (
             nx24047)) ;
    mux21_ni ix11779 (.Y (nx11778), .A0 (inputs_134__2), .A1 (inputs_135__2), .S0 (
             nx24047)) ;
    mux21_ni ix11811 (.Y (nx11810), .A0 (nx11794), .A1 (nx11806), .S0 (nx23451)
             ) ;
    mux21_ni ix11795 (.Y (nx11794), .A0 (inputs_148__2), .A1 (inputs_149__2), .S0 (
             nx24047)) ;
    mux21_ni ix11807 (.Y (nx11806), .A0 (inputs_150__2), .A1 (inputs_151__2), .S0 (
             nx24047)) ;
    nand04 ix10726 (.Y (nx10725), .A0 (nx22253), .A1 (nx23451), .A2 (nx24047), .A3 (
           nx11754)) ;
    mux21_ni ix11755 (.Y (nx11754), .A0 (inputs_131__2), .A1 (inputs_147__2), .S0 (
             nx22755)) ;
    mux21_ni ix11741 (.Y (nx11740), .A0 (nx11676), .A1 (nx11736), .S0 (nx22755)
             ) ;
    mux21_ni ix11677 (.Y (nx11676), .A0 (nx11644), .A1 (nx11672), .S0 (nx23215)
             ) ;
    mux21_ni ix11645 (.Y (nx11644), .A0 (nx11628), .A1 (nx11640), .S0 (nx23451)
             ) ;
    mux21_ni ix11629 (.Y (nx11628), .A0 (inputs_136__2), .A1 (inputs_137__2), .S0 (
             nx24047)) ;
    mux21_ni ix11641 (.Y (nx11640), .A0 (inputs_138__2), .A1 (inputs_139__2), .S0 (
             nx24049)) ;
    mux21_ni ix11673 (.Y (nx11672), .A0 (nx11656), .A1 (nx11668), .S0 (nx23451)
             ) ;
    mux21_ni ix11657 (.Y (nx11656), .A0 (inputs_140__2), .A1 (inputs_141__2), .S0 (
             nx24049)) ;
    mux21_ni ix11669 (.Y (nx11668), .A0 (inputs_142__2), .A1 (inputs_143__2), .S0 (
             nx24049)) ;
    mux21_ni ix11737 (.Y (nx11736), .A0 (nx11704), .A1 (nx11732), .S0 (nx23215)
             ) ;
    mux21_ni ix11705 (.Y (nx11704), .A0 (nx11688), .A1 (nx11700), .S0 (nx23451)
             ) ;
    mux21_ni ix11689 (.Y (nx11688), .A0 (inputs_152__2), .A1 (inputs_153__2), .S0 (
             nx24049)) ;
    mux21_ni ix11701 (.Y (nx11700), .A0 (inputs_154__2), .A1 (inputs_155__2), .S0 (
             nx24049)) ;
    mux21_ni ix11733 (.Y (nx11732), .A0 (nx11716), .A1 (nx11728), .S0 (nx23451)
             ) ;
    mux21_ni ix11717 (.Y (nx11716), .A0 (inputs_156__2), .A1 (inputs_157__2), .S0 (
             nx24049)) ;
    mux21_ni ix11729 (.Y (nx11728), .A0 (inputs_158__2), .A1 (inputs_159__2), .S0 (
             nx24049)) ;
    mux21_ni ix12033 (.Y (nx12032), .A0 (nx12026), .A1 (nx11948), .S0 (nx23129)
             ) ;
    oai21 ix12027 (.Y (nx12026), .A0 (nx22253), .A1 (nx10759), .B0 (nx10771)) ;
    mux21 ix10760 (.Y (nx10759), .A0 (nx11990), .A1 (nx12018), .S0 (nx22755)) ;
    mux21_ni ix11991 (.Y (nx11990), .A0 (nx11974), .A1 (nx11986), .S0 (nx23451)
             ) ;
    mux21_ni ix11975 (.Y (nx11974), .A0 (inputs_164__2), .A1 (inputs_165__2), .S0 (
             nx24051)) ;
    mux21_ni ix11987 (.Y (nx11986), .A0 (inputs_166__2), .A1 (inputs_167__2), .S0 (
             nx24051)) ;
    mux21_ni ix12019 (.Y (nx12018), .A0 (nx12002), .A1 (nx12014), .S0 (nx23453)
             ) ;
    mux21_ni ix12003 (.Y (nx12002), .A0 (inputs_180__2), .A1 (inputs_181__2), .S0 (
             nx24051)) ;
    mux21_ni ix12015 (.Y (nx12014), .A0 (inputs_182__2), .A1 (inputs_183__2), .S0 (
             nx24051)) ;
    nand04 ix10772 (.Y (nx10771), .A0 (nx22253), .A1 (nx23453), .A2 (nx24051), .A3 (
           nx11962)) ;
    mux21_ni ix11963 (.Y (nx11962), .A0 (inputs_163__2), .A1 (inputs_179__2), .S0 (
             nx22757)) ;
    mux21_ni ix11949 (.Y (nx11948), .A0 (nx11884), .A1 (nx11944), .S0 (nx22757)
             ) ;
    mux21_ni ix11885 (.Y (nx11884), .A0 (nx11852), .A1 (nx11880), .S0 (nx23215)
             ) ;
    mux21_ni ix11853 (.Y (nx11852), .A0 (nx11836), .A1 (nx11848), .S0 (nx23453)
             ) ;
    mux21_ni ix11837 (.Y (nx11836), .A0 (inputs_168__2), .A1 (inputs_169__2), .S0 (
             nx24051)) ;
    mux21_ni ix11849 (.Y (nx11848), .A0 (inputs_170__2), .A1 (inputs_171__2), .S0 (
             nx24051)) ;
    mux21_ni ix11881 (.Y (nx11880), .A0 (nx11864), .A1 (nx11876), .S0 (nx23453)
             ) ;
    mux21_ni ix11865 (.Y (nx11864), .A0 (inputs_172__2), .A1 (inputs_173__2), .S0 (
             nx24053)) ;
    mux21_ni ix11877 (.Y (nx11876), .A0 (inputs_174__2), .A1 (inputs_175__2), .S0 (
             nx24053)) ;
    mux21_ni ix11945 (.Y (nx11944), .A0 (nx11912), .A1 (nx11940), .S0 (nx23217)
             ) ;
    mux21_ni ix11913 (.Y (nx11912), .A0 (nx11896), .A1 (nx11908), .S0 (nx23453)
             ) ;
    mux21_ni ix11897 (.Y (nx11896), .A0 (inputs_184__2), .A1 (inputs_185__2), .S0 (
             nx24053)) ;
    mux21_ni ix11909 (.Y (nx11908), .A0 (inputs_186__2), .A1 (inputs_187__2), .S0 (
             nx24053)) ;
    mux21_ni ix11941 (.Y (nx11940), .A0 (nx11924), .A1 (nx11936), .S0 (nx23453)
             ) ;
    mux21_ni ix11925 (.Y (nx11924), .A0 (inputs_188__2), .A1 (inputs_189__2), .S0 (
             nx24053)) ;
    mux21_ni ix11937 (.Y (nx11936), .A0 (inputs_190__2), .A1 (inputs_191__2), .S0 (
             nx24053)) ;
    mux21_ni ix12457 (.Y (nx12456), .A0 (nx12244), .A1 (nx12452), .S0 (nx22553)
             ) ;
    mux21_ni ix12245 (.Y (nx12244), .A0 (nx12238), .A1 (nx12160), .S0 (nx23129)
             ) ;
    oai21 ix12239 (.Y (nx12238), .A0 (nx22253), .A1 (nx10803), .B0 (nx10815)) ;
    mux21 ix10804 (.Y (nx10803), .A0 (nx12202), .A1 (nx12230), .S0 (nx22757)) ;
    mux21_ni ix12203 (.Y (nx12202), .A0 (nx12186), .A1 (nx12198), .S0 (nx23453)
             ) ;
    mux21_ni ix12187 (.Y (nx12186), .A0 (inputs_196__2), .A1 (inputs_197__2), .S0 (
             nx24053)) ;
    mux21_ni ix12199 (.Y (nx12198), .A0 (inputs_198__2), .A1 (inputs_199__2), .S0 (
             nx24055)) ;
    mux21_ni ix12231 (.Y (nx12230), .A0 (nx12214), .A1 (nx12226), .S0 (nx23455)
             ) ;
    mux21_ni ix12215 (.Y (nx12214), .A0 (inputs_212__2), .A1 (inputs_213__2), .S0 (
             nx24055)) ;
    mux21_ni ix12227 (.Y (nx12226), .A0 (inputs_214__2), .A1 (inputs_215__2), .S0 (
             nx24055)) ;
    nand04 ix10816 (.Y (nx10815), .A0 (nx22253), .A1 (nx23455), .A2 (nx24055), .A3 (
           nx12174)) ;
    mux21_ni ix12175 (.Y (nx12174), .A0 (inputs_195__2), .A1 (inputs_211__2), .S0 (
             nx22757)) ;
    mux21_ni ix12161 (.Y (nx12160), .A0 (nx12096), .A1 (nx12156), .S0 (nx22757)
             ) ;
    mux21_ni ix12097 (.Y (nx12096), .A0 (nx12064), .A1 (nx12092), .S0 (nx23217)
             ) ;
    mux21_ni ix12065 (.Y (nx12064), .A0 (nx12048), .A1 (nx12060), .S0 (nx23455)
             ) ;
    mux21_ni ix12049 (.Y (nx12048), .A0 (inputs_200__2), .A1 (inputs_201__2), .S0 (
             nx24055)) ;
    mux21_ni ix12061 (.Y (nx12060), .A0 (inputs_202__2), .A1 (inputs_203__2), .S0 (
             nx24055)) ;
    mux21_ni ix12093 (.Y (nx12092), .A0 (nx12076), .A1 (nx12088), .S0 (nx23455)
             ) ;
    mux21_ni ix12077 (.Y (nx12076), .A0 (inputs_204__2), .A1 (inputs_205__2), .S0 (
             nx24055)) ;
    mux21_ni ix12089 (.Y (nx12088), .A0 (inputs_206__2), .A1 (inputs_207__2), .S0 (
             nx24057)) ;
    mux21_ni ix12157 (.Y (nx12156), .A0 (nx12124), .A1 (nx12152), .S0 (nx23217)
             ) ;
    mux21_ni ix12125 (.Y (nx12124), .A0 (nx12108), .A1 (nx12120), .S0 (nx23455)
             ) ;
    mux21_ni ix12109 (.Y (nx12108), .A0 (inputs_216__2), .A1 (inputs_217__2), .S0 (
             nx24057)) ;
    mux21_ni ix12121 (.Y (nx12120), .A0 (inputs_218__2), .A1 (inputs_219__2), .S0 (
             nx24057)) ;
    mux21_ni ix12153 (.Y (nx12152), .A0 (nx12136), .A1 (nx12148), .S0 (nx23455)
             ) ;
    mux21_ni ix12137 (.Y (nx12136), .A0 (inputs_220__2), .A1 (inputs_221__2), .S0 (
             nx24057)) ;
    mux21_ni ix12149 (.Y (nx12148), .A0 (inputs_222__2), .A1 (inputs_223__2), .S0 (
             nx24057)) ;
    mux21_ni ix12453 (.Y (nx12452), .A0 (nx12446), .A1 (nx12368), .S0 (nx23129)
             ) ;
    oai21 ix12447 (.Y (nx12446), .A0 (nx22253), .A1 (nx10847), .B0 (nx10859)) ;
    mux21 ix10848 (.Y (nx10847), .A0 (nx12410), .A1 (nx12438), .S0 (nx22757)) ;
    mux21_ni ix12411 (.Y (nx12410), .A0 (nx12394), .A1 (nx12406), .S0 (nx23455)
             ) ;
    mux21_ni ix12395 (.Y (nx12394), .A0 (inputs_228__2), .A1 (inputs_229__2), .S0 (
             nx24057)) ;
    mux21_ni ix12407 (.Y (nx12406), .A0 (inputs_230__2), .A1 (inputs_231__2), .S0 (
             nx24057)) ;
    mux21_ni ix12439 (.Y (nx12438), .A0 (nx12422), .A1 (nx12434), .S0 (nx23457)
             ) ;
    mux21_ni ix12423 (.Y (nx12422), .A0 (inputs_244__2), .A1 (inputs_245__2), .S0 (
             nx24059)) ;
    mux21_ni ix12435 (.Y (nx12434), .A0 (inputs_246__2), .A1 (inputs_247__2), .S0 (
             nx24059)) ;
    nand04 ix10860 (.Y (nx10859), .A0 (nx22255), .A1 (nx23457), .A2 (nx24059), .A3 (
           nx12382)) ;
    mux21_ni ix12383 (.Y (nx12382), .A0 (inputs_227__2), .A1 (inputs_243__2), .S0 (
             nx22757)) ;
    mux21_ni ix12369 (.Y (nx12368), .A0 (nx12304), .A1 (nx12364), .S0 (nx22759)
             ) ;
    mux21_ni ix12305 (.Y (nx12304), .A0 (nx12272), .A1 (nx12300), .S0 (nx23217)
             ) ;
    mux21_ni ix12273 (.Y (nx12272), .A0 (nx12256), .A1 (nx12268), .S0 (nx23457)
             ) ;
    mux21_ni ix12257 (.Y (nx12256), .A0 (inputs_232__2), .A1 (inputs_233__2), .S0 (
             nx24059)) ;
    mux21_ni ix12269 (.Y (nx12268), .A0 (inputs_234__2), .A1 (inputs_235__2), .S0 (
             nx24059)) ;
    mux21_ni ix12301 (.Y (nx12300), .A0 (nx12284), .A1 (nx12296), .S0 (nx23457)
             ) ;
    mux21_ni ix12285 (.Y (nx12284), .A0 (inputs_236__2), .A1 (inputs_237__2), .S0 (
             nx24059)) ;
    mux21_ni ix12297 (.Y (nx12296), .A0 (inputs_238__2), .A1 (inputs_239__2), .S0 (
             nx24059)) ;
    mux21_ni ix12365 (.Y (nx12364), .A0 (nx12332), .A1 (nx12360), .S0 (nx23217)
             ) ;
    mux21_ni ix12333 (.Y (nx12332), .A0 (nx12316), .A1 (nx12328), .S0 (nx23457)
             ) ;
    mux21_ni ix12317 (.Y (nx12316), .A0 (inputs_248__2), .A1 (inputs_249__2), .S0 (
             nx24061)) ;
    mux21_ni ix12329 (.Y (nx12328), .A0 (inputs_250__2), .A1 (inputs_251__2), .S0 (
             nx24061)) ;
    mux21_ni ix12361 (.Y (nx12360), .A0 (nx12344), .A1 (nx12356), .S0 (nx23457)
             ) ;
    mux21_ni ix12345 (.Y (nx12344), .A0 (inputs_252__2), .A1 (inputs_253__2), .S0 (
             nx24061)) ;
    mux21_ni ix12357 (.Y (nx12356), .A0 (inputs_254__2), .A1 (inputs_255__2), .S0 (
             nx24061)) ;
    oai21 ix16631 (.Y (\output [3]), .A0 (nx24851), .A1 (nx10887), .B0 (nx11241)
          ) ;
    mux21 ix10888 (.Y (nx10887), .A0 (nx13312), .A1 (nx14156), .S0 (nx22417)) ;
    mux21_ni ix13313 (.Y (nx13312), .A0 (nx12888), .A1 (nx13308), .S0 (nx22463)
             ) ;
    mux21_ni ix12889 (.Y (nx12888), .A0 (nx12676), .A1 (nx12884), .S0 (nx22553)
             ) ;
    mux21_ni ix12677 (.Y (nx12676), .A0 (nx12670), .A1 (nx12592), .S0 (nx23129)
             ) ;
    oai21 ix12671 (.Y (nx12670), .A0 (nx22255), .A1 (nx10897), .B0 (nx10907)) ;
    mux21 ix10898 (.Y (nx10897), .A0 (nx12634), .A1 (nx12662), .S0 (nx22759)) ;
    mux21_ni ix12635 (.Y (nx12634), .A0 (nx12618), .A1 (nx12630), .S0 (nx23457)
             ) ;
    mux21_ni ix12619 (.Y (nx12618), .A0 (inputs_260__3), .A1 (inputs_261__3), .S0 (
             nx24061)) ;
    mux21_ni ix12631 (.Y (nx12630), .A0 (inputs_262__3), .A1 (inputs_263__3), .S0 (
             nx24061)) ;
    mux21_ni ix12663 (.Y (nx12662), .A0 (nx12646), .A1 (nx12658), .S0 (nx23459)
             ) ;
    mux21_ni ix12647 (.Y (nx12646), .A0 (inputs_276__3), .A1 (inputs_277__3), .S0 (
             nx24061)) ;
    mux21_ni ix12659 (.Y (nx12658), .A0 (inputs_278__3), .A1 (inputs_279__3), .S0 (
             nx24063)) ;
    nand04 ix10908 (.Y (nx10907), .A0 (nx22255), .A1 (nx23459), .A2 (nx24063), .A3 (
           nx12606)) ;
    mux21_ni ix12607 (.Y (nx12606), .A0 (inputs_259__3), .A1 (inputs_275__3), .S0 (
             nx22759)) ;
    mux21_ni ix12593 (.Y (nx12592), .A0 (nx12528), .A1 (nx12588), .S0 (nx22759)
             ) ;
    mux21_ni ix12529 (.Y (nx12528), .A0 (nx12496), .A1 (nx12524), .S0 (nx23217)
             ) ;
    mux21_ni ix12497 (.Y (nx12496), .A0 (nx12480), .A1 (nx12492), .S0 (nx23459)
             ) ;
    mux21_ni ix12481 (.Y (nx12480), .A0 (inputs_264__3), .A1 (inputs_265__3), .S0 (
             nx24063)) ;
    mux21_ni ix12493 (.Y (nx12492), .A0 (inputs_266__3), .A1 (inputs_267__3), .S0 (
             nx24063)) ;
    mux21_ni ix12525 (.Y (nx12524), .A0 (nx12508), .A1 (nx12520), .S0 (nx23459)
             ) ;
    mux21_ni ix12509 (.Y (nx12508), .A0 (inputs_268__3), .A1 (inputs_269__3), .S0 (
             nx24063)) ;
    mux21_ni ix12521 (.Y (nx12520), .A0 (inputs_270__3), .A1 (inputs_271__3), .S0 (
             nx24063)) ;
    mux21_ni ix12589 (.Y (nx12588), .A0 (nx12556), .A1 (nx12584), .S0 (nx23217)
             ) ;
    mux21_ni ix12557 (.Y (nx12556), .A0 (nx12540), .A1 (nx12552), .S0 (nx23459)
             ) ;
    mux21_ni ix12541 (.Y (nx12540), .A0 (inputs_280__3), .A1 (inputs_281__3), .S0 (
             nx24063)) ;
    mux21_ni ix12553 (.Y (nx12552), .A0 (inputs_282__3), .A1 (inputs_283__3), .S0 (
             nx24065)) ;
    mux21_ni ix12585 (.Y (nx12584), .A0 (nx12568), .A1 (nx12580), .S0 (nx23459)
             ) ;
    mux21_ni ix12569 (.Y (nx12568), .A0 (inputs_284__3), .A1 (inputs_285__3), .S0 (
             nx24065)) ;
    mux21_ni ix12581 (.Y (nx12580), .A0 (inputs_286__3), .A1 (inputs_287__3), .S0 (
             nx24065)) ;
    mux21_ni ix12885 (.Y (nx12884), .A0 (nx12878), .A1 (nx12800), .S0 (nx23131)
             ) ;
    oai21 ix12879 (.Y (nx12878), .A0 (nx22255), .A1 (nx10939), .B0 (nx10949)) ;
    mux21 ix10940 (.Y (nx10939), .A0 (nx12842), .A1 (nx12870), .S0 (nx22759)) ;
    mux21_ni ix12843 (.Y (nx12842), .A0 (nx12826), .A1 (nx12838), .S0 (nx23459)
             ) ;
    mux21_ni ix12827 (.Y (nx12826), .A0 (inputs_292__3), .A1 (inputs_293__3), .S0 (
             nx24065)) ;
    mux21_ni ix12839 (.Y (nx12838), .A0 (inputs_294__3), .A1 (inputs_295__3), .S0 (
             nx24065)) ;
    mux21_ni ix12871 (.Y (nx12870), .A0 (nx12854), .A1 (nx12866), .S0 (nx23461)
             ) ;
    mux21_ni ix12855 (.Y (nx12854), .A0 (inputs_308__3), .A1 (inputs_309__3), .S0 (
             nx24065)) ;
    mux21_ni ix12867 (.Y (nx12866), .A0 (inputs_310__3), .A1 (inputs_311__3), .S0 (
             nx24065)) ;
    nand04 ix10950 (.Y (nx10949), .A0 (nx22255), .A1 (nx23461), .A2 (nx24067), .A3 (
           nx12814)) ;
    mux21_ni ix12815 (.Y (nx12814), .A0 (inputs_291__3), .A1 (inputs_307__3), .S0 (
             nx22759)) ;
    mux21_ni ix12801 (.Y (nx12800), .A0 (nx12736), .A1 (nx12796), .S0 (nx22759)
             ) ;
    mux21_ni ix12737 (.Y (nx12736), .A0 (nx12704), .A1 (nx12732), .S0 (nx23219)
             ) ;
    mux21_ni ix12705 (.Y (nx12704), .A0 (nx12688), .A1 (nx12700), .S0 (nx23461)
             ) ;
    mux21_ni ix12689 (.Y (nx12688), .A0 (inputs_296__3), .A1 (inputs_297__3), .S0 (
             nx24067)) ;
    mux21_ni ix12701 (.Y (nx12700), .A0 (inputs_298__3), .A1 (inputs_299__3), .S0 (
             nx24067)) ;
    mux21_ni ix12733 (.Y (nx12732), .A0 (nx12716), .A1 (nx12728), .S0 (nx23461)
             ) ;
    mux21_ni ix12717 (.Y (nx12716), .A0 (inputs_300__3), .A1 (inputs_301__3), .S0 (
             nx24067)) ;
    mux21_ni ix12729 (.Y (nx12728), .A0 (inputs_302__3), .A1 (inputs_303__3), .S0 (
             nx24067)) ;
    mux21_ni ix12797 (.Y (nx12796), .A0 (nx12764), .A1 (nx12792), .S0 (nx23219)
             ) ;
    mux21_ni ix12765 (.Y (nx12764), .A0 (nx12748), .A1 (nx12760), .S0 (nx23461)
             ) ;
    mux21_ni ix12749 (.Y (nx12748), .A0 (inputs_312__3), .A1 (inputs_313__3), .S0 (
             nx24067)) ;
    mux21_ni ix12761 (.Y (nx12760), .A0 (inputs_314__3), .A1 (inputs_315__3), .S0 (
             nx24067)) ;
    mux21_ni ix12793 (.Y (nx12792), .A0 (nx12776), .A1 (nx12788), .S0 (nx23461)
             ) ;
    mux21_ni ix12777 (.Y (nx12776), .A0 (inputs_316__3), .A1 (inputs_317__3), .S0 (
             nx24069)) ;
    mux21_ni ix12789 (.Y (nx12788), .A0 (inputs_318__3), .A1 (inputs_319__3), .S0 (
             nx24069)) ;
    mux21_ni ix13309 (.Y (nx13308), .A0 (nx13096), .A1 (nx13304), .S0 (nx22553)
             ) ;
    mux21_ni ix13097 (.Y (nx13096), .A0 (nx13090), .A1 (nx13012), .S0 (nx23131)
             ) ;
    oai21 ix13091 (.Y (nx13090), .A0 (nx22255), .A1 (nx10983), .B0 (nx10995)) ;
    mux21 ix10984 (.Y (nx10983), .A0 (nx13054), .A1 (nx13082), .S0 (nx22761)) ;
    mux21_ni ix13055 (.Y (nx13054), .A0 (nx13038), .A1 (nx13050), .S0 (nx23461)
             ) ;
    mux21_ni ix13039 (.Y (nx13038), .A0 (inputs_324__3), .A1 (inputs_325__3), .S0 (
             nx24069)) ;
    mux21_ni ix13051 (.Y (nx13050), .A0 (inputs_326__3), .A1 (inputs_327__3), .S0 (
             nx24069)) ;
    mux21_ni ix13083 (.Y (nx13082), .A0 (nx13066), .A1 (nx13078), .S0 (nx23463)
             ) ;
    mux21_ni ix13067 (.Y (nx13066), .A0 (inputs_340__3), .A1 (inputs_341__3), .S0 (
             nx24069)) ;
    mux21_ni ix13079 (.Y (nx13078), .A0 (inputs_342__3), .A1 (inputs_343__3), .S0 (
             nx24069)) ;
    nand04 ix10996 (.Y (nx10995), .A0 (nx22255), .A1 (nx23463), .A2 (nx24069), .A3 (
           nx13026)) ;
    mux21_ni ix13027 (.Y (nx13026), .A0 (inputs_323__3), .A1 (inputs_339__3), .S0 (
             nx22761)) ;
    mux21_ni ix13013 (.Y (nx13012), .A0 (nx12948), .A1 (nx13008), .S0 (nx22761)
             ) ;
    mux21_ni ix12949 (.Y (nx12948), .A0 (nx12916), .A1 (nx12944), .S0 (nx23219)
             ) ;
    mux21_ni ix12917 (.Y (nx12916), .A0 (nx12900), .A1 (nx12912), .S0 (nx23463)
             ) ;
    mux21_ni ix12901 (.Y (nx12900), .A0 (inputs_328__3), .A1 (inputs_329__3), .S0 (
             nx24071)) ;
    mux21_ni ix12913 (.Y (nx12912), .A0 (inputs_330__3), .A1 (inputs_331__3), .S0 (
             nx24071)) ;
    mux21_ni ix12945 (.Y (nx12944), .A0 (nx12928), .A1 (nx12940), .S0 (nx23463)
             ) ;
    mux21_ni ix12929 (.Y (nx12928), .A0 (inputs_332__3), .A1 (inputs_333__3), .S0 (
             nx24071)) ;
    mux21_ni ix12941 (.Y (nx12940), .A0 (inputs_334__3), .A1 (inputs_335__3), .S0 (
             nx24071)) ;
    mux21_ni ix13009 (.Y (nx13008), .A0 (nx12976), .A1 (nx13004), .S0 (nx23219)
             ) ;
    mux21_ni ix12977 (.Y (nx12976), .A0 (nx12960), .A1 (nx12972), .S0 (nx23463)
             ) ;
    mux21_ni ix12961 (.Y (nx12960), .A0 (inputs_344__3), .A1 (inputs_345__3), .S0 (
             nx24071)) ;
    mux21_ni ix12973 (.Y (nx12972), .A0 (inputs_346__3), .A1 (inputs_347__3), .S0 (
             nx24071)) ;
    mux21_ni ix13005 (.Y (nx13004), .A0 (nx12988), .A1 (nx13000), .S0 (nx23463)
             ) ;
    mux21_ni ix12989 (.Y (nx12988), .A0 (inputs_348__3), .A1 (inputs_349__3), .S0 (
             nx24071)) ;
    mux21_ni ix13001 (.Y (nx13000), .A0 (inputs_350__3), .A1 (inputs_351__3), .S0 (
             nx24073)) ;
    mux21_ni ix13305 (.Y (nx13304), .A0 (nx13298), .A1 (nx13220), .S0 (nx23131)
             ) ;
    oai21 ix13299 (.Y (nx13298), .A0 (nx22257), .A1 (nx11025), .B0 (nx11037)) ;
    mux21 ix11026 (.Y (nx11025), .A0 (nx13262), .A1 (nx13290), .S0 (nx22761)) ;
    mux21_ni ix13263 (.Y (nx13262), .A0 (nx13246), .A1 (nx13258), .S0 (nx23463)
             ) ;
    mux21_ni ix13247 (.Y (nx13246), .A0 (inputs_356__3), .A1 (inputs_357__3), .S0 (
             nx24073)) ;
    mux21_ni ix13259 (.Y (nx13258), .A0 (inputs_358__3), .A1 (inputs_359__3), .S0 (
             nx24073)) ;
    mux21_ni ix13291 (.Y (nx13290), .A0 (nx13274), .A1 (nx13286), .S0 (nx23465)
             ) ;
    mux21_ni ix13275 (.Y (nx13274), .A0 (inputs_372__3), .A1 (inputs_373__3), .S0 (
             nx24073)) ;
    mux21_ni ix13287 (.Y (nx13286), .A0 (inputs_374__3), .A1 (inputs_375__3), .S0 (
             nx24073)) ;
    nand04 ix11038 (.Y (nx11037), .A0 (nx22257), .A1 (nx23465), .A2 (nx24073), .A3 (
           nx13234)) ;
    mux21_ni ix13235 (.Y (nx13234), .A0 (inputs_355__3), .A1 (inputs_371__3), .S0 (
             nx22761)) ;
    mux21_ni ix13221 (.Y (nx13220), .A0 (nx13156), .A1 (nx13216), .S0 (nx22761)
             ) ;
    mux21_ni ix13157 (.Y (nx13156), .A0 (nx13124), .A1 (nx13152), .S0 (nx23219)
             ) ;
    mux21_ni ix13125 (.Y (nx13124), .A0 (nx13108), .A1 (nx13120), .S0 (nx23465)
             ) ;
    mux21_ni ix13109 (.Y (nx13108), .A0 (inputs_360__3), .A1 (inputs_361__3), .S0 (
             nx24073)) ;
    mux21_ni ix13121 (.Y (nx13120), .A0 (inputs_362__3), .A1 (inputs_363__3), .S0 (
             nx24075)) ;
    mux21_ni ix13153 (.Y (nx13152), .A0 (nx13136), .A1 (nx13148), .S0 (nx23465)
             ) ;
    mux21_ni ix13137 (.Y (nx13136), .A0 (inputs_364__3), .A1 (inputs_365__3), .S0 (
             nx24075)) ;
    mux21_ni ix13149 (.Y (nx13148), .A0 (inputs_366__3), .A1 (inputs_367__3), .S0 (
             nx24075)) ;
    mux21_ni ix13217 (.Y (nx13216), .A0 (nx13184), .A1 (nx13212), .S0 (nx23219)
             ) ;
    mux21_ni ix13185 (.Y (nx13184), .A0 (nx13168), .A1 (nx13180), .S0 (nx23465)
             ) ;
    mux21_ni ix13169 (.Y (nx13168), .A0 (inputs_376__3), .A1 (inputs_377__3), .S0 (
             nx24075)) ;
    mux21_ni ix13181 (.Y (nx13180), .A0 (inputs_378__3), .A1 (inputs_379__3), .S0 (
             nx24075)) ;
    mux21_ni ix13213 (.Y (nx13212), .A0 (nx13196), .A1 (nx13208), .S0 (nx23465)
             ) ;
    mux21_ni ix13197 (.Y (nx13196), .A0 (inputs_380__3), .A1 (inputs_381__3), .S0 (
             nx24075)) ;
    mux21_ni ix13209 (.Y (nx13208), .A0 (inputs_382__3), .A1 (inputs_383__3), .S0 (
             nx24075)) ;
    mux21_ni ix14157 (.Y (nx14156), .A0 (nx13732), .A1 (nx14152), .S0 (nx22465)
             ) ;
    mux21_ni ix13733 (.Y (nx13732), .A0 (nx13520), .A1 (nx13728), .S0 (nx22555)
             ) ;
    mux21_ni ix13521 (.Y (nx13520), .A0 (nx13514), .A1 (nx13436), .S0 (nx23131)
             ) ;
    oai21 ix13515 (.Y (nx13514), .A0 (nx22257), .A1 (nx11071), .B0 (nx11083)) ;
    mux21 ix11072 (.Y (nx11071), .A0 (nx13478), .A1 (nx13506), .S0 (nx22761)) ;
    mux21_ni ix13479 (.Y (nx13478), .A0 (nx13462), .A1 (nx13474), .S0 (nx23465)
             ) ;
    mux21_ni ix13463 (.Y (nx13462), .A0 (inputs_388__3), .A1 (inputs_389__3), .S0 (
             nx24077)) ;
    mux21_ni ix13475 (.Y (nx13474), .A0 (inputs_390__3), .A1 (inputs_391__3), .S0 (
             nx24077)) ;
    mux21_ni ix13507 (.Y (nx13506), .A0 (nx13490), .A1 (nx13502), .S0 (nx23467)
             ) ;
    mux21_ni ix13491 (.Y (nx13490), .A0 (inputs_404__3), .A1 (inputs_405__3), .S0 (
             nx24077)) ;
    mux21_ni ix13503 (.Y (nx13502), .A0 (inputs_406__3), .A1 (inputs_407__3), .S0 (
             nx24077)) ;
    nand04 ix11084 (.Y (nx11083), .A0 (nx22257), .A1 (nx23467), .A2 (nx24077), .A3 (
           nx13450)) ;
    mux21_ni ix13451 (.Y (nx13450), .A0 (inputs_387__3), .A1 (inputs_403__3), .S0 (
             nx22763)) ;
    mux21_ni ix13437 (.Y (nx13436), .A0 (nx13372), .A1 (nx13432), .S0 (nx22763)
             ) ;
    mux21_ni ix13373 (.Y (nx13372), .A0 (nx13340), .A1 (nx13368), .S0 (nx23219)
             ) ;
    mux21_ni ix13341 (.Y (nx13340), .A0 (nx13324), .A1 (nx13336), .S0 (nx23467)
             ) ;
    mux21_ni ix13325 (.Y (nx13324), .A0 (inputs_392__3), .A1 (inputs_393__3), .S0 (
             nx24077)) ;
    mux21_ni ix13337 (.Y (nx13336), .A0 (inputs_394__3), .A1 (inputs_395__3), .S0 (
             nx24077)) ;
    mux21_ni ix13369 (.Y (nx13368), .A0 (nx13352), .A1 (nx13364), .S0 (nx23467)
             ) ;
    mux21_ni ix13353 (.Y (nx13352), .A0 (inputs_396__3), .A1 (inputs_397__3), .S0 (
             nx24079)) ;
    mux21_ni ix13365 (.Y (nx13364), .A0 (inputs_398__3), .A1 (inputs_399__3), .S0 (
             nx24079)) ;
    mux21_ni ix13433 (.Y (nx13432), .A0 (nx13400), .A1 (nx13428), .S0 (nx23221)
             ) ;
    mux21_ni ix13401 (.Y (nx13400), .A0 (nx13384), .A1 (nx13396), .S0 (nx23467)
             ) ;
    mux21_ni ix13385 (.Y (nx13384), .A0 (inputs_408__3), .A1 (inputs_409__3), .S0 (
             nx24079)) ;
    mux21_ni ix13397 (.Y (nx13396), .A0 (inputs_410__3), .A1 (inputs_411__3), .S0 (
             nx24079)) ;
    mux21_ni ix13429 (.Y (nx13428), .A0 (nx13412), .A1 (nx13424), .S0 (nx23467)
             ) ;
    mux21_ni ix13413 (.Y (nx13412), .A0 (inputs_412__3), .A1 (inputs_413__3), .S0 (
             nx24079)) ;
    mux21_ni ix13425 (.Y (nx13424), .A0 (inputs_414__3), .A1 (inputs_415__3), .S0 (
             nx24079)) ;
    mux21_ni ix13729 (.Y (nx13728), .A0 (nx13722), .A1 (nx13644), .S0 (nx23131)
             ) ;
    oai21 ix13723 (.Y (nx13722), .A0 (nx22257), .A1 (nx11115), .B0 (nx11127)) ;
    mux21 ix11116 (.Y (nx11115), .A0 (nx13686), .A1 (nx13714), .S0 (nx22763)) ;
    mux21_ni ix13687 (.Y (nx13686), .A0 (nx13670), .A1 (nx13682), .S0 (nx23467)
             ) ;
    mux21_ni ix13671 (.Y (nx13670), .A0 (inputs_420__3), .A1 (inputs_421__3), .S0 (
             nx24079)) ;
    mux21_ni ix13683 (.Y (nx13682), .A0 (inputs_422__3), .A1 (inputs_423__3), .S0 (
             nx24081)) ;
    mux21_ni ix13715 (.Y (nx13714), .A0 (nx13698), .A1 (nx13710), .S0 (nx23469)
             ) ;
    mux21_ni ix13699 (.Y (nx13698), .A0 (inputs_436__3), .A1 (inputs_437__3), .S0 (
             nx24081)) ;
    mux21_ni ix13711 (.Y (nx13710), .A0 (inputs_438__3), .A1 (inputs_439__3), .S0 (
             nx24081)) ;
    nand04 ix11128 (.Y (nx11127), .A0 (nx22257), .A1 (nx23469), .A2 (nx24081), .A3 (
           nx13658)) ;
    mux21_ni ix13659 (.Y (nx13658), .A0 (inputs_419__3), .A1 (inputs_435__3), .S0 (
             nx22763)) ;
    mux21_ni ix13645 (.Y (nx13644), .A0 (nx13580), .A1 (nx13640), .S0 (nx22763)
             ) ;
    mux21_ni ix13581 (.Y (nx13580), .A0 (nx13548), .A1 (nx13576), .S0 (nx23221)
             ) ;
    mux21_ni ix13549 (.Y (nx13548), .A0 (nx13532), .A1 (nx13544), .S0 (nx23469)
             ) ;
    mux21_ni ix13533 (.Y (nx13532), .A0 (inputs_424__3), .A1 (inputs_425__3), .S0 (
             nx24081)) ;
    mux21_ni ix13545 (.Y (nx13544), .A0 (inputs_426__3), .A1 (inputs_427__3), .S0 (
             nx24081)) ;
    mux21_ni ix13577 (.Y (nx13576), .A0 (nx13560), .A1 (nx13572), .S0 (nx23469)
             ) ;
    mux21_ni ix13561 (.Y (nx13560), .A0 (inputs_428__3), .A1 (inputs_429__3), .S0 (
             nx24081)) ;
    mux21_ni ix13573 (.Y (nx13572), .A0 (inputs_430__3), .A1 (inputs_431__3), .S0 (
             nx24083)) ;
    mux21_ni ix13641 (.Y (nx13640), .A0 (nx13608), .A1 (nx13636), .S0 (nx23221)
             ) ;
    mux21_ni ix13609 (.Y (nx13608), .A0 (nx13592), .A1 (nx13604), .S0 (nx23469)
             ) ;
    mux21_ni ix13593 (.Y (nx13592), .A0 (inputs_440__3), .A1 (inputs_441__3), .S0 (
             nx24083)) ;
    mux21_ni ix13605 (.Y (nx13604), .A0 (inputs_442__3), .A1 (inputs_443__3), .S0 (
             nx24083)) ;
    mux21_ni ix13637 (.Y (nx13636), .A0 (nx13620), .A1 (nx13632), .S0 (nx23469)
             ) ;
    mux21_ni ix13621 (.Y (nx13620), .A0 (inputs_444__3), .A1 (inputs_445__3), .S0 (
             nx24083)) ;
    mux21_ni ix13633 (.Y (nx13632), .A0 (inputs_446__3), .A1 (inputs_447__3), .S0 (
             nx24083)) ;
    mux21_ni ix14153 (.Y (nx14152), .A0 (nx13940), .A1 (nx14148), .S0 (nx22555)
             ) ;
    mux21_ni ix13941 (.Y (nx13940), .A0 (nx13934), .A1 (nx13856), .S0 (nx23131)
             ) ;
    oai21 ix13935 (.Y (nx13934), .A0 (nx22257), .A1 (nx11159), .B0 (nx11169)) ;
    mux21 ix11160 (.Y (nx11159), .A0 (nx13898), .A1 (nx13926), .S0 (nx22763)) ;
    mux21_ni ix13899 (.Y (nx13898), .A0 (nx13882), .A1 (nx13894), .S0 (nx23469)
             ) ;
    mux21_ni ix13883 (.Y (nx13882), .A0 (inputs_452__3), .A1 (inputs_453__3), .S0 (
             nx24083)) ;
    mux21_ni ix13895 (.Y (nx13894), .A0 (inputs_454__3), .A1 (inputs_455__3), .S0 (
             nx24083)) ;
    mux21_ni ix13927 (.Y (nx13926), .A0 (nx13910), .A1 (nx13922), .S0 (nx23471)
             ) ;
    mux21_ni ix13911 (.Y (nx13910), .A0 (inputs_468__3), .A1 (inputs_469__3), .S0 (
             nx24085)) ;
    mux21_ni ix13923 (.Y (nx13922), .A0 (inputs_470__3), .A1 (inputs_471__3), .S0 (
             nx24085)) ;
    nand04 ix11170 (.Y (nx11169), .A0 (nx22259), .A1 (nx23471), .A2 (nx24085), .A3 (
           nx13870)) ;
    mux21_ni ix13871 (.Y (nx13870), .A0 (inputs_451__3), .A1 (inputs_467__3), .S0 (
             nx22763)) ;
    mux21_ni ix13857 (.Y (nx13856), .A0 (nx13792), .A1 (nx13852), .S0 (nx22765)
             ) ;
    mux21_ni ix13793 (.Y (nx13792), .A0 (nx13760), .A1 (nx13788), .S0 (nx23221)
             ) ;
    mux21_ni ix13761 (.Y (nx13760), .A0 (nx13744), .A1 (nx13756), .S0 (nx23471)
             ) ;
    mux21_ni ix13745 (.Y (nx13744), .A0 (inputs_456__3), .A1 (inputs_457__3), .S0 (
             nx24085)) ;
    mux21_ni ix13757 (.Y (nx13756), .A0 (inputs_458__3), .A1 (inputs_459__3), .S0 (
             nx24085)) ;
    mux21_ni ix13789 (.Y (nx13788), .A0 (nx13772), .A1 (nx13784), .S0 (nx23471)
             ) ;
    mux21_ni ix13773 (.Y (nx13772), .A0 (inputs_460__3), .A1 (inputs_461__3), .S0 (
             nx24085)) ;
    mux21_ni ix13785 (.Y (nx13784), .A0 (inputs_462__3), .A1 (inputs_463__3), .S0 (
             nx24085)) ;
    mux21_ni ix13853 (.Y (nx13852), .A0 (nx13820), .A1 (nx13848), .S0 (nx23221)
             ) ;
    mux21_ni ix13821 (.Y (nx13820), .A0 (nx13804), .A1 (nx13816), .S0 (nx23471)
             ) ;
    mux21_ni ix13805 (.Y (nx13804), .A0 (inputs_472__3), .A1 (inputs_473__3), .S0 (
             nx24087)) ;
    mux21_ni ix13817 (.Y (nx13816), .A0 (inputs_474__3), .A1 (inputs_475__3), .S0 (
             nx24087)) ;
    mux21_ni ix13849 (.Y (nx13848), .A0 (nx13832), .A1 (nx13844), .S0 (nx23471)
             ) ;
    mux21_ni ix13833 (.Y (nx13832), .A0 (inputs_476__3), .A1 (inputs_477__3), .S0 (
             nx24087)) ;
    mux21_ni ix13845 (.Y (nx13844), .A0 (inputs_478__3), .A1 (inputs_479__3), .S0 (
             nx24087)) ;
    mux21_ni ix14149 (.Y (nx14148), .A0 (nx14142), .A1 (nx14064), .S0 (nx23131)
             ) ;
    oai21 ix14143 (.Y (nx14142), .A0 (nx22259), .A1 (nx11201), .B0 (nx11213)) ;
    mux21 ix11202 (.Y (nx11201), .A0 (nx14106), .A1 (nx14134), .S0 (nx22765)) ;
    mux21_ni ix14107 (.Y (nx14106), .A0 (nx14090), .A1 (nx14102), .S0 (nx23471)
             ) ;
    mux21_ni ix14091 (.Y (nx14090), .A0 (inputs_484__3), .A1 (inputs_485__3), .S0 (
             nx24087)) ;
    mux21_ni ix14103 (.Y (nx14102), .A0 (inputs_486__3), .A1 (inputs_487__3), .S0 (
             nx24087)) ;
    mux21_ni ix14135 (.Y (nx14134), .A0 (nx14118), .A1 (nx14130), .S0 (nx23473)
             ) ;
    mux21_ni ix14119 (.Y (nx14118), .A0 (inputs_500__3), .A1 (inputs_501__3), .S0 (
             nx24087)) ;
    mux21_ni ix14131 (.Y (nx14130), .A0 (inputs_502__3), .A1 (inputs_503__3), .S0 (
             nx24089)) ;
    nand04 ix11214 (.Y (nx11213), .A0 (nx22259), .A1 (nx23473), .A2 (nx24089), .A3 (
           nx14078)) ;
    mux21_ni ix14079 (.Y (nx14078), .A0 (inputs_483__3), .A1 (inputs_499__3), .S0 (
             nx22765)) ;
    mux21_ni ix14065 (.Y (nx14064), .A0 (nx14000), .A1 (nx14060), .S0 (nx22765)
             ) ;
    mux21_ni ix14001 (.Y (nx14000), .A0 (nx13968), .A1 (nx13996), .S0 (nx23221)
             ) ;
    mux21_ni ix13969 (.Y (nx13968), .A0 (nx13952), .A1 (nx13964), .S0 (nx23473)
             ) ;
    mux21_ni ix13953 (.Y (nx13952), .A0 (inputs_488__3), .A1 (inputs_489__3), .S0 (
             nx24089)) ;
    mux21_ni ix13965 (.Y (nx13964), .A0 (inputs_490__3), .A1 (inputs_491__3), .S0 (
             nx24089)) ;
    mux21_ni ix13997 (.Y (nx13996), .A0 (nx13980), .A1 (nx13992), .S0 (nx23473)
             ) ;
    mux21_ni ix13981 (.Y (nx13980), .A0 (inputs_492__3), .A1 (inputs_493__3), .S0 (
             nx24089)) ;
    mux21_ni ix13993 (.Y (nx13992), .A0 (inputs_494__3), .A1 (inputs_495__3), .S0 (
             nx24089)) ;
    mux21_ni ix14061 (.Y (nx14060), .A0 (nx14028), .A1 (nx14056), .S0 (nx23221)
             ) ;
    mux21_ni ix14029 (.Y (nx14028), .A0 (nx14012), .A1 (nx14024), .S0 (nx23473)
             ) ;
    mux21_ni ix14013 (.Y (nx14012), .A0 (inputs_504__3), .A1 (inputs_505__3), .S0 (
             nx24089)) ;
    mux21_ni ix14025 (.Y (nx14024), .A0 (inputs_506__3), .A1 (inputs_507__3), .S0 (
             nx24091)) ;
    mux21_ni ix14057 (.Y (nx14056), .A0 (nx14040), .A1 (nx14052), .S0 (nx23473)
             ) ;
    mux21_ni ix14041 (.Y (nx14040), .A0 (inputs_508__3), .A1 (inputs_509__3), .S0 (
             nx24091)) ;
    mux21_ni ix14053 (.Y (nx14052), .A0 (inputs_510__3), .A1 (inputs_511__3), .S0 (
             nx24091)) ;
    aoi32 ix11242 (.Y (nx11241), .A0 (nx14926), .A1 (nx22385), .A2 (nx22259), .B0 (
          nx22219), .B1 (nx16622)) ;
    oai21 ix14927 (.Y (nx14926), .A0 (nx23473), .A1 (nx11245), .B0 (nx11347)) ;
    mux21 ix11246 (.Y (nx11245), .A0 (nx14664), .A1 (nx14916), .S0 (nx24091)) ;
    mux21_ni ix14665 (.Y (nx14664), .A0 (nx14536), .A1 (nx14660), .S0 (nx22395)
             ) ;
    mux21_ni ix14537 (.Y (nx14536), .A0 (nx14472), .A1 (nx14532), .S0 (nx22417)
             ) ;
    mux21_ni ix14473 (.Y (nx14472), .A0 (nx14440), .A1 (nx14468), .S0 (nx22465)
             ) ;
    mux21_ni ix14441 (.Y (nx14440), .A0 (nx14424), .A1 (nx14436), .S0 (nx22555)
             ) ;
    mux21_ni ix14425 (.Y (nx14424), .A0 (inputs_0__3), .A1 (inputs_16__3), .S0 (
             nx22765)) ;
    mux21_ni ix14437 (.Y (nx14436), .A0 (inputs_32__3), .A1 (inputs_48__3), .S0 (
             nx22765)) ;
    mux21_ni ix14469 (.Y (nx14468), .A0 (nx14452), .A1 (nx14464), .S0 (nx22555)
             ) ;
    mux21_ni ix14453 (.Y (nx14452), .A0 (inputs_64__3), .A1 (inputs_80__3), .S0 (
             nx22765)) ;
    mux21_ni ix14465 (.Y (nx14464), .A0 (inputs_96__3), .A1 (inputs_112__3), .S0 (
             nx22767)) ;
    mux21_ni ix14533 (.Y (nx14532), .A0 (nx14500), .A1 (nx14528), .S0 (nx22465)
             ) ;
    mux21_ni ix14501 (.Y (nx14500), .A0 (nx14484), .A1 (nx14496), .S0 (nx22555)
             ) ;
    mux21_ni ix14485 (.Y (nx14484), .A0 (inputs_128__3), .A1 (inputs_144__3), .S0 (
             nx22767)) ;
    mux21_ni ix14497 (.Y (nx14496), .A0 (inputs_160__3), .A1 (inputs_176__3), .S0 (
             nx22767)) ;
    mux21_ni ix14529 (.Y (nx14528), .A0 (nx14512), .A1 (nx14524), .S0 (nx22555)
             ) ;
    mux21_ni ix14513 (.Y (nx14512), .A0 (inputs_192__3), .A1 (inputs_208__3), .S0 (
             nx22767)) ;
    mux21_ni ix14525 (.Y (nx14524), .A0 (inputs_224__3), .A1 (inputs_240__3), .S0 (
             nx22767)) ;
    mux21_ni ix14661 (.Y (nx14660), .A0 (nx14596), .A1 (nx14656), .S0 (nx22417)
             ) ;
    mux21_ni ix14597 (.Y (nx14596), .A0 (nx14564), .A1 (nx14592), .S0 (nx22465)
             ) ;
    mux21_ni ix14565 (.Y (nx14564), .A0 (nx14548), .A1 (nx14560), .S0 (nx22555)
             ) ;
    mux21_ni ix14549 (.Y (nx14548), .A0 (inputs_256__3), .A1 (inputs_272__3), .S0 (
             nx22767)) ;
    mux21_ni ix14561 (.Y (nx14560), .A0 (inputs_288__3), .A1 (inputs_304__3), .S0 (
             nx22767)) ;
    mux21_ni ix14593 (.Y (nx14592), .A0 (nx14576), .A1 (nx14588), .S0 (nx22557)
             ) ;
    mux21_ni ix14577 (.Y (nx14576), .A0 (inputs_320__3), .A1 (inputs_336__3), .S0 (
             nx22769)) ;
    mux21_ni ix14589 (.Y (nx14588), .A0 (inputs_352__3), .A1 (inputs_368__3), .S0 (
             nx22769)) ;
    mux21_ni ix14657 (.Y (nx14656), .A0 (nx14624), .A1 (nx14652), .S0 (nx22465)
             ) ;
    mux21_ni ix14625 (.Y (nx14624), .A0 (nx14608), .A1 (nx14620), .S0 (nx22557)
             ) ;
    mux21_ni ix14609 (.Y (nx14608), .A0 (inputs_384__3), .A1 (inputs_400__3), .S0 (
             nx22769)) ;
    mux21_ni ix14621 (.Y (nx14620), .A0 (inputs_416__3), .A1 (inputs_432__3), .S0 (
             nx22769)) ;
    mux21_ni ix14653 (.Y (nx14652), .A0 (nx14636), .A1 (nx14648), .S0 (nx22557)
             ) ;
    mux21_ni ix14637 (.Y (nx14636), .A0 (inputs_448__3), .A1 (inputs_464__3), .S0 (
             nx22769)) ;
    mux21_ni ix14649 (.Y (nx14648), .A0 (inputs_480__3), .A1 (inputs_496__3), .S0 (
             nx22769)) ;
    mux21_ni ix14917 (.Y (nx14916), .A0 (nx14788), .A1 (nx14912), .S0 (nx22395)
             ) ;
    mux21_ni ix14789 (.Y (nx14788), .A0 (nx14724), .A1 (nx14784), .S0 (nx22417)
             ) ;
    mux21_ni ix14725 (.Y (nx14724), .A0 (nx14692), .A1 (nx14720), .S0 (nx22465)
             ) ;
    mux21_ni ix14693 (.Y (nx14692), .A0 (nx14676), .A1 (nx14688), .S0 (nx22557)
             ) ;
    mux21_ni ix14677 (.Y (nx14676), .A0 (inputs_1__3), .A1 (inputs_17__3), .S0 (
             nx22769)) ;
    mux21_ni ix14689 (.Y (nx14688), .A0 (inputs_33__3), .A1 (inputs_49__3), .S0 (
             nx22771)) ;
    mux21_ni ix14721 (.Y (nx14720), .A0 (nx14704), .A1 (nx14716), .S0 (nx22557)
             ) ;
    mux21_ni ix14705 (.Y (nx14704), .A0 (inputs_65__3), .A1 (inputs_81__3), .S0 (
             nx22771)) ;
    mux21_ni ix14717 (.Y (nx14716), .A0 (inputs_97__3), .A1 (inputs_113__3), .S0 (
             nx22771)) ;
    mux21_ni ix14785 (.Y (nx14784), .A0 (nx14752), .A1 (nx14780), .S0 (nx22465)
             ) ;
    mux21_ni ix14753 (.Y (nx14752), .A0 (nx14736), .A1 (nx14748), .S0 (nx22557)
             ) ;
    mux21_ni ix14737 (.Y (nx14736), .A0 (inputs_129__3), .A1 (inputs_145__3), .S0 (
             nx22771)) ;
    mux21_ni ix14749 (.Y (nx14748), .A0 (inputs_161__3), .A1 (inputs_177__3), .S0 (
             nx22771)) ;
    mux21_ni ix14781 (.Y (nx14780), .A0 (nx14764), .A1 (nx14776), .S0 (nx22557)
             ) ;
    mux21_ni ix14765 (.Y (nx14764), .A0 (inputs_193__3), .A1 (inputs_209__3), .S0 (
             nx22771)) ;
    mux21_ni ix14777 (.Y (nx14776), .A0 (inputs_225__3), .A1 (inputs_241__3), .S0 (
             nx22771)) ;
    mux21_ni ix14913 (.Y (nx14912), .A0 (nx14848), .A1 (nx14908), .S0 (nx22419)
             ) ;
    mux21_ni ix14849 (.Y (nx14848), .A0 (nx14816), .A1 (nx14844), .S0 (nx22467)
             ) ;
    mux21_ni ix14817 (.Y (nx14816), .A0 (nx14800), .A1 (nx14812), .S0 (nx22559)
             ) ;
    mux21_ni ix14801 (.Y (nx14800), .A0 (inputs_257__3), .A1 (inputs_273__3), .S0 (
             nx22773)) ;
    mux21_ni ix14813 (.Y (nx14812), .A0 (inputs_289__3), .A1 (inputs_305__3), .S0 (
             nx22773)) ;
    mux21_ni ix14845 (.Y (nx14844), .A0 (nx14828), .A1 (nx14840), .S0 (nx22559)
             ) ;
    mux21_ni ix14829 (.Y (nx14828), .A0 (inputs_321__3), .A1 (inputs_337__3), .S0 (
             nx22773)) ;
    mux21_ni ix14841 (.Y (nx14840), .A0 (inputs_353__3), .A1 (inputs_369__3), .S0 (
             nx22773)) ;
    mux21_ni ix14909 (.Y (nx14908), .A0 (nx14876), .A1 (nx14904), .S0 (nx22467)
             ) ;
    mux21_ni ix14877 (.Y (nx14876), .A0 (nx14860), .A1 (nx14872), .S0 (nx22559)
             ) ;
    mux21_ni ix14861 (.Y (nx14860), .A0 (inputs_385__3), .A1 (inputs_401__3), .S0 (
             nx22773)) ;
    mux21_ni ix14873 (.Y (nx14872), .A0 (inputs_417__3), .A1 (inputs_433__3), .S0 (
             nx22773)) ;
    mux21_ni ix14905 (.Y (nx14904), .A0 (nx14888), .A1 (nx14900), .S0 (nx22559)
             ) ;
    mux21_ni ix14889 (.Y (nx14888), .A0 (inputs_449__3), .A1 (inputs_465__3), .S0 (
             nx22773)) ;
    mux21_ni ix14901 (.Y (nx14900), .A0 (inputs_481__3), .A1 (inputs_497__3), .S0 (
             nx22775)) ;
    nand03 ix11348 (.Y (nx11347), .A0 (nx14410), .A1 (nx23475), .A2 (nx24879)) ;
    mux21_ni ix14411 (.Y (nx14410), .A0 (nx14282), .A1 (nx14406), .S0 (nx22395)
             ) ;
    mux21_ni ix14283 (.Y (nx14282), .A0 (nx14218), .A1 (nx14278), .S0 (nx22419)
             ) ;
    mux21_ni ix14219 (.Y (nx14218), .A0 (nx14186), .A1 (nx14214), .S0 (nx22467)
             ) ;
    mux21_ni ix14187 (.Y (nx14186), .A0 (nx14170), .A1 (nx14182), .S0 (nx22559)
             ) ;
    mux21_ni ix14171 (.Y (nx14170), .A0 (inputs_2__3), .A1 (inputs_18__3), .S0 (
             nx22775)) ;
    mux21_ni ix14183 (.Y (nx14182), .A0 (inputs_34__3), .A1 (inputs_50__3), .S0 (
             nx22775)) ;
    mux21_ni ix14215 (.Y (nx14214), .A0 (nx14198), .A1 (nx14210), .S0 (nx22559)
             ) ;
    mux21_ni ix14199 (.Y (nx14198), .A0 (inputs_66__3), .A1 (inputs_82__3), .S0 (
             nx22775)) ;
    mux21_ni ix14211 (.Y (nx14210), .A0 (inputs_98__3), .A1 (inputs_114__3), .S0 (
             nx22775)) ;
    mux21_ni ix14279 (.Y (nx14278), .A0 (nx14246), .A1 (nx14274), .S0 (nx22467)
             ) ;
    mux21_ni ix14247 (.Y (nx14246), .A0 (nx14230), .A1 (nx14242), .S0 (nx22559)
             ) ;
    mux21_ni ix14231 (.Y (nx14230), .A0 (inputs_130__3), .A1 (inputs_146__3), .S0 (
             nx22775)) ;
    mux21_ni ix14243 (.Y (nx14242), .A0 (inputs_162__3), .A1 (inputs_178__3), .S0 (
             nx22775)) ;
    mux21_ni ix14275 (.Y (nx14274), .A0 (nx14258), .A1 (nx14270), .S0 (nx22561)
             ) ;
    mux21_ni ix14259 (.Y (nx14258), .A0 (inputs_194__3), .A1 (inputs_210__3), .S0 (
             nx22777)) ;
    mux21_ni ix14271 (.Y (nx14270), .A0 (inputs_226__3), .A1 (inputs_242__3), .S0 (
             nx22777)) ;
    mux21_ni ix14407 (.Y (nx14406), .A0 (nx14342), .A1 (nx14402), .S0 (nx22419)
             ) ;
    mux21_ni ix14343 (.Y (nx14342), .A0 (nx14310), .A1 (nx14338), .S0 (nx22467)
             ) ;
    mux21_ni ix14311 (.Y (nx14310), .A0 (nx14294), .A1 (nx14306), .S0 (nx22561)
             ) ;
    mux21_ni ix14295 (.Y (nx14294), .A0 (inputs_258__3), .A1 (inputs_274__3), .S0 (
             nx22777)) ;
    mux21_ni ix14307 (.Y (nx14306), .A0 (inputs_290__3), .A1 (inputs_306__3), .S0 (
             nx22777)) ;
    mux21_ni ix14339 (.Y (nx14338), .A0 (nx14322), .A1 (nx14334), .S0 (nx22561)
             ) ;
    mux21_ni ix14323 (.Y (nx14322), .A0 (inputs_322__3), .A1 (inputs_338__3), .S0 (
             nx22777)) ;
    mux21_ni ix14335 (.Y (nx14334), .A0 (inputs_354__3), .A1 (inputs_370__3), .S0 (
             nx22777)) ;
    mux21_ni ix14403 (.Y (nx14402), .A0 (nx14370), .A1 (nx14398), .S0 (nx22467)
             ) ;
    mux21_ni ix14371 (.Y (nx14370), .A0 (nx14354), .A1 (nx14366), .S0 (nx22561)
             ) ;
    mux21_ni ix14355 (.Y (nx14354), .A0 (inputs_386__3), .A1 (inputs_402__3), .S0 (
             nx22777)) ;
    mux21_ni ix14367 (.Y (nx14366), .A0 (inputs_418__3), .A1 (inputs_434__3), .S0 (
             nx22779)) ;
    mux21_ni ix14399 (.Y (nx14398), .A0 (nx14382), .A1 (nx14394), .S0 (nx22561)
             ) ;
    mux21_ni ix14383 (.Y (nx14382), .A0 (inputs_450__3), .A1 (inputs_466__3), .S0 (
             nx22779)) ;
    mux21_ni ix14395 (.Y (nx14394), .A0 (inputs_482__3), .A1 (inputs_498__3), .S0 (
             nx22779)) ;
    mux21_ni ix16623 (.Y (nx16622), .A0 (nx15774), .A1 (nx16618), .S0 (nx22419)
             ) ;
    mux21_ni ix15775 (.Y (nx15774), .A0 (nx15350), .A1 (nx15770), .S0 (nx22467)
             ) ;
    mux21_ni ix15351 (.Y (nx15350), .A0 (nx15138), .A1 (nx15346), .S0 (nx22561)
             ) ;
    mux21_ni ix15139 (.Y (nx15138), .A0 (nx15132), .A1 (nx15054), .S0 (nx23133)
             ) ;
    oai21 ix15133 (.Y (nx15132), .A0 (nx22259), .A1 (nx11407), .B0 (nx11419)) ;
    mux21 ix11408 (.Y (nx11407), .A0 (nx15096), .A1 (nx15124), .S0 (nx22779)) ;
    mux21_ni ix15097 (.Y (nx15096), .A0 (nx15080), .A1 (nx15092), .S0 (nx23475)
             ) ;
    mux21_ni ix15081 (.Y (nx15080), .A0 (inputs_4__3), .A1 (inputs_5__3), .S0 (
             nx24091)) ;
    mux21_ni ix15093 (.Y (nx15092), .A0 (inputs_6__3), .A1 (inputs_7__3), .S0 (
             nx24091)) ;
    mux21_ni ix15125 (.Y (nx15124), .A0 (nx15108), .A1 (nx15120), .S0 (nx23475)
             ) ;
    mux21_ni ix15109 (.Y (nx15108), .A0 (inputs_20__3), .A1 (inputs_21__3), .S0 (
             nx24091)) ;
    mux21_ni ix15121 (.Y (nx15120), .A0 (inputs_22__3), .A1 (inputs_23__3), .S0 (
             nx24093)) ;
    nand04 ix11420 (.Y (nx11419), .A0 (nx22259), .A1 (nx23475), .A2 (nx24093), .A3 (
           nx15068)) ;
    mux21_ni ix15069 (.Y (nx15068), .A0 (inputs_3__3), .A1 (inputs_19__3), .S0 (
             nx22779)) ;
    mux21_ni ix15055 (.Y (nx15054), .A0 (nx14990), .A1 (nx15050), .S0 (nx22779)
             ) ;
    mux21_ni ix14991 (.Y (nx14990), .A0 (nx14958), .A1 (nx14986), .S0 (nx23223)
             ) ;
    mux21_ni ix14959 (.Y (nx14958), .A0 (nx14942), .A1 (nx14954), .S0 (nx23475)
             ) ;
    mux21_ni ix14943 (.Y (nx14942), .A0 (inputs_8__3), .A1 (inputs_9__3), .S0 (
             nx24093)) ;
    mux21_ni ix14955 (.Y (nx14954), .A0 (inputs_10__3), .A1 (inputs_11__3), .S0 (
             nx24093)) ;
    mux21_ni ix14987 (.Y (nx14986), .A0 (nx14970), .A1 (nx14982), .S0 (nx23475)
             ) ;
    mux21_ni ix14971 (.Y (nx14970), .A0 (inputs_12__3), .A1 (inputs_13__3), .S0 (
             nx24093)) ;
    mux21_ni ix14983 (.Y (nx14982), .A0 (inputs_14__3), .A1 (inputs_15__3), .S0 (
             nx24093)) ;
    mux21_ni ix15051 (.Y (nx15050), .A0 (nx15018), .A1 (nx15046), .S0 (nx23223)
             ) ;
    mux21_ni ix15019 (.Y (nx15018), .A0 (nx15002), .A1 (nx15014), .S0 (nx23475)
             ) ;
    mux21_ni ix15003 (.Y (nx15002), .A0 (inputs_24__3), .A1 (inputs_25__3), .S0 (
             nx24093)) ;
    mux21_ni ix15015 (.Y (nx15014), .A0 (inputs_26__3), .A1 (inputs_27__3), .S0 (
             nx24095)) ;
    mux21_ni ix15047 (.Y (nx15046), .A0 (nx15030), .A1 (nx15042), .S0 (nx23477)
             ) ;
    mux21_ni ix15031 (.Y (nx15030), .A0 (inputs_28__3), .A1 (inputs_29__3), .S0 (
             nx24095)) ;
    mux21_ni ix15043 (.Y (nx15042), .A0 (inputs_30__3), .A1 (inputs_31__3), .S0 (
             nx24095)) ;
    mux21_ni ix15347 (.Y (nx15346), .A0 (nx15340), .A1 (nx15262), .S0 (nx23133)
             ) ;
    oai21 ix15341 (.Y (nx15340), .A0 (nx22259), .A1 (nx11449), .B0 (nx11463)) ;
    mux21 ix11450 (.Y (nx11449), .A0 (nx15304), .A1 (nx15332), .S0 (nx22779)) ;
    mux21_ni ix15305 (.Y (nx15304), .A0 (nx15288), .A1 (nx15300), .S0 (nx23477)
             ) ;
    mux21_ni ix15289 (.Y (nx15288), .A0 (inputs_36__3), .A1 (inputs_37__3), .S0 (
             nx24095)) ;
    mux21_ni ix15301 (.Y (nx15300), .A0 (inputs_38__3), .A1 (inputs_39__3), .S0 (
             nx24095)) ;
    mux21_ni ix15333 (.Y (nx15332), .A0 (nx15316), .A1 (nx15328), .S0 (nx23477)
             ) ;
    mux21_ni ix15317 (.Y (nx15316), .A0 (inputs_52__3), .A1 (inputs_53__3), .S0 (
             nx24095)) ;
    mux21_ni ix15329 (.Y (nx15328), .A0 (inputs_54__3), .A1 (inputs_55__3), .S0 (
             nx24095)) ;
    nand04 ix11464 (.Y (nx11463), .A0 (nx22261), .A1 (nx23477), .A2 (nx24097), .A3 (
           nx15276)) ;
    mux21_ni ix15277 (.Y (nx15276), .A0 (inputs_35__3), .A1 (inputs_51__3), .S0 (
             nx22781)) ;
    mux21_ni ix15263 (.Y (nx15262), .A0 (nx15198), .A1 (nx15258), .S0 (nx22781)
             ) ;
    mux21_ni ix15199 (.Y (nx15198), .A0 (nx15166), .A1 (nx15194), .S0 (nx23223)
             ) ;
    mux21_ni ix15167 (.Y (nx15166), .A0 (nx15150), .A1 (nx15162), .S0 (nx23477)
             ) ;
    mux21_ni ix15151 (.Y (nx15150), .A0 (inputs_40__3), .A1 (inputs_41__3), .S0 (
             nx24097)) ;
    mux21_ni ix15163 (.Y (nx15162), .A0 (inputs_42__3), .A1 (inputs_43__3), .S0 (
             nx24097)) ;
    mux21_ni ix15195 (.Y (nx15194), .A0 (nx15178), .A1 (nx15190), .S0 (nx23477)
             ) ;
    mux21_ni ix15179 (.Y (nx15178), .A0 (inputs_44__3), .A1 (inputs_45__3), .S0 (
             nx24097)) ;
    mux21_ni ix15191 (.Y (nx15190), .A0 (inputs_46__3), .A1 (inputs_47__3), .S0 (
             nx24097)) ;
    mux21_ni ix15259 (.Y (nx15258), .A0 (nx15226), .A1 (nx15254), .S0 (nx23223)
             ) ;
    mux21_ni ix15227 (.Y (nx15226), .A0 (nx15210), .A1 (nx15222), .S0 (nx23477)
             ) ;
    mux21_ni ix15211 (.Y (nx15210), .A0 (inputs_56__3), .A1 (inputs_57__3), .S0 (
             nx24097)) ;
    mux21_ni ix15223 (.Y (nx15222), .A0 (inputs_58__3), .A1 (inputs_59__3), .S0 (
             nx24097)) ;
    mux21_ni ix15255 (.Y (nx15254), .A0 (nx15238), .A1 (nx15250), .S0 (nx23479)
             ) ;
    mux21_ni ix15239 (.Y (nx15238), .A0 (inputs_60__3), .A1 (inputs_61__3), .S0 (
             nx24099)) ;
    mux21_ni ix15251 (.Y (nx15250), .A0 (inputs_62__3), .A1 (inputs_63__3), .S0 (
             nx24099)) ;
    mux21_ni ix15771 (.Y (nx15770), .A0 (nx15558), .A1 (nx15766), .S0 (nx22561)
             ) ;
    mux21_ni ix15559 (.Y (nx15558), .A0 (nx15552), .A1 (nx15474), .S0 (nx23133)
             ) ;
    oai21 ix15553 (.Y (nx15552), .A0 (nx22261), .A1 (nx11495), .B0 (nx11507)) ;
    mux21 ix11496 (.Y (nx11495), .A0 (nx15516), .A1 (nx15544), .S0 (nx22781)) ;
    mux21_ni ix15517 (.Y (nx15516), .A0 (nx15500), .A1 (nx15512), .S0 (nx23479)
             ) ;
    mux21_ni ix15501 (.Y (nx15500), .A0 (inputs_68__3), .A1 (inputs_69__3), .S0 (
             nx24099)) ;
    mux21_ni ix15513 (.Y (nx15512), .A0 (inputs_70__3), .A1 (inputs_71__3), .S0 (
             nx24099)) ;
    mux21_ni ix15545 (.Y (nx15544), .A0 (nx15528), .A1 (nx15540), .S0 (nx23479)
             ) ;
    mux21_ni ix15529 (.Y (nx15528), .A0 (inputs_84__3), .A1 (inputs_85__3), .S0 (
             nx24099)) ;
    mux21_ni ix15541 (.Y (nx15540), .A0 (inputs_86__3), .A1 (inputs_87__3), .S0 (
             nx24099)) ;
    nand04 ix11508 (.Y (nx11507), .A0 (nx22261), .A1 (nx23479), .A2 (nx24099), .A3 (
           nx15488)) ;
    mux21_ni ix15489 (.Y (nx15488), .A0 (inputs_67__3), .A1 (inputs_83__3), .S0 (
             nx22781)) ;
    mux21_ni ix15475 (.Y (nx15474), .A0 (nx15410), .A1 (nx15470), .S0 (nx22781)
             ) ;
    mux21_ni ix15411 (.Y (nx15410), .A0 (nx15378), .A1 (nx15406), .S0 (nx23223)
             ) ;
    mux21_ni ix15379 (.Y (nx15378), .A0 (nx15362), .A1 (nx15374), .S0 (nx23479)
             ) ;
    mux21_ni ix15363 (.Y (nx15362), .A0 (inputs_72__3), .A1 (inputs_73__3), .S0 (
             nx24101)) ;
    mux21_ni ix15375 (.Y (nx15374), .A0 (inputs_74__3), .A1 (inputs_75__3), .S0 (
             nx24101)) ;
    mux21_ni ix15407 (.Y (nx15406), .A0 (nx15390), .A1 (nx15402), .S0 (nx23479)
             ) ;
    mux21_ni ix15391 (.Y (nx15390), .A0 (inputs_76__3), .A1 (inputs_77__3), .S0 (
             nx24101)) ;
    mux21_ni ix15403 (.Y (nx15402), .A0 (inputs_78__3), .A1 (inputs_79__3), .S0 (
             nx24101)) ;
    mux21_ni ix15471 (.Y (nx15470), .A0 (nx15438), .A1 (nx15466), .S0 (nx23223)
             ) ;
    mux21_ni ix15439 (.Y (nx15438), .A0 (nx15422), .A1 (nx15434), .S0 (nx23479)
             ) ;
    mux21_ni ix15423 (.Y (nx15422), .A0 (inputs_88__3), .A1 (inputs_89__3), .S0 (
             nx24101)) ;
    mux21_ni ix15435 (.Y (nx15434), .A0 (inputs_90__3), .A1 (inputs_91__3), .S0 (
             nx24101)) ;
    mux21_ni ix15467 (.Y (nx15466), .A0 (nx15450), .A1 (nx15462), .S0 (nx23481)
             ) ;
    mux21_ni ix15451 (.Y (nx15450), .A0 (inputs_92__3), .A1 (inputs_93__3), .S0 (
             nx24101)) ;
    mux21_ni ix15463 (.Y (nx15462), .A0 (inputs_94__3), .A1 (inputs_95__3), .S0 (
             nx24103)) ;
    mux21_ni ix15767 (.Y (nx15766), .A0 (nx15760), .A1 (nx15682), .S0 (nx23133)
             ) ;
    oai21 ix15761 (.Y (nx15760), .A0 (nx22261), .A1 (nx11541), .B0 (nx11553)) ;
    mux21 ix11542 (.Y (nx11541), .A0 (nx15724), .A1 (nx15752), .S0 (nx22781)) ;
    mux21_ni ix15725 (.Y (nx15724), .A0 (nx15708), .A1 (nx15720), .S0 (nx23481)
             ) ;
    mux21_ni ix15709 (.Y (nx15708), .A0 (inputs_100__3), .A1 (inputs_101__3), .S0 (
             nx24103)) ;
    mux21_ni ix15721 (.Y (nx15720), .A0 (inputs_102__3), .A1 (inputs_103__3), .S0 (
             nx24103)) ;
    mux21_ni ix15753 (.Y (nx15752), .A0 (nx15736), .A1 (nx15748), .S0 (nx23481)
             ) ;
    mux21_ni ix15737 (.Y (nx15736), .A0 (inputs_116__3), .A1 (inputs_117__3), .S0 (
             nx24103)) ;
    mux21_ni ix15749 (.Y (nx15748), .A0 (inputs_118__3), .A1 (inputs_119__3), .S0 (
             nx24103)) ;
    nand04 ix11554 (.Y (nx11553), .A0 (nx22261), .A1 (nx23481), .A2 (nx24103), .A3 (
           nx15696)) ;
    mux21_ni ix15697 (.Y (nx15696), .A0 (inputs_99__3), .A1 (inputs_115__3), .S0 (
             nx22781)) ;
    mux21_ni ix15683 (.Y (nx15682), .A0 (nx15618), .A1 (nx15678), .S0 (nx22783)
             ) ;
    mux21_ni ix15619 (.Y (nx15618), .A0 (nx15586), .A1 (nx15614), .S0 (nx23223)
             ) ;
    mux21_ni ix15587 (.Y (nx15586), .A0 (nx15570), .A1 (nx15582), .S0 (nx23481)
             ) ;
    mux21_ni ix15571 (.Y (nx15570), .A0 (inputs_104__3), .A1 (inputs_105__3), .S0 (
             nx24103)) ;
    mux21_ni ix15583 (.Y (nx15582), .A0 (inputs_106__3), .A1 (inputs_107__3), .S0 (
             nx24105)) ;
    mux21_ni ix15615 (.Y (nx15614), .A0 (nx15598), .A1 (nx15610), .S0 (nx23481)
             ) ;
    mux21_ni ix15599 (.Y (nx15598), .A0 (inputs_108__3), .A1 (inputs_109__3), .S0 (
             nx24105)) ;
    mux21_ni ix15611 (.Y (nx15610), .A0 (inputs_110__3), .A1 (inputs_111__3), .S0 (
             nx24105)) ;
    mux21_ni ix15679 (.Y (nx15678), .A0 (nx15646), .A1 (nx15674), .S0 (nx23225)
             ) ;
    mux21_ni ix15647 (.Y (nx15646), .A0 (nx15630), .A1 (nx15642), .S0 (nx23481)
             ) ;
    mux21_ni ix15631 (.Y (nx15630), .A0 (inputs_120__3), .A1 (inputs_121__3), .S0 (
             nx24105)) ;
    mux21_ni ix15643 (.Y (nx15642), .A0 (inputs_122__3), .A1 (inputs_123__3), .S0 (
             nx24105)) ;
    mux21_ni ix15675 (.Y (nx15674), .A0 (nx15658), .A1 (nx15670), .S0 (nx23483)
             ) ;
    mux21_ni ix15659 (.Y (nx15658), .A0 (inputs_124__3), .A1 (inputs_125__3), .S0 (
             nx24105)) ;
    mux21_ni ix15671 (.Y (nx15670), .A0 (inputs_126__3), .A1 (inputs_127__3), .S0 (
             nx24105)) ;
    mux21_ni ix16619 (.Y (nx16618), .A0 (nx16194), .A1 (nx16614), .S0 (nx22469)
             ) ;
    mux21_ni ix16195 (.Y (nx16194), .A0 (nx15982), .A1 (nx16190), .S0 (nx22563)
             ) ;
    mux21_ni ix15983 (.Y (nx15982), .A0 (nx15976), .A1 (nx15898), .S0 (nx23133)
             ) ;
    oai21 ix15977 (.Y (nx15976), .A0 (nx22261), .A1 (nx11587), .B0 (nx11601)) ;
    mux21 ix11588 (.Y (nx11587), .A0 (nx15940), .A1 (nx15968), .S0 (nx22783)) ;
    mux21_ni ix15941 (.Y (nx15940), .A0 (nx15924), .A1 (nx15936), .S0 (nx23483)
             ) ;
    mux21_ni ix15925 (.Y (nx15924), .A0 (inputs_132__3), .A1 (inputs_133__3), .S0 (
             nx24107)) ;
    mux21_ni ix15937 (.Y (nx15936), .A0 (inputs_134__3), .A1 (inputs_135__3), .S0 (
             nx24107)) ;
    mux21_ni ix15969 (.Y (nx15968), .A0 (nx15952), .A1 (nx15964), .S0 (nx23483)
             ) ;
    mux21_ni ix15953 (.Y (nx15952), .A0 (inputs_148__3), .A1 (inputs_149__3), .S0 (
             nx24107)) ;
    mux21_ni ix15965 (.Y (nx15964), .A0 (inputs_150__3), .A1 (inputs_151__3), .S0 (
             nx24107)) ;
    nand04 ix11602 (.Y (nx11601), .A0 (nx22261), .A1 (nx23483), .A2 (nx24107), .A3 (
           nx15912)) ;
    mux21_ni ix15913 (.Y (nx15912), .A0 (inputs_131__3), .A1 (inputs_147__3), .S0 (
             nx22783)) ;
    mux21_ni ix15899 (.Y (nx15898), .A0 (nx15834), .A1 (nx15894), .S0 (nx22783)
             ) ;
    mux21_ni ix15835 (.Y (nx15834), .A0 (nx15802), .A1 (nx15830), .S0 (nx23225)
             ) ;
    mux21_ni ix15803 (.Y (nx15802), .A0 (nx15786), .A1 (nx15798), .S0 (nx23483)
             ) ;
    mux21_ni ix15787 (.Y (nx15786), .A0 (inputs_136__3), .A1 (inputs_137__3), .S0 (
             nx24107)) ;
    mux21_ni ix15799 (.Y (nx15798), .A0 (inputs_138__3), .A1 (inputs_139__3), .S0 (
             nx24107)) ;
    mux21_ni ix15831 (.Y (nx15830), .A0 (nx15814), .A1 (nx15826), .S0 (nx23483)
             ) ;
    mux21_ni ix15815 (.Y (nx15814), .A0 (inputs_140__3), .A1 (inputs_141__3), .S0 (
             nx24109)) ;
    mux21_ni ix15827 (.Y (nx15826), .A0 (inputs_142__3), .A1 (inputs_143__3), .S0 (
             nx24109)) ;
    mux21_ni ix15895 (.Y (nx15894), .A0 (nx15862), .A1 (nx15890), .S0 (nx23225)
             ) ;
    mux21_ni ix15863 (.Y (nx15862), .A0 (nx15846), .A1 (nx15858), .S0 (nx23483)
             ) ;
    mux21_ni ix15847 (.Y (nx15846), .A0 (inputs_152__3), .A1 (inputs_153__3), .S0 (
             nx24109)) ;
    mux21_ni ix15859 (.Y (nx15858), .A0 (inputs_154__3), .A1 (inputs_155__3), .S0 (
             nx24109)) ;
    mux21_ni ix15891 (.Y (nx15890), .A0 (nx15874), .A1 (nx15886), .S0 (nx23485)
             ) ;
    mux21_ni ix15875 (.Y (nx15874), .A0 (inputs_156__3), .A1 (inputs_157__3), .S0 (
             nx24109)) ;
    mux21_ni ix15887 (.Y (nx15886), .A0 (inputs_158__3), .A1 (inputs_159__3), .S0 (
             nx24109)) ;
    mux21_ni ix16191 (.Y (nx16190), .A0 (nx16184), .A1 (nx16106), .S0 (nx23133)
             ) ;
    oai21 ix16185 (.Y (nx16184), .A0 (nx22263), .A1 (nx11633), .B0 (nx11645)) ;
    mux21 ix11634 (.Y (nx11633), .A0 (nx16148), .A1 (nx16176), .S0 (nx22783)) ;
    mux21_ni ix16149 (.Y (nx16148), .A0 (nx16132), .A1 (nx16144), .S0 (nx23485)
             ) ;
    mux21_ni ix16133 (.Y (nx16132), .A0 (inputs_164__3), .A1 (inputs_165__3), .S0 (
             nx24109)) ;
    mux21_ni ix16145 (.Y (nx16144), .A0 (inputs_166__3), .A1 (inputs_167__3), .S0 (
             nx24111)) ;
    mux21_ni ix16177 (.Y (nx16176), .A0 (nx16160), .A1 (nx16172), .S0 (nx23485)
             ) ;
    mux21_ni ix16161 (.Y (nx16160), .A0 (inputs_180__3), .A1 (inputs_181__3), .S0 (
             nx24111)) ;
    mux21_ni ix16173 (.Y (nx16172), .A0 (inputs_182__3), .A1 (inputs_183__3), .S0 (
             nx24111)) ;
    nand04 ix11646 (.Y (nx11645), .A0 (nx22263), .A1 (nx23485), .A2 (nx24111), .A3 (
           nx16120)) ;
    mux21_ni ix16121 (.Y (nx16120), .A0 (inputs_163__3), .A1 (inputs_179__3), .S0 (
             nx22783)) ;
    mux21_ni ix16107 (.Y (nx16106), .A0 (nx16042), .A1 (nx16102), .S0 (nx22783)
             ) ;
    mux21_ni ix16043 (.Y (nx16042), .A0 (nx16010), .A1 (nx16038), .S0 (nx23225)
             ) ;
    mux21_ni ix16011 (.Y (nx16010), .A0 (nx15994), .A1 (nx16006), .S0 (nx23485)
             ) ;
    mux21_ni ix15995 (.Y (nx15994), .A0 (inputs_168__3), .A1 (inputs_169__3), .S0 (
             nx24111)) ;
    mux21_ni ix16007 (.Y (nx16006), .A0 (inputs_170__3), .A1 (inputs_171__3), .S0 (
             nx24111)) ;
    mux21_ni ix16039 (.Y (nx16038), .A0 (nx16022), .A1 (nx16034), .S0 (nx23485)
             ) ;
    mux21_ni ix16023 (.Y (nx16022), .A0 (inputs_172__3), .A1 (inputs_173__3), .S0 (
             nx24111)) ;
    mux21_ni ix16035 (.Y (nx16034), .A0 (inputs_174__3), .A1 (inputs_175__3), .S0 (
             nx24113)) ;
    mux21_ni ix16103 (.Y (nx16102), .A0 (nx16070), .A1 (nx16098), .S0 (nx23225)
             ) ;
    mux21_ni ix16071 (.Y (nx16070), .A0 (nx16054), .A1 (nx16066), .S0 (nx23485)
             ) ;
    mux21_ni ix16055 (.Y (nx16054), .A0 (inputs_184__3), .A1 (inputs_185__3), .S0 (
             nx24113)) ;
    mux21_ni ix16067 (.Y (nx16066), .A0 (inputs_186__3), .A1 (inputs_187__3), .S0 (
             nx24113)) ;
    mux21_ni ix16099 (.Y (nx16098), .A0 (nx16082), .A1 (nx16094), .S0 (nx23487)
             ) ;
    mux21_ni ix16083 (.Y (nx16082), .A0 (inputs_188__3), .A1 (inputs_189__3), .S0 (
             nx24113)) ;
    mux21_ni ix16095 (.Y (nx16094), .A0 (inputs_190__3), .A1 (inputs_191__3), .S0 (
             nx24113)) ;
    mux21_ni ix16615 (.Y (nx16614), .A0 (nx16402), .A1 (nx16610), .S0 (nx22563)
             ) ;
    mux21_ni ix16403 (.Y (nx16402), .A0 (nx16396), .A1 (nx16318), .S0 (nx23133)
             ) ;
    oai21 ix16397 (.Y (nx16396), .A0 (nx22263), .A1 (nx11677), .B0 (nx11687)) ;
    mux21 ix11678 (.Y (nx11677), .A0 (nx16360), .A1 (nx16388), .S0 (nx22785)) ;
    mux21_ni ix16361 (.Y (nx16360), .A0 (nx16344), .A1 (nx16356), .S0 (nx23487)
             ) ;
    mux21_ni ix16345 (.Y (nx16344), .A0 (inputs_196__3), .A1 (inputs_197__3), .S0 (
             nx24113)) ;
    mux21_ni ix16357 (.Y (nx16356), .A0 (inputs_198__3), .A1 (inputs_199__3), .S0 (
             nx24113)) ;
    mux21_ni ix16389 (.Y (nx16388), .A0 (nx16372), .A1 (nx16384), .S0 (nx23487)
             ) ;
    mux21_ni ix16373 (.Y (nx16372), .A0 (inputs_212__3), .A1 (inputs_213__3), .S0 (
             nx24115)) ;
    mux21_ni ix16385 (.Y (nx16384), .A0 (inputs_214__3), .A1 (inputs_215__3), .S0 (
             nx24115)) ;
    nand04 ix11688 (.Y (nx11687), .A0 (nx22263), .A1 (nx23487), .A2 (nx24115), .A3 (
           nx16332)) ;
    mux21_ni ix16333 (.Y (nx16332), .A0 (inputs_195__3), .A1 (inputs_211__3), .S0 (
             nx22785)) ;
    mux21_ni ix16319 (.Y (nx16318), .A0 (nx16254), .A1 (nx16314), .S0 (nx22785)
             ) ;
    mux21_ni ix16255 (.Y (nx16254), .A0 (nx16222), .A1 (nx16250), .S0 (nx23225)
             ) ;
    mux21_ni ix16223 (.Y (nx16222), .A0 (nx16206), .A1 (nx16218), .S0 (nx23487)
             ) ;
    mux21_ni ix16207 (.Y (nx16206), .A0 (inputs_200__3), .A1 (inputs_201__3), .S0 (
             nx24115)) ;
    mux21_ni ix16219 (.Y (nx16218), .A0 (inputs_202__3), .A1 (inputs_203__3), .S0 (
             nx24115)) ;
    mux21_ni ix16251 (.Y (nx16250), .A0 (nx16234), .A1 (nx16246), .S0 (nx23487)
             ) ;
    mux21_ni ix16235 (.Y (nx16234), .A0 (inputs_204__3), .A1 (inputs_205__3), .S0 (
             nx24115)) ;
    mux21_ni ix16247 (.Y (nx16246), .A0 (inputs_206__3), .A1 (inputs_207__3), .S0 (
             nx24115)) ;
    mux21_ni ix16315 (.Y (nx16314), .A0 (nx16282), .A1 (nx16310), .S0 (nx23225)
             ) ;
    mux21_ni ix16283 (.Y (nx16282), .A0 (nx16266), .A1 (nx16278), .S0 (nx23487)
             ) ;
    mux21_ni ix16267 (.Y (nx16266), .A0 (inputs_216__3), .A1 (inputs_217__3), .S0 (
             nx24117)) ;
    mux21_ni ix16279 (.Y (nx16278), .A0 (inputs_218__3), .A1 (inputs_219__3), .S0 (
             nx24117)) ;
    mux21_ni ix16311 (.Y (nx16310), .A0 (nx16294), .A1 (nx16306), .S0 (nx23489)
             ) ;
    mux21_ni ix16295 (.Y (nx16294), .A0 (inputs_220__3), .A1 (inputs_221__3), .S0 (
             nx24117)) ;
    mux21_ni ix16307 (.Y (nx16306), .A0 (inputs_222__3), .A1 (inputs_223__3), .S0 (
             nx24117)) ;
    mux21_ni ix16611 (.Y (nx16610), .A0 (nx16604), .A1 (nx16526), .S0 (nx23135)
             ) ;
    oai21 ix16605 (.Y (nx16604), .A0 (nx22263), .A1 (nx11717), .B0 (nx11727)) ;
    mux21 ix11718 (.Y (nx11717), .A0 (nx16568), .A1 (nx16596), .S0 (nx22785)) ;
    mux21_ni ix16569 (.Y (nx16568), .A0 (nx16552), .A1 (nx16564), .S0 (nx23489)
             ) ;
    mux21_ni ix16553 (.Y (nx16552), .A0 (inputs_228__3), .A1 (inputs_229__3), .S0 (
             nx24117)) ;
    mux21_ni ix16565 (.Y (nx16564), .A0 (inputs_230__3), .A1 (inputs_231__3), .S0 (
             nx24117)) ;
    mux21_ni ix16597 (.Y (nx16596), .A0 (nx16580), .A1 (nx16592), .S0 (nx23489)
             ) ;
    mux21_ni ix16581 (.Y (nx16580), .A0 (inputs_244__3), .A1 (inputs_245__3), .S0 (
             nx24117)) ;
    mux21_ni ix16593 (.Y (nx16592), .A0 (inputs_246__3), .A1 (inputs_247__3), .S0 (
             nx24119)) ;
    nand04 ix11728 (.Y (nx11727), .A0 (nx22263), .A1 (nx23489), .A2 (nx24119), .A3 (
           nx16540)) ;
    mux21_ni ix16541 (.Y (nx16540), .A0 (inputs_227__3), .A1 (inputs_243__3), .S0 (
             nx22785)) ;
    mux21_ni ix16527 (.Y (nx16526), .A0 (nx16462), .A1 (nx16522), .S0 (nx22785)
             ) ;
    mux21_ni ix16463 (.Y (nx16462), .A0 (nx16430), .A1 (nx16458), .S0 (nx23227)
             ) ;
    mux21_ni ix16431 (.Y (nx16430), .A0 (nx16414), .A1 (nx16426), .S0 (nx23489)
             ) ;
    mux21_ni ix16415 (.Y (nx16414), .A0 (inputs_232__3), .A1 (inputs_233__3), .S0 (
             nx24119)) ;
    mux21_ni ix16427 (.Y (nx16426), .A0 (inputs_234__3), .A1 (inputs_235__3), .S0 (
             nx24119)) ;
    mux21_ni ix16459 (.Y (nx16458), .A0 (nx16442), .A1 (nx16454), .S0 (nx23489)
             ) ;
    mux21_ni ix16443 (.Y (nx16442), .A0 (inputs_236__3), .A1 (inputs_237__3), .S0 (
             nx24119)) ;
    mux21_ni ix16455 (.Y (nx16454), .A0 (inputs_238__3), .A1 (inputs_239__3), .S0 (
             nx24119)) ;
    mux21_ni ix16523 (.Y (nx16522), .A0 (nx16490), .A1 (nx16518), .S0 (nx23227)
             ) ;
    mux21_ni ix16491 (.Y (nx16490), .A0 (nx16474), .A1 (nx16486), .S0 (nx23489)
             ) ;
    mux21_ni ix16475 (.Y (nx16474), .A0 (inputs_248__3), .A1 (inputs_249__3), .S0 (
             nx24119)) ;
    mux21_ni ix16487 (.Y (nx16486), .A0 (inputs_250__3), .A1 (inputs_251__3), .S0 (
             nx24121)) ;
    mux21_ni ix16519 (.Y (nx16518), .A0 (nx16502), .A1 (nx16514), .S0 (nx23491)
             ) ;
    mux21_ni ix16503 (.Y (nx16502), .A0 (inputs_252__3), .A1 (inputs_253__3), .S0 (
             nx24121)) ;
    mux21_ni ix16515 (.Y (nx16514), .A0 (inputs_254__3), .A1 (inputs_255__3), .S0 (
             nx24121)) ;
    oai21 ix20789 (.Y (\output [4]), .A0 (nx22219), .A1 (nx11759), .B0 (nx12113)
          ) ;
    mux21 ix11760 (.Y (nx11759), .A0 (nx17470), .A1 (nx18314), .S0 (nx22419)) ;
    mux21_ni ix17471 (.Y (nx17470), .A0 (nx17046), .A1 (nx17466), .S0 (nx22469)
             ) ;
    mux21_ni ix17047 (.Y (nx17046), .A0 (nx16834), .A1 (nx17042), .S0 (nx22563)
             ) ;
    mux21_ni ix16835 (.Y (nx16834), .A0 (nx16828), .A1 (nx16750), .S0 (nx23135)
             ) ;
    oai21 ix16829 (.Y (nx16828), .A0 (nx22263), .A1 (nx11767), .B0 (nx11777)) ;
    mux21 ix11768 (.Y (nx11767), .A0 (nx16792), .A1 (nx16820), .S0 (nx22785)) ;
    mux21_ni ix16793 (.Y (nx16792), .A0 (nx16776), .A1 (nx16788), .S0 (nx23491)
             ) ;
    mux21_ni ix16777 (.Y (nx16776), .A0 (inputs_260__4), .A1 (inputs_261__4), .S0 (
             nx24121)) ;
    mux21_ni ix16789 (.Y (nx16788), .A0 (inputs_262__4), .A1 (inputs_263__4), .S0 (
             nx24121)) ;
    mux21_ni ix16821 (.Y (nx16820), .A0 (nx16804), .A1 (nx16816), .S0 (nx23491)
             ) ;
    mux21_ni ix16805 (.Y (nx16804), .A0 (inputs_276__4), .A1 (inputs_277__4), .S0 (
             nx24121)) ;
    mux21_ni ix16817 (.Y (nx16816), .A0 (inputs_278__4), .A1 (inputs_279__4), .S0 (
             nx24121)) ;
    nand04 ix11778 (.Y (nx11777), .A0 (nx22265), .A1 (nx23491), .A2 (nx24123), .A3 (
           nx16764)) ;
    mux21_ni ix16765 (.Y (nx16764), .A0 (inputs_259__4), .A1 (inputs_275__4), .S0 (
             nx22787)) ;
    mux21_ni ix16751 (.Y (nx16750), .A0 (nx16686), .A1 (nx16746), .S0 (nx22787)
             ) ;
    mux21_ni ix16687 (.Y (nx16686), .A0 (nx16654), .A1 (nx16682), .S0 (nx23227)
             ) ;
    mux21_ni ix16655 (.Y (nx16654), .A0 (nx16638), .A1 (nx16650), .S0 (nx23491)
             ) ;
    mux21_ni ix16639 (.Y (nx16638), .A0 (inputs_264__4), .A1 (inputs_265__4), .S0 (
             nx24123)) ;
    mux21_ni ix16651 (.Y (nx16650), .A0 (inputs_266__4), .A1 (inputs_267__4), .S0 (
             nx24123)) ;
    mux21_ni ix16683 (.Y (nx16682), .A0 (nx16666), .A1 (nx16678), .S0 (nx23491)
             ) ;
    mux21_ni ix16667 (.Y (nx16666), .A0 (inputs_268__4), .A1 (inputs_269__4), .S0 (
             nx24123)) ;
    mux21_ni ix16679 (.Y (nx16678), .A0 (inputs_270__4), .A1 (inputs_271__4), .S0 (
             nx24123)) ;
    mux21_ni ix16747 (.Y (nx16746), .A0 (nx16714), .A1 (nx16742), .S0 (nx23227)
             ) ;
    mux21_ni ix16715 (.Y (nx16714), .A0 (nx16698), .A1 (nx16710), .S0 (nx23491)
             ) ;
    mux21_ni ix16699 (.Y (nx16698), .A0 (inputs_280__4), .A1 (inputs_281__4), .S0 (
             nx24123)) ;
    mux21_ni ix16711 (.Y (nx16710), .A0 (inputs_282__4), .A1 (inputs_283__4), .S0 (
             nx24123)) ;
    mux21_ni ix16743 (.Y (nx16742), .A0 (nx16726), .A1 (nx16738), .S0 (nx23493)
             ) ;
    mux21_ni ix16727 (.Y (nx16726), .A0 (inputs_284__4), .A1 (inputs_285__4), .S0 (
             nx24125)) ;
    mux21_ni ix16739 (.Y (nx16738), .A0 (inputs_286__4), .A1 (inputs_287__4), .S0 (
             nx24125)) ;
    mux21_ni ix17043 (.Y (nx17042), .A0 (nx17036), .A1 (nx16958), .S0 (nx23135)
             ) ;
    oai21 ix17037 (.Y (nx17036), .A0 (nx22265), .A1 (nx11807), .B0 (nx11821)) ;
    mux21 ix11808 (.Y (nx11807), .A0 (nx17000), .A1 (nx17028), .S0 (nx22787)) ;
    mux21_ni ix17001 (.Y (nx17000), .A0 (nx16984), .A1 (nx16996), .S0 (nx23493)
             ) ;
    mux21_ni ix16985 (.Y (nx16984), .A0 (inputs_292__4), .A1 (inputs_293__4), .S0 (
             nx24125)) ;
    mux21_ni ix16997 (.Y (nx16996), .A0 (inputs_294__4), .A1 (inputs_295__4), .S0 (
             nx24125)) ;
    mux21_ni ix17029 (.Y (nx17028), .A0 (nx17012), .A1 (nx17024), .S0 (nx23493)
             ) ;
    mux21_ni ix17013 (.Y (nx17012), .A0 (inputs_308__4), .A1 (inputs_309__4), .S0 (
             nx24125)) ;
    mux21_ni ix17025 (.Y (nx17024), .A0 (inputs_310__4), .A1 (inputs_311__4), .S0 (
             nx24125)) ;
    nand04 ix11822 (.Y (nx11821), .A0 (nx22265), .A1 (nx23493), .A2 (nx24125), .A3 (
           nx16972)) ;
    mux21_ni ix16973 (.Y (nx16972), .A0 (inputs_291__4), .A1 (inputs_307__4), .S0 (
             nx22787)) ;
    mux21_ni ix16959 (.Y (nx16958), .A0 (nx16894), .A1 (nx16954), .S0 (nx22787)
             ) ;
    mux21_ni ix16895 (.Y (nx16894), .A0 (nx16862), .A1 (nx16890), .S0 (nx23227)
             ) ;
    mux21_ni ix16863 (.Y (nx16862), .A0 (nx16846), .A1 (nx16858), .S0 (nx23493)
             ) ;
    mux21_ni ix16847 (.Y (nx16846), .A0 (inputs_296__4), .A1 (inputs_297__4), .S0 (
             nx24127)) ;
    mux21_ni ix16859 (.Y (nx16858), .A0 (inputs_298__4), .A1 (inputs_299__4), .S0 (
             nx24127)) ;
    mux21_ni ix16891 (.Y (nx16890), .A0 (nx16874), .A1 (nx16886), .S0 (nx23493)
             ) ;
    mux21_ni ix16875 (.Y (nx16874), .A0 (inputs_300__4), .A1 (inputs_301__4), .S0 (
             nx24127)) ;
    mux21_ni ix16887 (.Y (nx16886), .A0 (inputs_302__4), .A1 (inputs_303__4), .S0 (
             nx24127)) ;
    mux21_ni ix16955 (.Y (nx16954), .A0 (nx16922), .A1 (nx16950), .S0 (nx23227)
             ) ;
    mux21_ni ix16923 (.Y (nx16922), .A0 (nx16906), .A1 (nx16918), .S0 (nx23493)
             ) ;
    mux21_ni ix16907 (.Y (nx16906), .A0 (inputs_312__4), .A1 (inputs_313__4), .S0 (
             nx24127)) ;
    mux21_ni ix16919 (.Y (nx16918), .A0 (inputs_314__4), .A1 (inputs_315__4), .S0 (
             nx24127)) ;
    mux21_ni ix16951 (.Y (nx16950), .A0 (nx16934), .A1 (nx16946), .S0 (nx23495)
             ) ;
    mux21_ni ix16935 (.Y (nx16934), .A0 (inputs_316__4), .A1 (inputs_317__4), .S0 (
             nx24127)) ;
    mux21_ni ix16947 (.Y (nx16946), .A0 (inputs_318__4), .A1 (inputs_319__4), .S0 (
             nx24129)) ;
    mux21_ni ix17467 (.Y (nx17466), .A0 (nx17254), .A1 (nx17462), .S0 (nx22563)
             ) ;
    mux21_ni ix17255 (.Y (nx17254), .A0 (nx17248), .A1 (nx17170), .S0 (nx23135)
             ) ;
    oai21 ix17249 (.Y (nx17248), .A0 (nx22265), .A1 (nx11853), .B0 (nx11863)) ;
    mux21 ix11854 (.Y (nx11853), .A0 (nx17212), .A1 (nx17240), .S0 (nx22787)) ;
    mux21_ni ix17213 (.Y (nx17212), .A0 (nx17196), .A1 (nx17208), .S0 (nx23495)
             ) ;
    mux21_ni ix17197 (.Y (nx17196), .A0 (inputs_324__4), .A1 (inputs_325__4), .S0 (
             nx24129)) ;
    mux21_ni ix17209 (.Y (nx17208), .A0 (inputs_326__4), .A1 (inputs_327__4), .S0 (
             nx24129)) ;
    mux21_ni ix17241 (.Y (nx17240), .A0 (nx17224), .A1 (nx17236), .S0 (nx23495)
             ) ;
    mux21_ni ix17225 (.Y (nx17224), .A0 (inputs_340__4), .A1 (inputs_341__4), .S0 (
             nx24129)) ;
    mux21_ni ix17237 (.Y (nx17236), .A0 (inputs_342__4), .A1 (inputs_343__4), .S0 (
             nx24129)) ;
    nand04 ix11864 (.Y (nx11863), .A0 (nx22265), .A1 (nx23495), .A2 (nx24129), .A3 (
           nx17184)) ;
    mux21_ni ix17185 (.Y (nx17184), .A0 (inputs_323__4), .A1 (inputs_339__4), .S0 (
             nx22787)) ;
    mux21_ni ix17171 (.Y (nx17170), .A0 (nx17106), .A1 (nx17166), .S0 (nx22789)
             ) ;
    mux21_ni ix17107 (.Y (nx17106), .A0 (nx17074), .A1 (nx17102), .S0 (nx23227)
             ) ;
    mux21_ni ix17075 (.Y (nx17074), .A0 (nx17058), .A1 (nx17070), .S0 (nx23495)
             ) ;
    mux21_ni ix17059 (.Y (nx17058), .A0 (inputs_328__4), .A1 (inputs_329__4), .S0 (
             nx24129)) ;
    mux21_ni ix17071 (.Y (nx17070), .A0 (inputs_330__4), .A1 (inputs_331__4), .S0 (
             nx24131)) ;
    mux21_ni ix17103 (.Y (nx17102), .A0 (nx17086), .A1 (nx17098), .S0 (nx23495)
             ) ;
    mux21_ni ix17087 (.Y (nx17086), .A0 (inputs_332__4), .A1 (inputs_333__4), .S0 (
             nx24131)) ;
    mux21_ni ix17099 (.Y (nx17098), .A0 (inputs_334__4), .A1 (inputs_335__4), .S0 (
             nx24131)) ;
    mux21_ni ix17167 (.Y (nx17166), .A0 (nx17134), .A1 (nx17162), .S0 (nx23229)
             ) ;
    mux21_ni ix17135 (.Y (nx17134), .A0 (nx17118), .A1 (nx17130), .S0 (nx23495)
             ) ;
    mux21_ni ix17119 (.Y (nx17118), .A0 (inputs_344__4), .A1 (inputs_345__4), .S0 (
             nx24131)) ;
    mux21_ni ix17131 (.Y (nx17130), .A0 (inputs_346__4), .A1 (inputs_347__4), .S0 (
             nx24131)) ;
    mux21_ni ix17163 (.Y (nx17162), .A0 (nx17146), .A1 (nx17158), .S0 (nx23497)
             ) ;
    mux21_ni ix17147 (.Y (nx17146), .A0 (inputs_348__4), .A1 (inputs_349__4), .S0 (
             nx24131)) ;
    mux21_ni ix17159 (.Y (nx17158), .A0 (inputs_350__4), .A1 (inputs_351__4), .S0 (
             nx24131)) ;
    mux21_ni ix17463 (.Y (nx17462), .A0 (nx17456), .A1 (nx17378), .S0 (nx23135)
             ) ;
    oai21 ix17457 (.Y (nx17456), .A0 (nx22265), .A1 (nx11893), .B0 (nx11905)) ;
    mux21 ix11894 (.Y (nx11893), .A0 (nx17420), .A1 (nx17448), .S0 (nx22789)) ;
    mux21_ni ix17421 (.Y (nx17420), .A0 (nx17404), .A1 (nx17416), .S0 (nx23497)
             ) ;
    mux21_ni ix17405 (.Y (nx17404), .A0 (inputs_356__4), .A1 (inputs_357__4), .S0 (
             nx24133)) ;
    mux21_ni ix17417 (.Y (nx17416), .A0 (inputs_358__4), .A1 (inputs_359__4), .S0 (
             nx24133)) ;
    mux21_ni ix17449 (.Y (nx17448), .A0 (nx17432), .A1 (nx17444), .S0 (nx23497)
             ) ;
    mux21_ni ix17433 (.Y (nx17432), .A0 (inputs_372__4), .A1 (inputs_373__4), .S0 (
             nx24133)) ;
    mux21_ni ix17445 (.Y (nx17444), .A0 (inputs_374__4), .A1 (inputs_375__4), .S0 (
             nx24133)) ;
    nand04 ix11906 (.Y (nx11905), .A0 (nx22265), .A1 (nx23497), .A2 (nx24133), .A3 (
           nx17392)) ;
    mux21_ni ix17393 (.Y (nx17392), .A0 (inputs_355__4), .A1 (inputs_371__4), .S0 (
             nx22789)) ;
    mux21_ni ix17379 (.Y (nx17378), .A0 (nx17314), .A1 (nx17374), .S0 (nx22789)
             ) ;
    mux21_ni ix17315 (.Y (nx17314), .A0 (nx17282), .A1 (nx17310), .S0 (nx23229)
             ) ;
    mux21_ni ix17283 (.Y (nx17282), .A0 (nx17266), .A1 (nx17278), .S0 (nx23497)
             ) ;
    mux21_ni ix17267 (.Y (nx17266), .A0 (inputs_360__4), .A1 (inputs_361__4), .S0 (
             nx24133)) ;
    mux21_ni ix17279 (.Y (nx17278), .A0 (inputs_362__4), .A1 (inputs_363__4), .S0 (
             nx24133)) ;
    mux21_ni ix17311 (.Y (nx17310), .A0 (nx17294), .A1 (nx17306), .S0 (nx23497)
             ) ;
    mux21_ni ix17295 (.Y (nx17294), .A0 (inputs_364__4), .A1 (inputs_365__4), .S0 (
             nx24135)) ;
    mux21_ni ix17307 (.Y (nx17306), .A0 (inputs_366__4), .A1 (inputs_367__4), .S0 (
             nx24135)) ;
    mux21_ni ix17375 (.Y (nx17374), .A0 (nx17342), .A1 (nx17370), .S0 (nx23229)
             ) ;
    mux21_ni ix17343 (.Y (nx17342), .A0 (nx17326), .A1 (nx17338), .S0 (nx23497)
             ) ;
    mux21_ni ix17327 (.Y (nx17326), .A0 (inputs_376__4), .A1 (inputs_377__4), .S0 (
             nx24135)) ;
    mux21_ni ix17339 (.Y (nx17338), .A0 (inputs_378__4), .A1 (inputs_379__4), .S0 (
             nx24135)) ;
    mux21_ni ix17371 (.Y (nx17370), .A0 (nx17354), .A1 (nx17366), .S0 (nx23499)
             ) ;
    mux21_ni ix17355 (.Y (nx17354), .A0 (inputs_380__4), .A1 (inputs_381__4), .S0 (
             nx24135)) ;
    mux21_ni ix17367 (.Y (nx17366), .A0 (inputs_382__4), .A1 (inputs_383__4), .S0 (
             nx24135)) ;
    mux21_ni ix18315 (.Y (nx18314), .A0 (nx17890), .A1 (nx18310), .S0 (nx22469)
             ) ;
    mux21_ni ix17891 (.Y (nx17890), .A0 (nx17678), .A1 (nx17886), .S0 (nx22563)
             ) ;
    mux21_ni ix17679 (.Y (nx17678), .A0 (nx17672), .A1 (nx17594), .S0 (nx23135)
             ) ;
    oai21 ix17673 (.Y (nx17672), .A0 (nx22267), .A1 (nx11939), .B0 (nx11953)) ;
    mux21 ix11940 (.Y (nx11939), .A0 (nx17636), .A1 (nx17664), .S0 (nx22789)) ;
    mux21_ni ix17637 (.Y (nx17636), .A0 (nx17620), .A1 (nx17632), .S0 (nx23499)
             ) ;
    mux21_ni ix17621 (.Y (nx17620), .A0 (inputs_388__4), .A1 (inputs_389__4), .S0 (
             nx24135)) ;
    mux21_ni ix17633 (.Y (nx17632), .A0 (inputs_390__4), .A1 (inputs_391__4), .S0 (
             nx24137)) ;
    mux21_ni ix17665 (.Y (nx17664), .A0 (nx17648), .A1 (nx17660), .S0 (nx23499)
             ) ;
    mux21_ni ix17649 (.Y (nx17648), .A0 (inputs_404__4), .A1 (inputs_405__4), .S0 (
             nx24137)) ;
    mux21_ni ix17661 (.Y (nx17660), .A0 (inputs_406__4), .A1 (inputs_407__4), .S0 (
             nx24137)) ;
    nand04 ix11954 (.Y (nx11953), .A0 (nx22267), .A1 (nx23499), .A2 (nx24137), .A3 (
           nx17608)) ;
    mux21_ni ix17609 (.Y (nx17608), .A0 (inputs_387__4), .A1 (inputs_403__4), .S0 (
             nx22789)) ;
    mux21_ni ix17595 (.Y (nx17594), .A0 (nx17530), .A1 (nx17590), .S0 (nx22789)
             ) ;
    mux21_ni ix17531 (.Y (nx17530), .A0 (nx17498), .A1 (nx17526), .S0 (nx23229)
             ) ;
    mux21_ni ix17499 (.Y (nx17498), .A0 (nx17482), .A1 (nx17494), .S0 (nx23499)
             ) ;
    mux21_ni ix17483 (.Y (nx17482), .A0 (inputs_392__4), .A1 (inputs_393__4), .S0 (
             nx24137)) ;
    mux21_ni ix17495 (.Y (nx17494), .A0 (inputs_394__4), .A1 (inputs_395__4), .S0 (
             nx24137)) ;
    mux21_ni ix17527 (.Y (nx17526), .A0 (nx17510), .A1 (nx17522), .S0 (nx23499)
             ) ;
    mux21_ni ix17511 (.Y (nx17510), .A0 (inputs_396__4), .A1 (inputs_397__4), .S0 (
             nx24137)) ;
    mux21_ni ix17523 (.Y (nx17522), .A0 (inputs_398__4), .A1 (inputs_399__4), .S0 (
             nx24139)) ;
    mux21_ni ix17591 (.Y (nx17590), .A0 (nx17558), .A1 (nx17586), .S0 (nx23229)
             ) ;
    mux21_ni ix17559 (.Y (nx17558), .A0 (nx17542), .A1 (nx17554), .S0 (nx23499)
             ) ;
    mux21_ni ix17543 (.Y (nx17542), .A0 (inputs_408__4), .A1 (inputs_409__4), .S0 (
             nx24139)) ;
    mux21_ni ix17555 (.Y (nx17554), .A0 (inputs_410__4), .A1 (inputs_411__4), .S0 (
             nx24139)) ;
    mux21_ni ix17587 (.Y (nx17586), .A0 (nx17570), .A1 (nx17582), .S0 (nx23501)
             ) ;
    mux21_ni ix17571 (.Y (nx17570), .A0 (inputs_412__4), .A1 (inputs_413__4), .S0 (
             nx24139)) ;
    mux21_ni ix17583 (.Y (nx17582), .A0 (inputs_414__4), .A1 (inputs_415__4), .S0 (
             nx24139)) ;
    mux21_ni ix17887 (.Y (nx17886), .A0 (nx17880), .A1 (nx17802), .S0 (nx23135)
             ) ;
    oai21 ix17881 (.Y (nx17880), .A0 (nx22267), .A1 (nx11983), .B0 (nx11995)) ;
    mux21 ix11984 (.Y (nx11983), .A0 (nx17844), .A1 (nx17872), .S0 (nx22791)) ;
    mux21_ni ix17845 (.Y (nx17844), .A0 (nx17828), .A1 (nx17840), .S0 (nx23501)
             ) ;
    mux21_ni ix17829 (.Y (nx17828), .A0 (inputs_420__4), .A1 (inputs_421__4), .S0 (
             nx24139)) ;
    mux21_ni ix17841 (.Y (nx17840), .A0 (inputs_422__4), .A1 (inputs_423__4), .S0 (
             nx24139)) ;
    mux21_ni ix17873 (.Y (nx17872), .A0 (nx17856), .A1 (nx17868), .S0 (nx23501)
             ) ;
    mux21_ni ix17857 (.Y (nx17856), .A0 (inputs_436__4), .A1 (inputs_437__4), .S0 (
             nx24141)) ;
    mux21_ni ix17869 (.Y (nx17868), .A0 (inputs_438__4), .A1 (inputs_439__4), .S0 (
             nx24141)) ;
    nand04 ix11996 (.Y (nx11995), .A0 (nx22267), .A1 (nx23501), .A2 (nx24141), .A3 (
           nx17816)) ;
    mux21_ni ix17817 (.Y (nx17816), .A0 (inputs_419__4), .A1 (inputs_435__4), .S0 (
             nx22791)) ;
    mux21_ni ix17803 (.Y (nx17802), .A0 (nx17738), .A1 (nx17798), .S0 (nx22791)
             ) ;
    mux21_ni ix17739 (.Y (nx17738), .A0 (nx17706), .A1 (nx17734), .S0 (nx23229)
             ) ;
    mux21_ni ix17707 (.Y (nx17706), .A0 (nx17690), .A1 (nx17702), .S0 (nx23501)
             ) ;
    mux21_ni ix17691 (.Y (nx17690), .A0 (inputs_424__4), .A1 (inputs_425__4), .S0 (
             nx24141)) ;
    mux21_ni ix17703 (.Y (nx17702), .A0 (inputs_426__4), .A1 (inputs_427__4), .S0 (
             nx24141)) ;
    mux21_ni ix17735 (.Y (nx17734), .A0 (nx17718), .A1 (nx17730), .S0 (nx23501)
             ) ;
    mux21_ni ix17719 (.Y (nx17718), .A0 (inputs_428__4), .A1 (inputs_429__4), .S0 (
             nx24141)) ;
    mux21_ni ix17731 (.Y (nx17730), .A0 (inputs_430__4), .A1 (inputs_431__4), .S0 (
             nx24141)) ;
    mux21_ni ix17799 (.Y (nx17798), .A0 (nx17766), .A1 (nx17794), .S0 (nx23229)
             ) ;
    mux21_ni ix17767 (.Y (nx17766), .A0 (nx17750), .A1 (nx17762), .S0 (nx23501)
             ) ;
    mux21_ni ix17751 (.Y (nx17750), .A0 (inputs_440__4), .A1 (inputs_441__4), .S0 (
             nx24143)) ;
    mux21_ni ix17763 (.Y (nx17762), .A0 (inputs_442__4), .A1 (inputs_443__4), .S0 (
             nx24143)) ;
    mux21_ni ix17795 (.Y (nx17794), .A0 (nx17778), .A1 (nx17790), .S0 (nx23503)
             ) ;
    mux21_ni ix17779 (.Y (nx17778), .A0 (inputs_444__4), .A1 (inputs_445__4), .S0 (
             nx24143)) ;
    mux21_ni ix17791 (.Y (nx17790), .A0 (inputs_446__4), .A1 (inputs_447__4), .S0 (
             nx24143)) ;
    mux21_ni ix18311 (.Y (nx18310), .A0 (nx18098), .A1 (nx18306), .S0 (nx22563)
             ) ;
    mux21_ni ix18099 (.Y (nx18098), .A0 (nx18092), .A1 (nx18014), .S0 (nx23137)
             ) ;
    oai21 ix18093 (.Y (nx18092), .A0 (nx22267), .A1 (nx12029), .B0 (nx12041)) ;
    mux21 ix12030 (.Y (nx12029), .A0 (nx18056), .A1 (nx18084), .S0 (nx22791)) ;
    mux21_ni ix18057 (.Y (nx18056), .A0 (nx18040), .A1 (nx18052), .S0 (nx23503)
             ) ;
    mux21_ni ix18041 (.Y (nx18040), .A0 (inputs_452__4), .A1 (inputs_453__4), .S0 (
             nx24143)) ;
    mux21_ni ix18053 (.Y (nx18052), .A0 (inputs_454__4), .A1 (inputs_455__4), .S0 (
             nx24143)) ;
    mux21_ni ix18085 (.Y (nx18084), .A0 (nx18068), .A1 (nx18080), .S0 (nx23503)
             ) ;
    mux21_ni ix18069 (.Y (nx18068), .A0 (inputs_468__4), .A1 (inputs_469__4), .S0 (
             nx24143)) ;
    mux21_ni ix18081 (.Y (nx18080), .A0 (inputs_470__4), .A1 (inputs_471__4), .S0 (
             nx24145)) ;
    nand04 ix12042 (.Y (nx12041), .A0 (nx22267), .A1 (nx23503), .A2 (nx24145), .A3 (
           nx18028)) ;
    mux21_ni ix18029 (.Y (nx18028), .A0 (inputs_451__4), .A1 (inputs_467__4), .S0 (
             nx22791)) ;
    mux21_ni ix18015 (.Y (nx18014), .A0 (nx17950), .A1 (nx18010), .S0 (nx22791)
             ) ;
    mux21_ni ix17951 (.Y (nx17950), .A0 (nx17918), .A1 (nx17946), .S0 (nx23231)
             ) ;
    mux21_ni ix17919 (.Y (nx17918), .A0 (nx17902), .A1 (nx17914), .S0 (nx23503)
             ) ;
    mux21_ni ix17903 (.Y (nx17902), .A0 (inputs_456__4), .A1 (inputs_457__4), .S0 (
             nx24145)) ;
    mux21_ni ix17915 (.Y (nx17914), .A0 (inputs_458__4), .A1 (inputs_459__4), .S0 (
             nx24145)) ;
    mux21_ni ix17947 (.Y (nx17946), .A0 (nx17930), .A1 (nx17942), .S0 (nx23503)
             ) ;
    mux21_ni ix17931 (.Y (nx17930), .A0 (inputs_460__4), .A1 (inputs_461__4), .S0 (
             nx24145)) ;
    mux21_ni ix17943 (.Y (nx17942), .A0 (inputs_462__4), .A1 (inputs_463__4), .S0 (
             nx24145)) ;
    mux21_ni ix18011 (.Y (nx18010), .A0 (nx17978), .A1 (nx18006), .S0 (nx23231)
             ) ;
    mux21_ni ix17979 (.Y (nx17978), .A0 (nx17962), .A1 (nx17974), .S0 (nx23503)
             ) ;
    mux21_ni ix17963 (.Y (nx17962), .A0 (inputs_472__4), .A1 (inputs_473__4), .S0 (
             nx24145)) ;
    mux21_ni ix17975 (.Y (nx17974), .A0 (inputs_474__4), .A1 (inputs_475__4), .S0 (
             nx24147)) ;
    mux21_ni ix18007 (.Y (nx18006), .A0 (nx17990), .A1 (nx18002), .S0 (nx23505)
             ) ;
    mux21_ni ix17991 (.Y (nx17990), .A0 (inputs_476__4), .A1 (inputs_477__4), .S0 (
             nx24147)) ;
    mux21_ni ix18003 (.Y (nx18002), .A0 (inputs_478__4), .A1 (inputs_479__4), .S0 (
             nx24147)) ;
    mux21_ni ix18307 (.Y (nx18306), .A0 (nx18300), .A1 (nx18222), .S0 (nx23137)
             ) ;
    oai21 ix18301 (.Y (nx18300), .A0 (nx22267), .A1 (nx12071), .B0 (nx12083)) ;
    mux21 ix12072 (.Y (nx12071), .A0 (nx18264), .A1 (nx18292), .S0 (nx22791)) ;
    mux21_ni ix18265 (.Y (nx18264), .A0 (nx18248), .A1 (nx18260), .S0 (nx23505)
             ) ;
    mux21_ni ix18249 (.Y (nx18248), .A0 (inputs_484__4), .A1 (inputs_485__4), .S0 (
             nx24147)) ;
    mux21_ni ix18261 (.Y (nx18260), .A0 (inputs_486__4), .A1 (inputs_487__4), .S0 (
             nx24147)) ;
    mux21_ni ix18293 (.Y (nx18292), .A0 (nx18276), .A1 (nx18288), .S0 (nx23505)
             ) ;
    mux21_ni ix18277 (.Y (nx18276), .A0 (inputs_500__4), .A1 (inputs_501__4), .S0 (
             nx24147)) ;
    mux21_ni ix18289 (.Y (nx18288), .A0 (inputs_502__4), .A1 (inputs_503__4), .S0 (
             nx24147)) ;
    nand04 ix12084 (.Y (nx12083), .A0 (nx22269), .A1 (nx23505), .A2 (nx24149), .A3 (
           nx18236)) ;
    mux21_ni ix18237 (.Y (nx18236), .A0 (inputs_483__4), .A1 (inputs_499__4), .S0 (
             nx22793)) ;
    mux21_ni ix18223 (.Y (nx18222), .A0 (nx18158), .A1 (nx18218), .S0 (nx22793)
             ) ;
    mux21_ni ix18159 (.Y (nx18158), .A0 (nx18126), .A1 (nx18154), .S0 (nx23231)
             ) ;
    mux21_ni ix18127 (.Y (nx18126), .A0 (nx18110), .A1 (nx18122), .S0 (nx23505)
             ) ;
    mux21_ni ix18111 (.Y (nx18110), .A0 (inputs_488__4), .A1 (inputs_489__4), .S0 (
             nx24149)) ;
    mux21_ni ix18123 (.Y (nx18122), .A0 (inputs_490__4), .A1 (inputs_491__4), .S0 (
             nx24149)) ;
    mux21_ni ix18155 (.Y (nx18154), .A0 (nx18138), .A1 (nx18150), .S0 (nx23505)
             ) ;
    mux21_ni ix18139 (.Y (nx18138), .A0 (inputs_492__4), .A1 (inputs_493__4), .S0 (
             nx24149)) ;
    mux21_ni ix18151 (.Y (nx18150), .A0 (inputs_494__4), .A1 (inputs_495__4), .S0 (
             nx24149)) ;
    mux21_ni ix18219 (.Y (nx18218), .A0 (nx18186), .A1 (nx18214), .S0 (nx23231)
             ) ;
    mux21_ni ix18187 (.Y (nx18186), .A0 (nx18170), .A1 (nx18182), .S0 (nx23505)
             ) ;
    mux21_ni ix18171 (.Y (nx18170), .A0 (inputs_504__4), .A1 (inputs_505__4), .S0 (
             nx24149)) ;
    mux21_ni ix18183 (.Y (nx18182), .A0 (inputs_506__4), .A1 (inputs_507__4), .S0 (
             nx24149)) ;
    mux21_ni ix18215 (.Y (nx18214), .A0 (nx18198), .A1 (nx18210), .S0 (nx23507)
             ) ;
    mux21_ni ix18199 (.Y (nx18198), .A0 (inputs_508__4), .A1 (inputs_509__4), .S0 (
             nx24151)) ;
    mux21_ni ix18211 (.Y (nx18210), .A0 (inputs_510__4), .A1 (inputs_511__4), .S0 (
             nx24151)) ;
    aoi32 ix12114 (.Y (nx12113), .A0 (nx19084), .A1 (nx22385), .A2 (nx22269), .B0 (
          nx22219), .B1 (nx20780)) ;
    oai21 ix19085 (.Y (nx19084), .A0 (nx23507), .A1 (nx12117), .B0 (nx12219)) ;
    mux21 ix12118 (.Y (nx12117), .A0 (nx18822), .A1 (nx19074), .S0 (nx24151)) ;
    mux21_ni ix18823 (.Y (nx18822), .A0 (nx18694), .A1 (nx18818), .S0 (nx22395)
             ) ;
    mux21_ni ix18695 (.Y (nx18694), .A0 (nx18630), .A1 (nx18690), .S0 (nx22419)
             ) ;
    mux21_ni ix18631 (.Y (nx18630), .A0 (nx18598), .A1 (nx18626), .S0 (nx22469)
             ) ;
    mux21_ni ix18599 (.Y (nx18598), .A0 (nx18582), .A1 (nx18594), .S0 (nx22563)
             ) ;
    mux21_ni ix18583 (.Y (nx18582), .A0 (inputs_0__4), .A1 (inputs_16__4), .S0 (
             nx22793)) ;
    mux21_ni ix18595 (.Y (nx18594), .A0 (inputs_32__4), .A1 (inputs_48__4), .S0 (
             nx22793)) ;
    mux21_ni ix18627 (.Y (nx18626), .A0 (nx18610), .A1 (nx18622), .S0 (nx22565)
             ) ;
    mux21_ni ix18611 (.Y (nx18610), .A0 (inputs_64__4), .A1 (inputs_80__4), .S0 (
             nx22793)) ;
    mux21_ni ix18623 (.Y (nx18622), .A0 (inputs_96__4), .A1 (inputs_112__4), .S0 (
             nx22793)) ;
    mux21_ni ix18691 (.Y (nx18690), .A0 (nx18658), .A1 (nx18686), .S0 (nx22469)
             ) ;
    mux21_ni ix18659 (.Y (nx18658), .A0 (nx18642), .A1 (nx18654), .S0 (nx22565)
             ) ;
    mux21_ni ix18643 (.Y (nx18642), .A0 (inputs_128__4), .A1 (inputs_144__4), .S0 (
             nx22793)) ;
    mux21_ni ix18655 (.Y (nx18654), .A0 (inputs_160__4), .A1 (inputs_176__4), .S0 (
             nx22795)) ;
    mux21_ni ix18687 (.Y (nx18686), .A0 (nx18670), .A1 (nx18682), .S0 (nx22565)
             ) ;
    mux21_ni ix18671 (.Y (nx18670), .A0 (inputs_192__4), .A1 (inputs_208__4), .S0 (
             nx22795)) ;
    mux21_ni ix18683 (.Y (nx18682), .A0 (inputs_224__4), .A1 (inputs_240__4), .S0 (
             nx22795)) ;
    mux21_ni ix18819 (.Y (nx18818), .A0 (nx18754), .A1 (nx18814), .S0 (nx22419)
             ) ;
    mux21_ni ix18755 (.Y (nx18754), .A0 (nx18722), .A1 (nx18750), .S0 (nx22469)
             ) ;
    mux21_ni ix18723 (.Y (nx18722), .A0 (nx18706), .A1 (nx18718), .S0 (nx22565)
             ) ;
    mux21_ni ix18707 (.Y (nx18706), .A0 (inputs_256__4), .A1 (inputs_272__4), .S0 (
             nx22795)) ;
    mux21_ni ix18719 (.Y (nx18718), .A0 (inputs_288__4), .A1 (inputs_304__4), .S0 (
             nx22795)) ;
    mux21_ni ix18751 (.Y (nx18750), .A0 (nx18734), .A1 (nx18746), .S0 (nx22565)
             ) ;
    mux21_ni ix18735 (.Y (nx18734), .A0 (inputs_320__4), .A1 (inputs_336__4), .S0 (
             nx22795)) ;
    mux21_ni ix18747 (.Y (nx18746), .A0 (inputs_352__4), .A1 (inputs_368__4), .S0 (
             nx22795)) ;
    mux21_ni ix18815 (.Y (nx18814), .A0 (nx18782), .A1 (nx18810), .S0 (nx22469)
             ) ;
    mux21_ni ix18783 (.Y (nx18782), .A0 (nx18766), .A1 (nx18778), .S0 (nx22565)
             ) ;
    mux21_ni ix18767 (.Y (nx18766), .A0 (inputs_384__4), .A1 (inputs_400__4), .S0 (
             nx22797)) ;
    mux21_ni ix18779 (.Y (nx18778), .A0 (inputs_416__4), .A1 (inputs_432__4), .S0 (
             nx22797)) ;
    mux21_ni ix18811 (.Y (nx18810), .A0 (nx18794), .A1 (nx18806), .S0 (nx22565)
             ) ;
    mux21_ni ix18795 (.Y (nx18794), .A0 (inputs_448__4), .A1 (inputs_464__4), .S0 (
             nx22797)) ;
    mux21_ni ix18807 (.Y (nx18806), .A0 (inputs_480__4), .A1 (inputs_496__4), .S0 (
             nx22797)) ;
    mux21_ni ix19075 (.Y (nx19074), .A0 (nx18946), .A1 (nx19070), .S0 (nx22395)
             ) ;
    mux21_ni ix18947 (.Y (nx18946), .A0 (nx18882), .A1 (nx18942), .S0 (nx22421)
             ) ;
    mux21_ni ix18883 (.Y (nx18882), .A0 (nx18850), .A1 (nx18878), .S0 (nx22471)
             ) ;
    mux21_ni ix18851 (.Y (nx18850), .A0 (nx18834), .A1 (nx18846), .S0 (nx22567)
             ) ;
    mux21_ni ix18835 (.Y (nx18834), .A0 (inputs_1__4), .A1 (inputs_17__4), .S0 (
             nx22797)) ;
    mux21_ni ix18847 (.Y (nx18846), .A0 (inputs_33__4), .A1 (inputs_49__4), .S0 (
             nx22797)) ;
    mux21_ni ix18879 (.Y (nx18878), .A0 (nx18862), .A1 (nx18874), .S0 (nx22567)
             ) ;
    mux21_ni ix18863 (.Y (nx18862), .A0 (inputs_65__4), .A1 (inputs_81__4), .S0 (
             nx22797)) ;
    mux21_ni ix18875 (.Y (nx18874), .A0 (inputs_97__4), .A1 (inputs_113__4), .S0 (
             nx22799)) ;
    mux21_ni ix18943 (.Y (nx18942), .A0 (nx18910), .A1 (nx18938), .S0 (nx22471)
             ) ;
    mux21_ni ix18911 (.Y (nx18910), .A0 (nx18894), .A1 (nx18906), .S0 (nx22567)
             ) ;
    mux21_ni ix18895 (.Y (nx18894), .A0 (inputs_129__4), .A1 (inputs_145__4), .S0 (
             nx22799)) ;
    mux21_ni ix18907 (.Y (nx18906), .A0 (inputs_161__4), .A1 (inputs_177__4), .S0 (
             nx22799)) ;
    mux21_ni ix18939 (.Y (nx18938), .A0 (nx18922), .A1 (nx18934), .S0 (nx22567)
             ) ;
    mux21_ni ix18923 (.Y (nx18922), .A0 (inputs_193__4), .A1 (inputs_209__4), .S0 (
             nx22799)) ;
    mux21_ni ix18935 (.Y (nx18934), .A0 (inputs_225__4), .A1 (inputs_241__4), .S0 (
             nx22799)) ;
    mux21_ni ix19071 (.Y (nx19070), .A0 (nx19006), .A1 (nx19066), .S0 (nx22421)
             ) ;
    mux21_ni ix19007 (.Y (nx19006), .A0 (nx18974), .A1 (nx19002), .S0 (nx22471)
             ) ;
    mux21_ni ix18975 (.Y (nx18974), .A0 (nx18958), .A1 (nx18970), .S0 (nx22567)
             ) ;
    mux21_ni ix18959 (.Y (nx18958), .A0 (inputs_257__4), .A1 (inputs_273__4), .S0 (
             nx22799)) ;
    mux21_ni ix18971 (.Y (nx18970), .A0 (inputs_289__4), .A1 (inputs_305__4), .S0 (
             nx22799)) ;
    mux21_ni ix19003 (.Y (nx19002), .A0 (nx18986), .A1 (nx18998), .S0 (nx22567)
             ) ;
    mux21_ni ix18987 (.Y (nx18986), .A0 (inputs_321__4), .A1 (inputs_337__4), .S0 (
             nx22801)) ;
    mux21_ni ix18999 (.Y (nx18998), .A0 (inputs_353__4), .A1 (inputs_369__4), .S0 (
             nx22801)) ;
    mux21_ni ix19067 (.Y (nx19066), .A0 (nx19034), .A1 (nx19062), .S0 (nx22471)
             ) ;
    mux21_ni ix19035 (.Y (nx19034), .A0 (nx19018), .A1 (nx19030), .S0 (nx22567)
             ) ;
    mux21_ni ix19019 (.Y (nx19018), .A0 (inputs_385__4), .A1 (inputs_401__4), .S0 (
             nx22801)) ;
    mux21_ni ix19031 (.Y (nx19030), .A0 (inputs_417__4), .A1 (inputs_433__4), .S0 (
             nx22801)) ;
    mux21_ni ix19063 (.Y (nx19062), .A0 (nx19046), .A1 (nx19058), .S0 (nx22569)
             ) ;
    mux21_ni ix19047 (.Y (nx19046), .A0 (inputs_449__4), .A1 (inputs_465__4), .S0 (
             nx22801)) ;
    mux21_ni ix19059 (.Y (nx19058), .A0 (inputs_481__4), .A1 (inputs_497__4), .S0 (
             nx22801)) ;
    nand03 ix12220 (.Y (nx12219), .A0 (nx18568), .A1 (nx23507), .A2 (nx24879)) ;
    mux21_ni ix18569 (.Y (nx18568), .A0 (nx18440), .A1 (nx18564), .S0 (nx22397)
             ) ;
    mux21_ni ix18441 (.Y (nx18440), .A0 (nx18376), .A1 (nx18436), .S0 (nx22421)
             ) ;
    mux21_ni ix18377 (.Y (nx18376), .A0 (nx18344), .A1 (nx18372), .S0 (nx22471)
             ) ;
    mux21_ni ix18345 (.Y (nx18344), .A0 (nx18328), .A1 (nx18340), .S0 (nx22569)
             ) ;
    mux21_ni ix18329 (.Y (nx18328), .A0 (inputs_2__4), .A1 (inputs_18__4), .S0 (
             nx22801)) ;
    mux21_ni ix18341 (.Y (nx18340), .A0 (inputs_34__4), .A1 (inputs_50__4), .S0 (
             nx22803)) ;
    mux21_ni ix18373 (.Y (nx18372), .A0 (nx18356), .A1 (nx18368), .S0 (nx22569)
             ) ;
    mux21_ni ix18357 (.Y (nx18356), .A0 (inputs_66__4), .A1 (inputs_82__4), .S0 (
             nx22803)) ;
    mux21_ni ix18369 (.Y (nx18368), .A0 (inputs_98__4), .A1 (inputs_114__4), .S0 (
             nx22803)) ;
    mux21_ni ix18437 (.Y (nx18436), .A0 (nx18404), .A1 (nx18432), .S0 (nx22471)
             ) ;
    mux21_ni ix18405 (.Y (nx18404), .A0 (nx18388), .A1 (nx18400), .S0 (nx22569)
             ) ;
    mux21_ni ix18389 (.Y (nx18388), .A0 (inputs_130__4), .A1 (inputs_146__4), .S0 (
             nx22803)) ;
    mux21_ni ix18401 (.Y (nx18400), .A0 (inputs_162__4), .A1 (inputs_178__4), .S0 (
             nx22803)) ;
    mux21_ni ix18433 (.Y (nx18432), .A0 (nx18416), .A1 (nx18428), .S0 (nx22569)
             ) ;
    mux21_ni ix18417 (.Y (nx18416), .A0 (inputs_194__4), .A1 (inputs_210__4), .S0 (
             nx22803)) ;
    mux21_ni ix18429 (.Y (nx18428), .A0 (inputs_226__4), .A1 (inputs_242__4), .S0 (
             nx22803)) ;
    mux21_ni ix18565 (.Y (nx18564), .A0 (nx18500), .A1 (nx18560), .S0 (nx22421)
             ) ;
    mux21_ni ix18501 (.Y (nx18500), .A0 (nx18468), .A1 (nx18496), .S0 (nx22471)
             ) ;
    mux21_ni ix18469 (.Y (nx18468), .A0 (nx18452), .A1 (nx18464), .S0 (nx22569)
             ) ;
    mux21_ni ix18453 (.Y (nx18452), .A0 (inputs_258__4), .A1 (inputs_274__4), .S0 (
             nx22805)) ;
    mux21_ni ix18465 (.Y (nx18464), .A0 (inputs_290__4), .A1 (inputs_306__4), .S0 (
             nx22805)) ;
    mux21_ni ix18497 (.Y (nx18496), .A0 (nx18480), .A1 (nx18492), .S0 (nx22569)
             ) ;
    mux21_ni ix18481 (.Y (nx18480), .A0 (inputs_322__4), .A1 (inputs_338__4), .S0 (
             nx22805)) ;
    mux21_ni ix18493 (.Y (nx18492), .A0 (inputs_354__4), .A1 (inputs_370__4), .S0 (
             nx22805)) ;
    mux21_ni ix18561 (.Y (nx18560), .A0 (nx18528), .A1 (nx18556), .S0 (nx22473)
             ) ;
    mux21_ni ix18529 (.Y (nx18528), .A0 (nx18512), .A1 (nx18524), .S0 (nx22571)
             ) ;
    mux21_ni ix18513 (.Y (nx18512), .A0 (inputs_386__4), .A1 (inputs_402__4), .S0 (
             nx22805)) ;
    mux21_ni ix18525 (.Y (nx18524), .A0 (inputs_418__4), .A1 (inputs_434__4), .S0 (
             nx22805)) ;
    mux21_ni ix18557 (.Y (nx18556), .A0 (nx18540), .A1 (nx18552), .S0 (nx22571)
             ) ;
    mux21_ni ix18541 (.Y (nx18540), .A0 (inputs_450__4), .A1 (inputs_466__4), .S0 (
             nx22805)) ;
    mux21_ni ix18553 (.Y (nx18552), .A0 (inputs_482__4), .A1 (inputs_498__4), .S0 (
             nx22807)) ;
    mux21_ni ix20781 (.Y (nx20780), .A0 (nx19932), .A1 (nx20776), .S0 (nx22421)
             ) ;
    mux21_ni ix19933 (.Y (nx19932), .A0 (nx19508), .A1 (nx19928), .S0 (nx22473)
             ) ;
    mux21_ni ix19509 (.Y (nx19508), .A0 (nx19296), .A1 (nx19504), .S0 (nx22571)
             ) ;
    mux21_ni ix19297 (.Y (nx19296), .A0 (nx19290), .A1 (nx19212), .S0 (nx23137)
             ) ;
    oai21 ix19291 (.Y (nx19290), .A0 (nx22269), .A1 (nx12279), .B0 (nx12291)) ;
    mux21 ix12280 (.Y (nx12279), .A0 (nx19254), .A1 (nx19282), .S0 (nx22807)) ;
    mux21_ni ix19255 (.Y (nx19254), .A0 (nx19238), .A1 (nx19250), .S0 (nx23507)
             ) ;
    mux21_ni ix19239 (.Y (nx19238), .A0 (inputs_4__4), .A1 (inputs_5__4), .S0 (
             nx24151)) ;
    mux21_ni ix19251 (.Y (nx19250), .A0 (inputs_6__4), .A1 (inputs_7__4), .S0 (
             nx24151)) ;
    mux21_ni ix19283 (.Y (nx19282), .A0 (nx19266), .A1 (nx19278), .S0 (nx23507)
             ) ;
    mux21_ni ix19267 (.Y (nx19266), .A0 (inputs_20__4), .A1 (inputs_21__4), .S0 (
             nx24151)) ;
    mux21_ni ix19279 (.Y (nx19278), .A0 (inputs_22__4), .A1 (inputs_23__4), .S0 (
             nx24151)) ;
    nand04 ix12292 (.Y (nx12291), .A0 (nx22269), .A1 (nx23507), .A2 (nx24153), .A3 (
           nx19226)) ;
    mux21_ni ix19227 (.Y (nx19226), .A0 (inputs_3__4), .A1 (inputs_19__4), .S0 (
             nx22807)) ;
    mux21_ni ix19213 (.Y (nx19212), .A0 (nx19148), .A1 (nx19208), .S0 (nx22807)
             ) ;
    mux21_ni ix19149 (.Y (nx19148), .A0 (nx19116), .A1 (nx19144), .S0 (nx23231)
             ) ;
    mux21_ni ix19117 (.Y (nx19116), .A0 (nx19100), .A1 (nx19112), .S0 (nx23507)
             ) ;
    mux21_ni ix19101 (.Y (nx19100), .A0 (inputs_8__4), .A1 (inputs_9__4), .S0 (
             nx24153)) ;
    mux21_ni ix19113 (.Y (nx19112), .A0 (inputs_10__4), .A1 (inputs_11__4), .S0 (
             nx24153)) ;
    mux21_ni ix19145 (.Y (nx19144), .A0 (nx19128), .A1 (nx19140), .S0 (nx23509)
             ) ;
    mux21_ni ix19129 (.Y (nx19128), .A0 (inputs_12__4), .A1 (inputs_13__4), .S0 (
             nx24153)) ;
    mux21_ni ix19141 (.Y (nx19140), .A0 (inputs_14__4), .A1 (inputs_15__4), .S0 (
             nx24153)) ;
    mux21_ni ix19209 (.Y (nx19208), .A0 (nx19176), .A1 (nx19204), .S0 (nx23231)
             ) ;
    mux21_ni ix19177 (.Y (nx19176), .A0 (nx19160), .A1 (nx19172), .S0 (nx23509)
             ) ;
    mux21_ni ix19161 (.Y (nx19160), .A0 (inputs_24__4), .A1 (inputs_25__4), .S0 (
             nx24153)) ;
    mux21_ni ix19173 (.Y (nx19172), .A0 (inputs_26__4), .A1 (inputs_27__4), .S0 (
             nx24153)) ;
    mux21_ni ix19205 (.Y (nx19204), .A0 (nx19188), .A1 (nx19200), .S0 (nx23509)
             ) ;
    mux21_ni ix19189 (.Y (nx19188), .A0 (inputs_28__4), .A1 (inputs_29__4), .S0 (
             nx24155)) ;
    mux21_ni ix19201 (.Y (nx19200), .A0 (inputs_30__4), .A1 (inputs_31__4), .S0 (
             nx24155)) ;
    mux21_ni ix19505 (.Y (nx19504), .A0 (nx19498), .A1 (nx19420), .S0 (nx23137)
             ) ;
    oai21 ix19499 (.Y (nx19498), .A0 (nx22269), .A1 (nx12323), .B0 (nx12337)) ;
    mux21 ix12324 (.Y (nx12323), .A0 (nx19462), .A1 (nx19490), .S0 (nx22807)) ;
    mux21_ni ix19463 (.Y (nx19462), .A0 (nx19446), .A1 (nx19458), .S0 (nx23509)
             ) ;
    mux21_ni ix19447 (.Y (nx19446), .A0 (inputs_36__4), .A1 (inputs_37__4), .S0 (
             nx24155)) ;
    mux21_ni ix19459 (.Y (nx19458), .A0 (inputs_38__4), .A1 (inputs_39__4), .S0 (
             nx24155)) ;
    mux21_ni ix19491 (.Y (nx19490), .A0 (nx19474), .A1 (nx19486), .S0 (nx23509)
             ) ;
    mux21_ni ix19475 (.Y (nx19474), .A0 (inputs_52__4), .A1 (inputs_53__4), .S0 (
             nx24155)) ;
    mux21_ni ix19487 (.Y (nx19486), .A0 (inputs_54__4), .A1 (inputs_55__4), .S0 (
             nx24155)) ;
    nand04 ix12338 (.Y (nx12337), .A0 (nx22269), .A1 (nx23509), .A2 (nx24155), .A3 (
           nx19434)) ;
    mux21_ni ix19435 (.Y (nx19434), .A0 (inputs_35__4), .A1 (inputs_51__4), .S0 (
             nx22807)) ;
    mux21_ni ix19421 (.Y (nx19420), .A0 (nx19356), .A1 (nx19416), .S0 (nx22807)
             ) ;
    mux21_ni ix19357 (.Y (nx19356), .A0 (nx19324), .A1 (nx19352), .S0 (nx23231)
             ) ;
    mux21_ni ix19325 (.Y (nx19324), .A0 (nx19308), .A1 (nx19320), .S0 (nx23509)
             ) ;
    mux21_ni ix19309 (.Y (nx19308), .A0 (inputs_40__4), .A1 (inputs_41__4), .S0 (
             nx24157)) ;
    mux21_ni ix19321 (.Y (nx19320), .A0 (inputs_42__4), .A1 (inputs_43__4), .S0 (
             nx24157)) ;
    mux21_ni ix19353 (.Y (nx19352), .A0 (nx19336), .A1 (nx19348), .S0 (nx23511)
             ) ;
    mux21_ni ix19337 (.Y (nx19336), .A0 (inputs_44__4), .A1 (inputs_45__4), .S0 (
             nx24157)) ;
    mux21_ni ix19349 (.Y (nx19348), .A0 (inputs_46__4), .A1 (inputs_47__4), .S0 (
             nx24157)) ;
    mux21_ni ix19417 (.Y (nx19416), .A0 (nx19384), .A1 (nx19412), .S0 (nx23233)
             ) ;
    mux21_ni ix19385 (.Y (nx19384), .A0 (nx19368), .A1 (nx19380), .S0 (nx23511)
             ) ;
    mux21_ni ix19369 (.Y (nx19368), .A0 (inputs_56__4), .A1 (inputs_57__4), .S0 (
             nx24157)) ;
    mux21_ni ix19381 (.Y (nx19380), .A0 (inputs_58__4), .A1 (inputs_59__4), .S0 (
             nx24157)) ;
    mux21_ni ix19413 (.Y (nx19412), .A0 (nx19396), .A1 (nx19408), .S0 (nx23511)
             ) ;
    mux21_ni ix19397 (.Y (nx19396), .A0 (inputs_60__4), .A1 (inputs_61__4), .S0 (
             nx24157)) ;
    mux21_ni ix19409 (.Y (nx19408), .A0 (inputs_62__4), .A1 (inputs_63__4), .S0 (
             nx24159)) ;
    mux21_ni ix19929 (.Y (nx19928), .A0 (nx19716), .A1 (nx19924), .S0 (nx22571)
             ) ;
    mux21_ni ix19717 (.Y (nx19716), .A0 (nx19710), .A1 (nx19632), .S0 (nx23137)
             ) ;
    oai21 ix19711 (.Y (nx19710), .A0 (nx22269), .A1 (nx12371), .B0 (nx12381)) ;
    mux21 ix12372 (.Y (nx12371), .A0 (nx19674), .A1 (nx19702), .S0 (nx22809)) ;
    mux21_ni ix19675 (.Y (nx19674), .A0 (nx19658), .A1 (nx19670), .S0 (nx23511)
             ) ;
    mux21_ni ix19659 (.Y (nx19658), .A0 (inputs_68__4), .A1 (inputs_69__4), .S0 (
             nx24159)) ;
    mux21_ni ix19671 (.Y (nx19670), .A0 (inputs_70__4), .A1 (inputs_71__4), .S0 (
             nx24159)) ;
    mux21_ni ix19703 (.Y (nx19702), .A0 (nx19686), .A1 (nx19698), .S0 (nx23511)
             ) ;
    mux21_ni ix19687 (.Y (nx19686), .A0 (inputs_84__4), .A1 (inputs_85__4), .S0 (
             nx24159)) ;
    mux21_ni ix19699 (.Y (nx19698), .A0 (inputs_86__4), .A1 (inputs_87__4), .S0 (
             nx24159)) ;
    nand04 ix12382 (.Y (nx12381), .A0 (nx22271), .A1 (nx23511), .A2 (nx24159), .A3 (
           nx19646)) ;
    mux21_ni ix19647 (.Y (nx19646), .A0 (inputs_67__4), .A1 (inputs_83__4), .S0 (
             nx22809)) ;
    mux21_ni ix19633 (.Y (nx19632), .A0 (nx19568), .A1 (nx19628), .S0 (nx22809)
             ) ;
    mux21_ni ix19569 (.Y (nx19568), .A0 (nx19536), .A1 (nx19564), .S0 (nx23233)
             ) ;
    mux21_ni ix19537 (.Y (nx19536), .A0 (nx19520), .A1 (nx19532), .S0 (nx23511)
             ) ;
    mux21_ni ix19521 (.Y (nx19520), .A0 (inputs_72__4), .A1 (inputs_73__4), .S0 (
             nx24159)) ;
    mux21_ni ix19533 (.Y (nx19532), .A0 (inputs_74__4), .A1 (inputs_75__4), .S0 (
             nx24161)) ;
    mux21_ni ix19565 (.Y (nx19564), .A0 (nx19548), .A1 (nx19560), .S0 (nx23513)
             ) ;
    mux21_ni ix19549 (.Y (nx19548), .A0 (inputs_76__4), .A1 (inputs_77__4), .S0 (
             nx24161)) ;
    mux21_ni ix19561 (.Y (nx19560), .A0 (inputs_78__4), .A1 (inputs_79__4), .S0 (
             nx24161)) ;
    mux21_ni ix19629 (.Y (nx19628), .A0 (nx19596), .A1 (nx19624), .S0 (nx23233)
             ) ;
    mux21_ni ix19597 (.Y (nx19596), .A0 (nx19580), .A1 (nx19592), .S0 (nx23513)
             ) ;
    mux21_ni ix19581 (.Y (nx19580), .A0 (inputs_88__4), .A1 (inputs_89__4), .S0 (
             nx24161)) ;
    mux21_ni ix19593 (.Y (nx19592), .A0 (inputs_90__4), .A1 (inputs_91__4), .S0 (
             nx24161)) ;
    mux21_ni ix19625 (.Y (nx19624), .A0 (nx19608), .A1 (nx19620), .S0 (nx23513)
             ) ;
    mux21_ni ix19609 (.Y (nx19608), .A0 (inputs_92__4), .A1 (inputs_93__4), .S0 (
             nx24161)) ;
    mux21_ni ix19621 (.Y (nx19620), .A0 (inputs_94__4), .A1 (inputs_95__4), .S0 (
             nx24161)) ;
    mux21_ni ix19925 (.Y (nx19924), .A0 (nx19918), .A1 (nx19840), .S0 (nx23137)
             ) ;
    oai21 ix19919 (.Y (nx19918), .A0 (nx22271), .A1 (nx12413), .B0 (nx12425)) ;
    mux21 ix12414 (.Y (nx12413), .A0 (nx19882), .A1 (nx19910), .S0 (nx22809)) ;
    mux21_ni ix19883 (.Y (nx19882), .A0 (nx19866), .A1 (nx19878), .S0 (nx23513)
             ) ;
    mux21_ni ix19867 (.Y (nx19866), .A0 (inputs_100__4), .A1 (inputs_101__4), .S0 (
             nx24163)) ;
    mux21_ni ix19879 (.Y (nx19878), .A0 (inputs_102__4), .A1 (inputs_103__4), .S0 (
             nx24163)) ;
    mux21_ni ix19911 (.Y (nx19910), .A0 (nx19894), .A1 (nx19906), .S0 (nx23513)
             ) ;
    mux21_ni ix19895 (.Y (nx19894), .A0 (inputs_116__4), .A1 (inputs_117__4), .S0 (
             nx24163)) ;
    mux21_ni ix19907 (.Y (nx19906), .A0 (inputs_118__4), .A1 (inputs_119__4), .S0 (
             nx24163)) ;
    nand04 ix12426 (.Y (nx12425), .A0 (nx22271), .A1 (nx23513), .A2 (nx24163), .A3 (
           nx19854)) ;
    mux21_ni ix19855 (.Y (nx19854), .A0 (inputs_99__4), .A1 (inputs_115__4), .S0 (
             nx22809)) ;
    mux21_ni ix19841 (.Y (nx19840), .A0 (nx19776), .A1 (nx19836), .S0 (nx22809)
             ) ;
    mux21_ni ix19777 (.Y (nx19776), .A0 (nx19744), .A1 (nx19772), .S0 (nx23233)
             ) ;
    mux21_ni ix19745 (.Y (nx19744), .A0 (nx19728), .A1 (nx19740), .S0 (nx23513)
             ) ;
    mux21_ni ix19729 (.Y (nx19728), .A0 (inputs_104__4), .A1 (inputs_105__4), .S0 (
             nx24163)) ;
    mux21_ni ix19741 (.Y (nx19740), .A0 (inputs_106__4), .A1 (inputs_107__4), .S0 (
             nx24163)) ;
    mux21_ni ix19773 (.Y (nx19772), .A0 (nx19756), .A1 (nx19768), .S0 (nx23515)
             ) ;
    mux21_ni ix19757 (.Y (nx19756), .A0 (inputs_108__4), .A1 (inputs_109__4), .S0 (
             nx24165)) ;
    mux21_ni ix19769 (.Y (nx19768), .A0 (inputs_110__4), .A1 (inputs_111__4), .S0 (
             nx24165)) ;
    mux21_ni ix19837 (.Y (nx19836), .A0 (nx19804), .A1 (nx19832), .S0 (nx23233)
             ) ;
    mux21_ni ix19805 (.Y (nx19804), .A0 (nx19788), .A1 (nx19800), .S0 (nx23515)
             ) ;
    mux21_ni ix19789 (.Y (nx19788), .A0 (inputs_120__4), .A1 (inputs_121__4), .S0 (
             nx24165)) ;
    mux21_ni ix19801 (.Y (nx19800), .A0 (inputs_122__4), .A1 (inputs_123__4), .S0 (
             nx24165)) ;
    mux21_ni ix19833 (.Y (nx19832), .A0 (nx19816), .A1 (nx19828), .S0 (nx23515)
             ) ;
    mux21_ni ix19817 (.Y (nx19816), .A0 (inputs_124__4), .A1 (inputs_125__4), .S0 (
             nx24165)) ;
    mux21_ni ix19829 (.Y (nx19828), .A0 (inputs_126__4), .A1 (inputs_127__4), .S0 (
             nx24165)) ;
    mux21_ni ix20777 (.Y (nx20776), .A0 (nx20352), .A1 (nx20772), .S0 (nx22473)
             ) ;
    mux21_ni ix20353 (.Y (nx20352), .A0 (nx20140), .A1 (nx20348), .S0 (nx22571)
             ) ;
    mux21_ni ix20141 (.Y (nx20140), .A0 (nx20134), .A1 (nx20056), .S0 (nx23137)
             ) ;
    oai21 ix20135 (.Y (nx20134), .A0 (nx22271), .A1 (nx12463), .B0 (nx12475)) ;
    mux21 ix12464 (.Y (nx12463), .A0 (nx20098), .A1 (nx20126), .S0 (nx22809)) ;
    mux21_ni ix20099 (.Y (nx20098), .A0 (nx20082), .A1 (nx20094), .S0 (nx23515)
             ) ;
    mux21_ni ix20083 (.Y (nx20082), .A0 (inputs_132__4), .A1 (inputs_133__4), .S0 (
             nx24165)) ;
    mux21_ni ix20095 (.Y (nx20094), .A0 (inputs_134__4), .A1 (inputs_135__4), .S0 (
             nx24167)) ;
    mux21_ni ix20127 (.Y (nx20126), .A0 (nx20110), .A1 (nx20122), .S0 (nx23515)
             ) ;
    mux21_ni ix20111 (.Y (nx20110), .A0 (inputs_148__4), .A1 (inputs_149__4), .S0 (
             nx24167)) ;
    mux21_ni ix20123 (.Y (nx20122), .A0 (inputs_150__4), .A1 (inputs_151__4), .S0 (
             nx24167)) ;
    nand04 ix12476 (.Y (nx12475), .A0 (nx22271), .A1 (nx23515), .A2 (nx24167), .A3 (
           nx20070)) ;
    mux21_ni ix20071 (.Y (nx20070), .A0 (inputs_131__4), .A1 (inputs_147__4), .S0 (
             nx22811)) ;
    mux21_ni ix20057 (.Y (nx20056), .A0 (nx19992), .A1 (nx20052), .S0 (nx22811)
             ) ;
    mux21_ni ix19993 (.Y (nx19992), .A0 (nx19960), .A1 (nx19988), .S0 (nx23233)
             ) ;
    mux21_ni ix19961 (.Y (nx19960), .A0 (nx19944), .A1 (nx19956), .S0 (nx23515)
             ) ;
    mux21_ni ix19945 (.Y (nx19944), .A0 (inputs_136__4), .A1 (inputs_137__4), .S0 (
             nx24167)) ;
    mux21_ni ix19957 (.Y (nx19956), .A0 (inputs_138__4), .A1 (inputs_139__4), .S0 (
             nx24167)) ;
    mux21_ni ix19989 (.Y (nx19988), .A0 (nx19972), .A1 (nx19984), .S0 (nx23517)
             ) ;
    mux21_ni ix19973 (.Y (nx19972), .A0 (inputs_140__4), .A1 (inputs_141__4), .S0 (
             nx24167)) ;
    mux21_ni ix19985 (.Y (nx19984), .A0 (inputs_142__4), .A1 (inputs_143__4), .S0 (
             nx24169)) ;
    mux21_ni ix20053 (.Y (nx20052), .A0 (nx20020), .A1 (nx20048), .S0 (nx23233)
             ) ;
    mux21_ni ix20021 (.Y (nx20020), .A0 (nx20004), .A1 (nx20016), .S0 (nx23517)
             ) ;
    mux21_ni ix20005 (.Y (nx20004), .A0 (inputs_152__4), .A1 (inputs_153__4), .S0 (
             nx24169)) ;
    mux21_ni ix20017 (.Y (nx20016), .A0 (inputs_154__4), .A1 (inputs_155__4), .S0 (
             nx24169)) ;
    mux21_ni ix20049 (.Y (nx20048), .A0 (nx20032), .A1 (nx20044), .S0 (nx23517)
             ) ;
    mux21_ni ix20033 (.Y (nx20032), .A0 (inputs_156__4), .A1 (inputs_157__4), .S0 (
             nx24169)) ;
    mux21_ni ix20045 (.Y (nx20044), .A0 (inputs_158__4), .A1 (inputs_159__4), .S0 (
             nx24169)) ;
    mux21_ni ix20349 (.Y (nx20348), .A0 (nx20342), .A1 (nx20264), .S0 (nx23139)
             ) ;
    oai21 ix20343 (.Y (nx20342), .A0 (nx22271), .A1 (nx12505), .B0 (nx12517)) ;
    mux21 ix12506 (.Y (nx12505), .A0 (nx20306), .A1 (nx20334), .S0 (nx22811)) ;
    mux21_ni ix20307 (.Y (nx20306), .A0 (nx20290), .A1 (nx20302), .S0 (nx23517)
             ) ;
    mux21_ni ix20291 (.Y (nx20290), .A0 (inputs_164__4), .A1 (inputs_165__4), .S0 (
             nx24169)) ;
    mux21_ni ix20303 (.Y (nx20302), .A0 (inputs_166__4), .A1 (inputs_167__4), .S0 (
             nx24169)) ;
    mux21_ni ix20335 (.Y (nx20334), .A0 (nx20318), .A1 (nx20330), .S0 (nx23517)
             ) ;
    mux21_ni ix20319 (.Y (nx20318), .A0 (inputs_180__4), .A1 (inputs_181__4), .S0 (
             nx24171)) ;
    mux21_ni ix20331 (.Y (nx20330), .A0 (inputs_182__4), .A1 (inputs_183__4), .S0 (
             nx24171)) ;
    nand04 ix12518 (.Y (nx12517), .A0 (nx22271), .A1 (nx23517), .A2 (nx24171), .A3 (
           nx20278)) ;
    mux21_ni ix20279 (.Y (nx20278), .A0 (inputs_163__4), .A1 (inputs_179__4), .S0 (
             nx22811)) ;
    mux21_ni ix20265 (.Y (nx20264), .A0 (nx20200), .A1 (nx20260), .S0 (nx22811)
             ) ;
    mux21_ni ix20201 (.Y (nx20200), .A0 (nx20168), .A1 (nx20196), .S0 (nx23235)
             ) ;
    mux21_ni ix20169 (.Y (nx20168), .A0 (nx20152), .A1 (nx20164), .S0 (nx23517)
             ) ;
    mux21_ni ix20153 (.Y (nx20152), .A0 (inputs_168__4), .A1 (inputs_169__4), .S0 (
             nx24171)) ;
    mux21_ni ix20165 (.Y (nx20164), .A0 (inputs_170__4), .A1 (inputs_171__4), .S0 (
             nx24171)) ;
    mux21_ni ix20197 (.Y (nx20196), .A0 (nx20180), .A1 (nx20192), .S0 (nx23519)
             ) ;
    mux21_ni ix20181 (.Y (nx20180), .A0 (inputs_172__4), .A1 (inputs_173__4), .S0 (
             nx24171)) ;
    mux21_ni ix20193 (.Y (nx20192), .A0 (inputs_174__4), .A1 (inputs_175__4), .S0 (
             nx24171)) ;
    mux21_ni ix20261 (.Y (nx20260), .A0 (nx20228), .A1 (nx20256), .S0 (nx23235)
             ) ;
    mux21_ni ix20229 (.Y (nx20228), .A0 (nx20212), .A1 (nx20224), .S0 (nx23519)
             ) ;
    mux21_ni ix20213 (.Y (nx20212), .A0 (inputs_184__4), .A1 (inputs_185__4), .S0 (
             nx24173)) ;
    mux21_ni ix20225 (.Y (nx20224), .A0 (inputs_186__4), .A1 (inputs_187__4), .S0 (
             nx24173)) ;
    mux21_ni ix20257 (.Y (nx20256), .A0 (nx20240), .A1 (nx20252), .S0 (nx23519)
             ) ;
    mux21_ni ix20241 (.Y (nx20240), .A0 (inputs_188__4), .A1 (inputs_189__4), .S0 (
             nx24173)) ;
    mux21_ni ix20253 (.Y (nx20252), .A0 (inputs_190__4), .A1 (inputs_191__4), .S0 (
             nx24173)) ;
    mux21_ni ix20773 (.Y (nx20772), .A0 (nx20560), .A1 (nx20768), .S0 (nx22571)
             ) ;
    mux21_ni ix20561 (.Y (nx20560), .A0 (nx20554), .A1 (nx20476), .S0 (nx23139)
             ) ;
    oai21 ix20555 (.Y (nx20554), .A0 (nx22273), .A1 (nx12549), .B0 (nx12561)) ;
    mux21 ix12550 (.Y (nx12549), .A0 (nx20518), .A1 (nx20546), .S0 (nx22811)) ;
    mux21_ni ix20519 (.Y (nx20518), .A0 (nx20502), .A1 (nx20514), .S0 (nx23519)
             ) ;
    mux21_ni ix20503 (.Y (nx20502), .A0 (inputs_196__4), .A1 (inputs_197__4), .S0 (
             nx24173)) ;
    mux21_ni ix20515 (.Y (nx20514), .A0 (inputs_198__4), .A1 (inputs_199__4), .S0 (
             nx24173)) ;
    mux21_ni ix20547 (.Y (nx20546), .A0 (nx20530), .A1 (nx20542), .S0 (nx23519)
             ) ;
    mux21_ni ix20531 (.Y (nx20530), .A0 (inputs_212__4), .A1 (inputs_213__4), .S0 (
             nx24173)) ;
    mux21_ni ix20543 (.Y (nx20542), .A0 (inputs_214__4), .A1 (inputs_215__4), .S0 (
             nx24175)) ;
    nand04 ix12562 (.Y (nx12561), .A0 (nx22273), .A1 (nx23519), .A2 (nx24175), .A3 (
           nx20490)) ;
    mux21_ni ix20491 (.Y (nx20490), .A0 (inputs_195__4), .A1 (inputs_211__4), .S0 (
             nx22811)) ;
    mux21_ni ix20477 (.Y (nx20476), .A0 (nx20412), .A1 (nx20472), .S0 (nx22813)
             ) ;
    mux21_ni ix20413 (.Y (nx20412), .A0 (nx20380), .A1 (nx20408), .S0 (nx23235)
             ) ;
    mux21_ni ix20381 (.Y (nx20380), .A0 (nx20364), .A1 (nx20376), .S0 (nx23519)
             ) ;
    mux21_ni ix20365 (.Y (nx20364), .A0 (inputs_200__4), .A1 (inputs_201__4), .S0 (
             nx24175)) ;
    mux21_ni ix20377 (.Y (nx20376), .A0 (inputs_202__4), .A1 (inputs_203__4), .S0 (
             nx24175)) ;
    mux21_ni ix20409 (.Y (nx20408), .A0 (nx20392), .A1 (nx20404), .S0 (nx23521)
             ) ;
    mux21_ni ix20393 (.Y (nx20392), .A0 (inputs_204__4), .A1 (inputs_205__4), .S0 (
             nx24175)) ;
    mux21_ni ix20405 (.Y (nx20404), .A0 (inputs_206__4), .A1 (inputs_207__4), .S0 (
             nx24175)) ;
    mux21_ni ix20473 (.Y (nx20472), .A0 (nx20440), .A1 (nx20468), .S0 (nx23235)
             ) ;
    mux21_ni ix20441 (.Y (nx20440), .A0 (nx20424), .A1 (nx20436), .S0 (nx23521)
             ) ;
    mux21_ni ix20425 (.Y (nx20424), .A0 (inputs_216__4), .A1 (inputs_217__4), .S0 (
             nx24175)) ;
    mux21_ni ix20437 (.Y (nx20436), .A0 (inputs_218__4), .A1 (inputs_219__4), .S0 (
             nx24177)) ;
    mux21_ni ix20469 (.Y (nx20468), .A0 (nx20452), .A1 (nx20464), .S0 (nx23521)
             ) ;
    mux21_ni ix20453 (.Y (nx20452), .A0 (inputs_220__4), .A1 (inputs_221__4), .S0 (
             nx24177)) ;
    mux21_ni ix20465 (.Y (nx20464), .A0 (inputs_222__4), .A1 (inputs_223__4), .S0 (
             nx24177)) ;
    mux21_ni ix20769 (.Y (nx20768), .A0 (nx20762), .A1 (nx20684), .S0 (nx23139)
             ) ;
    oai21 ix20763 (.Y (nx20762), .A0 (nx22273), .A1 (nx12593), .B0 (nx12603)) ;
    mux21 ix12594 (.Y (nx12593), .A0 (nx20726), .A1 (nx20754), .S0 (nx22813)) ;
    mux21_ni ix20727 (.Y (nx20726), .A0 (nx20710), .A1 (nx20722), .S0 (nx23521)
             ) ;
    mux21_ni ix20711 (.Y (nx20710), .A0 (inputs_228__4), .A1 (inputs_229__4), .S0 (
             nx24177)) ;
    mux21_ni ix20723 (.Y (nx20722), .A0 (inputs_230__4), .A1 (inputs_231__4), .S0 (
             nx24177)) ;
    mux21_ni ix20755 (.Y (nx20754), .A0 (nx20738), .A1 (nx20750), .S0 (nx23521)
             ) ;
    mux21_ni ix20739 (.Y (nx20738), .A0 (inputs_244__4), .A1 (inputs_245__4), .S0 (
             nx24177)) ;
    mux21_ni ix20751 (.Y (nx20750), .A0 (inputs_246__4), .A1 (inputs_247__4), .S0 (
             nx24177)) ;
    nand04 ix12604 (.Y (nx12603), .A0 (nx22273), .A1 (nx23521), .A2 (nx24179), .A3 (
           nx20698)) ;
    mux21_ni ix20699 (.Y (nx20698), .A0 (inputs_227__4), .A1 (inputs_243__4), .S0 (
             nx22813)) ;
    mux21_ni ix20685 (.Y (nx20684), .A0 (nx20620), .A1 (nx20680), .S0 (nx22813)
             ) ;
    mux21_ni ix20621 (.Y (nx20620), .A0 (nx20588), .A1 (nx20616), .S0 (nx23235)
             ) ;
    mux21_ni ix20589 (.Y (nx20588), .A0 (nx20572), .A1 (nx20584), .S0 (nx23521)
             ) ;
    mux21_ni ix20573 (.Y (nx20572), .A0 (inputs_232__4), .A1 (inputs_233__4), .S0 (
             nx24179)) ;
    mux21_ni ix20585 (.Y (nx20584), .A0 (inputs_234__4), .A1 (inputs_235__4), .S0 (
             nx24179)) ;
    mux21_ni ix20617 (.Y (nx20616), .A0 (nx20600), .A1 (nx20612), .S0 (nx23523)
             ) ;
    mux21_ni ix20601 (.Y (nx20600), .A0 (inputs_236__4), .A1 (inputs_237__4), .S0 (
             nx24179)) ;
    mux21_ni ix20613 (.Y (nx20612), .A0 (inputs_238__4), .A1 (inputs_239__4), .S0 (
             nx24179)) ;
    mux21_ni ix20681 (.Y (nx20680), .A0 (nx20648), .A1 (nx20676), .S0 (nx23235)
             ) ;
    mux21_ni ix20649 (.Y (nx20648), .A0 (nx20632), .A1 (nx20644), .S0 (nx23523)
             ) ;
    mux21_ni ix20633 (.Y (nx20632), .A0 (inputs_248__4), .A1 (inputs_249__4), .S0 (
             nx24179)) ;
    mux21_ni ix20645 (.Y (nx20644), .A0 (inputs_250__4), .A1 (inputs_251__4), .S0 (
             nx24179)) ;
    mux21_ni ix20677 (.Y (nx20676), .A0 (nx20660), .A1 (nx20672), .S0 (nx23523)
             ) ;
    mux21_ni ix20661 (.Y (nx20660), .A0 (inputs_252__4), .A1 (inputs_253__4), .S0 (
             nx24181)) ;
    mux21_ni ix20673 (.Y (nx20672), .A0 (inputs_254__4), .A1 (inputs_255__4), .S0 (
             nx24181)) ;
    oai21 ix24947 (.Y (\output [5]), .A0 (nx22219), .A1 (nx12633), .B0 (nx12993)
          ) ;
    mux21 ix12634 (.Y (nx12633), .A0 (nx21628), .A1 (nx22472), .S0 (nx22421)) ;
    mux21_ni ix21629 (.Y (nx21628), .A0 (nx21204), .A1 (nx21624), .S0 (nx22473)
             ) ;
    mux21_ni ix21205 (.Y (nx21204), .A0 (nx20992), .A1 (nx21200), .S0 (nx22571)
             ) ;
    mux21_ni ix20993 (.Y (nx20992), .A0 (nx20986), .A1 (nx20908), .S0 (nx23139)
             ) ;
    oai21 ix20987 (.Y (nx20986), .A0 (nx22273), .A1 (nx12641), .B0 (nx12653)) ;
    mux21 ix12642 (.Y (nx12641), .A0 (nx20950), .A1 (nx20978), .S0 (nx22813)) ;
    mux21_ni ix20951 (.Y (nx20950), .A0 (nx20934), .A1 (nx20946), .S0 (nx23523)
             ) ;
    mux21_ni ix20935 (.Y (nx20934), .A0 (inputs_260__5), .A1 (inputs_261__5), .S0 (
             nx24181)) ;
    mux21_ni ix20947 (.Y (nx20946), .A0 (inputs_262__5), .A1 (inputs_263__5), .S0 (
             nx24181)) ;
    mux21_ni ix20979 (.Y (nx20978), .A0 (nx20962), .A1 (nx20974), .S0 (nx23523)
             ) ;
    mux21_ni ix20963 (.Y (nx20962), .A0 (inputs_276__5), .A1 (inputs_277__5), .S0 (
             nx24181)) ;
    mux21_ni ix20975 (.Y (nx20974), .A0 (inputs_278__5), .A1 (inputs_279__5), .S0 (
             nx24181)) ;
    nand04 ix12654 (.Y (nx12653), .A0 (nx22273), .A1 (nx23523), .A2 (nx24181), .A3 (
           nx20922)) ;
    mux21_ni ix20923 (.Y (nx20922), .A0 (inputs_259__5), .A1 (inputs_275__5), .S0 (
             nx22813)) ;
    mux21_ni ix20909 (.Y (nx20908), .A0 (nx20844), .A1 (nx20904), .S0 (nx22813)
             ) ;
    mux21_ni ix20845 (.Y (nx20844), .A0 (nx20812), .A1 (nx20840), .S0 (nx23235)
             ) ;
    mux21_ni ix20813 (.Y (nx20812), .A0 (nx20796), .A1 (nx20808), .S0 (nx23523)
             ) ;
    mux21_ni ix20797 (.Y (nx20796), .A0 (inputs_264__5), .A1 (inputs_265__5), .S0 (
             nx24183)) ;
    mux21_ni ix20809 (.Y (nx20808), .A0 (inputs_266__5), .A1 (inputs_267__5), .S0 (
             nx24183)) ;
    mux21_ni ix20841 (.Y (nx20840), .A0 (nx20824), .A1 (nx20836), .S0 (nx23525)
             ) ;
    mux21_ni ix20825 (.Y (nx20824), .A0 (inputs_268__5), .A1 (inputs_269__5), .S0 (
             nx24183)) ;
    mux21_ni ix20837 (.Y (nx20836), .A0 (inputs_270__5), .A1 (inputs_271__5), .S0 (
             nx24183)) ;
    mux21_ni ix20905 (.Y (nx20904), .A0 (nx20872), .A1 (nx20900), .S0 (nx23237)
             ) ;
    mux21_ni ix20873 (.Y (nx20872), .A0 (nx20856), .A1 (nx20868), .S0 (nx23525)
             ) ;
    mux21_ni ix20857 (.Y (nx20856), .A0 (inputs_280__5), .A1 (inputs_281__5), .S0 (
             nx24183)) ;
    mux21_ni ix20869 (.Y (nx20868), .A0 (inputs_282__5), .A1 (inputs_283__5), .S0 (
             nx24183)) ;
    mux21_ni ix20901 (.Y (nx20900), .A0 (nx20884), .A1 (nx20896), .S0 (nx23525)
             ) ;
    mux21_ni ix20885 (.Y (nx20884), .A0 (inputs_284__5), .A1 (inputs_285__5), .S0 (
             nx24183)) ;
    mux21_ni ix20897 (.Y (nx20896), .A0 (inputs_286__5), .A1 (inputs_287__5), .S0 (
             nx24185)) ;
    mux21_ni ix21201 (.Y (nx21200), .A0 (nx21194), .A1 (nx21116), .S0 (nx23139)
             ) ;
    oai21 ix21195 (.Y (nx21194), .A0 (nx22273), .A1 (nx12685), .B0 (nx12697)) ;
    mux21 ix12686 (.Y (nx12685), .A0 (nx21158), .A1 (nx21186), .S0 (nx22815)) ;
    mux21_ni ix21159 (.Y (nx21158), .A0 (nx21142), .A1 (nx21154), .S0 (nx23525)
             ) ;
    mux21_ni ix21143 (.Y (nx21142), .A0 (inputs_292__5), .A1 (inputs_293__5), .S0 (
             nx24185)) ;
    mux21_ni ix21155 (.Y (nx21154), .A0 (inputs_294__5), .A1 (inputs_295__5), .S0 (
             nx24185)) ;
    mux21_ni ix21187 (.Y (nx21186), .A0 (nx21170), .A1 (nx21182), .S0 (nx23525)
             ) ;
    mux21_ni ix21171 (.Y (nx21170), .A0 (inputs_308__5), .A1 (inputs_309__5), .S0 (
             nx24185)) ;
    mux21_ni ix21183 (.Y (nx21182), .A0 (inputs_310__5), .A1 (inputs_311__5), .S0 (
             nx24185)) ;
    nand04 ix12698 (.Y (nx12697), .A0 (nx22275), .A1 (nx23525), .A2 (nx24185), .A3 (
           nx21130)) ;
    mux21_ni ix21131 (.Y (nx21130), .A0 (inputs_291__5), .A1 (inputs_307__5), .S0 (
             nx22815)) ;
    mux21_ni ix21117 (.Y (nx21116), .A0 (nx21052), .A1 (nx21112), .S0 (nx22815)
             ) ;
    mux21_ni ix21053 (.Y (nx21052), .A0 (nx21020), .A1 (nx21048), .S0 (nx23237)
             ) ;
    mux21_ni ix21021 (.Y (nx21020), .A0 (nx21004), .A1 (nx21016), .S0 (nx23525)
             ) ;
    mux21_ni ix21005 (.Y (nx21004), .A0 (inputs_296__5), .A1 (inputs_297__5), .S0 (
             nx24185)) ;
    mux21_ni ix21017 (.Y (nx21016), .A0 (inputs_298__5), .A1 (inputs_299__5), .S0 (
             nx24187)) ;
    mux21_ni ix21049 (.Y (nx21048), .A0 (nx21032), .A1 (nx21044), .S0 (nx23527)
             ) ;
    mux21_ni ix21033 (.Y (nx21032), .A0 (inputs_300__5), .A1 (inputs_301__5), .S0 (
             nx24187)) ;
    mux21_ni ix21045 (.Y (nx21044), .A0 (inputs_302__5), .A1 (inputs_303__5), .S0 (
             nx24187)) ;
    mux21_ni ix21113 (.Y (nx21112), .A0 (nx21080), .A1 (nx21108), .S0 (nx23237)
             ) ;
    mux21_ni ix21081 (.Y (nx21080), .A0 (nx21064), .A1 (nx21076), .S0 (nx23527)
             ) ;
    mux21_ni ix21065 (.Y (nx21064), .A0 (inputs_312__5), .A1 (inputs_313__5), .S0 (
             nx24187)) ;
    mux21_ni ix21077 (.Y (nx21076), .A0 (inputs_314__5), .A1 (inputs_315__5), .S0 (
             nx24187)) ;
    mux21_ni ix21109 (.Y (nx21108), .A0 (nx21092), .A1 (nx21104), .S0 (nx23527)
             ) ;
    mux21_ni ix21093 (.Y (nx21092), .A0 (inputs_316__5), .A1 (inputs_317__5), .S0 (
             nx24187)) ;
    mux21_ni ix21105 (.Y (nx21104), .A0 (inputs_318__5), .A1 (inputs_319__5), .S0 (
             nx24187)) ;
    mux21_ni ix21625 (.Y (nx21624), .A0 (nx21412), .A1 (nx21620), .S0 (nx22573)
             ) ;
    mux21_ni ix21413 (.Y (nx21412), .A0 (nx21406), .A1 (nx21328), .S0 (nx23139)
             ) ;
    oai21 ix21407 (.Y (nx21406), .A0 (nx22275), .A1 (nx12729), .B0 (nx12741)) ;
    mux21 ix12730 (.Y (nx12729), .A0 (nx21370), .A1 (nx21398), .S0 (nx22815)) ;
    mux21_ni ix21371 (.Y (nx21370), .A0 (nx21354), .A1 (nx21366), .S0 (nx23527)
             ) ;
    mux21_ni ix21355 (.Y (nx21354), .A0 (inputs_324__5), .A1 (inputs_325__5), .S0 (
             nx24189)) ;
    mux21_ni ix21367 (.Y (nx21366), .A0 (inputs_326__5), .A1 (inputs_327__5), .S0 (
             nx24189)) ;
    mux21_ni ix21399 (.Y (nx21398), .A0 (nx21382), .A1 (nx21394), .S0 (nx23527)
             ) ;
    mux21_ni ix21383 (.Y (nx21382), .A0 (inputs_340__5), .A1 (inputs_341__5), .S0 (
             nx24189)) ;
    mux21_ni ix21395 (.Y (nx21394), .A0 (inputs_342__5), .A1 (inputs_343__5), .S0 (
             nx24189)) ;
    nand04 ix12742 (.Y (nx12741), .A0 (nx22275), .A1 (nx23527), .A2 (nx24189), .A3 (
           nx21342)) ;
    mux21_ni ix21343 (.Y (nx21342), .A0 (inputs_323__5), .A1 (inputs_339__5), .S0 (
             nx22815)) ;
    mux21_ni ix21329 (.Y (nx21328), .A0 (nx21264), .A1 (nx21324), .S0 (nx22815)
             ) ;
    mux21_ni ix21265 (.Y (nx21264), .A0 (nx21232), .A1 (nx21260), .S0 (nx23237)
             ) ;
    mux21_ni ix21233 (.Y (nx21232), .A0 (nx21216), .A1 (nx21228), .S0 (nx23527)
             ) ;
    mux21_ni ix21217 (.Y (nx21216), .A0 (inputs_328__5), .A1 (inputs_329__5), .S0 (
             nx24189)) ;
    mux21_ni ix21229 (.Y (nx21228), .A0 (inputs_330__5), .A1 (inputs_331__5), .S0 (
             nx24189)) ;
    mux21_ni ix21261 (.Y (nx21260), .A0 (nx21244), .A1 (nx21256), .S0 (nx23529)
             ) ;
    mux21_ni ix21245 (.Y (nx21244), .A0 (inputs_332__5), .A1 (inputs_333__5), .S0 (
             nx24191)) ;
    mux21_ni ix21257 (.Y (nx21256), .A0 (inputs_334__5), .A1 (inputs_335__5), .S0 (
             nx24191)) ;
    mux21_ni ix21325 (.Y (nx21324), .A0 (nx21292), .A1 (nx21320), .S0 (nx23237)
             ) ;
    mux21_ni ix21293 (.Y (nx21292), .A0 (nx21276), .A1 (nx21288), .S0 (nx23529)
             ) ;
    mux21_ni ix21277 (.Y (nx21276), .A0 (inputs_344__5), .A1 (inputs_345__5), .S0 (
             nx24191)) ;
    mux21_ni ix21289 (.Y (nx21288), .A0 (inputs_346__5), .A1 (inputs_347__5), .S0 (
             nx24191)) ;
    mux21_ni ix21321 (.Y (nx21320), .A0 (nx21304), .A1 (nx21316), .S0 (nx23529)
             ) ;
    mux21_ni ix21305 (.Y (nx21304), .A0 (inputs_348__5), .A1 (inputs_349__5), .S0 (
             nx24191)) ;
    mux21_ni ix21317 (.Y (nx21316), .A0 (inputs_350__5), .A1 (inputs_351__5), .S0 (
             nx24191)) ;
    mux21_ni ix21621 (.Y (nx21620), .A0 (nx21614), .A1 (nx21536), .S0 (nx23139)
             ) ;
    oai21 ix21615 (.Y (nx21614), .A0 (nx22275), .A1 (nx12771), .B0 (nx12783)) ;
    mux21 ix12772 (.Y (nx12771), .A0 (nx21578), .A1 (nx21606), .S0 (nx22815)) ;
    mux21_ni ix21579 (.Y (nx21578), .A0 (nx21562), .A1 (nx21574), .S0 (nx23529)
             ) ;
    mux21_ni ix21563 (.Y (nx21562), .A0 (inputs_356__5), .A1 (inputs_357__5), .S0 (
             nx24191)) ;
    mux21_ni ix21575 (.Y (nx21574), .A0 (inputs_358__5), .A1 (inputs_359__5), .S0 (
             nx24193)) ;
    mux21_ni ix21607 (.Y (nx21606), .A0 (nx21590), .A1 (nx21602), .S0 (nx23529)
             ) ;
    mux21_ni ix21591 (.Y (nx21590), .A0 (inputs_372__5), .A1 (inputs_373__5), .S0 (
             nx24193)) ;
    mux21_ni ix21603 (.Y (nx21602), .A0 (inputs_374__5), .A1 (inputs_375__5), .S0 (
             nx24193)) ;
    nand04 ix12784 (.Y (nx12783), .A0 (nx22275), .A1 (nx23529), .A2 (nx24193), .A3 (
           nx21550)) ;
    mux21_ni ix21551 (.Y (nx21550), .A0 (inputs_355__5), .A1 (inputs_371__5), .S0 (
             nx22817)) ;
    mux21_ni ix21537 (.Y (nx21536), .A0 (nx21472), .A1 (nx21532), .S0 (nx22817)
             ) ;
    mux21_ni ix21473 (.Y (nx21472), .A0 (nx21440), .A1 (nx21468), .S0 (nx23237)
             ) ;
    mux21_ni ix21441 (.Y (nx21440), .A0 (nx21424), .A1 (nx21436), .S0 (nx23529)
             ) ;
    mux21_ni ix21425 (.Y (nx21424), .A0 (inputs_360__5), .A1 (inputs_361__5), .S0 (
             nx24193)) ;
    mux21_ni ix21437 (.Y (nx21436), .A0 (inputs_362__5), .A1 (inputs_363__5), .S0 (
             nx24193)) ;
    mux21_ni ix21469 (.Y (nx21468), .A0 (nx21452), .A1 (nx21464), .S0 (nx23531)
             ) ;
    mux21_ni ix21453 (.Y (nx21452), .A0 (inputs_364__5), .A1 (inputs_365__5), .S0 (
             nx24193)) ;
    mux21_ni ix21465 (.Y (nx21464), .A0 (inputs_366__5), .A1 (inputs_367__5), .S0 (
             nx24195)) ;
    mux21_ni ix21533 (.Y (nx21532), .A0 (nx21500), .A1 (nx21528), .S0 (nx23237)
             ) ;
    mux21_ni ix21501 (.Y (nx21500), .A0 (nx21484), .A1 (nx21496), .S0 (nx23531)
             ) ;
    mux21_ni ix21485 (.Y (nx21484), .A0 (inputs_376__5), .A1 (inputs_377__5), .S0 (
             nx24195)) ;
    mux21_ni ix21497 (.Y (nx21496), .A0 (inputs_378__5), .A1 (inputs_379__5), .S0 (
             nx24195)) ;
    mux21_ni ix21529 (.Y (nx21528), .A0 (nx21512), .A1 (nx21524), .S0 (nx23531)
             ) ;
    mux21_ni ix21513 (.Y (nx21512), .A0 (inputs_380__5), .A1 (inputs_381__5), .S0 (
             nx24195)) ;
    mux21_ni ix21525 (.Y (nx21524), .A0 (inputs_382__5), .A1 (inputs_383__5), .S0 (
             nx24195)) ;
    mux21_ni ix22473 (.Y (nx22472), .A0 (nx22048), .A1 (nx22468), .S0 (nx22473)
             ) ;
    mux21_ni ix22049 (.Y (nx22048), .A0 (nx21836), .A1 (nx22044), .S0 (nx22573)
             ) ;
    mux21_ni ix21837 (.Y (nx21836), .A0 (nx21830), .A1 (nx21752), .S0 (nx23141)
             ) ;
    oai21 ix21831 (.Y (nx21830), .A0 (nx22275), .A1 (nx12821), .B0 (nx12833)) ;
    mux21 ix12822 (.Y (nx12821), .A0 (nx21794), .A1 (nx21822), .S0 (nx22817)) ;
    mux21_ni ix21795 (.Y (nx21794), .A0 (nx21778), .A1 (nx21790), .S0 (nx23531)
             ) ;
    mux21_ni ix21779 (.Y (nx21778), .A0 (inputs_388__5), .A1 (inputs_389__5), .S0 (
             nx24195)) ;
    mux21_ni ix21791 (.Y (nx21790), .A0 (inputs_390__5), .A1 (inputs_391__5), .S0 (
             nx24195)) ;
    mux21_ni ix21823 (.Y (nx21822), .A0 (nx21806), .A1 (nx21818), .S0 (nx23531)
             ) ;
    mux21_ni ix21807 (.Y (nx21806), .A0 (inputs_404__5), .A1 (inputs_405__5), .S0 (
             nx24197)) ;
    mux21_ni ix21819 (.Y (nx21818), .A0 (inputs_406__5), .A1 (inputs_407__5), .S0 (
             nx24197)) ;
    nand04 ix12834 (.Y (nx12833), .A0 (nx22275), .A1 (nx23531), .A2 (nx24197), .A3 (
           nx21766)) ;
    mux21_ni ix21767 (.Y (nx21766), .A0 (inputs_387__5), .A1 (inputs_403__5), .S0 (
             nx22817)) ;
    mux21_ni ix21753 (.Y (nx21752), .A0 (nx21688), .A1 (nx21748), .S0 (nx22817)
             ) ;
    mux21_ni ix21689 (.Y (nx21688), .A0 (nx21656), .A1 (nx21684), .S0 (nx23239)
             ) ;
    mux21_ni ix21657 (.Y (nx21656), .A0 (nx21640), .A1 (nx21652), .S0 (nx23531)
             ) ;
    mux21_ni ix21641 (.Y (nx21640), .A0 (inputs_392__5), .A1 (inputs_393__5), .S0 (
             nx24197)) ;
    mux21_ni ix21653 (.Y (nx21652), .A0 (inputs_394__5), .A1 (inputs_395__5), .S0 (
             nx24197)) ;
    mux21_ni ix21685 (.Y (nx21684), .A0 (nx21668), .A1 (nx21680), .S0 (nx23533)
             ) ;
    mux21_ni ix21669 (.Y (nx21668), .A0 (inputs_396__5), .A1 (inputs_397__5), .S0 (
             nx24197)) ;
    mux21_ni ix21681 (.Y (nx21680), .A0 (inputs_398__5), .A1 (inputs_399__5), .S0 (
             nx24197)) ;
    mux21_ni ix21749 (.Y (nx21748), .A0 (nx21716), .A1 (nx21744), .S0 (nx23239)
             ) ;
    mux21_ni ix21717 (.Y (nx21716), .A0 (nx21700), .A1 (nx21712), .S0 (nx23533)
             ) ;
    mux21_ni ix21701 (.Y (nx21700), .A0 (inputs_408__5), .A1 (inputs_409__5), .S0 (
             nx24199)) ;
    mux21_ni ix21713 (.Y (nx21712), .A0 (inputs_410__5), .A1 (inputs_411__5), .S0 (
             nx24199)) ;
    mux21_ni ix21745 (.Y (nx21744), .A0 (nx21728), .A1 (nx21740), .S0 (nx23533)
             ) ;
    mux21_ni ix21729 (.Y (nx21728), .A0 (inputs_412__5), .A1 (inputs_413__5), .S0 (
             nx24199)) ;
    mux21_ni ix21741 (.Y (nx21740), .A0 (inputs_414__5), .A1 (inputs_415__5), .S0 (
             nx24199)) ;
    mux21_ni ix22045 (.Y (nx22044), .A0 (nx22038), .A1 (nx21960), .S0 (nx23141)
             ) ;
    oai21 ix22039 (.Y (nx22038), .A0 (nx22277), .A1 (nx12863), .B0 (nx12877)) ;
    mux21 ix12864 (.Y (nx12863), .A0 (nx22002), .A1 (nx22030), .S0 (nx22817)) ;
    mux21_ni ix22003 (.Y (nx22002), .A0 (nx21986), .A1 (nx21998), .S0 (nx23533)
             ) ;
    mux21_ni ix21987 (.Y (nx21986), .A0 (inputs_420__5), .A1 (inputs_421__5), .S0 (
             nx24199)) ;
    mux21_ni ix21999 (.Y (nx21998), .A0 (inputs_422__5), .A1 (inputs_423__5), .S0 (
             nx24199)) ;
    mux21_ni ix22031 (.Y (nx22030), .A0 (nx22014), .A1 (nx22026), .S0 (nx23533)
             ) ;
    mux21_ni ix22015 (.Y (nx22014), .A0 (inputs_436__5), .A1 (inputs_437__5), .S0 (
             nx24199)) ;
    mux21_ni ix22027 (.Y (nx22026), .A0 (inputs_438__5), .A1 (inputs_439__5), .S0 (
             nx24201)) ;
    nand04 ix12878 (.Y (nx12877), .A0 (nx22277), .A1 (nx23533), .A2 (nx24201), .A3 (
           nx21974)) ;
    mux21_ni ix21975 (.Y (nx21974), .A0 (inputs_419__5), .A1 (inputs_435__5), .S0 (
             nx22817)) ;
    mux21_ni ix21961 (.Y (nx21960), .A0 (nx21896), .A1 (nx21956), .S0 (nx22819)
             ) ;
    mux21_ni ix21897 (.Y (nx21896), .A0 (nx21864), .A1 (nx21892), .S0 (nx23239)
             ) ;
    mux21_ni ix21865 (.Y (nx21864), .A0 (nx21848), .A1 (nx21860), .S0 (nx23533)
             ) ;
    mux21_ni ix21849 (.Y (nx21848), .A0 (inputs_424__5), .A1 (inputs_425__5), .S0 (
             nx24201)) ;
    mux21_ni ix21861 (.Y (nx21860), .A0 (inputs_426__5), .A1 (inputs_427__5), .S0 (
             nx24201)) ;
    mux21_ni ix21893 (.Y (nx21892), .A0 (nx21876), .A1 (nx21888), .S0 (nx23535)
             ) ;
    mux21_ni ix21877 (.Y (nx21876), .A0 (inputs_428__5), .A1 (inputs_429__5), .S0 (
             nx24201)) ;
    mux21_ni ix21889 (.Y (nx21888), .A0 (inputs_430__5), .A1 (inputs_431__5), .S0 (
             nx24201)) ;
    mux21_ni ix21957 (.Y (nx21956), .A0 (nx21924), .A1 (nx21952), .S0 (nx23239)
             ) ;
    mux21_ni ix21925 (.Y (nx21924), .A0 (nx21908), .A1 (nx21920), .S0 (nx23535)
             ) ;
    mux21_ni ix21909 (.Y (nx21908), .A0 (inputs_440__5), .A1 (inputs_441__5), .S0 (
             nx24201)) ;
    mux21_ni ix21921 (.Y (nx21920), .A0 (inputs_442__5), .A1 (inputs_443__5), .S0 (
             nx24203)) ;
    mux21_ni ix21953 (.Y (nx21952), .A0 (nx21936), .A1 (nx21948), .S0 (nx23535)
             ) ;
    mux21_ni ix21937 (.Y (nx21936), .A0 (inputs_444__5), .A1 (inputs_445__5), .S0 (
             nx24203)) ;
    mux21_ni ix21949 (.Y (nx21948), .A0 (inputs_446__5), .A1 (inputs_447__5), .S0 (
             nx24203)) ;
    mux21_ni ix22469 (.Y (nx22468), .A0 (nx22256), .A1 (nx22464), .S0 (nx22573)
             ) ;
    mux21_ni ix22257 (.Y (nx22256), .A0 (nx22250), .A1 (nx22172), .S0 (nx23141)
             ) ;
    oai21 ix22251 (.Y (nx22250), .A0 (nx22277), .A1 (nx12909), .B0 (nx12921)) ;
    mux21 ix12910 (.Y (nx12909), .A0 (nx22214), .A1 (nx22242), .S0 (nx22819)) ;
    mux21_ni ix22215 (.Y (nx22214), .A0 (nx22198), .A1 (nx22210), .S0 (nx23535)
             ) ;
    mux21_ni ix22199 (.Y (nx22198), .A0 (inputs_452__5), .A1 (inputs_453__5), .S0 (
             nx24203)) ;
    mux21_ni ix22211 (.Y (nx22210), .A0 (inputs_454__5), .A1 (inputs_455__5), .S0 (
             nx24203)) ;
    mux21_ni ix22243 (.Y (nx22242), .A0 (nx22226), .A1 (nx22238), .S0 (nx23535)
             ) ;
    mux21_ni ix22227 (.Y (nx22226), .A0 (inputs_468__5), .A1 (inputs_469__5), .S0 (
             nx24203)) ;
    mux21_ni ix22239 (.Y (nx22238), .A0 (inputs_470__5), .A1 (inputs_471__5), .S0 (
             nx24203)) ;
    nand04 ix12922 (.Y (nx12921), .A0 (nx22277), .A1 (nx23535), .A2 (nx24205), .A3 (
           nx22186)) ;
    mux21_ni ix22187 (.Y (nx22186), .A0 (inputs_451__5), .A1 (inputs_467__5), .S0 (
             nx22819)) ;
    mux21_ni ix22173 (.Y (nx22172), .A0 (nx22108), .A1 (nx22168), .S0 (nx22819)
             ) ;
    mux21_ni ix22109 (.Y (nx22108), .A0 (nx22076), .A1 (nx22104), .S0 (nx23239)
             ) ;
    mux21_ni ix22077 (.Y (nx22076), .A0 (nx22060), .A1 (nx22072), .S0 (nx23535)
             ) ;
    mux21_ni ix22061 (.Y (nx22060), .A0 (inputs_456__5), .A1 (inputs_457__5), .S0 (
             nx24205)) ;
    mux21_ni ix22073 (.Y (nx22072), .A0 (inputs_458__5), .A1 (inputs_459__5), .S0 (
             nx24205)) ;
    mux21_ni ix22105 (.Y (nx22104), .A0 (nx22088), .A1 (nx22100), .S0 (nx23537)
             ) ;
    mux21_ni ix22089 (.Y (nx22088), .A0 (inputs_460__5), .A1 (inputs_461__5), .S0 (
             nx24205)) ;
    mux21_ni ix22101 (.Y (nx22100), .A0 (inputs_462__5), .A1 (inputs_463__5), .S0 (
             nx24205)) ;
    mux21_ni ix22169 (.Y (nx22168), .A0 (nx22136), .A1 (nx22164), .S0 (nx23239)
             ) ;
    mux21_ni ix22137 (.Y (nx22136), .A0 (nx22120), .A1 (nx22132), .S0 (nx23537)
             ) ;
    mux21_ni ix22121 (.Y (nx22120), .A0 (inputs_472__5), .A1 (inputs_473__5), .S0 (
             nx24205)) ;
    mux21_ni ix22133 (.Y (nx22132), .A0 (inputs_474__5), .A1 (inputs_475__5), .S0 (
             nx24205)) ;
    mux21_ni ix22165 (.Y (nx22164), .A0 (nx22148), .A1 (nx22160), .S0 (nx23537)
             ) ;
    mux21_ni ix22149 (.Y (nx22148), .A0 (inputs_476__5), .A1 (inputs_477__5), .S0 (
             nx24207)) ;
    mux21_ni ix22161 (.Y (nx22160), .A0 (inputs_478__5), .A1 (inputs_479__5), .S0 (
             nx24207)) ;
    mux21_ni ix22465 (.Y (nx22464), .A0 (nx22458), .A1 (nx22380), .S0 (nx23141)
             ) ;
    oai21 ix22459 (.Y (nx22458), .A0 (nx22277), .A1 (nx12953), .B0 (nx12965)) ;
    mux21 ix12954 (.Y (nx12953), .A0 (nx22422), .A1 (nx22450), .S0 (nx22819)) ;
    mux21_ni ix22423 (.Y (nx22422), .A0 (nx22406), .A1 (nx22418), .S0 (nx23537)
             ) ;
    mux21_ni ix22407 (.Y (nx22406), .A0 (inputs_484__5), .A1 (inputs_485__5), .S0 (
             nx24207)) ;
    mux21_ni ix22419 (.Y (nx22418), .A0 (inputs_486__5), .A1 (inputs_487__5), .S0 (
             nx24207)) ;
    mux21_ni ix22451 (.Y (nx22450), .A0 (nx22434), .A1 (nx22446), .S0 (nx23537)
             ) ;
    mux21_ni ix22435 (.Y (nx22434), .A0 (inputs_500__5), .A1 (inputs_501__5), .S0 (
             nx24207)) ;
    mux21_ni ix22447 (.Y (nx22446), .A0 (inputs_502__5), .A1 (inputs_503__5), .S0 (
             nx24207)) ;
    nand04 ix12966 (.Y (nx12965), .A0 (nx22277), .A1 (nx23537), .A2 (nx24207), .A3 (
           nx22394)) ;
    mux21_ni ix22395 (.Y (nx22394), .A0 (inputs_483__5), .A1 (inputs_499__5), .S0 (
             nx22819)) ;
    mux21_ni ix22381 (.Y (nx22380), .A0 (nx22316), .A1 (nx22376), .S0 (nx22819)
             ) ;
    mux21_ni ix22317 (.Y (nx22316), .A0 (nx22284), .A1 (nx22312), .S0 (nx23239)
             ) ;
    mux21_ni ix22285 (.Y (nx22284), .A0 (nx22268), .A1 (nx22280), .S0 (nx23537)
             ) ;
    mux21_ni ix22269 (.Y (nx22268), .A0 (inputs_488__5), .A1 (inputs_489__5), .S0 (
             nx24209)) ;
    mux21_ni ix22281 (.Y (nx22280), .A0 (inputs_490__5), .A1 (inputs_491__5), .S0 (
             nx24209)) ;
    mux21_ni ix22313 (.Y (nx22312), .A0 (nx22296), .A1 (nx22308), .S0 (nx23539)
             ) ;
    mux21_ni ix22297 (.Y (nx22296), .A0 (inputs_492__5), .A1 (inputs_493__5), .S0 (
             nx24209)) ;
    mux21_ni ix22309 (.Y (nx22308), .A0 (inputs_494__5), .A1 (inputs_495__5), .S0 (
             nx24209)) ;
    mux21_ni ix22377 (.Y (nx22376), .A0 (nx22344), .A1 (nx22372), .S0 (nx23241)
             ) ;
    mux21_ni ix22345 (.Y (nx22344), .A0 (nx22328), .A1 (nx22340), .S0 (nx23539)
             ) ;
    mux21_ni ix22329 (.Y (nx22328), .A0 (inputs_504__5), .A1 (inputs_505__5), .S0 (
             nx24209)) ;
    mux21_ni ix22341 (.Y (nx22340), .A0 (inputs_506__5), .A1 (inputs_507__5), .S0 (
             nx24209)) ;
    mux21_ni ix22373 (.Y (nx22372), .A0 (nx22356), .A1 (nx22368), .S0 (nx23539)
             ) ;
    mux21_ni ix22357 (.Y (nx22356), .A0 (inputs_508__5), .A1 (inputs_509__5), .S0 (
             nx24209)) ;
    mux21_ni ix22369 (.Y (nx22368), .A0 (inputs_510__5), .A1 (inputs_511__5), .S0 (
             nx24211)) ;
    aoi32 ix12994 (.Y (nx12993), .A0 (nx23242), .A1 (nx22385), .A2 (nx22277), .B0 (
          nx22219), .B1 (nx24938)) ;
    oai21 ix23243 (.Y (nx23242), .A0 (nx23539), .A1 (nx12997), .B0 (nx13101)) ;
    mux21 ix12998 (.Y (nx12997), .A0 (nx22980), .A1 (nx23232), .S0 (nx24211)) ;
    mux21_ni ix22981 (.Y (nx22980), .A0 (nx22852), .A1 (nx22976), .S0 (nx22397)
             ) ;
    mux21_ni ix22853 (.Y (nx22852), .A0 (nx22788), .A1 (nx22848), .S0 (nx22421)
             ) ;
    mux21_ni ix22789 (.Y (nx22788), .A0 (nx22756), .A1 (nx22784), .S0 (nx22473)
             ) ;
    mux21_ni ix22757 (.Y (nx22756), .A0 (nx22740), .A1 (nx22752), .S0 (nx22573)
             ) ;
    mux21_ni ix22741 (.Y (nx22740), .A0 (inputs_0__5), .A1 (inputs_16__5), .S0 (
             nx22821)) ;
    mux21_ni ix22753 (.Y (nx22752), .A0 (inputs_32__5), .A1 (inputs_48__5), .S0 (
             nx22821)) ;
    mux21_ni ix22785 (.Y (nx22784), .A0 (nx22768), .A1 (nx22780), .S0 (nx22573)
             ) ;
    mux21_ni ix22769 (.Y (nx22768), .A0 (inputs_64__5), .A1 (inputs_80__5), .S0 (
             nx22821)) ;
    mux21_ni ix22781 (.Y (nx22780), .A0 (inputs_96__5), .A1 (inputs_112__5), .S0 (
             nx22821)) ;
    mux21_ni ix22849 (.Y (nx22848), .A0 (nx22816), .A1 (nx22844), .S0 (nx22473)
             ) ;
    mux21_ni ix22817 (.Y (nx22816), .A0 (nx22800), .A1 (nx22812), .S0 (nx22573)
             ) ;
    mux21_ni ix22801 (.Y (nx22800), .A0 (inputs_128__5), .A1 (inputs_144__5), .S0 (
             nx22821)) ;
    mux21_ni ix22813 (.Y (nx22812), .A0 (inputs_160__5), .A1 (inputs_176__5), .S0 (
             nx22821)) ;
    mux21_ni ix22845 (.Y (nx22844), .A0 (nx22828), .A1 (nx22840), .S0 (nx22573)
             ) ;
    mux21_ni ix22829 (.Y (nx22828), .A0 (inputs_192__5), .A1 (inputs_208__5), .S0 (
             nx22821)) ;
    mux21_ni ix22841 (.Y (nx22840), .A0 (inputs_224__5), .A1 (inputs_240__5), .S0 (
             nx22823)) ;
    mux21_ni ix22977 (.Y (nx22976), .A0 (nx22912), .A1 (nx22972), .S0 (nx22423)
             ) ;
    mux21_ni ix22913 (.Y (nx22912), .A0 (nx22880), .A1 (nx22908), .S0 (nx22475)
             ) ;
    mux21_ni ix22881 (.Y (nx22880), .A0 (nx22864), .A1 (nx22876), .S0 (nx22575)
             ) ;
    mux21_ni ix22865 (.Y (nx22864), .A0 (inputs_256__5), .A1 (inputs_272__5), .S0 (
             nx22823)) ;
    mux21_ni ix22877 (.Y (nx22876), .A0 (inputs_288__5), .A1 (inputs_304__5), .S0 (
             nx22823)) ;
    mux21_ni ix22909 (.Y (nx22908), .A0 (nx22892), .A1 (nx22904), .S0 (nx22575)
             ) ;
    mux21_ni ix22893 (.Y (nx22892), .A0 (inputs_320__5), .A1 (inputs_336__5), .S0 (
             nx22823)) ;
    mux21_ni ix22905 (.Y (nx22904), .A0 (inputs_352__5), .A1 (inputs_368__5), .S0 (
             nx22823)) ;
    mux21_ni ix22973 (.Y (nx22972), .A0 (nx22940), .A1 (nx22968), .S0 (nx22475)
             ) ;
    mux21_ni ix22941 (.Y (nx22940), .A0 (nx22924), .A1 (nx22936), .S0 (nx22575)
             ) ;
    mux21_ni ix22925 (.Y (nx22924), .A0 (inputs_384__5), .A1 (inputs_400__5), .S0 (
             nx22823)) ;
    mux21_ni ix22937 (.Y (nx22936), .A0 (inputs_416__5), .A1 (inputs_432__5), .S0 (
             nx22823)) ;
    mux21_ni ix22969 (.Y (nx22968), .A0 (nx22952), .A1 (nx22964), .S0 (nx22575)
             ) ;
    mux21_ni ix22953 (.Y (nx22952), .A0 (inputs_448__5), .A1 (inputs_464__5), .S0 (
             nx22825)) ;
    mux21_ni ix22965 (.Y (nx22964), .A0 (inputs_480__5), .A1 (inputs_496__5), .S0 (
             nx22825)) ;
    mux21_ni ix23233 (.Y (nx23232), .A0 (nx23104), .A1 (nx23228), .S0 (nx22397)
             ) ;
    mux21_ni ix23105 (.Y (nx23104), .A0 (nx23040), .A1 (nx23100), .S0 (nx22423)
             ) ;
    mux21_ni ix23041 (.Y (nx23040), .A0 (nx23008), .A1 (nx23036), .S0 (nx22475)
             ) ;
    mux21_ni ix23009 (.Y (nx23008), .A0 (nx22992), .A1 (nx23004), .S0 (nx22575)
             ) ;
    mux21_ni ix22993 (.Y (nx22992), .A0 (inputs_1__5), .A1 (inputs_17__5), .S0 (
             nx22825)) ;
    mux21_ni ix23005 (.Y (nx23004), .A0 (inputs_33__5), .A1 (inputs_49__5), .S0 (
             nx22825)) ;
    mux21_ni ix23037 (.Y (nx23036), .A0 (nx23020), .A1 (nx23032), .S0 (nx22575)
             ) ;
    mux21_ni ix23021 (.Y (nx23020), .A0 (inputs_65__5), .A1 (inputs_81__5), .S0 (
             nx22825)) ;
    mux21_ni ix23033 (.Y (nx23032), .A0 (inputs_97__5), .A1 (inputs_113__5), .S0 (
             nx22825)) ;
    mux21_ni ix23101 (.Y (nx23100), .A0 (nx23068), .A1 (nx23096), .S0 (nx22475)
             ) ;
    mux21_ni ix23069 (.Y (nx23068), .A0 (nx23052), .A1 (nx23064), .S0 (nx22575)
             ) ;
    mux21_ni ix23053 (.Y (nx23052), .A0 (inputs_129__5), .A1 (inputs_145__5), .S0 (
             nx22825)) ;
    mux21_ni ix23065 (.Y (nx23064), .A0 (inputs_161__5), .A1 (inputs_177__5), .S0 (
             nx22827)) ;
    mux21_ni ix23097 (.Y (nx23096), .A0 (nx23080), .A1 (nx23092), .S0 (nx22577)
             ) ;
    mux21_ni ix23081 (.Y (nx23080), .A0 (inputs_193__5), .A1 (inputs_209__5), .S0 (
             nx22827)) ;
    mux21_ni ix23093 (.Y (nx23092), .A0 (inputs_225__5), .A1 (inputs_241__5), .S0 (
             nx22827)) ;
    mux21_ni ix23229 (.Y (nx23228), .A0 (nx23164), .A1 (nx23224), .S0 (nx22423)
             ) ;
    mux21_ni ix23165 (.Y (nx23164), .A0 (nx23132), .A1 (nx23160), .S0 (nx22475)
             ) ;
    mux21_ni ix23133 (.Y (nx23132), .A0 (nx23116), .A1 (nx23128), .S0 (nx22577)
             ) ;
    mux21_ni ix23117 (.Y (nx23116), .A0 (inputs_257__5), .A1 (inputs_273__5), .S0 (
             nx22827)) ;
    mux21_ni ix23129 (.Y (nx23128), .A0 (inputs_289__5), .A1 (inputs_305__5), .S0 (
             nx22827)) ;
    mux21_ni ix23161 (.Y (nx23160), .A0 (nx23144), .A1 (nx23156), .S0 (nx22577)
             ) ;
    mux21_ni ix23145 (.Y (nx23144), .A0 (inputs_321__5), .A1 (inputs_337__5), .S0 (
             nx22827)) ;
    mux21_ni ix23157 (.Y (nx23156), .A0 (inputs_353__5), .A1 (inputs_369__5), .S0 (
             nx22827)) ;
    mux21_ni ix23225 (.Y (nx23224), .A0 (nx23192), .A1 (nx23220), .S0 (nx22475)
             ) ;
    mux21_ni ix23193 (.Y (nx23192), .A0 (nx23176), .A1 (nx23188), .S0 (nx22577)
             ) ;
    mux21_ni ix23177 (.Y (nx23176), .A0 (inputs_385__5), .A1 (inputs_401__5), .S0 (
             nx22829)) ;
    mux21_ni ix23189 (.Y (nx23188), .A0 (inputs_417__5), .A1 (inputs_433__5), .S0 (
             nx22829)) ;
    mux21_ni ix23221 (.Y (nx23220), .A0 (nx23204), .A1 (nx23216), .S0 (nx22577)
             ) ;
    mux21_ni ix23205 (.Y (nx23204), .A0 (inputs_449__5), .A1 (inputs_465__5), .S0 (
             nx22829)) ;
    mux21_ni ix23217 (.Y (nx23216), .A0 (inputs_481__5), .A1 (inputs_497__5), .S0 (
             nx22829)) ;
    nand03 ix13102 (.Y (nx13101), .A0 (nx22726), .A1 (nx23539), .A2 (nx24879)) ;
    mux21_ni ix22727 (.Y (nx22726), .A0 (nx22598), .A1 (nx22722), .S0 (nx22397)
             ) ;
    mux21_ni ix22599 (.Y (nx22598), .A0 (nx22534), .A1 (nx22594), .S0 (nx22423)
             ) ;
    mux21_ni ix22535 (.Y (nx22534), .A0 (nx22502), .A1 (nx22530), .S0 (nx22475)
             ) ;
    mux21_ni ix22503 (.Y (nx22502), .A0 (nx22486), .A1 (nx22498), .S0 (nx22577)
             ) ;
    mux21_ni ix22487 (.Y (nx22486), .A0 (inputs_2__5), .A1 (inputs_18__5), .S0 (
             nx22829)) ;
    mux21_ni ix22499 (.Y (nx22498), .A0 (inputs_34__5), .A1 (inputs_50__5), .S0 (
             nx22829)) ;
    mux21_ni ix22531 (.Y (nx22530), .A0 (nx22514), .A1 (nx22526), .S0 (nx22577)
             ) ;
    mux21_ni ix22515 (.Y (nx22514), .A0 (inputs_66__5), .A1 (inputs_82__5), .S0 (
             nx22829)) ;
    mux21_ni ix22527 (.Y (nx22526), .A0 (inputs_98__5), .A1 (inputs_114__5), .S0 (
             nx22831)) ;
    mux21_ni ix22595 (.Y (nx22594), .A0 (nx22562), .A1 (nx22590), .S0 (nx22477)
             ) ;
    mux21_ni ix22563 (.Y (nx22562), .A0 (nx22546), .A1 (nx22558), .S0 (nx22579)
             ) ;
    mux21_ni ix22547 (.Y (nx22546), .A0 (inputs_130__5), .A1 (inputs_146__5), .S0 (
             nx22831)) ;
    mux21_ni ix22559 (.Y (nx22558), .A0 (inputs_162__5), .A1 (inputs_178__5), .S0 (
             nx22831)) ;
    mux21_ni ix22591 (.Y (nx22590), .A0 (nx22574), .A1 (nx22586), .S0 (nx22579)
             ) ;
    mux21_ni ix22575 (.Y (nx22574), .A0 (inputs_194__5), .A1 (inputs_210__5), .S0 (
             nx22831)) ;
    mux21_ni ix22587 (.Y (nx22586), .A0 (inputs_226__5), .A1 (inputs_242__5), .S0 (
             nx22831)) ;
    mux21_ni ix22723 (.Y (nx22722), .A0 (nx22658), .A1 (nx22718), .S0 (nx22423)
             ) ;
    mux21_ni ix22659 (.Y (nx22658), .A0 (nx22626), .A1 (nx22654), .S0 (nx22477)
             ) ;
    mux21_ni ix22627 (.Y (nx22626), .A0 (nx22610), .A1 (nx22622), .S0 (nx22579)
             ) ;
    mux21_ni ix22611 (.Y (nx22610), .A0 (inputs_258__5), .A1 (inputs_274__5), .S0 (
             nx22831)) ;
    mux21_ni ix22623 (.Y (nx22622), .A0 (inputs_290__5), .A1 (inputs_306__5), .S0 (
             nx22831)) ;
    mux21_ni ix22655 (.Y (nx22654), .A0 (nx22638), .A1 (nx22650), .S0 (nx22579)
             ) ;
    mux21_ni ix22639 (.Y (nx22638), .A0 (inputs_322__5), .A1 (inputs_338__5), .S0 (
             nx22833)) ;
    mux21_ni ix22651 (.Y (nx22650), .A0 (inputs_354__5), .A1 (inputs_370__5), .S0 (
             nx22833)) ;
    mux21_ni ix22719 (.Y (nx22718), .A0 (nx22686), .A1 (nx22714), .S0 (nx22477)
             ) ;
    mux21_ni ix22687 (.Y (nx22686), .A0 (nx22670), .A1 (nx22682), .S0 (nx22579)
             ) ;
    mux21_ni ix22671 (.Y (nx22670), .A0 (inputs_386__5), .A1 (inputs_402__5), .S0 (
             nx22833)) ;
    mux21_ni ix22683 (.Y (nx22682), .A0 (inputs_418__5), .A1 (inputs_434__5), .S0 (
             nx22833)) ;
    mux21_ni ix22715 (.Y (nx22714), .A0 (nx22698), .A1 (nx22710), .S0 (nx22579)
             ) ;
    mux21_ni ix22699 (.Y (nx22698), .A0 (inputs_450__5), .A1 (inputs_466__5), .S0 (
             nx22833)) ;
    mux21_ni ix22711 (.Y (nx22710), .A0 (inputs_482__5), .A1 (inputs_498__5), .S0 (
             nx22833)) ;
    mux21_ni ix24939 (.Y (nx24938), .A0 (nx24090), .A1 (nx24934), .S0 (nx22423)
             ) ;
    mux21_ni ix24091 (.Y (nx24090), .A0 (nx23666), .A1 (nx24086), .S0 (nx22477)
             ) ;
    mux21_ni ix23667 (.Y (nx23666), .A0 (nx23454), .A1 (nx23662), .S0 (nx22579)
             ) ;
    mux21_ni ix23455 (.Y (nx23454), .A0 (nx23448), .A1 (nx23370), .S0 (nx23141)
             ) ;
    oai21 ix23449 (.Y (nx23448), .A0 (nx22279), .A1 (nx13161), .B0 (nx13173)) ;
    mux21 ix13162 (.Y (nx13161), .A0 (nx23412), .A1 (nx23440), .S0 (nx22833)) ;
    mux21_ni ix23413 (.Y (nx23412), .A0 (nx23396), .A1 (nx23408), .S0 (nx23539)
             ) ;
    mux21_ni ix23397 (.Y (nx23396), .A0 (inputs_4__5), .A1 (inputs_5__5), .S0 (
             nx24211)) ;
    mux21_ni ix23409 (.Y (nx23408), .A0 (inputs_6__5), .A1 (inputs_7__5), .S0 (
             nx24211)) ;
    mux21_ni ix23441 (.Y (nx23440), .A0 (nx23424), .A1 (nx23436), .S0 (nx23539)
             ) ;
    mux21_ni ix23425 (.Y (nx23424), .A0 (inputs_20__5), .A1 (inputs_21__5), .S0 (
             nx24211)) ;
    mux21_ni ix23437 (.Y (nx23436), .A0 (inputs_22__5), .A1 (inputs_23__5), .S0 (
             nx24211)) ;
    nand04 ix13174 (.Y (nx13173), .A0 (nx22279), .A1 (nx23541), .A2 (nx24211), .A3 (
           nx23384)) ;
    mux21_ni ix23385 (.Y (nx23384), .A0 (inputs_3__5), .A1 (inputs_19__5), .S0 (
             nx22835)) ;
    mux21_ni ix23371 (.Y (nx23370), .A0 (nx23306), .A1 (nx23366), .S0 (nx22835)
             ) ;
    mux21_ni ix23307 (.Y (nx23306), .A0 (nx23274), .A1 (nx23302), .S0 (nx23241)
             ) ;
    mux21_ni ix23275 (.Y (nx23274), .A0 (nx23258), .A1 (nx23270), .S0 (nx23541)
             ) ;
    mux21_ni ix23259 (.Y (nx23258), .A0 (inputs_8__5), .A1 (inputs_9__5), .S0 (
             nx24213)) ;
    mux21_ni ix23271 (.Y (nx23270), .A0 (inputs_10__5), .A1 (inputs_11__5), .S0 (
             nx24213)) ;
    mux21_ni ix23303 (.Y (nx23302), .A0 (nx23286), .A1 (nx23298), .S0 (nx23541)
             ) ;
    mux21_ni ix23287 (.Y (nx23286), .A0 (inputs_12__5), .A1 (inputs_13__5), .S0 (
             nx24213)) ;
    mux21_ni ix23299 (.Y (nx23298), .A0 (inputs_14__5), .A1 (inputs_15__5), .S0 (
             nx24213)) ;
    mux21_ni ix23367 (.Y (nx23366), .A0 (nx23334), .A1 (nx23362), .S0 (nx23241)
             ) ;
    mux21_ni ix23335 (.Y (nx23334), .A0 (nx23318), .A1 (nx23330), .S0 (nx23541)
             ) ;
    mux21_ni ix23319 (.Y (nx23318), .A0 (inputs_24__5), .A1 (inputs_25__5), .S0 (
             nx24213)) ;
    mux21_ni ix23331 (.Y (nx23330), .A0 (inputs_26__5), .A1 (inputs_27__5), .S0 (
             nx24213)) ;
    mux21_ni ix23363 (.Y (nx23362), .A0 (nx23346), .A1 (nx23358), .S0 (nx23541)
             ) ;
    mux21_ni ix23347 (.Y (nx23346), .A0 (inputs_28__5), .A1 (inputs_29__5), .S0 (
             nx24213)) ;
    mux21_ni ix23359 (.Y (nx23358), .A0 (inputs_30__5), .A1 (inputs_31__5), .S0 (
             nx24215)) ;
    mux21_ni ix23663 (.Y (nx23662), .A0 (nx23656), .A1 (nx23578), .S0 (nx23141)
             ) ;
    oai21 ix23657 (.Y (nx23656), .A0 (nx22279), .A1 (nx13203), .B0 (nx13217)) ;
    mux21 ix13204 (.Y (nx13203), .A0 (nx23620), .A1 (nx23648), .S0 (nx22835)) ;
    mux21_ni ix23621 (.Y (nx23620), .A0 (nx23604), .A1 (nx23616), .S0 (nx23541)
             ) ;
    mux21_ni ix23605 (.Y (nx23604), .A0 (inputs_36__5), .A1 (inputs_37__5), .S0 (
             nx24215)) ;
    mux21_ni ix23617 (.Y (nx23616), .A0 (inputs_38__5), .A1 (inputs_39__5), .S0 (
             nx24215)) ;
    mux21_ni ix23649 (.Y (nx23648), .A0 (nx23632), .A1 (nx23644), .S0 (nx23541)
             ) ;
    mux21_ni ix23633 (.Y (nx23632), .A0 (inputs_52__5), .A1 (inputs_53__5), .S0 (
             nx24215)) ;
    mux21_ni ix23645 (.Y (nx23644), .A0 (inputs_54__5), .A1 (inputs_55__5), .S0 (
             nx24215)) ;
    nand04 ix13218 (.Y (nx13217), .A0 (nx22279), .A1 (nx23543), .A2 (nx24215), .A3 (
           nx23592)) ;
    mux21_ni ix23593 (.Y (nx23592), .A0 (inputs_35__5), .A1 (inputs_51__5), .S0 (
             nx22835)) ;
    mux21_ni ix23579 (.Y (nx23578), .A0 (nx23514), .A1 (nx23574), .S0 (nx22835)
             ) ;
    mux21_ni ix23515 (.Y (nx23514), .A0 (nx23482), .A1 (nx23510), .S0 (nx23241)
             ) ;
    mux21_ni ix23483 (.Y (nx23482), .A0 (nx23466), .A1 (nx23478), .S0 (nx23543)
             ) ;
    mux21_ni ix23467 (.Y (nx23466), .A0 (inputs_40__5), .A1 (inputs_41__5), .S0 (
             nx24215)) ;
    mux21_ni ix23479 (.Y (nx23478), .A0 (inputs_42__5), .A1 (inputs_43__5), .S0 (
             nx24217)) ;
    mux21_ni ix23511 (.Y (nx23510), .A0 (nx23494), .A1 (nx23506), .S0 (nx23543)
             ) ;
    mux21_ni ix23495 (.Y (nx23494), .A0 (inputs_44__5), .A1 (inputs_45__5), .S0 (
             nx24217)) ;
    mux21_ni ix23507 (.Y (nx23506), .A0 (inputs_46__5), .A1 (inputs_47__5), .S0 (
             nx24217)) ;
    mux21_ni ix23575 (.Y (nx23574), .A0 (nx23542), .A1 (nx23570), .S0 (nx23241)
             ) ;
    mux21_ni ix23543 (.Y (nx23542), .A0 (nx23526), .A1 (nx23538), .S0 (nx23543)
             ) ;
    mux21_ni ix23527 (.Y (nx23526), .A0 (inputs_56__5), .A1 (inputs_57__5), .S0 (
             nx24217)) ;
    mux21_ni ix23539 (.Y (nx23538), .A0 (inputs_58__5), .A1 (inputs_59__5), .S0 (
             nx24217)) ;
    mux21_ni ix23571 (.Y (nx23570), .A0 (nx23554), .A1 (nx23566), .S0 (nx23543)
             ) ;
    mux21_ni ix23555 (.Y (nx23554), .A0 (inputs_60__5), .A1 (inputs_61__5), .S0 (
             nx24217)) ;
    mux21_ni ix23567 (.Y (nx23566), .A0 (inputs_62__5), .A1 (inputs_63__5), .S0 (
             nx24217)) ;
    mux21_ni ix24087 (.Y (nx24086), .A0 (nx23874), .A1 (nx24082), .S0 (nx22581)
             ) ;
    mux21_ni ix23875 (.Y (nx23874), .A0 (nx23868), .A1 (nx23790), .S0 (nx23141)
             ) ;
    oai21 ix23869 (.Y (nx23868), .A0 (nx22279), .A1 (nx13251), .B0 (nx13263)) ;
    mux21 ix13252 (.Y (nx13251), .A0 (nx23832), .A1 (nx23860), .S0 (nx22835)) ;
    mux21_ni ix23833 (.Y (nx23832), .A0 (nx23816), .A1 (nx23828), .S0 (nx23543)
             ) ;
    mux21_ni ix23817 (.Y (nx23816), .A0 (inputs_68__5), .A1 (inputs_69__5), .S0 (
             nx24219)) ;
    mux21_ni ix23829 (.Y (nx23828), .A0 (inputs_70__5), .A1 (inputs_71__5), .S0 (
             nx24219)) ;
    mux21_ni ix23861 (.Y (nx23860), .A0 (nx23844), .A1 (nx23856), .S0 (nx23543)
             ) ;
    mux21_ni ix23845 (.Y (nx23844), .A0 (inputs_84__5), .A1 (inputs_85__5), .S0 (
             nx24219)) ;
    mux21_ni ix23857 (.Y (nx23856), .A0 (inputs_86__5), .A1 (inputs_87__5), .S0 (
             nx24219)) ;
    nand04 ix13264 (.Y (nx13263), .A0 (nx22279), .A1 (nx23545), .A2 (nx24219), .A3 (
           nx23804)) ;
    mux21_ni ix23805 (.Y (nx23804), .A0 (inputs_67__5), .A1 (inputs_83__5), .S0 (
             nx22835)) ;
    mux21_ni ix23791 (.Y (nx23790), .A0 (nx23726), .A1 (nx23786), .S0 (nx22837)
             ) ;
    mux21_ni ix23727 (.Y (nx23726), .A0 (nx23694), .A1 (nx23722), .S0 (nx23241)
             ) ;
    mux21_ni ix23695 (.Y (nx23694), .A0 (nx23678), .A1 (nx23690), .S0 (nx23545)
             ) ;
    mux21_ni ix23679 (.Y (nx23678), .A0 (inputs_72__5), .A1 (inputs_73__5), .S0 (
             nx24219)) ;
    mux21_ni ix23691 (.Y (nx23690), .A0 (inputs_74__5), .A1 (inputs_75__5), .S0 (
             nx24219)) ;
    mux21_ni ix23723 (.Y (nx23722), .A0 (nx23706), .A1 (nx23718), .S0 (nx23545)
             ) ;
    mux21_ni ix23707 (.Y (nx23706), .A0 (inputs_76__5), .A1 (inputs_77__5), .S0 (
             nx24221)) ;
    mux21_ni ix23719 (.Y (nx23718), .A0 (inputs_78__5), .A1 (inputs_79__5), .S0 (
             nx24221)) ;
    mux21_ni ix23787 (.Y (nx23786), .A0 (nx23754), .A1 (nx23782), .S0 (nx23241)
             ) ;
    mux21_ni ix23755 (.Y (nx23754), .A0 (nx23738), .A1 (nx23750), .S0 (nx23545)
             ) ;
    mux21_ni ix23739 (.Y (nx23738), .A0 (inputs_88__5), .A1 (inputs_89__5), .S0 (
             nx24221)) ;
    mux21_ni ix23751 (.Y (nx23750), .A0 (inputs_90__5), .A1 (inputs_91__5), .S0 (
             nx24221)) ;
    mux21_ni ix23783 (.Y (nx23782), .A0 (nx23766), .A1 (nx23778), .S0 (nx23545)
             ) ;
    mux21_ni ix23767 (.Y (nx23766), .A0 (inputs_92__5), .A1 (inputs_93__5), .S0 (
             nx24221)) ;
    mux21_ni ix23779 (.Y (nx23778), .A0 (inputs_94__5), .A1 (inputs_95__5), .S0 (
             nx24221)) ;
    mux21_ni ix24083 (.Y (nx24082), .A0 (nx24076), .A1 (nx23998), .S0 (nx23143)
             ) ;
    oai21 ix24077 (.Y (nx24076), .A0 (nx22279), .A1 (nx13293), .B0 (nx13305)) ;
    mux21 ix13294 (.Y (nx13293), .A0 (nx24040), .A1 (nx24068), .S0 (nx22837)) ;
    mux21_ni ix24041 (.Y (nx24040), .A0 (nx24024), .A1 (nx24036), .S0 (nx23545)
             ) ;
    mux21_ni ix24025 (.Y (nx24024), .A0 (inputs_100__5), .A1 (inputs_101__5), .S0 (
             nx24221)) ;
    mux21_ni ix24037 (.Y (nx24036), .A0 (inputs_102__5), .A1 (inputs_103__5), .S0 (
             nx24223)) ;
    mux21_ni ix24069 (.Y (nx24068), .A0 (nx24052), .A1 (nx24064), .S0 (nx23545)
             ) ;
    mux21_ni ix24053 (.Y (nx24052), .A0 (inputs_116__5), .A1 (inputs_117__5), .S0 (
             nx24223)) ;
    mux21_ni ix24065 (.Y (nx24064), .A0 (inputs_118__5), .A1 (inputs_119__5), .S0 (
             nx24223)) ;
    nand04 ix13306 (.Y (nx13305), .A0 (nx22281), .A1 (nx23547), .A2 (nx24223), .A3 (
           nx24012)) ;
    mux21_ni ix24013 (.Y (nx24012), .A0 (inputs_99__5), .A1 (inputs_115__5), .S0 (
             nx22837)) ;
    mux21_ni ix23999 (.Y (nx23998), .A0 (nx23934), .A1 (nx23994), .S0 (nx22837)
             ) ;
    mux21_ni ix23935 (.Y (nx23934), .A0 (nx23902), .A1 (nx23930), .S0 (nx23243)
             ) ;
    mux21_ni ix23903 (.Y (nx23902), .A0 (nx23886), .A1 (nx23898), .S0 (nx23547)
             ) ;
    mux21_ni ix23887 (.Y (nx23886), .A0 (inputs_104__5), .A1 (inputs_105__5), .S0 (
             nx24223)) ;
    mux21_ni ix23899 (.Y (nx23898), .A0 (inputs_106__5), .A1 (inputs_107__5), .S0 (
             nx24223)) ;
    mux21_ni ix23931 (.Y (nx23930), .A0 (nx23914), .A1 (nx23926), .S0 (nx23547)
             ) ;
    mux21_ni ix23915 (.Y (nx23914), .A0 (inputs_108__5), .A1 (inputs_109__5), .S0 (
             nx24223)) ;
    mux21_ni ix23927 (.Y (nx23926), .A0 (inputs_110__5), .A1 (inputs_111__5), .S0 (
             nx24225)) ;
    mux21_ni ix23995 (.Y (nx23994), .A0 (nx23962), .A1 (nx23990), .S0 (nx23243)
             ) ;
    mux21_ni ix23963 (.Y (nx23962), .A0 (nx23946), .A1 (nx23958), .S0 (nx23547)
             ) ;
    mux21_ni ix23947 (.Y (nx23946), .A0 (inputs_120__5), .A1 (inputs_121__5), .S0 (
             nx24225)) ;
    mux21_ni ix23959 (.Y (nx23958), .A0 (inputs_122__5), .A1 (inputs_123__5), .S0 (
             nx24225)) ;
    mux21_ni ix23991 (.Y (nx23990), .A0 (nx23974), .A1 (nx23986), .S0 (nx23547)
             ) ;
    mux21_ni ix23975 (.Y (nx23974), .A0 (inputs_124__5), .A1 (inputs_125__5), .S0 (
             nx24225)) ;
    mux21_ni ix23987 (.Y (nx23986), .A0 (inputs_126__5), .A1 (inputs_127__5), .S0 (
             nx24225)) ;
    mux21_ni ix24935 (.Y (nx24934), .A0 (nx24510), .A1 (nx24930), .S0 (nx22477)
             ) ;
    mux21_ni ix24511 (.Y (nx24510), .A0 (nx24298), .A1 (nx24506), .S0 (nx22581)
             ) ;
    mux21_ni ix24299 (.Y (nx24298), .A0 (nx24292), .A1 (nx24214), .S0 (nx23143)
             ) ;
    oai21 ix24293 (.Y (nx24292), .A0 (nx22281), .A1 (nx13339), .B0 (nx13349)) ;
    mux21 ix13340 (.Y (nx13339), .A0 (nx24256), .A1 (nx24284), .S0 (nx22837)) ;
    mux21_ni ix24257 (.Y (nx24256), .A0 (nx24240), .A1 (nx24252), .S0 (nx23547)
             ) ;
    mux21_ni ix24241 (.Y (nx24240), .A0 (inputs_132__5), .A1 (inputs_133__5), .S0 (
             nx24225)) ;
    mux21_ni ix24253 (.Y (nx24252), .A0 (inputs_134__5), .A1 (inputs_135__5), .S0 (
             nx24225)) ;
    mux21_ni ix24285 (.Y (nx24284), .A0 (nx24268), .A1 (nx24280), .S0 (nx23547)
             ) ;
    mux21_ni ix24269 (.Y (nx24268), .A0 (inputs_148__5), .A1 (inputs_149__5), .S0 (
             nx24227)) ;
    mux21_ni ix24281 (.Y (nx24280), .A0 (inputs_150__5), .A1 (inputs_151__5), .S0 (
             nx24227)) ;
    nand04 ix13350 (.Y (nx13349), .A0 (nx22281), .A1 (nx23549), .A2 (nx24227), .A3 (
           nx24228)) ;
    mux21_ni ix24229 (.Y (nx24228), .A0 (inputs_131__5), .A1 (inputs_147__5), .S0 (
             nx22837)) ;
    mux21_ni ix24215 (.Y (nx24214), .A0 (nx24150), .A1 (nx24210), .S0 (nx22837)
             ) ;
    mux21_ni ix24151 (.Y (nx24150), .A0 (nx24118), .A1 (nx24146), .S0 (nx23243)
             ) ;
    mux21_ni ix24119 (.Y (nx24118), .A0 (nx24102), .A1 (nx24114), .S0 (nx23549)
             ) ;
    mux21_ni ix24103 (.Y (nx24102), .A0 (inputs_136__5), .A1 (inputs_137__5), .S0 (
             nx24227)) ;
    mux21_ni ix24115 (.Y (nx24114), .A0 (inputs_138__5), .A1 (inputs_139__5), .S0 (
             nx24227)) ;
    mux21_ni ix24147 (.Y (nx24146), .A0 (nx24130), .A1 (nx24142), .S0 (nx23549)
             ) ;
    mux21_ni ix24131 (.Y (nx24130), .A0 (inputs_140__5), .A1 (inputs_141__5), .S0 (
             nx24227)) ;
    mux21_ni ix24143 (.Y (nx24142), .A0 (inputs_142__5), .A1 (inputs_143__5), .S0 (
             nx24227)) ;
    mux21_ni ix24211 (.Y (nx24210), .A0 (nx24178), .A1 (nx24206), .S0 (nx23243)
             ) ;
    mux21_ni ix24179 (.Y (nx24178), .A0 (nx24162), .A1 (nx24174), .S0 (nx23549)
             ) ;
    mux21_ni ix24163 (.Y (nx24162), .A0 (inputs_152__5), .A1 (inputs_153__5), .S0 (
             nx24229)) ;
    mux21_ni ix24175 (.Y (nx24174), .A0 (inputs_154__5), .A1 (inputs_155__5), .S0 (
             nx24229)) ;
    mux21_ni ix24207 (.Y (nx24206), .A0 (nx24190), .A1 (nx24202), .S0 (nx23549)
             ) ;
    mux21_ni ix24191 (.Y (nx24190), .A0 (inputs_156__5), .A1 (inputs_157__5), .S0 (
             nx24229)) ;
    mux21_ni ix24203 (.Y (nx24202), .A0 (inputs_158__5), .A1 (inputs_159__5), .S0 (
             nx24229)) ;
    mux21_ni ix24507 (.Y (nx24506), .A0 (nx24500), .A1 (nx24422), .S0 (nx23143)
             ) ;
    oai21 ix24501 (.Y (nx24500), .A0 (nx22281), .A1 (nx13381), .B0 (nx13393)) ;
    mux21 ix13382 (.Y (nx13381), .A0 (nx24464), .A1 (nx24492), .S0 (nx22839)) ;
    mux21_ni ix24465 (.Y (nx24464), .A0 (nx24448), .A1 (nx24460), .S0 (nx23549)
             ) ;
    mux21_ni ix24449 (.Y (nx24448), .A0 (inputs_164__5), .A1 (inputs_165__5), .S0 (
             nx24229)) ;
    mux21_ni ix24461 (.Y (nx24460), .A0 (inputs_166__5), .A1 (inputs_167__5), .S0 (
             nx24229)) ;
    mux21_ni ix24493 (.Y (nx24492), .A0 (nx24476), .A1 (nx24488), .S0 (nx23549)
             ) ;
    mux21_ni ix24477 (.Y (nx24476), .A0 (inputs_180__5), .A1 (inputs_181__5), .S0 (
             nx24229)) ;
    mux21_ni ix24489 (.Y (nx24488), .A0 (inputs_182__5), .A1 (inputs_183__5), .S0 (
             nx24231)) ;
    nand04 ix13394 (.Y (nx13393), .A0 (nx22281), .A1 (nx23551), .A2 (nx24231), .A3 (
           nx24436)) ;
    mux21_ni ix24437 (.Y (nx24436), .A0 (inputs_163__5), .A1 (inputs_179__5), .S0 (
             nx22839)) ;
    mux21_ni ix24423 (.Y (nx24422), .A0 (nx24358), .A1 (nx24418), .S0 (nx22839)
             ) ;
    mux21_ni ix24359 (.Y (nx24358), .A0 (nx24326), .A1 (nx24354), .S0 (nx23243)
             ) ;
    mux21_ni ix24327 (.Y (nx24326), .A0 (nx24310), .A1 (nx24322), .S0 (nx23551)
             ) ;
    mux21_ni ix24311 (.Y (nx24310), .A0 (inputs_168__5), .A1 (inputs_169__5), .S0 (
             nx24231)) ;
    mux21_ni ix24323 (.Y (nx24322), .A0 (inputs_170__5), .A1 (inputs_171__5), .S0 (
             nx24231)) ;
    mux21_ni ix24355 (.Y (nx24354), .A0 (nx24338), .A1 (nx24350), .S0 (nx23551)
             ) ;
    mux21_ni ix24339 (.Y (nx24338), .A0 (inputs_172__5), .A1 (inputs_173__5), .S0 (
             nx24231)) ;
    mux21_ni ix24351 (.Y (nx24350), .A0 (inputs_174__5), .A1 (inputs_175__5), .S0 (
             nx24231)) ;
    mux21_ni ix24419 (.Y (nx24418), .A0 (nx24386), .A1 (nx24414), .S0 (nx23243)
             ) ;
    mux21_ni ix24387 (.Y (nx24386), .A0 (nx24370), .A1 (nx24382), .S0 (nx23551)
             ) ;
    mux21_ni ix24371 (.Y (nx24370), .A0 (inputs_184__5), .A1 (inputs_185__5), .S0 (
             nx24231)) ;
    mux21_ni ix24383 (.Y (nx24382), .A0 (inputs_186__5), .A1 (inputs_187__5), .S0 (
             nx24233)) ;
    mux21_ni ix24415 (.Y (nx24414), .A0 (nx24398), .A1 (nx24410), .S0 (nx23551)
             ) ;
    mux21_ni ix24399 (.Y (nx24398), .A0 (inputs_188__5), .A1 (inputs_189__5), .S0 (
             nx24233)) ;
    mux21_ni ix24411 (.Y (nx24410), .A0 (inputs_190__5), .A1 (inputs_191__5), .S0 (
             nx24233)) ;
    mux21_ni ix24931 (.Y (nx24930), .A0 (nx24718), .A1 (nx24926), .S0 (nx22581)
             ) ;
    mux21_ni ix24719 (.Y (nx24718), .A0 (nx24712), .A1 (nx24634), .S0 (nx23143)
             ) ;
    oai21 ix24713 (.Y (nx24712), .A0 (nx22281), .A1 (nx13425), .B0 (nx13439)) ;
    mux21 ix13426 (.Y (nx13425), .A0 (nx24676), .A1 (nx24704), .S0 (nx22839)) ;
    mux21_ni ix24677 (.Y (nx24676), .A0 (nx24660), .A1 (nx24672), .S0 (nx23551)
             ) ;
    mux21_ni ix24661 (.Y (nx24660), .A0 (inputs_196__5), .A1 (inputs_197__5), .S0 (
             nx24233)) ;
    mux21_ni ix24673 (.Y (nx24672), .A0 (inputs_198__5), .A1 (inputs_199__5), .S0 (
             nx24233)) ;
    mux21_ni ix24705 (.Y (nx24704), .A0 (nx24688), .A1 (nx24700), .S0 (nx23551)
             ) ;
    mux21_ni ix24689 (.Y (nx24688), .A0 (inputs_212__5), .A1 (inputs_213__5), .S0 (
             nx24233)) ;
    mux21_ni ix24701 (.Y (nx24700), .A0 (inputs_214__5), .A1 (inputs_215__5), .S0 (
             nx24233)) ;
    nand04 ix13440 (.Y (nx13439), .A0 (nx22281), .A1 (nx23553), .A2 (nx24235), .A3 (
           nx24648)) ;
    mux21_ni ix24649 (.Y (nx24648), .A0 (inputs_195__5), .A1 (inputs_211__5), .S0 (
             nx22839)) ;
    mux21_ni ix24635 (.Y (nx24634), .A0 (nx24570), .A1 (nx24630), .S0 (nx22839)
             ) ;
    mux21_ni ix24571 (.Y (nx24570), .A0 (nx24538), .A1 (nx24566), .S0 (nx23243)
             ) ;
    mux21_ni ix24539 (.Y (nx24538), .A0 (nx24522), .A1 (nx24534), .S0 (nx23553)
             ) ;
    mux21_ni ix24523 (.Y (nx24522), .A0 (inputs_200__5), .A1 (inputs_201__5), .S0 (
             nx24235)) ;
    mux21_ni ix24535 (.Y (nx24534), .A0 (inputs_202__5), .A1 (inputs_203__5), .S0 (
             nx24235)) ;
    mux21_ni ix24567 (.Y (nx24566), .A0 (nx24550), .A1 (nx24562), .S0 (nx23553)
             ) ;
    mux21_ni ix24551 (.Y (nx24550), .A0 (inputs_204__5), .A1 (inputs_205__5), .S0 (
             nx24235)) ;
    mux21_ni ix24563 (.Y (nx24562), .A0 (inputs_206__5), .A1 (inputs_207__5), .S0 (
             nx24235)) ;
    mux21_ni ix24631 (.Y (nx24630), .A0 (nx24598), .A1 (nx24626), .S0 (nx23245)
             ) ;
    mux21_ni ix24599 (.Y (nx24598), .A0 (nx24582), .A1 (nx24594), .S0 (nx23553)
             ) ;
    mux21_ni ix24583 (.Y (nx24582), .A0 (inputs_216__5), .A1 (inputs_217__5), .S0 (
             nx24235)) ;
    mux21_ni ix24595 (.Y (nx24594), .A0 (inputs_218__5), .A1 (inputs_219__5), .S0 (
             nx24235)) ;
    mux21_ni ix24627 (.Y (nx24626), .A0 (nx24610), .A1 (nx24622), .S0 (nx23553)
             ) ;
    mux21_ni ix24611 (.Y (nx24610), .A0 (inputs_220__5), .A1 (inputs_221__5), .S0 (
             nx24237)) ;
    mux21_ni ix24623 (.Y (nx24622), .A0 (inputs_222__5), .A1 (inputs_223__5), .S0 (
             nx24237)) ;
    mux21_ni ix24927 (.Y (nx24926), .A0 (nx24920), .A1 (nx24842), .S0 (nx23143)
             ) ;
    oai21 ix24921 (.Y (nx24920), .A0 (nx22283), .A1 (nx13469), .B0 (nx13483)) ;
    mux21 ix13470 (.Y (nx13469), .A0 (nx24884), .A1 (nx24912), .S0 (nx22839)) ;
    mux21_ni ix24885 (.Y (nx24884), .A0 (nx24868), .A1 (nx24880), .S0 (nx23553)
             ) ;
    mux21_ni ix24869 (.Y (nx24868), .A0 (inputs_228__5), .A1 (inputs_229__5), .S0 (
             nx24237)) ;
    mux21_ni ix24881 (.Y (nx24880), .A0 (inputs_230__5), .A1 (inputs_231__5), .S0 (
             nx24237)) ;
    mux21_ni ix24913 (.Y (nx24912), .A0 (nx24896), .A1 (nx24908), .S0 (nx23553)
             ) ;
    mux21_ni ix24897 (.Y (nx24896), .A0 (inputs_244__5), .A1 (inputs_245__5), .S0 (
             nx24237)) ;
    mux21_ni ix24909 (.Y (nx24908), .A0 (inputs_246__5), .A1 (inputs_247__5), .S0 (
             nx24237)) ;
    nand04 ix13484 (.Y (nx13483), .A0 (nx22283), .A1 (nx23555), .A2 (nx24237), .A3 (
           nx24856)) ;
    mux21_ni ix24857 (.Y (nx24856), .A0 (inputs_227__5), .A1 (inputs_243__5), .S0 (
             nx22841)) ;
    mux21_ni ix24843 (.Y (nx24842), .A0 (nx24778), .A1 (nx24838), .S0 (nx22841)
             ) ;
    mux21_ni ix24779 (.Y (nx24778), .A0 (nx24746), .A1 (nx24774), .S0 (nx23245)
             ) ;
    mux21_ni ix24747 (.Y (nx24746), .A0 (nx24730), .A1 (nx24742), .S0 (nx23555)
             ) ;
    mux21_ni ix24731 (.Y (nx24730), .A0 (inputs_232__5), .A1 (inputs_233__5), .S0 (
             nx24239)) ;
    mux21_ni ix24743 (.Y (nx24742), .A0 (inputs_234__5), .A1 (inputs_235__5), .S0 (
             nx24239)) ;
    mux21_ni ix24775 (.Y (nx24774), .A0 (nx24758), .A1 (nx24770), .S0 (nx23555)
             ) ;
    mux21_ni ix24759 (.Y (nx24758), .A0 (inputs_236__5), .A1 (inputs_237__5), .S0 (
             nx24239)) ;
    mux21_ni ix24771 (.Y (nx24770), .A0 (inputs_238__5), .A1 (inputs_239__5), .S0 (
             nx24239)) ;
    mux21_ni ix24839 (.Y (nx24838), .A0 (nx24806), .A1 (nx24834), .S0 (nx23245)
             ) ;
    mux21_ni ix24807 (.Y (nx24806), .A0 (nx24790), .A1 (nx24802), .S0 (nx23555)
             ) ;
    mux21_ni ix24791 (.Y (nx24790), .A0 (inputs_248__5), .A1 (inputs_249__5), .S0 (
             nx24239)) ;
    mux21_ni ix24803 (.Y (nx24802), .A0 (inputs_250__5), .A1 (inputs_251__5), .S0 (
             nx24239)) ;
    mux21_ni ix24835 (.Y (nx24834), .A0 (nx24818), .A1 (nx24830), .S0 (nx23555)
             ) ;
    mux21_ni ix24819 (.Y (nx24818), .A0 (inputs_252__5), .A1 (inputs_253__5), .S0 (
             nx24239)) ;
    mux21_ni ix24831 (.Y (nx24830), .A0 (inputs_254__5), .A1 (inputs_255__5), .S0 (
             nx24241)) ;
    oai21 ix29105 (.Y (\output [6]), .A0 (nx22219), .A1 (nx13513), .B0 (nx13869)
          ) ;
    mux21 ix13514 (.Y (nx13513), .A0 (nx25786), .A1 (nx26630), .S0 (nx22423)) ;
    mux21_ni ix25787 (.Y (nx25786), .A0 (nx25362), .A1 (nx25782), .S0 (nx22477)
             ) ;
    mux21_ni ix25363 (.Y (nx25362), .A0 (nx25150), .A1 (nx25358), .S0 (nx22581)
             ) ;
    mux21_ni ix25151 (.Y (nx25150), .A0 (nx25144), .A1 (nx25066), .S0 (nx23143)
             ) ;
    oai21 ix25145 (.Y (nx25144), .A0 (nx22283), .A1 (nx13521), .B0 (nx13531)) ;
    mux21 ix13522 (.Y (nx13521), .A0 (nx25108), .A1 (nx25136), .S0 (nx22841)) ;
    mux21_ni ix25109 (.Y (nx25108), .A0 (nx25092), .A1 (nx25104), .S0 (nx23555)
             ) ;
    mux21_ni ix25093 (.Y (nx25092), .A0 (inputs_260__6), .A1 (inputs_261__6), .S0 (
             nx24241)) ;
    mux21_ni ix25105 (.Y (nx25104), .A0 (inputs_262__6), .A1 (inputs_263__6), .S0 (
             nx24241)) ;
    mux21_ni ix25137 (.Y (nx25136), .A0 (nx25120), .A1 (nx25132), .S0 (nx23555)
             ) ;
    mux21_ni ix25121 (.Y (nx25120), .A0 (inputs_276__6), .A1 (inputs_277__6), .S0 (
             nx24241)) ;
    mux21_ni ix25133 (.Y (nx25132), .A0 (inputs_278__6), .A1 (inputs_279__6), .S0 (
             nx24241)) ;
    nand04 ix13532 (.Y (nx13531), .A0 (nx22283), .A1 (nx23557), .A2 (nx24241), .A3 (
           nx25080)) ;
    mux21_ni ix25081 (.Y (nx25080), .A0 (inputs_259__6), .A1 (inputs_275__6), .S0 (
             nx22841)) ;
    mux21_ni ix25067 (.Y (nx25066), .A0 (nx25002), .A1 (nx25062), .S0 (nx22841)
             ) ;
    mux21_ni ix25003 (.Y (nx25002), .A0 (nx24970), .A1 (nx24998), .S0 (nx23245)
             ) ;
    mux21_ni ix24971 (.Y (nx24970), .A0 (nx24954), .A1 (nx24966), .S0 (nx23557)
             ) ;
    mux21_ni ix24955 (.Y (nx24954), .A0 (inputs_264__6), .A1 (inputs_265__6), .S0 (
             nx24241)) ;
    mux21_ni ix24967 (.Y (nx24966), .A0 (inputs_266__6), .A1 (inputs_267__6), .S0 (
             nx24243)) ;
    mux21_ni ix24999 (.Y (nx24998), .A0 (nx24982), .A1 (nx24994), .S0 (nx23557)
             ) ;
    mux21_ni ix24983 (.Y (nx24982), .A0 (inputs_268__6), .A1 (inputs_269__6), .S0 (
             nx24243)) ;
    mux21_ni ix24995 (.Y (nx24994), .A0 (inputs_270__6), .A1 (inputs_271__6), .S0 (
             nx24243)) ;
    mux21_ni ix25063 (.Y (nx25062), .A0 (nx25030), .A1 (nx25058), .S0 (nx23245)
             ) ;
    mux21_ni ix25031 (.Y (nx25030), .A0 (nx25014), .A1 (nx25026), .S0 (nx23557)
             ) ;
    mux21_ni ix25015 (.Y (nx25014), .A0 (inputs_280__6), .A1 (inputs_281__6), .S0 (
             nx24243)) ;
    mux21_ni ix25027 (.Y (nx25026), .A0 (inputs_282__6), .A1 (inputs_283__6), .S0 (
             nx24243)) ;
    mux21_ni ix25059 (.Y (nx25058), .A0 (nx25042), .A1 (nx25054), .S0 (nx23557)
             ) ;
    mux21_ni ix25043 (.Y (nx25042), .A0 (inputs_284__6), .A1 (inputs_285__6), .S0 (
             nx24243)) ;
    mux21_ni ix25055 (.Y (nx25054), .A0 (inputs_286__6), .A1 (inputs_287__6), .S0 (
             nx24243)) ;
    mux21_ni ix25359 (.Y (nx25358), .A0 (nx25352), .A1 (nx25274), .S0 (nx23143)
             ) ;
    oai21 ix25353 (.Y (nx25352), .A0 (nx22283), .A1 (nx13561), .B0 (nx13571)) ;
    mux21 ix13562 (.Y (nx13561), .A0 (nx25316), .A1 (nx25344), .S0 (nx22841)) ;
    mux21_ni ix25317 (.Y (nx25316), .A0 (nx25300), .A1 (nx25312), .S0 (nx23557)
             ) ;
    mux21_ni ix25301 (.Y (nx25300), .A0 (inputs_292__6), .A1 (inputs_293__6), .S0 (
             nx24245)) ;
    mux21_ni ix25313 (.Y (nx25312), .A0 (inputs_294__6), .A1 (inputs_295__6), .S0 (
             nx24245)) ;
    mux21_ni ix25345 (.Y (nx25344), .A0 (nx25328), .A1 (nx25340), .S0 (nx23557)
             ) ;
    mux21_ni ix25329 (.Y (nx25328), .A0 (inputs_308__6), .A1 (inputs_309__6), .S0 (
             nx24245)) ;
    mux21_ni ix25341 (.Y (nx25340), .A0 (inputs_310__6), .A1 (inputs_311__6), .S0 (
             nx24245)) ;
    nand04 ix13572 (.Y (nx13571), .A0 (nx22283), .A1 (nx23559), .A2 (nx24245), .A3 (
           nx25288)) ;
    mux21_ni ix25289 (.Y (nx25288), .A0 (inputs_291__6), .A1 (inputs_307__6), .S0 (
             nx22841)) ;
    mux21_ni ix25275 (.Y (nx25274), .A0 (nx25210), .A1 (nx25270), .S0 (nx22843)
             ) ;
    mux21_ni ix25211 (.Y (nx25210), .A0 (nx25178), .A1 (nx25206), .S0 (nx23245)
             ) ;
    mux21_ni ix25179 (.Y (nx25178), .A0 (nx25162), .A1 (nx25174), .S0 (nx23559)
             ) ;
    mux21_ni ix25163 (.Y (nx25162), .A0 (inputs_296__6), .A1 (inputs_297__6), .S0 (
             nx24245)) ;
    mux21_ni ix25175 (.Y (nx25174), .A0 (inputs_298__6), .A1 (inputs_299__6), .S0 (
             nx24245)) ;
    mux21_ni ix25207 (.Y (nx25206), .A0 (nx25190), .A1 (nx25202), .S0 (nx23559)
             ) ;
    mux21_ni ix25191 (.Y (nx25190), .A0 (inputs_300__6), .A1 (inputs_301__6), .S0 (
             nx24247)) ;
    mux21_ni ix25203 (.Y (nx25202), .A0 (inputs_302__6), .A1 (inputs_303__6), .S0 (
             nx24247)) ;
    mux21_ni ix25271 (.Y (nx25270), .A0 (nx25238), .A1 (nx25266), .S0 (nx23245)
             ) ;
    mux21_ni ix25239 (.Y (nx25238), .A0 (nx25222), .A1 (nx25234), .S0 (nx23559)
             ) ;
    mux21_ni ix25223 (.Y (nx25222), .A0 (inputs_312__6), .A1 (inputs_313__6), .S0 (
             nx24247)) ;
    mux21_ni ix25235 (.Y (nx25234), .A0 (inputs_314__6), .A1 (inputs_315__6), .S0 (
             nx24247)) ;
    mux21_ni ix25267 (.Y (nx25266), .A0 (nx25250), .A1 (nx25262), .S0 (nx23559)
             ) ;
    mux21_ni ix25251 (.Y (nx25250), .A0 (inputs_316__6), .A1 (inputs_317__6), .S0 (
             nx24247)) ;
    mux21_ni ix25263 (.Y (nx25262), .A0 (inputs_318__6), .A1 (inputs_319__6), .S0 (
             nx24247)) ;
    mux21_ni ix25783 (.Y (nx25782), .A0 (nx25570), .A1 (nx25778), .S0 (nx22581)
             ) ;
    mux21_ni ix25571 (.Y (nx25570), .A0 (nx25564), .A1 (nx25486), .S0 (nx23145)
             ) ;
    oai21 ix25565 (.Y (nx25564), .A0 (nx22283), .A1 (nx13603), .B0 (nx13615)) ;
    mux21 ix13604 (.Y (nx13603), .A0 (nx25528), .A1 (nx25556), .S0 (nx22843)) ;
    mux21_ni ix25529 (.Y (nx25528), .A0 (nx25512), .A1 (nx25524), .S0 (nx23559)
             ) ;
    mux21_ni ix25513 (.Y (nx25512), .A0 (inputs_324__6), .A1 (inputs_325__6), .S0 (
             nx24247)) ;
    mux21_ni ix25525 (.Y (nx25524), .A0 (inputs_326__6), .A1 (inputs_327__6), .S0 (
             nx24249)) ;
    mux21_ni ix25557 (.Y (nx25556), .A0 (nx25540), .A1 (nx25552), .S0 (nx23559)
             ) ;
    mux21_ni ix25541 (.Y (nx25540), .A0 (inputs_340__6), .A1 (inputs_341__6), .S0 (
             nx24249)) ;
    mux21_ni ix25553 (.Y (nx25552), .A0 (inputs_342__6), .A1 (inputs_343__6), .S0 (
             nx24249)) ;
    nand04 ix13616 (.Y (nx13615), .A0 (nx22285), .A1 (nx23561), .A2 (nx24249), .A3 (
           nx25500)) ;
    mux21_ni ix25501 (.Y (nx25500), .A0 (inputs_323__6), .A1 (inputs_339__6), .S0 (
             nx22843)) ;
    mux21_ni ix25487 (.Y (nx25486), .A0 (nx25422), .A1 (nx25482), .S0 (nx22843)
             ) ;
    mux21_ni ix25423 (.Y (nx25422), .A0 (nx25390), .A1 (nx25418), .S0 (nx23247)
             ) ;
    mux21_ni ix25391 (.Y (nx25390), .A0 (nx25374), .A1 (nx25386), .S0 (nx23561)
             ) ;
    mux21_ni ix25375 (.Y (nx25374), .A0 (inputs_328__6), .A1 (inputs_329__6), .S0 (
             nx24249)) ;
    mux21_ni ix25387 (.Y (nx25386), .A0 (inputs_330__6), .A1 (inputs_331__6), .S0 (
             nx24249)) ;
    mux21_ni ix25419 (.Y (nx25418), .A0 (nx25402), .A1 (nx25414), .S0 (nx23561)
             ) ;
    mux21_ni ix25403 (.Y (nx25402), .A0 (inputs_332__6), .A1 (inputs_333__6), .S0 (
             nx24249)) ;
    mux21_ni ix25415 (.Y (nx25414), .A0 (inputs_334__6), .A1 (inputs_335__6), .S0 (
             nx24251)) ;
    mux21_ni ix25483 (.Y (nx25482), .A0 (nx25450), .A1 (nx25478), .S0 (nx23247)
             ) ;
    mux21_ni ix25451 (.Y (nx25450), .A0 (nx25434), .A1 (nx25446), .S0 (nx23561)
             ) ;
    mux21_ni ix25435 (.Y (nx25434), .A0 (inputs_344__6), .A1 (inputs_345__6), .S0 (
             nx24251)) ;
    mux21_ni ix25447 (.Y (nx25446), .A0 (inputs_346__6), .A1 (inputs_347__6), .S0 (
             nx24251)) ;
    mux21_ni ix25479 (.Y (nx25478), .A0 (nx25462), .A1 (nx25474), .S0 (nx23561)
             ) ;
    mux21_ni ix25463 (.Y (nx25462), .A0 (inputs_348__6), .A1 (inputs_349__6), .S0 (
             nx24251)) ;
    mux21_ni ix25475 (.Y (nx25474), .A0 (inputs_350__6), .A1 (inputs_351__6), .S0 (
             nx24251)) ;
    mux21_ni ix25779 (.Y (nx25778), .A0 (nx25772), .A1 (nx25694), .S0 (nx23145)
             ) ;
    oai21 ix25773 (.Y (nx25772), .A0 (nx22285), .A1 (nx13649), .B0 (nx13661)) ;
    mux21 ix13650 (.Y (nx13649), .A0 (nx25736), .A1 (nx25764), .S0 (nx22843)) ;
    mux21_ni ix25737 (.Y (nx25736), .A0 (nx25720), .A1 (nx25732), .S0 (nx23561)
             ) ;
    mux21_ni ix25721 (.Y (nx25720), .A0 (inputs_356__6), .A1 (inputs_357__6), .S0 (
             nx24251)) ;
    mux21_ni ix25733 (.Y (nx25732), .A0 (inputs_358__6), .A1 (inputs_359__6), .S0 (
             nx24251)) ;
    mux21_ni ix25765 (.Y (nx25764), .A0 (nx25748), .A1 (nx25760), .S0 (nx23561)
             ) ;
    mux21_ni ix25749 (.Y (nx25748), .A0 (inputs_372__6), .A1 (inputs_373__6), .S0 (
             nx24253)) ;
    mux21_ni ix25761 (.Y (nx25760), .A0 (inputs_374__6), .A1 (inputs_375__6), .S0 (
             nx24253)) ;
    nand04 ix13662 (.Y (nx13661), .A0 (nx22285), .A1 (nx23563), .A2 (nx24253), .A3 (
           nx25708)) ;
    mux21_ni ix25709 (.Y (nx25708), .A0 (inputs_355__6), .A1 (inputs_371__6), .S0 (
             nx22843)) ;
    mux21_ni ix25695 (.Y (nx25694), .A0 (nx25630), .A1 (nx25690), .S0 (nx22843)
             ) ;
    mux21_ni ix25631 (.Y (nx25630), .A0 (nx25598), .A1 (nx25626), .S0 (nx23247)
             ) ;
    mux21_ni ix25599 (.Y (nx25598), .A0 (nx25582), .A1 (nx25594), .S0 (nx23563)
             ) ;
    mux21_ni ix25583 (.Y (nx25582), .A0 (inputs_360__6), .A1 (inputs_361__6), .S0 (
             nx24253)) ;
    mux21_ni ix25595 (.Y (nx25594), .A0 (inputs_362__6), .A1 (inputs_363__6), .S0 (
             nx24253)) ;
    mux21_ni ix25627 (.Y (nx25626), .A0 (nx25610), .A1 (nx25622), .S0 (nx23563)
             ) ;
    mux21_ni ix25611 (.Y (nx25610), .A0 (inputs_364__6), .A1 (inputs_365__6), .S0 (
             nx24253)) ;
    mux21_ni ix25623 (.Y (nx25622), .A0 (inputs_366__6), .A1 (inputs_367__6), .S0 (
             nx24253)) ;
    mux21_ni ix25691 (.Y (nx25690), .A0 (nx25658), .A1 (nx25686), .S0 (nx23247)
             ) ;
    mux21_ni ix25659 (.Y (nx25658), .A0 (nx25642), .A1 (nx25654), .S0 (nx23563)
             ) ;
    mux21_ni ix25643 (.Y (nx25642), .A0 (inputs_376__6), .A1 (inputs_377__6), .S0 (
             nx24255)) ;
    mux21_ni ix25655 (.Y (nx25654), .A0 (inputs_378__6), .A1 (inputs_379__6), .S0 (
             nx24255)) ;
    mux21_ni ix25687 (.Y (nx25686), .A0 (nx25670), .A1 (nx25682), .S0 (nx23563)
             ) ;
    mux21_ni ix25671 (.Y (nx25670), .A0 (inputs_380__6), .A1 (inputs_381__6), .S0 (
             nx24255)) ;
    mux21_ni ix25683 (.Y (nx25682), .A0 (inputs_382__6), .A1 (inputs_383__6), .S0 (
             nx24255)) ;
    mux21_ni ix26631 (.Y (nx26630), .A0 (nx26206), .A1 (nx26626), .S0 (nx22477)
             ) ;
    mux21_ni ix26207 (.Y (nx26206), .A0 (nx25994), .A1 (nx26202), .S0 (nx22581)
             ) ;
    mux21_ni ix25995 (.Y (nx25994), .A0 (nx25988), .A1 (nx25910), .S0 (nx23145)
             ) ;
    oai21 ix25989 (.Y (nx25988), .A0 (nx22285), .A1 (nx13695), .B0 (nx13707)) ;
    mux21 ix13696 (.Y (nx13695), .A0 (nx25952), .A1 (nx25980), .S0 (nx22845)) ;
    mux21_ni ix25953 (.Y (nx25952), .A0 (nx25936), .A1 (nx25948), .S0 (nx23563)
             ) ;
    mux21_ni ix25937 (.Y (nx25936), .A0 (inputs_388__6), .A1 (inputs_389__6), .S0 (
             nx24255)) ;
    mux21_ni ix25949 (.Y (nx25948), .A0 (inputs_390__6), .A1 (inputs_391__6), .S0 (
             nx24255)) ;
    mux21_ni ix25981 (.Y (nx25980), .A0 (nx25964), .A1 (nx25976), .S0 (nx23563)
             ) ;
    mux21_ni ix25965 (.Y (nx25964), .A0 (inputs_404__6), .A1 (inputs_405__6), .S0 (
             nx24255)) ;
    mux21_ni ix25977 (.Y (nx25976), .A0 (inputs_406__6), .A1 (inputs_407__6), .S0 (
             nx24257)) ;
    nand04 ix13708 (.Y (nx13707), .A0 (nx22285), .A1 (nx23565), .A2 (nx24257), .A3 (
           nx25924)) ;
    mux21_ni ix25925 (.Y (nx25924), .A0 (inputs_387__6), .A1 (inputs_403__6), .S0 (
             nx22845)) ;
    mux21_ni ix25911 (.Y (nx25910), .A0 (nx25846), .A1 (nx25906), .S0 (nx22845)
             ) ;
    mux21_ni ix25847 (.Y (nx25846), .A0 (nx25814), .A1 (nx25842), .S0 (nx23247)
             ) ;
    mux21_ni ix25815 (.Y (nx25814), .A0 (nx25798), .A1 (nx25810), .S0 (nx23565)
             ) ;
    mux21_ni ix25799 (.Y (nx25798), .A0 (inputs_392__6), .A1 (inputs_393__6), .S0 (
             nx24257)) ;
    mux21_ni ix25811 (.Y (nx25810), .A0 (inputs_394__6), .A1 (inputs_395__6), .S0 (
             nx24257)) ;
    mux21_ni ix25843 (.Y (nx25842), .A0 (nx25826), .A1 (nx25838), .S0 (nx23565)
             ) ;
    mux21_ni ix25827 (.Y (nx25826), .A0 (inputs_396__6), .A1 (inputs_397__6), .S0 (
             nx24257)) ;
    mux21_ni ix25839 (.Y (nx25838), .A0 (inputs_398__6), .A1 (inputs_399__6), .S0 (
             nx24257)) ;
    mux21_ni ix25907 (.Y (nx25906), .A0 (nx25874), .A1 (nx25902), .S0 (nx23247)
             ) ;
    mux21_ni ix25875 (.Y (nx25874), .A0 (nx25858), .A1 (nx25870), .S0 (nx23565)
             ) ;
    mux21_ni ix25859 (.Y (nx25858), .A0 (inputs_408__6), .A1 (inputs_409__6), .S0 (
             nx24257)) ;
    mux21_ni ix25871 (.Y (nx25870), .A0 (inputs_410__6), .A1 (inputs_411__6), .S0 (
             nx24259)) ;
    mux21_ni ix25903 (.Y (nx25902), .A0 (nx25886), .A1 (nx25898), .S0 (nx23565)
             ) ;
    mux21_ni ix25887 (.Y (nx25886), .A0 (inputs_412__6), .A1 (inputs_413__6), .S0 (
             nx24259)) ;
    mux21_ni ix25899 (.Y (nx25898), .A0 (inputs_414__6), .A1 (inputs_415__6), .S0 (
             nx24259)) ;
    mux21_ni ix26203 (.Y (nx26202), .A0 (nx26196), .A1 (nx26118), .S0 (nx23145)
             ) ;
    oai21 ix26197 (.Y (nx26196), .A0 (nx22285), .A1 (nx13741), .B0 (nx13753)) ;
    mux21 ix13742 (.Y (nx13741), .A0 (nx26160), .A1 (nx26188), .S0 (nx22845)) ;
    mux21_ni ix26161 (.Y (nx26160), .A0 (nx26144), .A1 (nx26156), .S0 (nx23565)
             ) ;
    mux21_ni ix26145 (.Y (nx26144), .A0 (inputs_420__6), .A1 (inputs_421__6), .S0 (
             nx24259)) ;
    mux21_ni ix26157 (.Y (nx26156), .A0 (inputs_422__6), .A1 (inputs_423__6), .S0 (
             nx24259)) ;
    mux21_ni ix26189 (.Y (nx26188), .A0 (nx26172), .A1 (nx26184), .S0 (nx23565)
             ) ;
    mux21_ni ix26173 (.Y (nx26172), .A0 (inputs_436__6), .A1 (inputs_437__6), .S0 (
             nx24259)) ;
    mux21_ni ix26185 (.Y (nx26184), .A0 (inputs_438__6), .A1 (inputs_439__6), .S0 (
             nx24259)) ;
    nand04 ix13754 (.Y (nx13753), .A0 (nx22285), .A1 (nx23567), .A2 (nx24261), .A3 (
           nx26132)) ;
    mux21_ni ix26133 (.Y (nx26132), .A0 (inputs_419__6), .A1 (inputs_435__6), .S0 (
             nx22845)) ;
    mux21_ni ix26119 (.Y (nx26118), .A0 (nx26054), .A1 (nx26114), .S0 (nx22845)
             ) ;
    mux21_ni ix26055 (.Y (nx26054), .A0 (nx26022), .A1 (nx26050), .S0 (nx23247)
             ) ;
    mux21_ni ix26023 (.Y (nx26022), .A0 (nx26006), .A1 (nx26018), .S0 (nx23567)
             ) ;
    mux21_ni ix26007 (.Y (nx26006), .A0 (inputs_424__6), .A1 (inputs_425__6), .S0 (
             nx24261)) ;
    mux21_ni ix26019 (.Y (nx26018), .A0 (inputs_426__6), .A1 (inputs_427__6), .S0 (
             nx24261)) ;
    mux21_ni ix26051 (.Y (nx26050), .A0 (nx26034), .A1 (nx26046), .S0 (nx23567)
             ) ;
    mux21_ni ix26035 (.Y (nx26034), .A0 (inputs_428__6), .A1 (inputs_429__6), .S0 (
             nx24261)) ;
    mux21_ni ix26047 (.Y (nx26046), .A0 (inputs_430__6), .A1 (inputs_431__6), .S0 (
             nx24261)) ;
    mux21_ni ix26115 (.Y (nx26114), .A0 (nx26082), .A1 (nx26110), .S0 (nx23249)
             ) ;
    mux21_ni ix26083 (.Y (nx26082), .A0 (nx26066), .A1 (nx26078), .S0 (nx23567)
             ) ;
    mux21_ni ix26067 (.Y (nx26066), .A0 (inputs_440__6), .A1 (inputs_441__6), .S0 (
             nx24261)) ;
    mux21_ni ix26079 (.Y (nx26078), .A0 (inputs_442__6), .A1 (inputs_443__6), .S0 (
             nx24261)) ;
    mux21_ni ix26111 (.Y (nx26110), .A0 (nx26094), .A1 (nx26106), .S0 (nx23567)
             ) ;
    mux21_ni ix26095 (.Y (nx26094), .A0 (inputs_444__6), .A1 (inputs_445__6), .S0 (
             nx24263)) ;
    mux21_ni ix26107 (.Y (nx26106), .A0 (inputs_446__6), .A1 (inputs_447__6), .S0 (
             nx24263)) ;
    mux21_ni ix26627 (.Y (nx26626), .A0 (nx26414), .A1 (nx26622), .S0 (nx22581)
             ) ;
    mux21_ni ix26415 (.Y (nx26414), .A0 (nx26408), .A1 (nx26330), .S0 (nx23145)
             ) ;
    oai21 ix26409 (.Y (nx26408), .A0 (nx22287), .A1 (nx13785), .B0 (nx13797)) ;
    mux21 ix13786 (.Y (nx13785), .A0 (nx26372), .A1 (nx26400), .S0 (nx22845)) ;
    mux21_ni ix26373 (.Y (nx26372), .A0 (nx26356), .A1 (nx26368), .S0 (nx23567)
             ) ;
    mux21_ni ix26357 (.Y (nx26356), .A0 (inputs_452__6), .A1 (inputs_453__6), .S0 (
             nx24263)) ;
    mux21_ni ix26369 (.Y (nx26368), .A0 (inputs_454__6), .A1 (inputs_455__6), .S0 (
             nx24263)) ;
    mux21_ni ix26401 (.Y (nx26400), .A0 (nx26384), .A1 (nx26396), .S0 (nx23567)
             ) ;
    mux21_ni ix26385 (.Y (nx26384), .A0 (inputs_468__6), .A1 (inputs_469__6), .S0 (
             nx24263)) ;
    mux21_ni ix26397 (.Y (nx26396), .A0 (inputs_470__6), .A1 (inputs_471__6), .S0 (
             nx24263)) ;
    nand04 ix13798 (.Y (nx13797), .A0 (nx22287), .A1 (nx23569), .A2 (nx24263), .A3 (
           nx26344)) ;
    mux21_ni ix26345 (.Y (nx26344), .A0 (inputs_451__6), .A1 (inputs_467__6), .S0 (
             nx22847)) ;
    mux21_ni ix26331 (.Y (nx26330), .A0 (nx26266), .A1 (nx26326), .S0 (nx22847)
             ) ;
    mux21_ni ix26267 (.Y (nx26266), .A0 (nx26234), .A1 (nx26262), .S0 (nx23249)
             ) ;
    mux21_ni ix26235 (.Y (nx26234), .A0 (nx26218), .A1 (nx26230), .S0 (nx23569)
             ) ;
    mux21_ni ix26219 (.Y (nx26218), .A0 (inputs_456__6), .A1 (inputs_457__6), .S0 (
             nx24265)) ;
    mux21_ni ix26231 (.Y (nx26230), .A0 (inputs_458__6), .A1 (inputs_459__6), .S0 (
             nx24265)) ;
    mux21_ni ix26263 (.Y (nx26262), .A0 (nx26246), .A1 (nx26258), .S0 (nx23569)
             ) ;
    mux21_ni ix26247 (.Y (nx26246), .A0 (inputs_460__6), .A1 (inputs_461__6), .S0 (
             nx24265)) ;
    mux21_ni ix26259 (.Y (nx26258), .A0 (inputs_462__6), .A1 (inputs_463__6), .S0 (
             nx24265)) ;
    mux21_ni ix26327 (.Y (nx26326), .A0 (nx26294), .A1 (nx26322), .S0 (nx23249)
             ) ;
    mux21_ni ix26295 (.Y (nx26294), .A0 (nx26278), .A1 (nx26290), .S0 (nx23569)
             ) ;
    mux21_ni ix26279 (.Y (nx26278), .A0 (inputs_472__6), .A1 (inputs_473__6), .S0 (
             nx24265)) ;
    mux21_ni ix26291 (.Y (nx26290), .A0 (inputs_474__6), .A1 (inputs_475__6), .S0 (
             nx24265)) ;
    mux21_ni ix26323 (.Y (nx26322), .A0 (nx26306), .A1 (nx26318), .S0 (nx23569)
             ) ;
    mux21_ni ix26307 (.Y (nx26306), .A0 (inputs_476__6), .A1 (inputs_477__6), .S0 (
             nx24265)) ;
    mux21_ni ix26319 (.Y (nx26318), .A0 (inputs_478__6), .A1 (inputs_479__6), .S0 (
             nx24267)) ;
    mux21_ni ix26623 (.Y (nx26622), .A0 (nx26616), .A1 (nx26538), .S0 (nx23145)
             ) ;
    oai21 ix26617 (.Y (nx26616), .A0 (nx22287), .A1 (nx13827), .B0 (nx13839)) ;
    mux21 ix13828 (.Y (nx13827), .A0 (nx26580), .A1 (nx26608), .S0 (nx22847)) ;
    mux21_ni ix26581 (.Y (nx26580), .A0 (nx26564), .A1 (nx26576), .S0 (nx23569)
             ) ;
    mux21_ni ix26565 (.Y (nx26564), .A0 (inputs_484__6), .A1 (inputs_485__6), .S0 (
             nx24267)) ;
    mux21_ni ix26577 (.Y (nx26576), .A0 (inputs_486__6), .A1 (inputs_487__6), .S0 (
             nx24267)) ;
    mux21_ni ix26609 (.Y (nx26608), .A0 (nx26592), .A1 (nx26604), .S0 (nx23569)
             ) ;
    mux21_ni ix26593 (.Y (nx26592), .A0 (inputs_500__6), .A1 (inputs_501__6), .S0 (
             nx24267)) ;
    mux21_ni ix26605 (.Y (nx26604), .A0 (inputs_502__6), .A1 (inputs_503__6), .S0 (
             nx24267)) ;
    nand04 ix13840 (.Y (nx13839), .A0 (nx22287), .A1 (nx23571), .A2 (nx24267), .A3 (
           nx26552)) ;
    mux21_ni ix26553 (.Y (nx26552), .A0 (inputs_483__6), .A1 (inputs_499__6), .S0 (
             nx22847)) ;
    mux21_ni ix26539 (.Y (nx26538), .A0 (nx26474), .A1 (nx26534), .S0 (nx22847)
             ) ;
    mux21_ni ix26475 (.Y (nx26474), .A0 (nx26442), .A1 (nx26470), .S0 (nx23249)
             ) ;
    mux21_ni ix26443 (.Y (nx26442), .A0 (nx26426), .A1 (nx26438), .S0 (nx23571)
             ) ;
    mux21_ni ix26427 (.Y (nx26426), .A0 (inputs_488__6), .A1 (inputs_489__6), .S0 (
             nx24267)) ;
    mux21_ni ix26439 (.Y (nx26438), .A0 (inputs_490__6), .A1 (inputs_491__6), .S0 (
             nx24269)) ;
    mux21_ni ix26471 (.Y (nx26470), .A0 (nx26454), .A1 (nx26466), .S0 (nx23571)
             ) ;
    mux21_ni ix26455 (.Y (nx26454), .A0 (inputs_492__6), .A1 (inputs_493__6), .S0 (
             nx24269)) ;
    mux21_ni ix26467 (.Y (nx26466), .A0 (inputs_494__6), .A1 (inputs_495__6), .S0 (
             nx24269)) ;
    mux21_ni ix26535 (.Y (nx26534), .A0 (nx26502), .A1 (nx26530), .S0 (nx23249)
             ) ;
    mux21_ni ix26503 (.Y (nx26502), .A0 (nx26486), .A1 (nx26498), .S0 (nx23571)
             ) ;
    mux21_ni ix26487 (.Y (nx26486), .A0 (inputs_504__6), .A1 (inputs_505__6), .S0 (
             nx24269)) ;
    mux21_ni ix26499 (.Y (nx26498), .A0 (inputs_506__6), .A1 (inputs_507__6), .S0 (
             nx24269)) ;
    mux21_ni ix26531 (.Y (nx26530), .A0 (nx26514), .A1 (nx26526), .S0 (nx23571)
             ) ;
    mux21_ni ix26515 (.Y (nx26514), .A0 (inputs_508__6), .A1 (inputs_509__6), .S0 (
             nx24269)) ;
    mux21_ni ix26527 (.Y (nx26526), .A0 (inputs_510__6), .A1 (inputs_511__6), .S0 (
             nx24269)) ;
    aoi32 ix13870 (.Y (nx13869), .A0 (nx27400), .A1 (nx22387), .A2 (nx22287), .B0 (
          nx22219), .B1 (nx29096)) ;
    oai21 ix27401 (.Y (nx27400), .A0 (nx23571), .A1 (nx13873), .B0 (nx13973)) ;
    mux21 ix13874 (.Y (nx13873), .A0 (nx27138), .A1 (nx27390), .S0 (nx24271)) ;
    mux21_ni ix27139 (.Y (nx27138), .A0 (nx27010), .A1 (nx27134), .S0 (nx22397)
             ) ;
    mux21_ni ix27011 (.Y (nx27010), .A0 (nx26946), .A1 (nx27006), .S0 (nx22425)
             ) ;
    mux21_ni ix26947 (.Y (nx26946), .A0 (nx26914), .A1 (nx26942), .S0 (nx22479)
             ) ;
    mux21_ni ix26915 (.Y (nx26914), .A0 (nx26898), .A1 (nx26910), .S0 (nx22583)
             ) ;
    mux21_ni ix26899 (.Y (nx26898), .A0 (inputs_0__6), .A1 (inputs_16__6), .S0 (
             nx22847)) ;
    mux21_ni ix26911 (.Y (nx26910), .A0 (inputs_32__6), .A1 (inputs_48__6), .S0 (
             nx22847)) ;
    mux21_ni ix26943 (.Y (nx26942), .A0 (nx26926), .A1 (nx26938), .S0 (nx22583)
             ) ;
    mux21_ni ix26927 (.Y (nx26926), .A0 (inputs_64__6), .A1 (inputs_80__6), .S0 (
             nx22849)) ;
    mux21_ni ix26939 (.Y (nx26938), .A0 (inputs_96__6), .A1 (inputs_112__6), .S0 (
             nx22849)) ;
    mux21_ni ix27007 (.Y (nx27006), .A0 (nx26974), .A1 (nx27002), .S0 (nx22479)
             ) ;
    mux21_ni ix26975 (.Y (nx26974), .A0 (nx26958), .A1 (nx26970), .S0 (nx22583)
             ) ;
    mux21_ni ix26959 (.Y (nx26958), .A0 (inputs_128__6), .A1 (inputs_144__6), .S0 (
             nx22849)) ;
    mux21_ni ix26971 (.Y (nx26970), .A0 (inputs_160__6), .A1 (inputs_176__6), .S0 (
             nx22849)) ;
    mux21_ni ix27003 (.Y (nx27002), .A0 (nx26986), .A1 (nx26998), .S0 (nx22583)
             ) ;
    mux21_ni ix26987 (.Y (nx26986), .A0 (inputs_192__6), .A1 (inputs_208__6), .S0 (
             nx22849)) ;
    mux21_ni ix26999 (.Y (nx26998), .A0 (inputs_224__6), .A1 (inputs_240__6), .S0 (
             nx22849)) ;
    mux21_ni ix27135 (.Y (nx27134), .A0 (nx27070), .A1 (nx27130), .S0 (nx22425)
             ) ;
    mux21_ni ix27071 (.Y (nx27070), .A0 (nx27038), .A1 (nx27066), .S0 (nx22479)
             ) ;
    mux21_ni ix27039 (.Y (nx27038), .A0 (nx27022), .A1 (nx27034), .S0 (nx22583)
             ) ;
    mux21_ni ix27023 (.Y (nx27022), .A0 (inputs_256__6), .A1 (inputs_272__6), .S0 (
             nx22849)) ;
    mux21_ni ix27035 (.Y (nx27034), .A0 (inputs_288__6), .A1 (inputs_304__6), .S0 (
             nx22851)) ;
    mux21_ni ix27067 (.Y (nx27066), .A0 (nx27050), .A1 (nx27062), .S0 (nx22583)
             ) ;
    mux21_ni ix27051 (.Y (nx27050), .A0 (inputs_320__6), .A1 (inputs_336__6), .S0 (
             nx22851)) ;
    mux21_ni ix27063 (.Y (nx27062), .A0 (inputs_352__6), .A1 (inputs_368__6), .S0 (
             nx22851)) ;
    mux21_ni ix27131 (.Y (nx27130), .A0 (nx27098), .A1 (nx27126), .S0 (nx22479)
             ) ;
    mux21_ni ix27099 (.Y (nx27098), .A0 (nx27082), .A1 (nx27094), .S0 (nx22583)
             ) ;
    mux21_ni ix27083 (.Y (nx27082), .A0 (inputs_384__6), .A1 (inputs_400__6), .S0 (
             nx22851)) ;
    mux21_ni ix27095 (.Y (nx27094), .A0 (inputs_416__6), .A1 (inputs_432__6), .S0 (
             nx22851)) ;
    mux21_ni ix27127 (.Y (nx27126), .A0 (nx27110), .A1 (nx27122), .S0 (nx22585)
             ) ;
    mux21_ni ix27111 (.Y (nx27110), .A0 (inputs_448__6), .A1 (inputs_464__6), .S0 (
             nx22851)) ;
    mux21_ni ix27123 (.Y (nx27122), .A0 (inputs_480__6), .A1 (inputs_496__6), .S0 (
             nx22851)) ;
    mux21_ni ix27391 (.Y (nx27390), .A0 (nx27262), .A1 (nx27386), .S0 (nx22397)
             ) ;
    mux21_ni ix27263 (.Y (nx27262), .A0 (nx27198), .A1 (nx27258), .S0 (nx22425)
             ) ;
    mux21_ni ix27199 (.Y (nx27198), .A0 (nx27166), .A1 (nx27194), .S0 (nx22479)
             ) ;
    mux21_ni ix27167 (.Y (nx27166), .A0 (nx27150), .A1 (nx27162), .S0 (nx22585)
             ) ;
    mux21_ni ix27151 (.Y (nx27150), .A0 (inputs_1__6), .A1 (inputs_17__6), .S0 (
             nx22853)) ;
    mux21_ni ix27163 (.Y (nx27162), .A0 (inputs_33__6), .A1 (inputs_49__6), .S0 (
             nx22853)) ;
    mux21_ni ix27195 (.Y (nx27194), .A0 (nx27178), .A1 (nx27190), .S0 (nx22585)
             ) ;
    mux21_ni ix27179 (.Y (nx27178), .A0 (inputs_65__6), .A1 (inputs_81__6), .S0 (
             nx22853)) ;
    mux21_ni ix27191 (.Y (nx27190), .A0 (inputs_97__6), .A1 (inputs_113__6), .S0 (
             nx22853)) ;
    mux21_ni ix27259 (.Y (nx27258), .A0 (nx27226), .A1 (nx27254), .S0 (nx22479)
             ) ;
    mux21_ni ix27227 (.Y (nx27226), .A0 (nx27210), .A1 (nx27222), .S0 (nx22585)
             ) ;
    mux21_ni ix27211 (.Y (nx27210), .A0 (inputs_129__6), .A1 (inputs_145__6), .S0 (
             nx22853)) ;
    mux21_ni ix27223 (.Y (nx27222), .A0 (inputs_161__6), .A1 (inputs_177__6), .S0 (
             nx22853)) ;
    mux21_ni ix27255 (.Y (nx27254), .A0 (nx27238), .A1 (nx27250), .S0 (nx22585)
             ) ;
    mux21_ni ix27239 (.Y (nx27238), .A0 (inputs_193__6), .A1 (inputs_209__6), .S0 (
             nx22853)) ;
    mux21_ni ix27251 (.Y (nx27250), .A0 (inputs_225__6), .A1 (inputs_241__6), .S0 (
             nx22855)) ;
    mux21_ni ix27387 (.Y (nx27386), .A0 (nx27322), .A1 (nx27382), .S0 (nx22425)
             ) ;
    mux21_ni ix27323 (.Y (nx27322), .A0 (nx27290), .A1 (nx27318), .S0 (nx22479)
             ) ;
    mux21_ni ix27291 (.Y (nx27290), .A0 (nx27274), .A1 (nx27286), .S0 (nx22585)
             ) ;
    mux21_ni ix27275 (.Y (nx27274), .A0 (inputs_257__6), .A1 (inputs_273__6), .S0 (
             nx22855)) ;
    mux21_ni ix27287 (.Y (nx27286), .A0 (inputs_289__6), .A1 (inputs_305__6), .S0 (
             nx22855)) ;
    mux21_ni ix27319 (.Y (nx27318), .A0 (nx27302), .A1 (nx27314), .S0 (nx22585)
             ) ;
    mux21_ni ix27303 (.Y (nx27302), .A0 (inputs_321__6), .A1 (inputs_337__6), .S0 (
             nx22855)) ;
    mux21_ni ix27315 (.Y (nx27314), .A0 (inputs_353__6), .A1 (inputs_369__6), .S0 (
             nx22855)) ;
    mux21_ni ix27383 (.Y (nx27382), .A0 (nx27350), .A1 (nx27378), .S0 (nx22481)
             ) ;
    mux21_ni ix27351 (.Y (nx27350), .A0 (nx27334), .A1 (nx27346), .S0 (nx22587)
             ) ;
    mux21_ni ix27335 (.Y (nx27334), .A0 (inputs_385__6), .A1 (inputs_401__6), .S0 (
             nx22855)) ;
    mux21_ni ix27347 (.Y (nx27346), .A0 (inputs_417__6), .A1 (inputs_433__6), .S0 (
             nx22855)) ;
    mux21_ni ix27379 (.Y (nx27378), .A0 (nx27362), .A1 (nx27374), .S0 (nx22587)
             ) ;
    mux21_ni ix27363 (.Y (nx27362), .A0 (inputs_449__6), .A1 (inputs_465__6), .S0 (
             nx22857)) ;
    mux21_ni ix27375 (.Y (nx27374), .A0 (inputs_481__6), .A1 (inputs_497__6), .S0 (
             nx22857)) ;
    nand03 ix13974 (.Y (nx13973), .A0 (nx26884), .A1 (nx23571), .A2 (nx24879)) ;
    mux21_ni ix26885 (.Y (nx26884), .A0 (nx26756), .A1 (nx26880), .S0 (nx22397)
             ) ;
    mux21_ni ix26757 (.Y (nx26756), .A0 (nx26692), .A1 (nx26752), .S0 (nx22425)
             ) ;
    mux21_ni ix26693 (.Y (nx26692), .A0 (nx26660), .A1 (nx26688), .S0 (nx22481)
             ) ;
    mux21_ni ix26661 (.Y (nx26660), .A0 (nx26644), .A1 (nx26656), .S0 (nx22587)
             ) ;
    mux21_ni ix26645 (.Y (nx26644), .A0 (inputs_2__6), .A1 (inputs_18__6), .S0 (
             nx22857)) ;
    mux21_ni ix26657 (.Y (nx26656), .A0 (inputs_34__6), .A1 (inputs_50__6), .S0 (
             nx22857)) ;
    mux21_ni ix26689 (.Y (nx26688), .A0 (nx26672), .A1 (nx26684), .S0 (nx22587)
             ) ;
    mux21_ni ix26673 (.Y (nx26672), .A0 (inputs_66__6), .A1 (inputs_82__6), .S0 (
             nx22857)) ;
    mux21_ni ix26685 (.Y (nx26684), .A0 (inputs_98__6), .A1 (inputs_114__6), .S0 (
             nx22857)) ;
    mux21_ni ix26753 (.Y (nx26752), .A0 (nx26720), .A1 (nx26748), .S0 (nx22481)
             ) ;
    mux21_ni ix26721 (.Y (nx26720), .A0 (nx26704), .A1 (nx26716), .S0 (nx22587)
             ) ;
    mux21_ni ix26705 (.Y (nx26704), .A0 (inputs_130__6), .A1 (inputs_146__6), .S0 (
             nx22857)) ;
    mux21_ni ix26717 (.Y (nx26716), .A0 (inputs_162__6), .A1 (inputs_178__6), .S0 (
             nx22859)) ;
    mux21_ni ix26749 (.Y (nx26748), .A0 (nx26732), .A1 (nx26744), .S0 (nx22587)
             ) ;
    mux21_ni ix26733 (.Y (nx26732), .A0 (inputs_194__6), .A1 (inputs_210__6), .S0 (
             nx22859)) ;
    mux21_ni ix26745 (.Y (nx26744), .A0 (inputs_226__6), .A1 (inputs_242__6), .S0 (
             nx22859)) ;
    mux21_ni ix26881 (.Y (nx26880), .A0 (nx26816), .A1 (nx26876), .S0 (nx22425)
             ) ;
    mux21_ni ix26817 (.Y (nx26816), .A0 (nx26784), .A1 (nx26812), .S0 (nx22481)
             ) ;
    mux21_ni ix26785 (.Y (nx26784), .A0 (nx26768), .A1 (nx26780), .S0 (nx22587)
             ) ;
    mux21_ni ix26769 (.Y (nx26768), .A0 (inputs_258__6), .A1 (inputs_274__6), .S0 (
             nx22859)) ;
    mux21_ni ix26781 (.Y (nx26780), .A0 (inputs_290__6), .A1 (inputs_306__6), .S0 (
             nx22859)) ;
    mux21_ni ix26813 (.Y (nx26812), .A0 (nx26796), .A1 (nx26808), .S0 (nx22589)
             ) ;
    mux21_ni ix26797 (.Y (nx26796), .A0 (inputs_322__6), .A1 (inputs_338__6), .S0 (
             nx22859)) ;
    mux21_ni ix26809 (.Y (nx26808), .A0 (inputs_354__6), .A1 (inputs_370__6), .S0 (
             nx22859)) ;
    mux21_ni ix26877 (.Y (nx26876), .A0 (nx26844), .A1 (nx26872), .S0 (nx22481)
             ) ;
    mux21_ni ix26845 (.Y (nx26844), .A0 (nx26828), .A1 (nx26840), .S0 (nx22589)
             ) ;
    mux21_ni ix26829 (.Y (nx26828), .A0 (inputs_386__6), .A1 (inputs_402__6), .S0 (
             nx22861)) ;
    mux21_ni ix26841 (.Y (nx26840), .A0 (inputs_418__6), .A1 (inputs_434__6), .S0 (
             nx22861)) ;
    mux21_ni ix26873 (.Y (nx26872), .A0 (nx26856), .A1 (nx26868), .S0 (nx22589)
             ) ;
    mux21_ni ix26857 (.Y (nx26856), .A0 (inputs_450__6), .A1 (inputs_466__6), .S0 (
             nx22861)) ;
    mux21_ni ix26869 (.Y (nx26868), .A0 (inputs_482__6), .A1 (inputs_498__6), .S0 (
             nx22861)) ;
    mux21_ni ix29097 (.Y (nx29096), .A0 (nx28248), .A1 (nx29092), .S0 (nx22425)
             ) ;
    mux21_ni ix28249 (.Y (nx28248), .A0 (nx27824), .A1 (nx28244), .S0 (nx22481)
             ) ;
    mux21_ni ix27825 (.Y (nx27824), .A0 (nx27612), .A1 (nx27820), .S0 (nx22589)
             ) ;
    mux21_ni ix27613 (.Y (nx27612), .A0 (nx27606), .A1 (nx27528), .S0 (nx23145)
             ) ;
    oai21 ix27607 (.Y (nx27606), .A0 (nx22287), .A1 (nx14033), .B0 (nx14045)) ;
    mux21 ix14034 (.Y (nx14033), .A0 (nx27570), .A1 (nx27598), .S0 (nx22861)) ;
    mux21_ni ix27571 (.Y (nx27570), .A0 (nx27554), .A1 (nx27566), .S0 (nx23573)
             ) ;
    mux21_ni ix27555 (.Y (nx27554), .A0 (inputs_4__6), .A1 (inputs_5__6), .S0 (
             nx24271)) ;
    mux21_ni ix27567 (.Y (nx27566), .A0 (inputs_6__6), .A1 (inputs_7__6), .S0 (
             nx24271)) ;
    mux21_ni ix27599 (.Y (nx27598), .A0 (nx27582), .A1 (nx27594), .S0 (nx23573)
             ) ;
    mux21_ni ix27583 (.Y (nx27582), .A0 (inputs_20__6), .A1 (inputs_21__6), .S0 (
             nx24271)) ;
    mux21_ni ix27595 (.Y (nx27594), .A0 (inputs_22__6), .A1 (inputs_23__6), .S0 (
             nx24271)) ;
    nand04 ix14046 (.Y (nx14045), .A0 (nx22287), .A1 (nx23573), .A2 (nx24271), .A3 (
           nx27542)) ;
    mux21_ni ix27543 (.Y (nx27542), .A0 (inputs_3__6), .A1 (inputs_19__6), .S0 (
             nx22861)) ;
    mux21_ni ix27529 (.Y (nx27528), .A0 (nx27464), .A1 (nx27524), .S0 (nx22861)
             ) ;
    mux21_ni ix27465 (.Y (nx27464), .A0 (nx27432), .A1 (nx27460), .S0 (nx23249)
             ) ;
    mux21_ni ix27433 (.Y (nx27432), .A0 (nx27416), .A1 (nx27428), .S0 (nx23573)
             ) ;
    mux21_ni ix27417 (.Y (nx27416), .A0 (inputs_8__6), .A1 (inputs_9__6), .S0 (
             nx24271)) ;
    mux21_ni ix27429 (.Y (nx27428), .A0 (inputs_10__6), .A1 (inputs_11__6), .S0 (
             nx24273)) ;
    mux21_ni ix27461 (.Y (nx27460), .A0 (nx27444), .A1 (nx27456), .S0 (nx23573)
             ) ;
    mux21_ni ix27445 (.Y (nx27444), .A0 (inputs_12__6), .A1 (inputs_13__6), .S0 (
             nx24273)) ;
    mux21_ni ix27457 (.Y (nx27456), .A0 (inputs_14__6), .A1 (inputs_15__6), .S0 (
             nx24273)) ;
    mux21_ni ix27525 (.Y (nx27524), .A0 (nx27492), .A1 (nx27520), .S0 (nx23249)
             ) ;
    mux21_ni ix27493 (.Y (nx27492), .A0 (nx27476), .A1 (nx27488), .S0 (nx23573)
             ) ;
    mux21_ni ix27477 (.Y (nx27476), .A0 (inputs_24__6), .A1 (inputs_25__6), .S0 (
             nx24273)) ;
    mux21_ni ix27489 (.Y (nx27488), .A0 (inputs_26__6), .A1 (inputs_27__6), .S0 (
             nx24273)) ;
    mux21_ni ix27521 (.Y (nx27520), .A0 (nx27504), .A1 (nx27516), .S0 (nx23573)
             ) ;
    mux21_ni ix27505 (.Y (nx27504), .A0 (inputs_28__6), .A1 (inputs_29__6), .S0 (
             nx24273)) ;
    mux21_ni ix27517 (.Y (nx27516), .A0 (inputs_30__6), .A1 (inputs_31__6), .S0 (
             nx24273)) ;
    mux21_ni ix27821 (.Y (nx27820), .A0 (nx27814), .A1 (nx27736), .S0 (nx23147)
             ) ;
    oai21 ix27815 (.Y (nx27814), .A0 (nx22289), .A1 (nx14077), .B0 (nx14089)) ;
    mux21 ix14078 (.Y (nx14077), .A0 (nx27778), .A1 (nx27806), .S0 (nx22863)) ;
    mux21_ni ix27779 (.Y (nx27778), .A0 (nx27762), .A1 (nx27774), .S0 (nx23575)
             ) ;
    mux21_ni ix27763 (.Y (nx27762), .A0 (inputs_36__6), .A1 (inputs_37__6), .S0 (
             nx24275)) ;
    mux21_ni ix27775 (.Y (nx27774), .A0 (inputs_38__6), .A1 (inputs_39__6), .S0 (
             nx24275)) ;
    mux21_ni ix27807 (.Y (nx27806), .A0 (nx27790), .A1 (nx27802), .S0 (nx23575)
             ) ;
    mux21_ni ix27791 (.Y (nx27790), .A0 (inputs_52__6), .A1 (inputs_53__6), .S0 (
             nx24275)) ;
    mux21_ni ix27803 (.Y (nx27802), .A0 (inputs_54__6), .A1 (inputs_55__6), .S0 (
             nx24275)) ;
    nand04 ix14090 (.Y (nx14089), .A0 (nx22289), .A1 (nx23575), .A2 (nx24275), .A3 (
           nx27750)) ;
    mux21_ni ix27751 (.Y (nx27750), .A0 (inputs_35__6), .A1 (inputs_51__6), .S0 (
             nx22863)) ;
    mux21_ni ix27737 (.Y (nx27736), .A0 (nx27672), .A1 (nx27732), .S0 (nx22863)
             ) ;
    mux21_ni ix27673 (.Y (nx27672), .A0 (nx27640), .A1 (nx27668), .S0 (nx23251)
             ) ;
    mux21_ni ix27641 (.Y (nx27640), .A0 (nx27624), .A1 (nx27636), .S0 (nx23575)
             ) ;
    mux21_ni ix27625 (.Y (nx27624), .A0 (inputs_40__6), .A1 (inputs_41__6), .S0 (
             nx24275)) ;
    mux21_ni ix27637 (.Y (nx27636), .A0 (inputs_42__6), .A1 (inputs_43__6), .S0 (
             nx24275)) ;
    mux21_ni ix27669 (.Y (nx27668), .A0 (nx27652), .A1 (nx27664), .S0 (nx23575)
             ) ;
    mux21_ni ix27653 (.Y (nx27652), .A0 (inputs_44__6), .A1 (inputs_45__6), .S0 (
             nx24277)) ;
    mux21_ni ix27665 (.Y (nx27664), .A0 (inputs_46__6), .A1 (inputs_47__6), .S0 (
             nx24277)) ;
    mux21_ni ix27733 (.Y (nx27732), .A0 (nx27700), .A1 (nx27728), .S0 (nx23251)
             ) ;
    mux21_ni ix27701 (.Y (nx27700), .A0 (nx27684), .A1 (nx27696), .S0 (nx23575)
             ) ;
    mux21_ni ix27685 (.Y (nx27684), .A0 (inputs_56__6), .A1 (inputs_57__6), .S0 (
             nx24277)) ;
    mux21_ni ix27697 (.Y (nx27696), .A0 (inputs_58__6), .A1 (inputs_59__6), .S0 (
             nx24277)) ;
    mux21_ni ix27729 (.Y (nx27728), .A0 (nx27712), .A1 (nx27724), .S0 (nx23575)
             ) ;
    mux21_ni ix27713 (.Y (nx27712), .A0 (inputs_60__6), .A1 (inputs_61__6), .S0 (
             nx24277)) ;
    mux21_ni ix27725 (.Y (nx27724), .A0 (inputs_62__6), .A1 (inputs_63__6), .S0 (
             nx24277)) ;
    mux21_ni ix28245 (.Y (nx28244), .A0 (nx28032), .A1 (nx28240), .S0 (nx22589)
             ) ;
    mux21_ni ix28033 (.Y (nx28032), .A0 (nx28026), .A1 (nx27948), .S0 (nx23147)
             ) ;
    oai21 ix28027 (.Y (nx28026), .A0 (nx22289), .A1 (nx14121), .B0 (nx14133)) ;
    mux21 ix14122 (.Y (nx14121), .A0 (nx27990), .A1 (nx28018), .S0 (nx22863)) ;
    mux21_ni ix27991 (.Y (nx27990), .A0 (nx27974), .A1 (nx27986), .S0 (nx23577)
             ) ;
    mux21_ni ix27975 (.Y (nx27974), .A0 (inputs_68__6), .A1 (inputs_69__6), .S0 (
             nx24277)) ;
    mux21_ni ix27987 (.Y (nx27986), .A0 (inputs_70__6), .A1 (inputs_71__6), .S0 (
             nx24279)) ;
    mux21_ni ix28019 (.Y (nx28018), .A0 (nx28002), .A1 (nx28014), .S0 (nx23577)
             ) ;
    mux21_ni ix28003 (.Y (nx28002), .A0 (inputs_84__6), .A1 (inputs_85__6), .S0 (
             nx24279)) ;
    mux21_ni ix28015 (.Y (nx28014), .A0 (inputs_86__6), .A1 (inputs_87__6), .S0 (
             nx24279)) ;
    nand04 ix14134 (.Y (nx14133), .A0 (nx22289), .A1 (nx23577), .A2 (nx24279), .A3 (
           nx27962)) ;
    mux21_ni ix27963 (.Y (nx27962), .A0 (inputs_67__6), .A1 (inputs_83__6), .S0 (
             nx22863)) ;
    mux21_ni ix27949 (.Y (nx27948), .A0 (nx27884), .A1 (nx27944), .S0 (nx22863)
             ) ;
    mux21_ni ix27885 (.Y (nx27884), .A0 (nx27852), .A1 (nx27880), .S0 (nx23251)
             ) ;
    mux21_ni ix27853 (.Y (nx27852), .A0 (nx27836), .A1 (nx27848), .S0 (nx23577)
             ) ;
    mux21_ni ix27837 (.Y (nx27836), .A0 (inputs_72__6), .A1 (inputs_73__6), .S0 (
             nx24279)) ;
    mux21_ni ix27849 (.Y (nx27848), .A0 (inputs_74__6), .A1 (inputs_75__6), .S0 (
             nx24279)) ;
    mux21_ni ix27881 (.Y (nx27880), .A0 (nx27864), .A1 (nx27876), .S0 (nx23577)
             ) ;
    mux21_ni ix27865 (.Y (nx27864), .A0 (inputs_76__6), .A1 (inputs_77__6), .S0 (
             nx24279)) ;
    mux21_ni ix27877 (.Y (nx27876), .A0 (inputs_78__6), .A1 (inputs_79__6), .S0 (
             nx24281)) ;
    mux21_ni ix27945 (.Y (nx27944), .A0 (nx27912), .A1 (nx27940), .S0 (nx23251)
             ) ;
    mux21_ni ix27913 (.Y (nx27912), .A0 (nx27896), .A1 (nx27908), .S0 (nx23577)
             ) ;
    mux21_ni ix27897 (.Y (nx27896), .A0 (inputs_88__6), .A1 (inputs_89__6), .S0 (
             nx24281)) ;
    mux21_ni ix27909 (.Y (nx27908), .A0 (inputs_90__6), .A1 (inputs_91__6), .S0 (
             nx24281)) ;
    mux21_ni ix27941 (.Y (nx27940), .A0 (nx27924), .A1 (nx27936), .S0 (nx23577)
             ) ;
    mux21_ni ix27925 (.Y (nx27924), .A0 (inputs_92__6), .A1 (inputs_93__6), .S0 (
             nx24281)) ;
    mux21_ni ix27937 (.Y (nx27936), .A0 (inputs_94__6), .A1 (inputs_95__6), .S0 (
             nx24281)) ;
    mux21_ni ix28241 (.Y (nx28240), .A0 (nx28234), .A1 (nx28156), .S0 (nx23147)
             ) ;
    oai21 ix28235 (.Y (nx28234), .A0 (nx22289), .A1 (nx14167), .B0 (nx14179)) ;
    mux21 ix14168 (.Y (nx14167), .A0 (nx28198), .A1 (nx28226), .S0 (nx22863)) ;
    mux21_ni ix28199 (.Y (nx28198), .A0 (nx28182), .A1 (nx28194), .S0 (nx23579)
             ) ;
    mux21_ni ix28183 (.Y (nx28182), .A0 (inputs_100__6), .A1 (inputs_101__6), .S0 (
             nx24281)) ;
    mux21_ni ix28195 (.Y (nx28194), .A0 (inputs_102__6), .A1 (inputs_103__6), .S0 (
             nx24281)) ;
    mux21_ni ix28227 (.Y (nx28226), .A0 (nx28210), .A1 (nx28222), .S0 (nx23579)
             ) ;
    mux21_ni ix28211 (.Y (nx28210), .A0 (inputs_116__6), .A1 (inputs_117__6), .S0 (
             nx24283)) ;
    mux21_ni ix28223 (.Y (nx28222), .A0 (inputs_118__6), .A1 (inputs_119__6), .S0 (
             nx24283)) ;
    nand04 ix14180 (.Y (nx14179), .A0 (nx22289), .A1 (nx23579), .A2 (nx24283), .A3 (
           nx28170)) ;
    mux21_ni ix28171 (.Y (nx28170), .A0 (inputs_99__6), .A1 (inputs_115__6), .S0 (
             nx22865)) ;
    mux21_ni ix28157 (.Y (nx28156), .A0 (nx28092), .A1 (nx28152), .S0 (nx22865)
             ) ;
    mux21_ni ix28093 (.Y (nx28092), .A0 (nx28060), .A1 (nx28088), .S0 (nx23251)
             ) ;
    mux21_ni ix28061 (.Y (nx28060), .A0 (nx28044), .A1 (nx28056), .S0 (nx23579)
             ) ;
    mux21_ni ix28045 (.Y (nx28044), .A0 (inputs_104__6), .A1 (inputs_105__6), .S0 (
             nx24283)) ;
    mux21_ni ix28057 (.Y (nx28056), .A0 (inputs_106__6), .A1 (inputs_107__6), .S0 (
             nx24283)) ;
    mux21_ni ix28089 (.Y (nx28088), .A0 (nx28072), .A1 (nx28084), .S0 (nx23579)
             ) ;
    mux21_ni ix28073 (.Y (nx28072), .A0 (inputs_108__6), .A1 (inputs_109__6), .S0 (
             nx24283)) ;
    mux21_ni ix28085 (.Y (nx28084), .A0 (inputs_110__6), .A1 (inputs_111__6), .S0 (
             nx24283)) ;
    mux21_ni ix28153 (.Y (nx28152), .A0 (nx28120), .A1 (nx28148), .S0 (nx23251)
             ) ;
    mux21_ni ix28121 (.Y (nx28120), .A0 (nx28104), .A1 (nx28116), .S0 (nx23579)
             ) ;
    mux21_ni ix28105 (.Y (nx28104), .A0 (inputs_120__6), .A1 (inputs_121__6), .S0 (
             nx24285)) ;
    mux21_ni ix28117 (.Y (nx28116), .A0 (inputs_122__6), .A1 (inputs_123__6), .S0 (
             nx24285)) ;
    mux21_ni ix28149 (.Y (nx28148), .A0 (nx28132), .A1 (nx28144), .S0 (nx23579)
             ) ;
    mux21_ni ix28133 (.Y (nx28132), .A0 (inputs_124__6), .A1 (inputs_125__6), .S0 (
             nx24285)) ;
    mux21_ni ix28145 (.Y (nx28144), .A0 (inputs_126__6), .A1 (inputs_127__6), .S0 (
             nx24285)) ;
    mux21_ni ix29093 (.Y (nx29092), .A0 (nx28668), .A1 (nx29088), .S0 (nx22481)
             ) ;
    mux21_ni ix28669 (.Y (nx28668), .A0 (nx28456), .A1 (nx28664), .S0 (nx22589)
             ) ;
    mux21_ni ix28457 (.Y (nx28456), .A0 (nx28450), .A1 (nx28372), .S0 (nx23147)
             ) ;
    oai21 ix28451 (.Y (nx28450), .A0 (nx22289), .A1 (nx14213), .B0 (nx14225)) ;
    mux21 ix14214 (.Y (nx14213), .A0 (nx28414), .A1 (nx28442), .S0 (nx22865)) ;
    mux21_ni ix28415 (.Y (nx28414), .A0 (nx28398), .A1 (nx28410), .S0 (nx23581)
             ) ;
    mux21_ni ix28399 (.Y (nx28398), .A0 (inputs_132__6), .A1 (inputs_133__6), .S0 (
             nx24285)) ;
    mux21_ni ix28411 (.Y (nx28410), .A0 (inputs_134__6), .A1 (inputs_135__6), .S0 (
             nx24285)) ;
    mux21_ni ix28443 (.Y (nx28442), .A0 (nx28426), .A1 (nx28438), .S0 (nx23581)
             ) ;
    mux21_ni ix28427 (.Y (nx28426), .A0 (inputs_148__6), .A1 (inputs_149__6), .S0 (
             nx24285)) ;
    mux21_ni ix28439 (.Y (nx28438), .A0 (inputs_150__6), .A1 (inputs_151__6), .S0 (
             nx24287)) ;
    nand04 ix14226 (.Y (nx14225), .A0 (nx22291), .A1 (nx23581), .A2 (nx24287), .A3 (
           nx28386)) ;
    mux21_ni ix28387 (.Y (nx28386), .A0 (inputs_131__6), .A1 (inputs_147__6), .S0 (
             nx22865)) ;
    mux21_ni ix28373 (.Y (nx28372), .A0 (nx28308), .A1 (nx28368), .S0 (nx22865)
             ) ;
    mux21_ni ix28309 (.Y (nx28308), .A0 (nx28276), .A1 (nx28304), .S0 (nx23251)
             ) ;
    mux21_ni ix28277 (.Y (nx28276), .A0 (nx28260), .A1 (nx28272), .S0 (nx23581)
             ) ;
    mux21_ni ix28261 (.Y (nx28260), .A0 (inputs_136__6), .A1 (inputs_137__6), .S0 (
             nx24287)) ;
    mux21_ni ix28273 (.Y (nx28272), .A0 (inputs_138__6), .A1 (inputs_139__6), .S0 (
             nx24287)) ;
    mux21_ni ix28305 (.Y (nx28304), .A0 (nx28288), .A1 (nx28300), .S0 (nx23581)
             ) ;
    mux21_ni ix28289 (.Y (nx28288), .A0 (inputs_140__6), .A1 (inputs_141__6), .S0 (
             nx24287)) ;
    mux21_ni ix28301 (.Y (nx28300), .A0 (inputs_142__6), .A1 (inputs_143__6), .S0 (
             nx24287)) ;
    mux21_ni ix28369 (.Y (nx28368), .A0 (nx28336), .A1 (nx28364), .S0 (nx23253)
             ) ;
    mux21_ni ix28337 (.Y (nx28336), .A0 (nx28320), .A1 (nx28332), .S0 (nx23581)
             ) ;
    mux21_ni ix28321 (.Y (nx28320), .A0 (inputs_152__6), .A1 (inputs_153__6), .S0 (
             nx24287)) ;
    mux21_ni ix28333 (.Y (nx28332), .A0 (inputs_154__6), .A1 (inputs_155__6), .S0 (
             nx24289)) ;
    mux21_ni ix28365 (.Y (nx28364), .A0 (nx28348), .A1 (nx28360), .S0 (nx23581)
             ) ;
    mux21_ni ix28349 (.Y (nx28348), .A0 (inputs_156__6), .A1 (inputs_157__6), .S0 (
             nx24289)) ;
    mux21_ni ix28361 (.Y (nx28360), .A0 (inputs_158__6), .A1 (inputs_159__6), .S0 (
             nx24289)) ;
    mux21_ni ix28665 (.Y (nx28664), .A0 (nx28658), .A1 (nx28580), .S0 (nx23147)
             ) ;
    oai21 ix28659 (.Y (nx28658), .A0 (nx22291), .A1 (nx14255), .B0 (nx14267)) ;
    mux21 ix14256 (.Y (nx14255), .A0 (nx28622), .A1 (nx28650), .S0 (nx22865)) ;
    mux21_ni ix28623 (.Y (nx28622), .A0 (nx28606), .A1 (nx28618), .S0 (nx23583)
             ) ;
    mux21_ni ix28607 (.Y (nx28606), .A0 (inputs_164__6), .A1 (inputs_165__6), .S0 (
             nx24289)) ;
    mux21_ni ix28619 (.Y (nx28618), .A0 (inputs_166__6), .A1 (inputs_167__6), .S0 (
             nx24289)) ;
    mux21_ni ix28651 (.Y (nx28650), .A0 (nx28634), .A1 (nx28646), .S0 (nx23583)
             ) ;
    mux21_ni ix28635 (.Y (nx28634), .A0 (inputs_180__6), .A1 (inputs_181__6), .S0 (
             nx24289)) ;
    mux21_ni ix28647 (.Y (nx28646), .A0 (inputs_182__6), .A1 (inputs_183__6), .S0 (
             nx24289)) ;
    nand04 ix14268 (.Y (nx14267), .A0 (nx22291), .A1 (nx23583), .A2 (nx24291), .A3 (
           nx28594)) ;
    mux21_ni ix28595 (.Y (nx28594), .A0 (inputs_163__6), .A1 (inputs_179__6), .S0 (
             nx22865)) ;
    mux21_ni ix28581 (.Y (nx28580), .A0 (nx28516), .A1 (nx28576), .S0 (nx22867)
             ) ;
    mux21_ni ix28517 (.Y (nx28516), .A0 (nx28484), .A1 (nx28512), .S0 (nx23253)
             ) ;
    mux21_ni ix28485 (.Y (nx28484), .A0 (nx28468), .A1 (nx28480), .S0 (nx23583)
             ) ;
    mux21_ni ix28469 (.Y (nx28468), .A0 (inputs_168__6), .A1 (inputs_169__6), .S0 (
             nx24291)) ;
    mux21_ni ix28481 (.Y (nx28480), .A0 (inputs_170__6), .A1 (inputs_171__6), .S0 (
             nx24291)) ;
    mux21_ni ix28513 (.Y (nx28512), .A0 (nx28496), .A1 (nx28508), .S0 (nx23583)
             ) ;
    mux21_ni ix28497 (.Y (nx28496), .A0 (inputs_172__6), .A1 (inputs_173__6), .S0 (
             nx24291)) ;
    mux21_ni ix28509 (.Y (nx28508), .A0 (inputs_174__6), .A1 (inputs_175__6), .S0 (
             nx24291)) ;
    mux21_ni ix28577 (.Y (nx28576), .A0 (nx28544), .A1 (nx28572), .S0 (nx23253)
             ) ;
    mux21_ni ix28545 (.Y (nx28544), .A0 (nx28528), .A1 (nx28540), .S0 (nx23583)
             ) ;
    mux21_ni ix28529 (.Y (nx28528), .A0 (inputs_184__6), .A1 (inputs_185__6), .S0 (
             nx24291)) ;
    mux21_ni ix28541 (.Y (nx28540), .A0 (inputs_186__6), .A1 (inputs_187__6), .S0 (
             nx24291)) ;
    mux21_ni ix28573 (.Y (nx28572), .A0 (nx28556), .A1 (nx28568), .S0 (nx23583)
             ) ;
    mux21_ni ix28557 (.Y (nx28556), .A0 (inputs_188__6), .A1 (inputs_189__6), .S0 (
             nx24293)) ;
    mux21_ni ix28569 (.Y (nx28568), .A0 (inputs_190__6), .A1 (inputs_191__6), .S0 (
             nx24293)) ;
    mux21_ni ix29089 (.Y (nx29088), .A0 (nx28876), .A1 (nx29084), .S0 (nx22589)
             ) ;
    mux21_ni ix28877 (.Y (nx28876), .A0 (nx28870), .A1 (nx28792), .S0 (nx23147)
             ) ;
    oai21 ix28871 (.Y (nx28870), .A0 (nx22291), .A1 (nx14301), .B0 (nx14315)) ;
    mux21 ix14302 (.Y (nx14301), .A0 (nx28834), .A1 (nx28862), .S0 (nx22867)) ;
    mux21_ni ix28835 (.Y (nx28834), .A0 (nx28818), .A1 (nx28830), .S0 (nx23585)
             ) ;
    mux21_ni ix28819 (.Y (nx28818), .A0 (inputs_196__6), .A1 (inputs_197__6), .S0 (
             nx24293)) ;
    mux21_ni ix28831 (.Y (nx28830), .A0 (inputs_198__6), .A1 (inputs_199__6), .S0 (
             nx24293)) ;
    mux21_ni ix28863 (.Y (nx28862), .A0 (nx28846), .A1 (nx28858), .S0 (nx23585)
             ) ;
    mux21_ni ix28847 (.Y (nx28846), .A0 (inputs_212__6), .A1 (inputs_213__6), .S0 (
             nx24293)) ;
    mux21_ni ix28859 (.Y (nx28858), .A0 (inputs_214__6), .A1 (inputs_215__6), .S0 (
             nx24293)) ;
    nand04 ix14316 (.Y (nx14315), .A0 (nx22291), .A1 (nx23585), .A2 (nx24293), .A3 (
           nx28806)) ;
    mux21_ni ix28807 (.Y (nx28806), .A0 (inputs_195__6), .A1 (inputs_211__6), .S0 (
             nx22867)) ;
    mux21_ni ix28793 (.Y (nx28792), .A0 (nx28728), .A1 (nx28788), .S0 (nx22867)
             ) ;
    mux21_ni ix28729 (.Y (nx28728), .A0 (nx28696), .A1 (nx28724), .S0 (nx23253)
             ) ;
    mux21_ni ix28697 (.Y (nx28696), .A0 (nx28680), .A1 (nx28692), .S0 (nx23585)
             ) ;
    mux21_ni ix28681 (.Y (nx28680), .A0 (inputs_200__6), .A1 (inputs_201__6), .S0 (
             nx24295)) ;
    mux21_ni ix28693 (.Y (nx28692), .A0 (inputs_202__6), .A1 (inputs_203__6), .S0 (
             nx24295)) ;
    mux21_ni ix28725 (.Y (nx28724), .A0 (nx28708), .A1 (nx28720), .S0 (nx23585)
             ) ;
    mux21_ni ix28709 (.Y (nx28708), .A0 (inputs_204__6), .A1 (inputs_205__6), .S0 (
             nx24295)) ;
    mux21_ni ix28721 (.Y (nx28720), .A0 (inputs_206__6), .A1 (inputs_207__6), .S0 (
             nx24295)) ;
    mux21_ni ix28789 (.Y (nx28788), .A0 (nx28756), .A1 (nx28784), .S0 (nx23253)
             ) ;
    mux21_ni ix28757 (.Y (nx28756), .A0 (nx28740), .A1 (nx28752), .S0 (nx23585)
             ) ;
    mux21_ni ix28741 (.Y (nx28740), .A0 (inputs_216__6), .A1 (inputs_217__6), .S0 (
             nx24295)) ;
    mux21_ni ix28753 (.Y (nx28752), .A0 (inputs_218__6), .A1 (inputs_219__6), .S0 (
             nx24295)) ;
    mux21_ni ix28785 (.Y (nx28784), .A0 (nx28768), .A1 (nx28780), .S0 (nx23585)
             ) ;
    mux21_ni ix28769 (.Y (nx28768), .A0 (inputs_220__6), .A1 (inputs_221__6), .S0 (
             nx24295)) ;
    mux21_ni ix28781 (.Y (nx28780), .A0 (inputs_222__6), .A1 (inputs_223__6), .S0 (
             nx24297)) ;
    mux21_ni ix29085 (.Y (nx29084), .A0 (nx29078), .A1 (nx29000), .S0 (nx23147)
             ) ;
    oai21 ix29079 (.Y (nx29078), .A0 (nx22291), .A1 (nx14347), .B0 (nx14359)) ;
    mux21 ix14348 (.Y (nx14347), .A0 (nx29042), .A1 (nx29070), .S0 (nx22867)) ;
    mux21_ni ix29043 (.Y (nx29042), .A0 (nx29026), .A1 (nx29038), .S0 (nx23587)
             ) ;
    mux21_ni ix29027 (.Y (nx29026), .A0 (inputs_228__6), .A1 (inputs_229__6), .S0 (
             nx24297)) ;
    mux21_ni ix29039 (.Y (nx29038), .A0 (inputs_230__6), .A1 (inputs_231__6), .S0 (
             nx24297)) ;
    mux21_ni ix29071 (.Y (nx29070), .A0 (nx29054), .A1 (nx29066), .S0 (nx23587)
             ) ;
    mux21_ni ix29055 (.Y (nx29054), .A0 (inputs_244__6), .A1 (inputs_245__6), .S0 (
             nx24297)) ;
    mux21_ni ix29067 (.Y (nx29066), .A0 (inputs_246__6), .A1 (inputs_247__6), .S0 (
             nx24297)) ;
    nand04 ix14360 (.Y (nx14359), .A0 (nx22291), .A1 (nx23587), .A2 (nx24297), .A3 (
           nx29014)) ;
    mux21_ni ix29015 (.Y (nx29014), .A0 (inputs_227__6), .A1 (inputs_243__6), .S0 (
             nx22867)) ;
    mux21_ni ix29001 (.Y (nx29000), .A0 (nx28936), .A1 (nx28996), .S0 (nx22867)
             ) ;
    mux21_ni ix28937 (.Y (nx28936), .A0 (nx28904), .A1 (nx28932), .S0 (nx23253)
             ) ;
    mux21_ni ix28905 (.Y (nx28904), .A0 (nx28888), .A1 (nx28900), .S0 (nx23587)
             ) ;
    mux21_ni ix28889 (.Y (nx28888), .A0 (inputs_232__6), .A1 (inputs_233__6), .S0 (
             nx24297)) ;
    mux21_ni ix28901 (.Y (nx28900), .A0 (inputs_234__6), .A1 (inputs_235__6), .S0 (
             nx24299)) ;
    mux21_ni ix28933 (.Y (nx28932), .A0 (nx28916), .A1 (nx28928), .S0 (nx23587)
             ) ;
    mux21_ni ix28917 (.Y (nx28916), .A0 (inputs_236__6), .A1 (inputs_237__6), .S0 (
             nx24299)) ;
    mux21_ni ix28929 (.Y (nx28928), .A0 (inputs_238__6), .A1 (inputs_239__6), .S0 (
             nx24299)) ;
    mux21_ni ix28997 (.Y (nx28996), .A0 (nx28964), .A1 (nx28992), .S0 (nx23253)
             ) ;
    mux21_ni ix28965 (.Y (nx28964), .A0 (nx28948), .A1 (nx28960), .S0 (nx23587)
             ) ;
    mux21_ni ix28949 (.Y (nx28948), .A0 (inputs_248__6), .A1 (inputs_249__6), .S0 (
             nx24299)) ;
    mux21_ni ix28961 (.Y (nx28960), .A0 (inputs_250__6), .A1 (inputs_251__6), .S0 (
             nx24299)) ;
    mux21_ni ix28993 (.Y (nx28992), .A0 (nx28976), .A1 (nx28988), .S0 (nx23587)
             ) ;
    mux21_ni ix28977 (.Y (nx28976), .A0 (inputs_252__6), .A1 (inputs_253__6), .S0 (
             nx24299)) ;
    mux21_ni ix28989 (.Y (nx28988), .A0 (inputs_254__6), .A1 (inputs_255__6), .S0 (
             nx24299)) ;
    oai21 ix33263 (.Y (\output [7]), .A0 (nx22221), .A1 (nx14387), .B0 (nx14741)
          ) ;
    mux21 ix14388 (.Y (nx14387), .A0 (nx29944), .A1 (nx30788), .S0 (nx22427)) ;
    mux21_ni ix29945 (.Y (nx29944), .A0 (nx29520), .A1 (nx29940), .S0 (nx22483)
             ) ;
    mux21_ni ix29521 (.Y (nx29520), .A0 (nx29308), .A1 (nx29516), .S0 (nx22591)
             ) ;
    mux21_ni ix29309 (.Y (nx29308), .A0 (nx29302), .A1 (nx29224), .S0 (nx23149)
             ) ;
    oai21 ix29303 (.Y (nx29302), .A0 (nx22293), .A1 (nx14395), .B0 (nx14409)) ;
    mux21 ix14396 (.Y (nx14395), .A0 (nx29266), .A1 (nx29294), .S0 (nx22869)) ;
    mux21_ni ix29267 (.Y (nx29266), .A0 (nx29250), .A1 (nx29262), .S0 (nx23589)
             ) ;
    mux21_ni ix29251 (.Y (nx29250), .A0 (inputs_260__7), .A1 (inputs_261__7), .S0 (
             nx24301)) ;
    mux21_ni ix29263 (.Y (nx29262), .A0 (inputs_262__7), .A1 (inputs_263__7), .S0 (
             nx24301)) ;
    mux21_ni ix29295 (.Y (nx29294), .A0 (nx29278), .A1 (nx29290), .S0 (nx23589)
             ) ;
    mux21_ni ix29279 (.Y (nx29278), .A0 (inputs_276__7), .A1 (inputs_277__7), .S0 (
             nx24301)) ;
    mux21_ni ix29291 (.Y (nx29290), .A0 (inputs_278__7), .A1 (inputs_279__7), .S0 (
             nx24301)) ;
    nand04 ix14410 (.Y (nx14409), .A0 (nx22293), .A1 (nx23589), .A2 (nx24301), .A3 (
           nx29238)) ;
    mux21_ni ix29239 (.Y (nx29238), .A0 (inputs_259__7), .A1 (inputs_275__7), .S0 (
             nx22869)) ;
    mux21_ni ix29225 (.Y (nx29224), .A0 (nx29160), .A1 (nx29220), .S0 (nx22869)
             ) ;
    mux21_ni ix29161 (.Y (nx29160), .A0 (nx29128), .A1 (nx29156), .S0 (nx23255)
             ) ;
    mux21_ni ix29129 (.Y (nx29128), .A0 (nx29112), .A1 (nx29124), .S0 (nx23589)
             ) ;
    mux21_ni ix29113 (.Y (nx29112), .A0 (inputs_264__7), .A1 (inputs_265__7), .S0 (
             nx24301)) ;
    mux21_ni ix29125 (.Y (nx29124), .A0 (inputs_266__7), .A1 (inputs_267__7), .S0 (
             nx24301)) ;
    mux21_ni ix29157 (.Y (nx29156), .A0 (nx29140), .A1 (nx29152), .S0 (nx23589)
             ) ;
    mux21_ni ix29141 (.Y (nx29140), .A0 (inputs_268__7), .A1 (inputs_269__7), .S0 (
             nx24303)) ;
    mux21_ni ix29153 (.Y (nx29152), .A0 (inputs_270__7), .A1 (inputs_271__7), .S0 (
             nx24303)) ;
    mux21_ni ix29221 (.Y (nx29220), .A0 (nx29188), .A1 (nx29216), .S0 (nx23255)
             ) ;
    mux21_ni ix29189 (.Y (nx29188), .A0 (nx29172), .A1 (nx29184), .S0 (nx23589)
             ) ;
    mux21_ni ix29173 (.Y (nx29172), .A0 (inputs_280__7), .A1 (inputs_281__7), .S0 (
             nx24303)) ;
    mux21_ni ix29185 (.Y (nx29184), .A0 (inputs_282__7), .A1 (inputs_283__7), .S0 (
             nx24303)) ;
    mux21_ni ix29217 (.Y (nx29216), .A0 (nx29200), .A1 (nx29212), .S0 (nx23589)
             ) ;
    mux21_ni ix29201 (.Y (nx29200), .A0 (inputs_284__7), .A1 (inputs_285__7), .S0 (
             nx24303)) ;
    mux21_ni ix29213 (.Y (nx29212), .A0 (inputs_286__7), .A1 (inputs_287__7), .S0 (
             nx24303)) ;
    mux21_ni ix29517 (.Y (nx29516), .A0 (nx29510), .A1 (nx29432), .S0 (nx23149)
             ) ;
    oai21 ix29511 (.Y (nx29510), .A0 (nx22293), .A1 (nx14439), .B0 (nx14449)) ;
    mux21 ix14440 (.Y (nx14439), .A0 (nx29474), .A1 (nx29502), .S0 (nx22869)) ;
    mux21_ni ix29475 (.Y (nx29474), .A0 (nx29458), .A1 (nx29470), .S0 (nx23591)
             ) ;
    mux21_ni ix29459 (.Y (nx29458), .A0 (inputs_292__7), .A1 (inputs_293__7), .S0 (
             nx24303)) ;
    mux21_ni ix29471 (.Y (nx29470), .A0 (inputs_294__7), .A1 (inputs_295__7), .S0 (
             nx24305)) ;
    mux21_ni ix29503 (.Y (nx29502), .A0 (nx29486), .A1 (nx29498), .S0 (nx23591)
             ) ;
    mux21_ni ix29487 (.Y (nx29486), .A0 (inputs_308__7), .A1 (inputs_309__7), .S0 (
             nx24305)) ;
    mux21_ni ix29499 (.Y (nx29498), .A0 (inputs_310__7), .A1 (inputs_311__7), .S0 (
             nx24305)) ;
    nand04 ix14450 (.Y (nx14449), .A0 (nx22293), .A1 (nx23591), .A2 (nx24305), .A3 (
           nx29446)) ;
    mux21_ni ix29447 (.Y (nx29446), .A0 (inputs_291__7), .A1 (inputs_307__7), .S0 (
             nx22869)) ;
    mux21_ni ix29433 (.Y (nx29432), .A0 (nx29368), .A1 (nx29428), .S0 (nx22869)
             ) ;
    mux21_ni ix29369 (.Y (nx29368), .A0 (nx29336), .A1 (nx29364), .S0 (nx23255)
             ) ;
    mux21_ni ix29337 (.Y (nx29336), .A0 (nx29320), .A1 (nx29332), .S0 (nx23591)
             ) ;
    mux21_ni ix29321 (.Y (nx29320), .A0 (inputs_296__7), .A1 (inputs_297__7), .S0 (
             nx24305)) ;
    mux21_ni ix29333 (.Y (nx29332), .A0 (inputs_298__7), .A1 (inputs_299__7), .S0 (
             nx24305)) ;
    mux21_ni ix29365 (.Y (nx29364), .A0 (nx29348), .A1 (nx29360), .S0 (nx23591)
             ) ;
    mux21_ni ix29349 (.Y (nx29348), .A0 (inputs_300__7), .A1 (inputs_301__7), .S0 (
             nx24305)) ;
    mux21_ni ix29361 (.Y (nx29360), .A0 (inputs_302__7), .A1 (inputs_303__7), .S0 (
             nx24307)) ;
    mux21_ni ix29429 (.Y (nx29428), .A0 (nx29396), .A1 (nx29424), .S0 (nx23255)
             ) ;
    mux21_ni ix29397 (.Y (nx29396), .A0 (nx29380), .A1 (nx29392), .S0 (nx23591)
             ) ;
    mux21_ni ix29381 (.Y (nx29380), .A0 (inputs_312__7), .A1 (inputs_313__7), .S0 (
             nx24307)) ;
    mux21_ni ix29393 (.Y (nx29392), .A0 (inputs_314__7), .A1 (inputs_315__7), .S0 (
             nx24307)) ;
    mux21_ni ix29425 (.Y (nx29424), .A0 (nx29408), .A1 (nx29420), .S0 (nx23591)
             ) ;
    mux21_ni ix29409 (.Y (nx29408), .A0 (inputs_316__7), .A1 (inputs_317__7), .S0 (
             nx24307)) ;
    mux21_ni ix29421 (.Y (nx29420), .A0 (inputs_318__7), .A1 (inputs_319__7), .S0 (
             nx24307)) ;
    mux21_ni ix29941 (.Y (nx29940), .A0 (nx29728), .A1 (nx29936), .S0 (nx22591)
             ) ;
    mux21_ni ix29729 (.Y (nx29728), .A0 (nx29722), .A1 (nx29644), .S0 (nx23149)
             ) ;
    oai21 ix29723 (.Y (nx29722), .A0 (nx22293), .A1 (nx14481), .B0 (nx14493)) ;
    mux21 ix14482 (.Y (nx14481), .A0 (nx29686), .A1 (nx29714), .S0 (nx22869)) ;
    mux21_ni ix29687 (.Y (nx29686), .A0 (nx29670), .A1 (nx29682), .S0 (nx23593)
             ) ;
    mux21_ni ix29671 (.Y (nx29670), .A0 (inputs_324__7), .A1 (inputs_325__7), .S0 (
             nx24307)) ;
    mux21_ni ix29683 (.Y (nx29682), .A0 (inputs_326__7), .A1 (inputs_327__7), .S0 (
             nx24307)) ;
    mux21_ni ix29715 (.Y (nx29714), .A0 (nx29698), .A1 (nx29710), .S0 (nx23593)
             ) ;
    mux21_ni ix29699 (.Y (nx29698), .A0 (inputs_340__7), .A1 (inputs_341__7), .S0 (
             nx24309)) ;
    mux21_ni ix29711 (.Y (nx29710), .A0 (inputs_342__7), .A1 (inputs_343__7), .S0 (
             nx24309)) ;
    nand04 ix14494 (.Y (nx14493), .A0 (nx22293), .A1 (nx23593), .A2 (nx24309), .A3 (
           nx29658)) ;
    mux21_ni ix29659 (.Y (nx29658), .A0 (inputs_323__7), .A1 (inputs_339__7), .S0 (
             nx22871)) ;
    mux21_ni ix29645 (.Y (nx29644), .A0 (nx29580), .A1 (nx29640), .S0 (nx22871)
             ) ;
    mux21_ni ix29581 (.Y (nx29580), .A0 (nx29548), .A1 (nx29576), .S0 (nx23255)
             ) ;
    mux21_ni ix29549 (.Y (nx29548), .A0 (nx29532), .A1 (nx29544), .S0 (nx23593)
             ) ;
    mux21_ni ix29533 (.Y (nx29532), .A0 (inputs_328__7), .A1 (inputs_329__7), .S0 (
             nx24309)) ;
    mux21_ni ix29545 (.Y (nx29544), .A0 (inputs_330__7), .A1 (inputs_331__7), .S0 (
             nx24309)) ;
    mux21_ni ix29577 (.Y (nx29576), .A0 (nx29560), .A1 (nx29572), .S0 (nx23593)
             ) ;
    mux21_ni ix29561 (.Y (nx29560), .A0 (inputs_332__7), .A1 (inputs_333__7), .S0 (
             nx24309)) ;
    mux21_ni ix29573 (.Y (nx29572), .A0 (inputs_334__7), .A1 (inputs_335__7), .S0 (
             nx24309)) ;
    mux21_ni ix29641 (.Y (nx29640), .A0 (nx29608), .A1 (nx29636), .S0 (nx23255)
             ) ;
    mux21_ni ix29609 (.Y (nx29608), .A0 (nx29592), .A1 (nx29604), .S0 (nx23593)
             ) ;
    mux21_ni ix29593 (.Y (nx29592), .A0 (inputs_344__7), .A1 (inputs_345__7), .S0 (
             nx24311)) ;
    mux21_ni ix29605 (.Y (nx29604), .A0 (inputs_346__7), .A1 (inputs_347__7), .S0 (
             nx24311)) ;
    mux21_ni ix29637 (.Y (nx29636), .A0 (nx29620), .A1 (nx29632), .S0 (nx23593)
             ) ;
    mux21_ni ix29621 (.Y (nx29620), .A0 (inputs_348__7), .A1 (inputs_349__7), .S0 (
             nx24311)) ;
    mux21_ni ix29633 (.Y (nx29632), .A0 (inputs_350__7), .A1 (inputs_351__7), .S0 (
             nx24311)) ;
    mux21_ni ix29937 (.Y (nx29936), .A0 (nx29930), .A1 (nx29852), .S0 (nx23149)
             ) ;
    oai21 ix29931 (.Y (nx29930), .A0 (nx22293), .A1 (nx14523), .B0 (nx14537)) ;
    mux21 ix14524 (.Y (nx14523), .A0 (nx29894), .A1 (nx29922), .S0 (nx22871)) ;
    mux21_ni ix29895 (.Y (nx29894), .A0 (nx29878), .A1 (nx29890), .S0 (nx23595)
             ) ;
    mux21_ni ix29879 (.Y (nx29878), .A0 (inputs_356__7), .A1 (inputs_357__7), .S0 (
             nx24311)) ;
    mux21_ni ix29891 (.Y (nx29890), .A0 (inputs_358__7), .A1 (inputs_359__7), .S0 (
             nx24311)) ;
    mux21_ni ix29923 (.Y (nx29922), .A0 (nx29906), .A1 (nx29918), .S0 (nx23595)
             ) ;
    mux21_ni ix29907 (.Y (nx29906), .A0 (inputs_372__7), .A1 (inputs_373__7), .S0 (
             nx24311)) ;
    mux21_ni ix29919 (.Y (nx29918), .A0 (inputs_374__7), .A1 (inputs_375__7), .S0 (
             nx24313)) ;
    nand04 ix14538 (.Y (nx14537), .A0 (nx22295), .A1 (nx23595), .A2 (nx24313), .A3 (
           nx29866)) ;
    mux21_ni ix29867 (.Y (nx29866), .A0 (inputs_355__7), .A1 (inputs_371__7), .S0 (
             nx22871)) ;
    mux21_ni ix29853 (.Y (nx29852), .A0 (nx29788), .A1 (nx29848), .S0 (nx22871)
             ) ;
    mux21_ni ix29789 (.Y (nx29788), .A0 (nx29756), .A1 (nx29784), .S0 (nx23255)
             ) ;
    mux21_ni ix29757 (.Y (nx29756), .A0 (nx29740), .A1 (nx29752), .S0 (nx23595)
             ) ;
    mux21_ni ix29741 (.Y (nx29740), .A0 (inputs_360__7), .A1 (inputs_361__7), .S0 (
             nx24313)) ;
    mux21_ni ix29753 (.Y (nx29752), .A0 (inputs_362__7), .A1 (inputs_363__7), .S0 (
             nx24313)) ;
    mux21_ni ix29785 (.Y (nx29784), .A0 (nx29768), .A1 (nx29780), .S0 (nx23595)
             ) ;
    mux21_ni ix29769 (.Y (nx29768), .A0 (inputs_364__7), .A1 (inputs_365__7), .S0 (
             nx24313)) ;
    mux21_ni ix29781 (.Y (nx29780), .A0 (inputs_366__7), .A1 (inputs_367__7), .S0 (
             nx24313)) ;
    mux21_ni ix29849 (.Y (nx29848), .A0 (nx29816), .A1 (nx29844), .S0 (nx23257)
             ) ;
    mux21_ni ix29817 (.Y (nx29816), .A0 (nx29800), .A1 (nx29812), .S0 (nx23595)
             ) ;
    mux21_ni ix29801 (.Y (nx29800), .A0 (inputs_376__7), .A1 (inputs_377__7), .S0 (
             nx24313)) ;
    mux21_ni ix29813 (.Y (nx29812), .A0 (inputs_378__7), .A1 (inputs_379__7), .S0 (
             nx24315)) ;
    mux21_ni ix29845 (.Y (nx29844), .A0 (nx29828), .A1 (nx29840), .S0 (nx23595)
             ) ;
    mux21_ni ix29829 (.Y (nx29828), .A0 (inputs_380__7), .A1 (inputs_381__7), .S0 (
             nx24315)) ;
    mux21_ni ix29841 (.Y (nx29840), .A0 (inputs_382__7), .A1 (inputs_383__7), .S0 (
             nx24315)) ;
    mux21_ni ix30789 (.Y (nx30788), .A0 (nx30364), .A1 (nx30784), .S0 (nx22483)
             ) ;
    mux21_ni ix30365 (.Y (nx30364), .A0 (nx30152), .A1 (nx30360), .S0 (nx22591)
             ) ;
    mux21_ni ix30153 (.Y (nx30152), .A0 (nx30146), .A1 (nx30068), .S0 (nx23149)
             ) ;
    oai21 ix30147 (.Y (nx30146), .A0 (nx22295), .A1 (nx14569), .B0 (nx14581)) ;
    mux21 ix14570 (.Y (nx14569), .A0 (nx30110), .A1 (nx30138), .S0 (nx22871)) ;
    mux21_ni ix30111 (.Y (nx30110), .A0 (nx30094), .A1 (nx30106), .S0 (nx23597)
             ) ;
    mux21_ni ix30095 (.Y (nx30094), .A0 (inputs_388__7), .A1 (inputs_389__7), .S0 (
             nx24315)) ;
    mux21_ni ix30107 (.Y (nx30106), .A0 (inputs_390__7), .A1 (inputs_391__7), .S0 (
             nx24315)) ;
    mux21_ni ix30139 (.Y (nx30138), .A0 (nx30122), .A1 (nx30134), .S0 (nx23597)
             ) ;
    mux21_ni ix30123 (.Y (nx30122), .A0 (inputs_404__7), .A1 (inputs_405__7), .S0 (
             nx24315)) ;
    mux21_ni ix30135 (.Y (nx30134), .A0 (inputs_406__7), .A1 (inputs_407__7), .S0 (
             nx24315)) ;
    nand04 ix14582 (.Y (nx14581), .A0 (nx22295), .A1 (nx23597), .A2 (nx24317), .A3 (
           nx30082)) ;
    mux21_ni ix30083 (.Y (nx30082), .A0 (inputs_387__7), .A1 (inputs_403__7), .S0 (
             nx22871)) ;
    mux21_ni ix30069 (.Y (nx30068), .A0 (nx30004), .A1 (nx30064), .S0 (nx22873)
             ) ;
    mux21_ni ix30005 (.Y (nx30004), .A0 (nx29972), .A1 (nx30000), .S0 (nx23257)
             ) ;
    mux21_ni ix29973 (.Y (nx29972), .A0 (nx29956), .A1 (nx29968), .S0 (nx23597)
             ) ;
    mux21_ni ix29957 (.Y (nx29956), .A0 (inputs_392__7), .A1 (inputs_393__7), .S0 (
             nx24317)) ;
    mux21_ni ix29969 (.Y (nx29968), .A0 (inputs_394__7), .A1 (inputs_395__7), .S0 (
             nx24317)) ;
    mux21_ni ix30001 (.Y (nx30000), .A0 (nx29984), .A1 (nx29996), .S0 (nx23597)
             ) ;
    mux21_ni ix29985 (.Y (nx29984), .A0 (inputs_396__7), .A1 (inputs_397__7), .S0 (
             nx24317)) ;
    mux21_ni ix29997 (.Y (nx29996), .A0 (inputs_398__7), .A1 (inputs_399__7), .S0 (
             nx24317)) ;
    mux21_ni ix30065 (.Y (nx30064), .A0 (nx30032), .A1 (nx30060), .S0 (nx23257)
             ) ;
    mux21_ni ix30033 (.Y (nx30032), .A0 (nx30016), .A1 (nx30028), .S0 (nx23597)
             ) ;
    mux21_ni ix30017 (.Y (nx30016), .A0 (inputs_408__7), .A1 (inputs_409__7), .S0 (
             nx24317)) ;
    mux21_ni ix30029 (.Y (nx30028), .A0 (inputs_410__7), .A1 (inputs_411__7), .S0 (
             nx24317)) ;
    mux21_ni ix30061 (.Y (nx30060), .A0 (nx30044), .A1 (nx30056), .S0 (nx23597)
             ) ;
    mux21_ni ix30045 (.Y (nx30044), .A0 (inputs_412__7), .A1 (inputs_413__7), .S0 (
             nx24319)) ;
    mux21_ni ix30057 (.Y (nx30056), .A0 (inputs_414__7), .A1 (inputs_415__7), .S0 (
             nx24319)) ;
    mux21_ni ix30361 (.Y (nx30360), .A0 (nx30354), .A1 (nx30276), .S0 (nx23149)
             ) ;
    oai21 ix30355 (.Y (nx30354), .A0 (nx22295), .A1 (nx14613), .B0 (nx14625)) ;
    mux21 ix14614 (.Y (nx14613), .A0 (nx30318), .A1 (nx30346), .S0 (nx22873)) ;
    mux21_ni ix30319 (.Y (nx30318), .A0 (nx30302), .A1 (nx30314), .S0 (nx23599)
             ) ;
    mux21_ni ix30303 (.Y (nx30302), .A0 (inputs_420__7), .A1 (inputs_421__7), .S0 (
             nx24319)) ;
    mux21_ni ix30315 (.Y (nx30314), .A0 (inputs_422__7), .A1 (inputs_423__7), .S0 (
             nx24319)) ;
    mux21_ni ix30347 (.Y (nx30346), .A0 (nx30330), .A1 (nx30342), .S0 (nx23599)
             ) ;
    mux21_ni ix30331 (.Y (nx30330), .A0 (inputs_436__7), .A1 (inputs_437__7), .S0 (
             nx24319)) ;
    mux21_ni ix30343 (.Y (nx30342), .A0 (inputs_438__7), .A1 (inputs_439__7), .S0 (
             nx24319)) ;
    nand04 ix14626 (.Y (nx14625), .A0 (nx22295), .A1 (nx23599), .A2 (nx24319), .A3 (
           nx30290)) ;
    mux21_ni ix30291 (.Y (nx30290), .A0 (inputs_419__7), .A1 (inputs_435__7), .S0 (
             nx22873)) ;
    mux21_ni ix30277 (.Y (nx30276), .A0 (nx30212), .A1 (nx30272), .S0 (nx22873)
             ) ;
    mux21_ni ix30213 (.Y (nx30212), .A0 (nx30180), .A1 (nx30208), .S0 (nx23257)
             ) ;
    mux21_ni ix30181 (.Y (nx30180), .A0 (nx30164), .A1 (nx30176), .S0 (nx23599)
             ) ;
    mux21_ni ix30165 (.Y (nx30164), .A0 (inputs_424__7), .A1 (inputs_425__7), .S0 (
             nx24321)) ;
    mux21_ni ix30177 (.Y (nx30176), .A0 (inputs_426__7), .A1 (inputs_427__7), .S0 (
             nx24321)) ;
    mux21_ni ix30209 (.Y (nx30208), .A0 (nx30192), .A1 (nx30204), .S0 (nx23599)
             ) ;
    mux21_ni ix30193 (.Y (nx30192), .A0 (inputs_428__7), .A1 (inputs_429__7), .S0 (
             nx24321)) ;
    mux21_ni ix30205 (.Y (nx30204), .A0 (inputs_430__7), .A1 (inputs_431__7), .S0 (
             nx24321)) ;
    mux21_ni ix30273 (.Y (nx30272), .A0 (nx30240), .A1 (nx30268), .S0 (nx23257)
             ) ;
    mux21_ni ix30241 (.Y (nx30240), .A0 (nx30224), .A1 (nx30236), .S0 (nx23599)
             ) ;
    mux21_ni ix30225 (.Y (nx30224), .A0 (inputs_440__7), .A1 (inputs_441__7), .S0 (
             nx24321)) ;
    mux21_ni ix30237 (.Y (nx30236), .A0 (inputs_442__7), .A1 (inputs_443__7), .S0 (
             nx24321)) ;
    mux21_ni ix30269 (.Y (nx30268), .A0 (nx30252), .A1 (nx30264), .S0 (nx23599)
             ) ;
    mux21_ni ix30253 (.Y (nx30252), .A0 (inputs_444__7), .A1 (inputs_445__7), .S0 (
             nx24321)) ;
    mux21_ni ix30265 (.Y (nx30264), .A0 (inputs_446__7), .A1 (inputs_447__7), .S0 (
             nx24323)) ;
    mux21_ni ix30785 (.Y (nx30784), .A0 (nx30572), .A1 (nx30780), .S0 (nx22591)
             ) ;
    mux21_ni ix30573 (.Y (nx30572), .A0 (nx30566), .A1 (nx30488), .S0 (nx23149)
             ) ;
    oai21 ix30567 (.Y (nx30566), .A0 (nx22295), .A1 (nx14657), .B0 (nx14669)) ;
    mux21 ix14658 (.Y (nx14657), .A0 (nx30530), .A1 (nx30558), .S0 (nx22873)) ;
    mux21_ni ix30531 (.Y (nx30530), .A0 (nx30514), .A1 (nx30526), .S0 (nx23601)
             ) ;
    mux21_ni ix30515 (.Y (nx30514), .A0 (inputs_452__7), .A1 (inputs_453__7), .S0 (
             nx24323)) ;
    mux21_ni ix30527 (.Y (nx30526), .A0 (inputs_454__7), .A1 (inputs_455__7), .S0 (
             nx24323)) ;
    mux21_ni ix30559 (.Y (nx30558), .A0 (nx30542), .A1 (nx30554), .S0 (nx23601)
             ) ;
    mux21_ni ix30543 (.Y (nx30542), .A0 (inputs_468__7), .A1 (inputs_469__7), .S0 (
             nx24323)) ;
    mux21_ni ix30555 (.Y (nx30554), .A0 (inputs_470__7), .A1 (inputs_471__7), .S0 (
             nx24323)) ;
    nand04 ix14670 (.Y (nx14669), .A0 (nx22295), .A1 (nx23601), .A2 (nx24323), .A3 (
           nx30502)) ;
    mux21_ni ix30503 (.Y (nx30502), .A0 (inputs_451__7), .A1 (inputs_467__7), .S0 (
             nx22873)) ;
    mux21_ni ix30489 (.Y (nx30488), .A0 (nx30424), .A1 (nx30484), .S0 (nx22873)
             ) ;
    mux21_ni ix30425 (.Y (nx30424), .A0 (nx30392), .A1 (nx30420), .S0 (nx23257)
             ) ;
    mux21_ni ix30393 (.Y (nx30392), .A0 (nx30376), .A1 (nx30388), .S0 (nx23601)
             ) ;
    mux21_ni ix30377 (.Y (nx30376), .A0 (inputs_456__7), .A1 (inputs_457__7), .S0 (
             nx24323)) ;
    mux21_ni ix30389 (.Y (nx30388), .A0 (inputs_458__7), .A1 (inputs_459__7), .S0 (
             nx24325)) ;
    mux21_ni ix30421 (.Y (nx30420), .A0 (nx30404), .A1 (nx30416), .S0 (nx23601)
             ) ;
    mux21_ni ix30405 (.Y (nx30404), .A0 (inputs_460__7), .A1 (inputs_461__7), .S0 (
             nx24325)) ;
    mux21_ni ix30417 (.Y (nx30416), .A0 (inputs_462__7), .A1 (inputs_463__7), .S0 (
             nx24325)) ;
    mux21_ni ix30485 (.Y (nx30484), .A0 (nx30452), .A1 (nx30480), .S0 (nx23257)
             ) ;
    mux21_ni ix30453 (.Y (nx30452), .A0 (nx30436), .A1 (nx30448), .S0 (nx23601)
             ) ;
    mux21_ni ix30437 (.Y (nx30436), .A0 (inputs_472__7), .A1 (inputs_473__7), .S0 (
             nx24325)) ;
    mux21_ni ix30449 (.Y (nx30448), .A0 (inputs_474__7), .A1 (inputs_475__7), .S0 (
             nx24325)) ;
    mux21_ni ix30481 (.Y (nx30480), .A0 (nx30464), .A1 (nx30476), .S0 (nx23601)
             ) ;
    mux21_ni ix30465 (.Y (nx30464), .A0 (inputs_476__7), .A1 (inputs_477__7), .S0 (
             nx24325)) ;
    mux21_ni ix30477 (.Y (nx30476), .A0 (inputs_478__7), .A1 (inputs_479__7), .S0 (
             nx24325)) ;
    mux21_ni ix30781 (.Y (nx30780), .A0 (nx30774), .A1 (nx30696), .S0 (nx23151)
             ) ;
    oai21 ix30775 (.Y (nx30774), .A0 (nx22297), .A1 (nx14699), .B0 (nx14711)) ;
    mux21 ix14700 (.Y (nx14699), .A0 (nx30738), .A1 (nx30766), .S0 (nx22875)) ;
    mux21_ni ix30739 (.Y (nx30738), .A0 (nx30722), .A1 (nx30734), .S0 (nx23603)
             ) ;
    mux21_ni ix30723 (.Y (nx30722), .A0 (inputs_484__7), .A1 (inputs_485__7), .S0 (
             nx24327)) ;
    mux21_ni ix30735 (.Y (nx30734), .A0 (inputs_486__7), .A1 (inputs_487__7), .S0 (
             nx24327)) ;
    mux21_ni ix30767 (.Y (nx30766), .A0 (nx30750), .A1 (nx30762), .S0 (nx23603)
             ) ;
    mux21_ni ix30751 (.Y (nx30750), .A0 (inputs_500__7), .A1 (inputs_501__7), .S0 (
             nx24327)) ;
    mux21_ni ix30763 (.Y (nx30762), .A0 (inputs_502__7), .A1 (inputs_503__7), .S0 (
             nx24327)) ;
    nand04 ix14712 (.Y (nx14711), .A0 (nx22297), .A1 (nx23603), .A2 (nx24327), .A3 (
           nx30710)) ;
    mux21_ni ix30711 (.Y (nx30710), .A0 (inputs_483__7), .A1 (inputs_499__7), .S0 (
             nx22875)) ;
    mux21_ni ix30697 (.Y (nx30696), .A0 (nx30632), .A1 (nx30692), .S0 (nx22875)
             ) ;
    mux21_ni ix30633 (.Y (nx30632), .A0 (nx30600), .A1 (nx30628), .S0 (nx23259)
             ) ;
    mux21_ni ix30601 (.Y (nx30600), .A0 (nx30584), .A1 (nx30596), .S0 (nx23603)
             ) ;
    mux21_ni ix30585 (.Y (nx30584), .A0 (inputs_488__7), .A1 (inputs_489__7), .S0 (
             nx24327)) ;
    mux21_ni ix30597 (.Y (nx30596), .A0 (inputs_490__7), .A1 (inputs_491__7), .S0 (
             nx24327)) ;
    mux21_ni ix30629 (.Y (nx30628), .A0 (nx30612), .A1 (nx30624), .S0 (nx23603)
             ) ;
    mux21_ni ix30613 (.Y (nx30612), .A0 (inputs_492__7), .A1 (inputs_493__7), .S0 (
             nx24329)) ;
    mux21_ni ix30625 (.Y (nx30624), .A0 (inputs_494__7), .A1 (inputs_495__7), .S0 (
             nx24329)) ;
    mux21_ni ix30693 (.Y (nx30692), .A0 (nx30660), .A1 (nx30688), .S0 (nx23259)
             ) ;
    mux21_ni ix30661 (.Y (nx30660), .A0 (nx30644), .A1 (nx30656), .S0 (nx23603)
             ) ;
    mux21_ni ix30645 (.Y (nx30644), .A0 (inputs_504__7), .A1 (inputs_505__7), .S0 (
             nx24329)) ;
    mux21_ni ix30657 (.Y (nx30656), .A0 (inputs_506__7), .A1 (inputs_507__7), .S0 (
             nx24329)) ;
    mux21_ni ix30689 (.Y (nx30688), .A0 (nx30672), .A1 (nx30684), .S0 (nx23603)
             ) ;
    mux21_ni ix30673 (.Y (nx30672), .A0 (inputs_508__7), .A1 (inputs_509__7), .S0 (
             nx24329)) ;
    mux21_ni ix30685 (.Y (nx30684), .A0 (inputs_510__7), .A1 (inputs_511__7), .S0 (
             nx24329)) ;
    aoi32 ix14742 (.Y (nx14741), .A0 (nx31558), .A1 (nx22387), .A2 (nx22297), .B0 (
          nx22221), .B1 (nx33254)) ;
    oai21 ix31559 (.Y (nx31558), .A0 (nx23605), .A1 (nx14745), .B0 (nx14847)) ;
    mux21 ix14746 (.Y (nx14745), .A0 (nx31296), .A1 (nx31548), .S0 (nx24329)) ;
    mux21_ni ix31297 (.Y (nx31296), .A0 (nx31168), .A1 (nx31292), .S0 (nx22399)
             ) ;
    mux21_ni ix31169 (.Y (nx31168), .A0 (nx31104), .A1 (nx31164), .S0 (nx22427)
             ) ;
    mux21_ni ix31105 (.Y (nx31104), .A0 (nx31072), .A1 (nx31100), .S0 (nx22483)
             ) ;
    mux21_ni ix31073 (.Y (nx31072), .A0 (nx31056), .A1 (nx31068), .S0 (nx22591)
             ) ;
    mux21_ni ix31057 (.Y (nx31056), .A0 (inputs_0__7), .A1 (inputs_16__7), .S0 (
             nx22875)) ;
    mux21_ni ix31069 (.Y (nx31068), .A0 (inputs_32__7), .A1 (inputs_48__7), .S0 (
             nx22875)) ;
    mux21_ni ix31101 (.Y (nx31100), .A0 (nx31084), .A1 (nx31096), .S0 (nx22591)
             ) ;
    mux21_ni ix31085 (.Y (nx31084), .A0 (inputs_64__7), .A1 (inputs_80__7), .S0 (
             nx22875)) ;
    mux21_ni ix31097 (.Y (nx31096), .A0 (inputs_96__7), .A1 (inputs_112__7), .S0 (
             nx22875)) ;
    mux21_ni ix31165 (.Y (nx31164), .A0 (nx31132), .A1 (nx31160), .S0 (nx22483)
             ) ;
    mux21_ni ix31133 (.Y (nx31132), .A0 (nx31116), .A1 (nx31128), .S0 (nx22591)
             ) ;
    mux21_ni ix31117 (.Y (nx31116), .A0 (inputs_128__7), .A1 (inputs_144__7), .S0 (
             nx22877)) ;
    mux21_ni ix31129 (.Y (nx31128), .A0 (inputs_160__7), .A1 (inputs_176__7), .S0 (
             nx22877)) ;
    mux21_ni ix31161 (.Y (nx31160), .A0 (nx31144), .A1 (nx31156), .S0 (nx22593)
             ) ;
    mux21_ni ix31145 (.Y (nx31144), .A0 (inputs_192__7), .A1 (inputs_208__7), .S0 (
             nx22877)) ;
    mux21_ni ix31157 (.Y (nx31156), .A0 (inputs_224__7), .A1 (inputs_240__7), .S0 (
             nx22877)) ;
    mux21_ni ix31293 (.Y (nx31292), .A0 (nx31228), .A1 (nx31288), .S0 (nx22427)
             ) ;
    mux21_ni ix31229 (.Y (nx31228), .A0 (nx31196), .A1 (nx31224), .S0 (nx22483)
             ) ;
    mux21_ni ix31197 (.Y (nx31196), .A0 (nx31180), .A1 (nx31192), .S0 (nx22593)
             ) ;
    mux21_ni ix31181 (.Y (nx31180), .A0 (inputs_256__7), .A1 (inputs_272__7), .S0 (
             nx22877)) ;
    mux21_ni ix31193 (.Y (nx31192), .A0 (inputs_288__7), .A1 (inputs_304__7), .S0 (
             nx22877)) ;
    mux21_ni ix31225 (.Y (nx31224), .A0 (nx31208), .A1 (nx31220), .S0 (nx22593)
             ) ;
    mux21_ni ix31209 (.Y (nx31208), .A0 (inputs_320__7), .A1 (inputs_336__7), .S0 (
             nx22877)) ;
    mux21_ni ix31221 (.Y (nx31220), .A0 (inputs_352__7), .A1 (inputs_368__7), .S0 (
             nx22879)) ;
    mux21_ni ix31289 (.Y (nx31288), .A0 (nx31256), .A1 (nx31284), .S0 (nx22483)
             ) ;
    mux21_ni ix31257 (.Y (nx31256), .A0 (nx31240), .A1 (nx31252), .S0 (nx22593)
             ) ;
    mux21_ni ix31241 (.Y (nx31240), .A0 (inputs_384__7), .A1 (inputs_400__7), .S0 (
             nx22879)) ;
    mux21_ni ix31253 (.Y (nx31252), .A0 (inputs_416__7), .A1 (inputs_432__7), .S0 (
             nx22879)) ;
    mux21_ni ix31285 (.Y (nx31284), .A0 (nx31268), .A1 (nx31280), .S0 (nx22593)
             ) ;
    mux21_ni ix31269 (.Y (nx31268), .A0 (inputs_448__7), .A1 (inputs_464__7), .S0 (
             nx22879)) ;
    mux21_ni ix31281 (.Y (nx31280), .A0 (inputs_480__7), .A1 (inputs_496__7), .S0 (
             nx22879)) ;
    mux21_ni ix31549 (.Y (nx31548), .A0 (nx31420), .A1 (nx31544), .S0 (nx22399)
             ) ;
    mux21_ni ix31421 (.Y (nx31420), .A0 (nx31356), .A1 (nx31416), .S0 (nx22427)
             ) ;
    mux21_ni ix31357 (.Y (nx31356), .A0 (nx31324), .A1 (nx31352), .S0 (nx22483)
             ) ;
    mux21_ni ix31325 (.Y (nx31324), .A0 (nx31308), .A1 (nx31320), .S0 (nx22593)
             ) ;
    mux21_ni ix31309 (.Y (nx31308), .A0 (inputs_1__7), .A1 (inputs_17__7), .S0 (
             nx22879)) ;
    mux21_ni ix31321 (.Y (nx31320), .A0 (inputs_33__7), .A1 (inputs_49__7), .S0 (
             nx22879)) ;
    mux21_ni ix31353 (.Y (nx31352), .A0 (nx31336), .A1 (nx31348), .S0 (nx22593)
             ) ;
    mux21_ni ix31337 (.Y (nx31336), .A0 (inputs_65__7), .A1 (inputs_81__7), .S0 (
             nx22881)) ;
    mux21_ni ix31349 (.Y (nx31348), .A0 (inputs_97__7), .A1 (inputs_113__7), .S0 (
             nx22881)) ;
    mux21_ni ix31417 (.Y (nx31416), .A0 (nx31384), .A1 (nx31412), .S0 (nx22485)
             ) ;
    mux21_ni ix31385 (.Y (nx31384), .A0 (nx31368), .A1 (nx31380), .S0 (nx22595)
             ) ;
    mux21_ni ix31369 (.Y (nx31368), .A0 (inputs_129__7), .A1 (inputs_145__7), .S0 (
             nx22881)) ;
    mux21_ni ix31381 (.Y (nx31380), .A0 (inputs_161__7), .A1 (inputs_177__7), .S0 (
             nx22881)) ;
    mux21_ni ix31413 (.Y (nx31412), .A0 (nx31396), .A1 (nx31408), .S0 (nx22595)
             ) ;
    mux21_ni ix31397 (.Y (nx31396), .A0 (inputs_193__7), .A1 (inputs_209__7), .S0 (
             nx22881)) ;
    mux21_ni ix31409 (.Y (nx31408), .A0 (inputs_225__7), .A1 (inputs_241__7), .S0 (
             nx22881)) ;
    mux21_ni ix31545 (.Y (nx31544), .A0 (nx31480), .A1 (nx31540), .S0 (nx22427)
             ) ;
    mux21_ni ix31481 (.Y (nx31480), .A0 (nx31448), .A1 (nx31476), .S0 (nx22485)
             ) ;
    mux21_ni ix31449 (.Y (nx31448), .A0 (nx31432), .A1 (nx31444), .S0 (nx22595)
             ) ;
    mux21_ni ix31433 (.Y (nx31432), .A0 (inputs_257__7), .A1 (inputs_273__7), .S0 (
             nx22881)) ;
    mux21_ni ix31445 (.Y (nx31444), .A0 (inputs_289__7), .A1 (inputs_305__7), .S0 (
             nx22883)) ;
    mux21_ni ix31477 (.Y (nx31476), .A0 (nx31460), .A1 (nx31472), .S0 (nx22595)
             ) ;
    mux21_ni ix31461 (.Y (nx31460), .A0 (inputs_321__7), .A1 (inputs_337__7), .S0 (
             nx22883)) ;
    mux21_ni ix31473 (.Y (nx31472), .A0 (inputs_353__7), .A1 (inputs_369__7), .S0 (
             nx22883)) ;
    mux21_ni ix31541 (.Y (nx31540), .A0 (nx31508), .A1 (nx31536), .S0 (nx22485)
             ) ;
    mux21_ni ix31509 (.Y (nx31508), .A0 (nx31492), .A1 (nx31504), .S0 (nx22595)
             ) ;
    mux21_ni ix31493 (.Y (nx31492), .A0 (inputs_385__7), .A1 (inputs_401__7), .S0 (
             nx22883)) ;
    mux21_ni ix31505 (.Y (nx31504), .A0 (inputs_417__7), .A1 (inputs_433__7), .S0 (
             nx22883)) ;
    mux21_ni ix31537 (.Y (nx31536), .A0 (nx31520), .A1 (nx31532), .S0 (nx22595)
             ) ;
    mux21_ni ix31521 (.Y (nx31520), .A0 (inputs_449__7), .A1 (inputs_465__7), .S0 (
             nx22883)) ;
    mux21_ni ix31533 (.Y (nx31532), .A0 (inputs_481__7), .A1 (inputs_497__7), .S0 (
             nx22883)) ;
    nand03 ix14848 (.Y (nx14847), .A0 (nx31042), .A1 (nx23605), .A2 (nx22381)) ;
    mux21_ni ix31043 (.Y (nx31042), .A0 (nx30914), .A1 (nx31038), .S0 (nx22399)
             ) ;
    mux21_ni ix30915 (.Y (nx30914), .A0 (nx30850), .A1 (nx30910), .S0 (nx22427)
             ) ;
    mux21_ni ix30851 (.Y (nx30850), .A0 (nx30818), .A1 (nx30846), .S0 (nx22485)
             ) ;
    mux21_ni ix30819 (.Y (nx30818), .A0 (nx30802), .A1 (nx30814), .S0 (nx22595)
             ) ;
    mux21_ni ix30803 (.Y (nx30802), .A0 (inputs_2__7), .A1 (inputs_18__7), .S0 (
             nx22885)) ;
    mux21_ni ix30815 (.Y (nx30814), .A0 (inputs_34__7), .A1 (inputs_50__7), .S0 (
             nx22885)) ;
    mux21_ni ix30847 (.Y (nx30846), .A0 (nx30830), .A1 (nx30842), .S0 (nx22597)
             ) ;
    mux21_ni ix30831 (.Y (nx30830), .A0 (inputs_66__7), .A1 (inputs_82__7), .S0 (
             nx22885)) ;
    mux21_ni ix30843 (.Y (nx30842), .A0 (inputs_98__7), .A1 (inputs_114__7), .S0 (
             nx22885)) ;
    mux21_ni ix30911 (.Y (nx30910), .A0 (nx30878), .A1 (nx30906), .S0 (nx22485)
             ) ;
    mux21_ni ix30879 (.Y (nx30878), .A0 (nx30862), .A1 (nx30874), .S0 (nx22597)
             ) ;
    mux21_ni ix30863 (.Y (nx30862), .A0 (inputs_130__7), .A1 (inputs_146__7), .S0 (
             nx22885)) ;
    mux21_ni ix30875 (.Y (nx30874), .A0 (inputs_162__7), .A1 (inputs_178__7), .S0 (
             nx22885)) ;
    mux21_ni ix30907 (.Y (nx30906), .A0 (nx30890), .A1 (nx30902), .S0 (nx22597)
             ) ;
    mux21_ni ix30891 (.Y (nx30890), .A0 (inputs_194__7), .A1 (inputs_210__7), .S0 (
             nx22885)) ;
    mux21_ni ix30903 (.Y (nx30902), .A0 (inputs_226__7), .A1 (inputs_242__7), .S0 (
             nx22887)) ;
    mux21_ni ix31039 (.Y (nx31038), .A0 (nx30974), .A1 (nx31034), .S0 (nx22427)
             ) ;
    mux21_ni ix30975 (.Y (nx30974), .A0 (nx30942), .A1 (nx30970), .S0 (nx22485)
             ) ;
    mux21_ni ix30943 (.Y (nx30942), .A0 (nx30926), .A1 (nx30938), .S0 (nx22597)
             ) ;
    mux21_ni ix30927 (.Y (nx30926), .A0 (inputs_258__7), .A1 (inputs_274__7), .S0 (
             nx22887)) ;
    mux21_ni ix30939 (.Y (nx30938), .A0 (inputs_290__7), .A1 (inputs_306__7), .S0 (
             nx22887)) ;
    mux21_ni ix30971 (.Y (nx30970), .A0 (nx30954), .A1 (nx30966), .S0 (nx22597)
             ) ;
    mux21_ni ix30955 (.Y (nx30954), .A0 (inputs_322__7), .A1 (inputs_338__7), .S0 (
             nx22887)) ;
    mux21_ni ix30967 (.Y (nx30966), .A0 (inputs_354__7), .A1 (inputs_370__7), .S0 (
             nx22887)) ;
    mux21_ni ix31035 (.Y (nx31034), .A0 (nx31002), .A1 (nx31030), .S0 (nx22485)
             ) ;
    mux21_ni ix31003 (.Y (nx31002), .A0 (nx30986), .A1 (nx30998), .S0 (nx22597)
             ) ;
    mux21_ni ix30987 (.Y (nx30986), .A0 (inputs_386__7), .A1 (inputs_402__7), .S0 (
             nx22887)) ;
    mux21_ni ix30999 (.Y (nx30998), .A0 (inputs_418__7), .A1 (inputs_434__7), .S0 (
             nx22887)) ;
    mux21_ni ix31031 (.Y (nx31030), .A0 (nx31014), .A1 (nx31026), .S0 (nx22597)
             ) ;
    mux21_ni ix31015 (.Y (nx31014), .A0 (inputs_450__7), .A1 (inputs_466__7), .S0 (
             nx22889)) ;
    mux21_ni ix31027 (.Y (nx31026), .A0 (inputs_482__7), .A1 (inputs_498__7), .S0 (
             nx22889)) ;
    mux21_ni ix33255 (.Y (nx33254), .A0 (nx32406), .A1 (nx33250), .S0 (nx22429)
             ) ;
    mux21_ni ix32407 (.Y (nx32406), .A0 (nx31982), .A1 (nx32402), .S0 (nx22487)
             ) ;
    mux21_ni ix31983 (.Y (nx31982), .A0 (nx31770), .A1 (nx31978), .S0 (nx22599)
             ) ;
    mux21_ni ix31771 (.Y (nx31770), .A0 (nx31764), .A1 (nx31686), .S0 (nx23151)
             ) ;
    oai21 ix31765 (.Y (nx31764), .A0 (nx22297), .A1 (nx14905), .B0 (nx14919)) ;
    mux21 ix14906 (.Y (nx14905), .A0 (nx31728), .A1 (nx31756), .S0 (nx22889)) ;
    mux21_ni ix31729 (.Y (nx31728), .A0 (nx31712), .A1 (nx31724), .S0 (nx23605)
             ) ;
    mux21_ni ix31713 (.Y (nx31712), .A0 (inputs_4__7), .A1 (inputs_5__7), .S0 (
             nx24331)) ;
    mux21_ni ix31725 (.Y (nx31724), .A0 (inputs_6__7), .A1 (inputs_7__7), .S0 (
             nx24331)) ;
    mux21_ni ix31757 (.Y (nx31756), .A0 (nx31740), .A1 (nx31752), .S0 (nx23605)
             ) ;
    mux21_ni ix31741 (.Y (nx31740), .A0 (inputs_20__7), .A1 (inputs_21__7), .S0 (
             nx24331)) ;
    mux21_ni ix31753 (.Y (nx31752), .A0 (inputs_22__7), .A1 (inputs_23__7), .S0 (
             nx24331)) ;
    nand04 ix14920 (.Y (nx14919), .A0 (nx22297), .A1 (nx23605), .A2 (nx24331), .A3 (
           nx31700)) ;
    mux21_ni ix31701 (.Y (nx31700), .A0 (inputs_3__7), .A1 (inputs_19__7), .S0 (
             nx22889)) ;
    mux21_ni ix31687 (.Y (nx31686), .A0 (nx31622), .A1 (nx31682), .S0 (nx22889)
             ) ;
    mux21_ni ix31623 (.Y (nx31622), .A0 (nx31590), .A1 (nx31618), .S0 (nx23259)
             ) ;
    mux21_ni ix31591 (.Y (nx31590), .A0 (nx31574), .A1 (nx31586), .S0 (nx23605)
             ) ;
    mux21_ni ix31575 (.Y (nx31574), .A0 (inputs_8__7), .A1 (inputs_9__7), .S0 (
             nx24331)) ;
    mux21_ni ix31587 (.Y (nx31586), .A0 (inputs_10__7), .A1 (inputs_11__7), .S0 (
             nx24331)) ;
    mux21_ni ix31619 (.Y (nx31618), .A0 (nx31602), .A1 (nx31614), .S0 (nx23605)
             ) ;
    mux21_ni ix31603 (.Y (nx31602), .A0 (inputs_12__7), .A1 (inputs_13__7), .S0 (
             nx24333)) ;
    mux21_ni ix31615 (.Y (nx31614), .A0 (inputs_14__7), .A1 (inputs_15__7), .S0 (
             nx24333)) ;
    mux21_ni ix31683 (.Y (nx31682), .A0 (nx31650), .A1 (nx31678), .S0 (nx23259)
             ) ;
    mux21_ni ix31651 (.Y (nx31650), .A0 (nx31634), .A1 (nx31646), .S0 (nx23607)
             ) ;
    mux21_ni ix31635 (.Y (nx31634), .A0 (inputs_24__7), .A1 (inputs_25__7), .S0 (
             nx24333)) ;
    mux21_ni ix31647 (.Y (nx31646), .A0 (inputs_26__7), .A1 (inputs_27__7), .S0 (
             nx24333)) ;
    mux21_ni ix31679 (.Y (nx31678), .A0 (nx31662), .A1 (nx31674), .S0 (nx23607)
             ) ;
    mux21_ni ix31663 (.Y (nx31662), .A0 (inputs_28__7), .A1 (inputs_29__7), .S0 (
             nx24333)) ;
    mux21_ni ix31675 (.Y (nx31674), .A0 (inputs_30__7), .A1 (inputs_31__7), .S0 (
             nx24333)) ;
    mux21_ni ix31979 (.Y (nx31978), .A0 (nx31972), .A1 (nx31894), .S0 (nx23151)
             ) ;
    oai21 ix31973 (.Y (nx31972), .A0 (nx22297), .A1 (nx14947), .B0 (nx14959)) ;
    mux21 ix14948 (.Y (nx14947), .A0 (nx31936), .A1 (nx31964), .S0 (nx22889)) ;
    mux21_ni ix31937 (.Y (nx31936), .A0 (nx31920), .A1 (nx31932), .S0 (nx23607)
             ) ;
    mux21_ni ix31921 (.Y (nx31920), .A0 (inputs_36__7), .A1 (inputs_37__7), .S0 (
             nx24333)) ;
    mux21_ni ix31933 (.Y (nx31932), .A0 (inputs_38__7), .A1 (inputs_39__7), .S0 (
             nx24335)) ;
    mux21_ni ix31965 (.Y (nx31964), .A0 (nx31948), .A1 (nx31960), .S0 (nx23607)
             ) ;
    mux21_ni ix31949 (.Y (nx31948), .A0 (inputs_52__7), .A1 (inputs_53__7), .S0 (
             nx24335)) ;
    mux21_ni ix31961 (.Y (nx31960), .A0 (inputs_54__7), .A1 (inputs_55__7), .S0 (
             nx24335)) ;
    nand04 ix14960 (.Y (nx14959), .A0 (nx22297), .A1 (nx23607), .A2 (nx24335), .A3 (
           nx31908)) ;
    mux21_ni ix31909 (.Y (nx31908), .A0 (inputs_35__7), .A1 (inputs_51__7), .S0 (
             nx22889)) ;
    mux21_ni ix31895 (.Y (nx31894), .A0 (nx31830), .A1 (nx31890), .S0 (nx22891)
             ) ;
    mux21_ni ix31831 (.Y (nx31830), .A0 (nx31798), .A1 (nx31826), .S0 (nx23259)
             ) ;
    mux21_ni ix31799 (.Y (nx31798), .A0 (nx31782), .A1 (nx31794), .S0 (nx23607)
             ) ;
    mux21_ni ix31783 (.Y (nx31782), .A0 (inputs_40__7), .A1 (inputs_41__7), .S0 (
             nx24335)) ;
    mux21_ni ix31795 (.Y (nx31794), .A0 (inputs_42__7), .A1 (inputs_43__7), .S0 (
             nx24335)) ;
    mux21_ni ix31827 (.Y (nx31826), .A0 (nx31810), .A1 (nx31822), .S0 (nx23607)
             ) ;
    mux21_ni ix31811 (.Y (nx31810), .A0 (inputs_44__7), .A1 (inputs_45__7), .S0 (
             nx24335)) ;
    mux21_ni ix31823 (.Y (nx31822), .A0 (inputs_46__7), .A1 (inputs_47__7), .S0 (
             nx24337)) ;
    mux21_ni ix31891 (.Y (nx31890), .A0 (nx31858), .A1 (nx31886), .S0 (nx23259)
             ) ;
    mux21_ni ix31859 (.Y (nx31858), .A0 (nx31842), .A1 (nx31854), .S0 (nx23609)
             ) ;
    mux21_ni ix31843 (.Y (nx31842), .A0 (inputs_56__7), .A1 (inputs_57__7), .S0 (
             nx24337)) ;
    mux21_ni ix31855 (.Y (nx31854), .A0 (inputs_58__7), .A1 (inputs_59__7), .S0 (
             nx24337)) ;
    mux21_ni ix31887 (.Y (nx31886), .A0 (nx31870), .A1 (nx31882), .S0 (nx23609)
             ) ;
    mux21_ni ix31871 (.Y (nx31870), .A0 (inputs_60__7), .A1 (inputs_61__7), .S0 (
             nx24337)) ;
    mux21_ni ix31883 (.Y (nx31882), .A0 (inputs_62__7), .A1 (inputs_63__7), .S0 (
             nx24337)) ;
    mux21_ni ix32403 (.Y (nx32402), .A0 (nx32190), .A1 (nx32398), .S0 (nx22599)
             ) ;
    mux21_ni ix32191 (.Y (nx32190), .A0 (nx32184), .A1 (nx32106), .S0 (nx23151)
             ) ;
    oai21 ix32185 (.Y (nx32184), .A0 (nx22299), .A1 (nx14991), .B0 (nx15001)) ;
    mux21 ix14992 (.Y (nx14991), .A0 (nx32148), .A1 (nx32176), .S0 (nx22891)) ;
    mux21_ni ix32149 (.Y (nx32148), .A0 (nx32132), .A1 (nx32144), .S0 (nx23609)
             ) ;
    mux21_ni ix32133 (.Y (nx32132), .A0 (inputs_68__7), .A1 (inputs_69__7), .S0 (
             nx24337)) ;
    mux21_ni ix32145 (.Y (nx32144), .A0 (inputs_70__7), .A1 (inputs_71__7), .S0 (
             nx24337)) ;
    mux21_ni ix32177 (.Y (nx32176), .A0 (nx32160), .A1 (nx32172), .S0 (nx23609)
             ) ;
    mux21_ni ix32161 (.Y (nx32160), .A0 (inputs_84__7), .A1 (inputs_85__7), .S0 (
             nx24339)) ;
    mux21_ni ix32173 (.Y (nx32172), .A0 (inputs_86__7), .A1 (inputs_87__7), .S0 (
             nx24339)) ;
    nand04 ix15002 (.Y (nx15001), .A0 (nx22299), .A1 (nx23609), .A2 (nx24339), .A3 (
           nx32120)) ;
    mux21_ni ix32121 (.Y (nx32120), .A0 (inputs_67__7), .A1 (inputs_83__7), .S0 (
             nx22891)) ;
    mux21_ni ix32107 (.Y (nx32106), .A0 (nx32042), .A1 (nx32102), .S0 (nx22891)
             ) ;
    mux21_ni ix32043 (.Y (nx32042), .A0 (nx32010), .A1 (nx32038), .S0 (nx23259)
             ) ;
    mux21_ni ix32011 (.Y (nx32010), .A0 (nx31994), .A1 (nx32006), .S0 (nx23609)
             ) ;
    mux21_ni ix31995 (.Y (nx31994), .A0 (inputs_72__7), .A1 (inputs_73__7), .S0 (
             nx24339)) ;
    mux21_ni ix32007 (.Y (nx32006), .A0 (inputs_74__7), .A1 (inputs_75__7), .S0 (
             nx24339)) ;
    mux21_ni ix32039 (.Y (nx32038), .A0 (nx32022), .A1 (nx32034), .S0 (nx23609)
             ) ;
    mux21_ni ix32023 (.Y (nx32022), .A0 (inputs_76__7), .A1 (inputs_77__7), .S0 (
             nx24339)) ;
    mux21_ni ix32035 (.Y (nx32034), .A0 (inputs_78__7), .A1 (inputs_79__7), .S0 (
             nx24339)) ;
    mux21_ni ix32103 (.Y (nx32102), .A0 (nx32070), .A1 (nx32098), .S0 (nx23261)
             ) ;
    mux21_ni ix32071 (.Y (nx32070), .A0 (nx32054), .A1 (nx32066), .S0 (nx23611)
             ) ;
    mux21_ni ix32055 (.Y (nx32054), .A0 (inputs_88__7), .A1 (inputs_89__7), .S0 (
             nx24341)) ;
    mux21_ni ix32067 (.Y (nx32066), .A0 (inputs_90__7), .A1 (inputs_91__7), .S0 (
             nx24341)) ;
    mux21_ni ix32099 (.Y (nx32098), .A0 (nx32082), .A1 (nx32094), .S0 (nx23611)
             ) ;
    mux21_ni ix32083 (.Y (nx32082), .A0 (inputs_92__7), .A1 (inputs_93__7), .S0 (
             nx24341)) ;
    mux21_ni ix32095 (.Y (nx32094), .A0 (inputs_94__7), .A1 (inputs_95__7), .S0 (
             nx24341)) ;
    mux21_ni ix32399 (.Y (nx32398), .A0 (nx32392), .A1 (nx32314), .S0 (nx23151)
             ) ;
    oai21 ix32393 (.Y (nx32392), .A0 (nx22299), .A1 (nx15031), .B0 (nx15041)) ;
    mux21 ix15032 (.Y (nx15031), .A0 (nx32356), .A1 (nx32384), .S0 (nx22891)) ;
    mux21_ni ix32357 (.Y (nx32356), .A0 (nx32340), .A1 (nx32352), .S0 (nx23611)
             ) ;
    mux21_ni ix32341 (.Y (nx32340), .A0 (inputs_100__7), .A1 (inputs_101__7), .S0 (
             nx24341)) ;
    mux21_ni ix32353 (.Y (nx32352), .A0 (inputs_102__7), .A1 (inputs_103__7), .S0 (
             nx24341)) ;
    mux21_ni ix32385 (.Y (nx32384), .A0 (nx32368), .A1 (nx32380), .S0 (nx23611)
             ) ;
    mux21_ni ix32369 (.Y (nx32368), .A0 (inputs_116__7), .A1 (inputs_117__7), .S0 (
             nx24341)) ;
    mux21_ni ix32381 (.Y (nx32380), .A0 (inputs_118__7), .A1 (inputs_119__7), .S0 (
             nx24343)) ;
    nand04 ix15042 (.Y (nx15041), .A0 (nx22299), .A1 (nx23611), .A2 (nx24343), .A3 (
           nx32328)) ;
    mux21_ni ix32329 (.Y (nx32328), .A0 (inputs_99__7), .A1 (inputs_115__7), .S0 (
             nx22891)) ;
    mux21_ni ix32315 (.Y (nx32314), .A0 (nx32250), .A1 (nx32310), .S0 (nx22891)
             ) ;
    mux21_ni ix32251 (.Y (nx32250), .A0 (nx32218), .A1 (nx32246), .S0 (nx23261)
             ) ;
    mux21_ni ix32219 (.Y (nx32218), .A0 (nx32202), .A1 (nx32214), .S0 (nx23611)
             ) ;
    mux21_ni ix32203 (.Y (nx32202), .A0 (inputs_104__7), .A1 (inputs_105__7), .S0 (
             nx24343)) ;
    mux21_ni ix32215 (.Y (nx32214), .A0 (inputs_106__7), .A1 (inputs_107__7), .S0 (
             nx24343)) ;
    mux21_ni ix32247 (.Y (nx32246), .A0 (nx32230), .A1 (nx32242), .S0 (nx23611)
             ) ;
    mux21_ni ix32231 (.Y (nx32230), .A0 (inputs_108__7), .A1 (inputs_109__7), .S0 (
             nx24343)) ;
    mux21_ni ix32243 (.Y (nx32242), .A0 (inputs_110__7), .A1 (inputs_111__7), .S0 (
             nx24343)) ;
    mux21_ni ix32311 (.Y (nx32310), .A0 (nx32278), .A1 (nx32306), .S0 (nx23261)
             ) ;
    mux21_ni ix32279 (.Y (nx32278), .A0 (nx32262), .A1 (nx32274), .S0 (nx23613)
             ) ;
    mux21_ni ix32263 (.Y (nx32262), .A0 (inputs_120__7), .A1 (inputs_121__7), .S0 (
             nx24343)) ;
    mux21_ni ix32275 (.Y (nx32274), .A0 (inputs_122__7), .A1 (inputs_123__7), .S0 (
             nx24345)) ;
    mux21_ni ix32307 (.Y (nx32306), .A0 (nx32290), .A1 (nx32302), .S0 (nx23613)
             ) ;
    mux21_ni ix32291 (.Y (nx32290), .A0 (inputs_124__7), .A1 (inputs_125__7), .S0 (
             nx24345)) ;
    mux21_ni ix32303 (.Y (nx32302), .A0 (inputs_126__7), .A1 (inputs_127__7), .S0 (
             nx24345)) ;
    mux21_ni ix33251 (.Y (nx33250), .A0 (nx32826), .A1 (nx33246), .S0 (nx22487)
             ) ;
    mux21_ni ix32827 (.Y (nx32826), .A0 (nx32614), .A1 (nx32822), .S0 (nx22599)
             ) ;
    mux21_ni ix32615 (.Y (nx32614), .A0 (nx32608), .A1 (nx32530), .S0 (nx23151)
             ) ;
    oai21 ix32609 (.Y (nx32608), .A0 (nx22299), .A1 (nx15077), .B0 (nx15089)) ;
    mux21 ix15078 (.Y (nx15077), .A0 (nx32572), .A1 (nx32600), .S0 (nx22893)) ;
    mux21_ni ix32573 (.Y (nx32572), .A0 (nx32556), .A1 (nx32568), .S0 (nx23613)
             ) ;
    mux21_ni ix32557 (.Y (nx32556), .A0 (inputs_132__7), .A1 (inputs_133__7), .S0 (
             nx24345)) ;
    mux21_ni ix32569 (.Y (nx32568), .A0 (inputs_134__7), .A1 (inputs_135__7), .S0 (
             nx24345)) ;
    mux21_ni ix32601 (.Y (nx32600), .A0 (nx32584), .A1 (nx32596), .S0 (nx23613)
             ) ;
    mux21_ni ix32585 (.Y (nx32584), .A0 (inputs_148__7), .A1 (inputs_149__7), .S0 (
             nx24345)) ;
    mux21_ni ix32597 (.Y (nx32596), .A0 (inputs_150__7), .A1 (inputs_151__7), .S0 (
             nx24345)) ;
    nand04 ix15090 (.Y (nx15089), .A0 (nx22299), .A1 (nx23613), .A2 (nx24347), .A3 (
           nx32544)) ;
    mux21_ni ix32545 (.Y (nx32544), .A0 (inputs_131__7), .A1 (inputs_147__7), .S0 (
             nx22893)) ;
    mux21_ni ix32531 (.Y (nx32530), .A0 (nx32466), .A1 (nx32526), .S0 (nx22893)
             ) ;
    mux21_ni ix32467 (.Y (nx32466), .A0 (nx32434), .A1 (nx32462), .S0 (nx23261)
             ) ;
    mux21_ni ix32435 (.Y (nx32434), .A0 (nx32418), .A1 (nx32430), .S0 (nx23613)
             ) ;
    mux21_ni ix32419 (.Y (nx32418), .A0 (inputs_136__7), .A1 (inputs_137__7), .S0 (
             nx24347)) ;
    mux21_ni ix32431 (.Y (nx32430), .A0 (inputs_138__7), .A1 (inputs_139__7), .S0 (
             nx24347)) ;
    mux21_ni ix32463 (.Y (nx32462), .A0 (nx32446), .A1 (nx32458), .S0 (nx23613)
             ) ;
    mux21_ni ix32447 (.Y (nx32446), .A0 (inputs_140__7), .A1 (inputs_141__7), .S0 (
             nx24347)) ;
    mux21_ni ix32459 (.Y (nx32458), .A0 (inputs_142__7), .A1 (inputs_143__7), .S0 (
             nx24347)) ;
    mux21_ni ix32527 (.Y (nx32526), .A0 (nx32494), .A1 (nx32522), .S0 (nx23261)
             ) ;
    mux21_ni ix32495 (.Y (nx32494), .A0 (nx32478), .A1 (nx32490), .S0 (nx23615)
             ) ;
    mux21_ni ix32479 (.Y (nx32478), .A0 (inputs_152__7), .A1 (inputs_153__7), .S0 (
             nx24347)) ;
    mux21_ni ix32491 (.Y (nx32490), .A0 (inputs_154__7), .A1 (inputs_155__7), .S0 (
             nx24347)) ;
    mux21_ni ix32523 (.Y (nx32522), .A0 (nx32506), .A1 (nx32518), .S0 (nx23615)
             ) ;
    mux21_ni ix32507 (.Y (nx32506), .A0 (inputs_156__7), .A1 (inputs_157__7), .S0 (
             nx24349)) ;
    mux21_ni ix32519 (.Y (nx32518), .A0 (inputs_158__7), .A1 (inputs_159__7), .S0 (
             nx24349)) ;
    mux21_ni ix32823 (.Y (nx32822), .A0 (nx32816), .A1 (nx32738), .S0 (nx23151)
             ) ;
    oai21 ix32817 (.Y (nx32816), .A0 (nx22299), .A1 (nx15119), .B0 (nx15133)) ;
    mux21 ix15120 (.Y (nx15119), .A0 (nx32780), .A1 (nx32808), .S0 (nx22893)) ;
    mux21_ni ix32781 (.Y (nx32780), .A0 (nx32764), .A1 (nx32776), .S0 (nx23615)
             ) ;
    mux21_ni ix32765 (.Y (nx32764), .A0 (inputs_164__7), .A1 (inputs_165__7), .S0 (
             nx24349)) ;
    mux21_ni ix32777 (.Y (nx32776), .A0 (inputs_166__7), .A1 (inputs_167__7), .S0 (
             nx24349)) ;
    mux21_ni ix32809 (.Y (nx32808), .A0 (nx32792), .A1 (nx32804), .S0 (nx23615)
             ) ;
    mux21_ni ix32793 (.Y (nx32792), .A0 (inputs_180__7), .A1 (inputs_181__7), .S0 (
             nx24349)) ;
    mux21_ni ix32805 (.Y (nx32804), .A0 (inputs_182__7), .A1 (inputs_183__7), .S0 (
             nx24349)) ;
    nand04 ix15134 (.Y (nx15133), .A0 (nx22301), .A1 (nx23615), .A2 (nx24349), .A3 (
           nx32752)) ;
    mux21_ni ix32753 (.Y (nx32752), .A0 (inputs_163__7), .A1 (inputs_179__7), .S0 (
             nx22893)) ;
    mux21_ni ix32739 (.Y (nx32738), .A0 (nx32674), .A1 (nx32734), .S0 (nx22893)
             ) ;
    mux21_ni ix32675 (.Y (nx32674), .A0 (nx32642), .A1 (nx32670), .S0 (nx23261)
             ) ;
    mux21_ni ix32643 (.Y (nx32642), .A0 (nx32626), .A1 (nx32638), .S0 (nx23615)
             ) ;
    mux21_ni ix32627 (.Y (nx32626), .A0 (inputs_168__7), .A1 (inputs_169__7), .S0 (
             nx24351)) ;
    mux21_ni ix32639 (.Y (nx32638), .A0 (inputs_170__7), .A1 (inputs_171__7), .S0 (
             nx24351)) ;
    mux21_ni ix32671 (.Y (nx32670), .A0 (nx32654), .A1 (nx32666), .S0 (nx23615)
             ) ;
    mux21_ni ix32655 (.Y (nx32654), .A0 (inputs_172__7), .A1 (inputs_173__7), .S0 (
             nx24351)) ;
    mux21_ni ix32667 (.Y (nx32666), .A0 (inputs_174__7), .A1 (inputs_175__7), .S0 (
             nx24351)) ;
    mux21_ni ix32735 (.Y (nx32734), .A0 (nx32702), .A1 (nx32730), .S0 (nx23261)
             ) ;
    mux21_ni ix32703 (.Y (nx32702), .A0 (nx32686), .A1 (nx32698), .S0 (nx23617)
             ) ;
    mux21_ni ix32687 (.Y (nx32686), .A0 (inputs_184__7), .A1 (inputs_185__7), .S0 (
             nx24351)) ;
    mux21_ni ix32699 (.Y (nx32698), .A0 (inputs_186__7), .A1 (inputs_187__7), .S0 (
             nx24351)) ;
    mux21_ni ix32731 (.Y (nx32730), .A0 (nx32714), .A1 (nx32726), .S0 (nx23617)
             ) ;
    mux21_ni ix32715 (.Y (nx32714), .A0 (inputs_188__7), .A1 (inputs_189__7), .S0 (
             nx24351)) ;
    mux21_ni ix32727 (.Y (nx32726), .A0 (inputs_190__7), .A1 (inputs_191__7), .S0 (
             nx24353)) ;
    mux21_ni ix33247 (.Y (nx33246), .A0 (nx33034), .A1 (nx33242), .S0 (nx22599)
             ) ;
    mux21_ni ix33035 (.Y (nx33034), .A0 (nx33028), .A1 (nx32950), .S0 (nx23153)
             ) ;
    oai21 ix33029 (.Y (nx33028), .A0 (nx22301), .A1 (nx15163), .B0 (nx15175)) ;
    mux21 ix15164 (.Y (nx15163), .A0 (nx32992), .A1 (nx33020), .S0 (nx22893)) ;
    mux21_ni ix32993 (.Y (nx32992), .A0 (nx32976), .A1 (nx32988), .S0 (nx23617)
             ) ;
    mux21_ni ix32977 (.Y (nx32976), .A0 (inputs_196__7), .A1 (inputs_197__7), .S0 (
             nx24353)) ;
    mux21_ni ix32989 (.Y (nx32988), .A0 (inputs_198__7), .A1 (inputs_199__7), .S0 (
             nx24353)) ;
    mux21_ni ix33021 (.Y (nx33020), .A0 (nx33004), .A1 (nx33016), .S0 (nx23617)
             ) ;
    mux21_ni ix33005 (.Y (nx33004), .A0 (inputs_212__7), .A1 (inputs_213__7), .S0 (
             nx24353)) ;
    mux21_ni ix33017 (.Y (nx33016), .A0 (inputs_214__7), .A1 (inputs_215__7), .S0 (
             nx24353)) ;
    nand04 ix15176 (.Y (nx15175), .A0 (nx22301), .A1 (nx23617), .A2 (nx24353), .A3 (
           nx32964)) ;
    mux21_ni ix32965 (.Y (nx32964), .A0 (inputs_195__7), .A1 (inputs_211__7), .S0 (
             nx22895)) ;
    mux21_ni ix32951 (.Y (nx32950), .A0 (nx32886), .A1 (nx32946), .S0 (nx22895)
             ) ;
    mux21_ni ix32887 (.Y (nx32886), .A0 (nx32854), .A1 (nx32882), .S0 (nx23263)
             ) ;
    mux21_ni ix32855 (.Y (nx32854), .A0 (nx32838), .A1 (nx32850), .S0 (nx23617)
             ) ;
    mux21_ni ix32839 (.Y (nx32838), .A0 (inputs_200__7), .A1 (inputs_201__7), .S0 (
             nx24353)) ;
    mux21_ni ix32851 (.Y (nx32850), .A0 (inputs_202__7), .A1 (inputs_203__7), .S0 (
             nx24355)) ;
    mux21_ni ix32883 (.Y (nx32882), .A0 (nx32866), .A1 (nx32878), .S0 (nx23617)
             ) ;
    mux21_ni ix32867 (.Y (nx32866), .A0 (inputs_204__7), .A1 (inputs_205__7), .S0 (
             nx24355)) ;
    mux21_ni ix32879 (.Y (nx32878), .A0 (inputs_206__7), .A1 (inputs_207__7), .S0 (
             nx24355)) ;
    mux21_ni ix32947 (.Y (nx32946), .A0 (nx32914), .A1 (nx32942), .S0 (nx23263)
             ) ;
    mux21_ni ix32915 (.Y (nx32914), .A0 (nx32898), .A1 (nx32910), .S0 (nx23619)
             ) ;
    mux21_ni ix32899 (.Y (nx32898), .A0 (inputs_216__7), .A1 (inputs_217__7), .S0 (
             nx24355)) ;
    mux21_ni ix32911 (.Y (nx32910), .A0 (inputs_218__7), .A1 (inputs_219__7), .S0 (
             nx24355)) ;
    mux21_ni ix32943 (.Y (nx32942), .A0 (nx32926), .A1 (nx32938), .S0 (nx23619)
             ) ;
    mux21_ni ix32927 (.Y (nx32926), .A0 (inputs_220__7), .A1 (inputs_221__7), .S0 (
             nx24355)) ;
    mux21_ni ix32939 (.Y (nx32938), .A0 (inputs_222__7), .A1 (inputs_223__7), .S0 (
             nx24355)) ;
    mux21_ni ix33243 (.Y (nx33242), .A0 (nx33236), .A1 (nx33158), .S0 (nx23153)
             ) ;
    oai21 ix33237 (.Y (nx33236), .A0 (nx22301), .A1 (nx15207), .B0 (nx15219)) ;
    mux21 ix15208 (.Y (nx15207), .A0 (nx33200), .A1 (nx33228), .S0 (nx22895)) ;
    mux21_ni ix33201 (.Y (nx33200), .A0 (nx33184), .A1 (nx33196), .S0 (nx23619)
             ) ;
    mux21_ni ix33185 (.Y (nx33184), .A0 (inputs_228__7), .A1 (inputs_229__7), .S0 (
             nx24357)) ;
    mux21_ni ix33197 (.Y (nx33196), .A0 (inputs_230__7), .A1 (inputs_231__7), .S0 (
             nx24357)) ;
    mux21_ni ix33229 (.Y (nx33228), .A0 (nx33212), .A1 (nx33224), .S0 (nx23619)
             ) ;
    mux21_ni ix33213 (.Y (nx33212), .A0 (inputs_244__7), .A1 (inputs_245__7), .S0 (
             nx24357)) ;
    mux21_ni ix33225 (.Y (nx33224), .A0 (inputs_246__7), .A1 (inputs_247__7), .S0 (
             nx24357)) ;
    nand04 ix15220 (.Y (nx15219), .A0 (nx22301), .A1 (nx23619), .A2 (nx24357), .A3 (
           nx33172)) ;
    mux21_ni ix33173 (.Y (nx33172), .A0 (inputs_227__7), .A1 (inputs_243__7), .S0 (
             nx22895)) ;
    mux21_ni ix33159 (.Y (nx33158), .A0 (nx33094), .A1 (nx33154), .S0 (nx22895)
             ) ;
    mux21_ni ix33095 (.Y (nx33094), .A0 (nx33062), .A1 (nx33090), .S0 (nx23263)
             ) ;
    mux21_ni ix33063 (.Y (nx33062), .A0 (nx33046), .A1 (nx33058), .S0 (nx23619)
             ) ;
    mux21_ni ix33047 (.Y (nx33046), .A0 (inputs_232__7), .A1 (inputs_233__7), .S0 (
             nx24357)) ;
    mux21_ni ix33059 (.Y (nx33058), .A0 (inputs_234__7), .A1 (inputs_235__7), .S0 (
             nx24357)) ;
    mux21_ni ix33091 (.Y (nx33090), .A0 (nx33074), .A1 (nx33086), .S0 (nx23619)
             ) ;
    mux21_ni ix33075 (.Y (nx33074), .A0 (inputs_236__7), .A1 (inputs_237__7), .S0 (
             nx24359)) ;
    mux21_ni ix33087 (.Y (nx33086), .A0 (inputs_238__7), .A1 (inputs_239__7), .S0 (
             nx24359)) ;
    mux21_ni ix33155 (.Y (nx33154), .A0 (nx33122), .A1 (nx33150), .S0 (nx23263)
             ) ;
    mux21_ni ix33123 (.Y (nx33122), .A0 (nx33106), .A1 (nx33118), .S0 (nx23621)
             ) ;
    mux21_ni ix33107 (.Y (nx33106), .A0 (inputs_248__7), .A1 (inputs_249__7), .S0 (
             nx24359)) ;
    mux21_ni ix33119 (.Y (nx33118), .A0 (inputs_250__7), .A1 (inputs_251__7), .S0 (
             nx24359)) ;
    mux21_ni ix33151 (.Y (nx33150), .A0 (nx33134), .A1 (nx33146), .S0 (nx23621)
             ) ;
    mux21_ni ix33135 (.Y (nx33134), .A0 (inputs_252__7), .A1 (inputs_253__7), .S0 (
             nx24359)) ;
    mux21_ni ix33147 (.Y (nx33146), .A0 (inputs_254__7), .A1 (inputs_255__7), .S0 (
             nx24359)) ;
    oai21 ix37421 (.Y (\output [8]), .A0 (nx22221), .A1 (nx15247), .B0 (nx15607)
          ) ;
    mux21 ix15248 (.Y (nx15247), .A0 (nx34102), .A1 (nx34946), .S0 (nx22429)) ;
    mux21_ni ix34103 (.Y (nx34102), .A0 (nx33678), .A1 (nx34098), .S0 (nx22487)
             ) ;
    mux21_ni ix33679 (.Y (nx33678), .A0 (nx33466), .A1 (nx33674), .S0 (nx22599)
             ) ;
    mux21_ni ix33467 (.Y (nx33466), .A0 (nx33460), .A1 (nx33382), .S0 (nx23153)
             ) ;
    oai21 ix33461 (.Y (nx33460), .A0 (nx22301), .A1 (nx15257), .B0 (nx15269)) ;
    mux21 ix15258 (.Y (nx15257), .A0 (nx33424), .A1 (nx33452), .S0 (nx22895)) ;
    mux21_ni ix33425 (.Y (nx33424), .A0 (nx33408), .A1 (nx33420), .S0 (nx23621)
             ) ;
    mux21_ni ix33409 (.Y (nx33408), .A0 (inputs_260__8), .A1 (inputs_261__8), .S0 (
             nx24359)) ;
    mux21_ni ix33421 (.Y (nx33420), .A0 (inputs_262__8), .A1 (inputs_263__8), .S0 (
             nx24361)) ;
    mux21_ni ix33453 (.Y (nx33452), .A0 (nx33436), .A1 (nx33448), .S0 (nx23621)
             ) ;
    mux21_ni ix33437 (.Y (nx33436), .A0 (inputs_276__8), .A1 (inputs_277__8), .S0 (
             nx24361)) ;
    mux21_ni ix33449 (.Y (nx33448), .A0 (inputs_278__8), .A1 (inputs_279__8), .S0 (
             nx24361)) ;
    nand04 ix15270 (.Y (nx15269), .A0 (nx22301), .A1 (nx23621), .A2 (nx24361), .A3 (
           nx33396)) ;
    mux21_ni ix33397 (.Y (nx33396), .A0 (inputs_259__8), .A1 (inputs_275__8), .S0 (
             nx22895)) ;
    mux21_ni ix33383 (.Y (nx33382), .A0 (nx33318), .A1 (nx33378), .S0 (nx22897)
             ) ;
    mux21_ni ix33319 (.Y (nx33318), .A0 (nx33286), .A1 (nx33314), .S0 (nx23263)
             ) ;
    mux21_ni ix33287 (.Y (nx33286), .A0 (nx33270), .A1 (nx33282), .S0 (nx23621)
             ) ;
    mux21_ni ix33271 (.Y (nx33270), .A0 (inputs_264__8), .A1 (inputs_265__8), .S0 (
             nx24361)) ;
    mux21_ni ix33283 (.Y (nx33282), .A0 (inputs_266__8), .A1 (inputs_267__8), .S0 (
             nx24361)) ;
    mux21_ni ix33315 (.Y (nx33314), .A0 (nx33298), .A1 (nx33310), .S0 (nx23621)
             ) ;
    mux21_ni ix33299 (.Y (nx33298), .A0 (inputs_268__8), .A1 (inputs_269__8), .S0 (
             nx24361)) ;
    mux21_ni ix33311 (.Y (nx33310), .A0 (inputs_270__8), .A1 (inputs_271__8), .S0 (
             nx24363)) ;
    mux21_ni ix33379 (.Y (nx33378), .A0 (nx33346), .A1 (nx33374), .S0 (nx23263)
             ) ;
    mux21_ni ix33347 (.Y (nx33346), .A0 (nx33330), .A1 (nx33342), .S0 (nx23623)
             ) ;
    mux21_ni ix33331 (.Y (nx33330), .A0 (inputs_280__8), .A1 (inputs_281__8), .S0 (
             nx24363)) ;
    mux21_ni ix33343 (.Y (nx33342), .A0 (inputs_282__8), .A1 (inputs_283__8), .S0 (
             nx24363)) ;
    mux21_ni ix33375 (.Y (nx33374), .A0 (nx33358), .A1 (nx33370), .S0 (nx23623)
             ) ;
    mux21_ni ix33359 (.Y (nx33358), .A0 (inputs_284__8), .A1 (inputs_285__8), .S0 (
             nx24363)) ;
    mux21_ni ix33371 (.Y (nx33370), .A0 (inputs_286__8), .A1 (inputs_287__8), .S0 (
             nx24363)) ;
    mux21_ni ix33675 (.Y (nx33674), .A0 (nx33668), .A1 (nx33590), .S0 (nx23153)
             ) ;
    oai21 ix33669 (.Y (nx33668), .A0 (nx22303), .A1 (nx15299), .B0 (nx15311)) ;
    mux21 ix15300 (.Y (nx15299), .A0 (nx33632), .A1 (nx33660), .S0 (nx22897)) ;
    mux21_ni ix33633 (.Y (nx33632), .A0 (nx33616), .A1 (nx33628), .S0 (nx23623)
             ) ;
    mux21_ni ix33617 (.Y (nx33616), .A0 (inputs_292__8), .A1 (inputs_293__8), .S0 (
             nx24363)) ;
    mux21_ni ix33629 (.Y (nx33628), .A0 (inputs_294__8), .A1 (inputs_295__8), .S0 (
             nx24363)) ;
    mux21_ni ix33661 (.Y (nx33660), .A0 (nx33644), .A1 (nx33656), .S0 (nx23623)
             ) ;
    mux21_ni ix33645 (.Y (nx33644), .A0 (inputs_308__8), .A1 (inputs_309__8), .S0 (
             nx24365)) ;
    mux21_ni ix33657 (.Y (nx33656), .A0 (inputs_310__8), .A1 (inputs_311__8), .S0 (
             nx24365)) ;
    nand04 ix15312 (.Y (nx15311), .A0 (nx22303), .A1 (nx23623), .A2 (nx24365), .A3 (
           nx33604)) ;
    mux21_ni ix33605 (.Y (nx33604), .A0 (inputs_291__8), .A1 (inputs_307__8), .S0 (
             nx22897)) ;
    mux21_ni ix33591 (.Y (nx33590), .A0 (nx33526), .A1 (nx33586), .S0 (nx22897)
             ) ;
    mux21_ni ix33527 (.Y (nx33526), .A0 (nx33494), .A1 (nx33522), .S0 (nx23263)
             ) ;
    mux21_ni ix33495 (.Y (nx33494), .A0 (nx33478), .A1 (nx33490), .S0 (nx23623)
             ) ;
    mux21_ni ix33479 (.Y (nx33478), .A0 (inputs_296__8), .A1 (inputs_297__8), .S0 (
             nx24365)) ;
    mux21_ni ix33491 (.Y (nx33490), .A0 (inputs_298__8), .A1 (inputs_299__8), .S0 (
             nx24365)) ;
    mux21_ni ix33523 (.Y (nx33522), .A0 (nx33506), .A1 (nx33518), .S0 (nx23623)
             ) ;
    mux21_ni ix33507 (.Y (nx33506), .A0 (inputs_300__8), .A1 (inputs_301__8), .S0 (
             nx24365)) ;
    mux21_ni ix33519 (.Y (nx33518), .A0 (inputs_302__8), .A1 (inputs_303__8), .S0 (
             nx24365)) ;
    mux21_ni ix33587 (.Y (nx33586), .A0 (nx33554), .A1 (nx33582), .S0 (nx23265)
             ) ;
    mux21_ni ix33555 (.Y (nx33554), .A0 (nx33538), .A1 (nx33550), .S0 (nx23625)
             ) ;
    mux21_ni ix33539 (.Y (nx33538), .A0 (inputs_312__8), .A1 (inputs_313__8), .S0 (
             nx24367)) ;
    mux21_ni ix33551 (.Y (nx33550), .A0 (inputs_314__8), .A1 (inputs_315__8), .S0 (
             nx24367)) ;
    mux21_ni ix33583 (.Y (nx33582), .A0 (nx33566), .A1 (nx33578), .S0 (nx23625)
             ) ;
    mux21_ni ix33567 (.Y (nx33566), .A0 (inputs_316__8), .A1 (inputs_317__8), .S0 (
             nx24367)) ;
    mux21_ni ix33579 (.Y (nx33578), .A0 (inputs_318__8), .A1 (inputs_319__8), .S0 (
             nx24367)) ;
    mux21_ni ix34099 (.Y (nx34098), .A0 (nx33886), .A1 (nx34094), .S0 (nx22599)
             ) ;
    mux21_ni ix33887 (.Y (nx33886), .A0 (nx33880), .A1 (nx33802), .S0 (nx23153)
             ) ;
    oai21 ix33881 (.Y (nx33880), .A0 (nx22303), .A1 (nx15345), .B0 (nx15357)) ;
    mux21 ix15346 (.Y (nx15345), .A0 (nx33844), .A1 (nx33872), .S0 (nx22897)) ;
    mux21_ni ix33845 (.Y (nx33844), .A0 (nx33828), .A1 (nx33840), .S0 (nx23625)
             ) ;
    mux21_ni ix33829 (.Y (nx33828), .A0 (inputs_324__8), .A1 (inputs_325__8), .S0 (
             nx24367)) ;
    mux21_ni ix33841 (.Y (nx33840), .A0 (inputs_326__8), .A1 (inputs_327__8), .S0 (
             nx24367)) ;
    mux21_ni ix33873 (.Y (nx33872), .A0 (nx33856), .A1 (nx33868), .S0 (nx23625)
             ) ;
    mux21_ni ix33857 (.Y (nx33856), .A0 (inputs_340__8), .A1 (inputs_341__8), .S0 (
             nx24367)) ;
    mux21_ni ix33869 (.Y (nx33868), .A0 (inputs_342__8), .A1 (inputs_343__8), .S0 (
             nx24369)) ;
    nand04 ix15358 (.Y (nx15357), .A0 (nx22303), .A1 (nx23625), .A2 (nx24369), .A3 (
           nx33816)) ;
    mux21_ni ix33817 (.Y (nx33816), .A0 (inputs_323__8), .A1 (inputs_339__8), .S0 (
             nx22897)) ;
    mux21_ni ix33803 (.Y (nx33802), .A0 (nx33738), .A1 (nx33798), .S0 (nx22897)
             ) ;
    mux21_ni ix33739 (.Y (nx33738), .A0 (nx33706), .A1 (nx33734), .S0 (nx23265)
             ) ;
    mux21_ni ix33707 (.Y (nx33706), .A0 (nx33690), .A1 (nx33702), .S0 (nx23625)
             ) ;
    mux21_ni ix33691 (.Y (nx33690), .A0 (inputs_328__8), .A1 (inputs_329__8), .S0 (
             nx24369)) ;
    mux21_ni ix33703 (.Y (nx33702), .A0 (inputs_330__8), .A1 (inputs_331__8), .S0 (
             nx24369)) ;
    mux21_ni ix33735 (.Y (nx33734), .A0 (nx33718), .A1 (nx33730), .S0 (nx23625)
             ) ;
    mux21_ni ix33719 (.Y (nx33718), .A0 (inputs_332__8), .A1 (inputs_333__8), .S0 (
             nx24369)) ;
    mux21_ni ix33731 (.Y (nx33730), .A0 (inputs_334__8), .A1 (inputs_335__8), .S0 (
             nx24369)) ;
    mux21_ni ix33799 (.Y (nx33798), .A0 (nx33766), .A1 (nx33794), .S0 (nx23265)
             ) ;
    mux21_ni ix33767 (.Y (nx33766), .A0 (nx33750), .A1 (nx33762), .S0 (nx23627)
             ) ;
    mux21_ni ix33751 (.Y (nx33750), .A0 (inputs_344__8), .A1 (inputs_345__8), .S0 (
             nx24369)) ;
    mux21_ni ix33763 (.Y (nx33762), .A0 (inputs_346__8), .A1 (inputs_347__8), .S0 (
             nx24371)) ;
    mux21_ni ix33795 (.Y (nx33794), .A0 (nx33778), .A1 (nx33790), .S0 (nx23627)
             ) ;
    mux21_ni ix33779 (.Y (nx33778), .A0 (inputs_348__8), .A1 (inputs_349__8), .S0 (
             nx24371)) ;
    mux21_ni ix33791 (.Y (nx33790), .A0 (inputs_350__8), .A1 (inputs_351__8), .S0 (
             nx24371)) ;
    mux21_ni ix34095 (.Y (nx34094), .A0 (nx34088), .A1 (nx34010), .S0 (nx23153)
             ) ;
    oai21 ix34089 (.Y (nx34088), .A0 (nx22303), .A1 (nx15387), .B0 (nx15399)) ;
    mux21 ix15388 (.Y (nx15387), .A0 (nx34052), .A1 (nx34080), .S0 (nx22899)) ;
    mux21_ni ix34053 (.Y (nx34052), .A0 (nx34036), .A1 (nx34048), .S0 (nx23627)
             ) ;
    mux21_ni ix34037 (.Y (nx34036), .A0 (inputs_356__8), .A1 (inputs_357__8), .S0 (
             nx24371)) ;
    mux21_ni ix34049 (.Y (nx34048), .A0 (inputs_358__8), .A1 (inputs_359__8), .S0 (
             nx24371)) ;
    mux21_ni ix34081 (.Y (nx34080), .A0 (nx34064), .A1 (nx34076), .S0 (nx23627)
             ) ;
    mux21_ni ix34065 (.Y (nx34064), .A0 (inputs_372__8), .A1 (inputs_373__8), .S0 (
             nx24371)) ;
    mux21_ni ix34077 (.Y (nx34076), .A0 (inputs_374__8), .A1 (inputs_375__8), .S0 (
             nx24371)) ;
    nand04 ix15400 (.Y (nx15399), .A0 (nx22303), .A1 (nx23627), .A2 (nx24373), .A3 (
           nx34024)) ;
    mux21_ni ix34025 (.Y (nx34024), .A0 (inputs_355__8), .A1 (inputs_371__8), .S0 (
             nx22899)) ;
    mux21_ni ix34011 (.Y (nx34010), .A0 (nx33946), .A1 (nx34006), .S0 (nx22899)
             ) ;
    mux21_ni ix33947 (.Y (nx33946), .A0 (nx33914), .A1 (nx33942), .S0 (nx23265)
             ) ;
    mux21_ni ix33915 (.Y (nx33914), .A0 (nx33898), .A1 (nx33910), .S0 (nx23627)
             ) ;
    mux21_ni ix33899 (.Y (nx33898), .A0 (inputs_360__8), .A1 (inputs_361__8), .S0 (
             nx24373)) ;
    mux21_ni ix33911 (.Y (nx33910), .A0 (inputs_362__8), .A1 (inputs_363__8), .S0 (
             nx24373)) ;
    mux21_ni ix33943 (.Y (nx33942), .A0 (nx33926), .A1 (nx33938), .S0 (nx23627)
             ) ;
    mux21_ni ix33927 (.Y (nx33926), .A0 (inputs_364__8), .A1 (inputs_365__8), .S0 (
             nx24373)) ;
    mux21_ni ix33939 (.Y (nx33938), .A0 (inputs_366__8), .A1 (inputs_367__8), .S0 (
             nx24373)) ;
    mux21_ni ix34007 (.Y (nx34006), .A0 (nx33974), .A1 (nx34002), .S0 (nx23265)
             ) ;
    mux21_ni ix33975 (.Y (nx33974), .A0 (nx33958), .A1 (nx33970), .S0 (nx23629)
             ) ;
    mux21_ni ix33959 (.Y (nx33958), .A0 (inputs_376__8), .A1 (inputs_377__8), .S0 (
             nx24373)) ;
    mux21_ni ix33971 (.Y (nx33970), .A0 (inputs_378__8), .A1 (inputs_379__8), .S0 (
             nx24373)) ;
    mux21_ni ix34003 (.Y (nx34002), .A0 (nx33986), .A1 (nx33998), .S0 (nx23629)
             ) ;
    mux21_ni ix33987 (.Y (nx33986), .A0 (inputs_380__8), .A1 (inputs_381__8), .S0 (
             nx24375)) ;
    mux21_ni ix33999 (.Y (nx33998), .A0 (inputs_382__8), .A1 (inputs_383__8), .S0 (
             nx24375)) ;
    mux21_ni ix34947 (.Y (nx34946), .A0 (nx34522), .A1 (nx34942), .S0 (nx22487)
             ) ;
    mux21_ni ix34523 (.Y (nx34522), .A0 (nx34310), .A1 (nx34518), .S0 (nx22599)
             ) ;
    mux21_ni ix34311 (.Y (nx34310), .A0 (nx34304), .A1 (nx34226), .S0 (nx23153)
             ) ;
    oai21 ix34305 (.Y (nx34304), .A0 (nx22303), .A1 (nx15433), .B0 (nx15445)) ;
    mux21 ix15434 (.Y (nx15433), .A0 (nx34268), .A1 (nx34296), .S0 (nx22899)) ;
    mux21_ni ix34269 (.Y (nx34268), .A0 (nx34252), .A1 (nx34264), .S0 (nx23629)
             ) ;
    mux21_ni ix34253 (.Y (nx34252), .A0 (inputs_388__8), .A1 (inputs_389__8), .S0 (
             nx24375)) ;
    mux21_ni ix34265 (.Y (nx34264), .A0 (inputs_390__8), .A1 (inputs_391__8), .S0 (
             nx24375)) ;
    mux21_ni ix34297 (.Y (nx34296), .A0 (nx34280), .A1 (nx34292), .S0 (nx23629)
             ) ;
    mux21_ni ix34281 (.Y (nx34280), .A0 (inputs_404__8), .A1 (inputs_405__8), .S0 (
             nx24375)) ;
    mux21_ni ix34293 (.Y (nx34292), .A0 (inputs_406__8), .A1 (inputs_407__8), .S0 (
             nx24375)) ;
    nand04 ix15446 (.Y (nx15445), .A0 (nx22305), .A1 (nx23629), .A2 (nx24375), .A3 (
           nx34240)) ;
    mux21_ni ix34241 (.Y (nx34240), .A0 (inputs_387__8), .A1 (inputs_403__8), .S0 (
             nx22899)) ;
    mux21_ni ix34227 (.Y (nx34226), .A0 (nx34162), .A1 (nx34222), .S0 (nx22899)
             ) ;
    mux21_ni ix34163 (.Y (nx34162), .A0 (nx34130), .A1 (nx34158), .S0 (nx23265)
             ) ;
    mux21_ni ix34131 (.Y (nx34130), .A0 (nx34114), .A1 (nx34126), .S0 (nx23629)
             ) ;
    mux21_ni ix34115 (.Y (nx34114), .A0 (inputs_392__8), .A1 (inputs_393__8), .S0 (
             nx24377)) ;
    mux21_ni ix34127 (.Y (nx34126), .A0 (inputs_394__8), .A1 (inputs_395__8), .S0 (
             nx24377)) ;
    mux21_ni ix34159 (.Y (nx34158), .A0 (nx34142), .A1 (nx34154), .S0 (nx23629)
             ) ;
    mux21_ni ix34143 (.Y (nx34142), .A0 (inputs_396__8), .A1 (inputs_397__8), .S0 (
             nx24377)) ;
    mux21_ni ix34155 (.Y (nx34154), .A0 (inputs_398__8), .A1 (inputs_399__8), .S0 (
             nx24377)) ;
    mux21_ni ix34223 (.Y (nx34222), .A0 (nx34190), .A1 (nx34218), .S0 (nx23265)
             ) ;
    mux21_ni ix34191 (.Y (nx34190), .A0 (nx34174), .A1 (nx34186), .S0 (nx23631)
             ) ;
    mux21_ni ix34175 (.Y (nx34174), .A0 (inputs_408__8), .A1 (inputs_409__8), .S0 (
             nx24377)) ;
    mux21_ni ix34187 (.Y (nx34186), .A0 (inputs_410__8), .A1 (inputs_411__8), .S0 (
             nx24377)) ;
    mux21_ni ix34219 (.Y (nx34218), .A0 (nx34202), .A1 (nx34214), .S0 (nx23631)
             ) ;
    mux21_ni ix34203 (.Y (nx34202), .A0 (inputs_412__8), .A1 (inputs_413__8), .S0 (
             nx24377)) ;
    mux21_ni ix34215 (.Y (nx34214), .A0 (inputs_414__8), .A1 (inputs_415__8), .S0 (
             nx24379)) ;
    mux21_ni ix34519 (.Y (nx34518), .A0 (nx34512), .A1 (nx34434), .S0 (nx23155)
             ) ;
    oai21 ix34513 (.Y (nx34512), .A0 (nx22305), .A1 (nx15479), .B0 (nx15491)) ;
    mux21 ix15480 (.Y (nx15479), .A0 (nx34476), .A1 (nx34504), .S0 (nx22899)) ;
    mux21_ni ix34477 (.Y (nx34476), .A0 (nx34460), .A1 (nx34472), .S0 (nx23631)
             ) ;
    mux21_ni ix34461 (.Y (nx34460), .A0 (inputs_420__8), .A1 (inputs_421__8), .S0 (
             nx24379)) ;
    mux21_ni ix34473 (.Y (nx34472), .A0 (inputs_422__8), .A1 (inputs_423__8), .S0 (
             nx24379)) ;
    mux21_ni ix34505 (.Y (nx34504), .A0 (nx34488), .A1 (nx34500), .S0 (nx23631)
             ) ;
    mux21_ni ix34489 (.Y (nx34488), .A0 (inputs_436__8), .A1 (inputs_437__8), .S0 (
             nx24379)) ;
    mux21_ni ix34501 (.Y (nx34500), .A0 (inputs_438__8), .A1 (inputs_439__8), .S0 (
             nx24379)) ;
    nand04 ix15492 (.Y (nx15491), .A0 (nx22305), .A1 (nx23631), .A2 (nx24379), .A3 (
           nx34448)) ;
    mux21_ni ix34449 (.Y (nx34448), .A0 (inputs_419__8), .A1 (inputs_435__8), .S0 (
             nx22901)) ;
    mux21_ni ix34435 (.Y (nx34434), .A0 (nx34370), .A1 (nx34430), .S0 (nx22901)
             ) ;
    mux21_ni ix34371 (.Y (nx34370), .A0 (nx34338), .A1 (nx34366), .S0 (nx23267)
             ) ;
    mux21_ni ix34339 (.Y (nx34338), .A0 (nx34322), .A1 (nx34334), .S0 (nx23631)
             ) ;
    mux21_ni ix34323 (.Y (nx34322), .A0 (inputs_424__8), .A1 (inputs_425__8), .S0 (
             nx24379)) ;
    mux21_ni ix34335 (.Y (nx34334), .A0 (inputs_426__8), .A1 (inputs_427__8), .S0 (
             nx24381)) ;
    mux21_ni ix34367 (.Y (nx34366), .A0 (nx34350), .A1 (nx34362), .S0 (nx23631)
             ) ;
    mux21_ni ix34351 (.Y (nx34350), .A0 (inputs_428__8), .A1 (inputs_429__8), .S0 (
             nx24381)) ;
    mux21_ni ix34363 (.Y (nx34362), .A0 (inputs_430__8), .A1 (inputs_431__8), .S0 (
             nx24381)) ;
    mux21_ni ix34431 (.Y (nx34430), .A0 (nx34398), .A1 (nx34426), .S0 (nx23267)
             ) ;
    mux21_ni ix34399 (.Y (nx34398), .A0 (nx34382), .A1 (nx34394), .S0 (nx23633)
             ) ;
    mux21_ni ix34383 (.Y (nx34382), .A0 (inputs_440__8), .A1 (inputs_441__8), .S0 (
             nx24381)) ;
    mux21_ni ix34395 (.Y (nx34394), .A0 (inputs_442__8), .A1 (inputs_443__8), .S0 (
             nx24381)) ;
    mux21_ni ix34427 (.Y (nx34426), .A0 (nx34410), .A1 (nx34422), .S0 (nx23633)
             ) ;
    mux21_ni ix34411 (.Y (nx34410), .A0 (inputs_444__8), .A1 (inputs_445__8), .S0 (
             nx24381)) ;
    mux21_ni ix34423 (.Y (nx34422), .A0 (inputs_446__8), .A1 (inputs_447__8), .S0 (
             nx24381)) ;
    mux21_ni ix34943 (.Y (nx34942), .A0 (nx34730), .A1 (nx34938), .S0 (nx22601)
             ) ;
    mux21_ni ix34731 (.Y (nx34730), .A0 (nx34724), .A1 (nx34646), .S0 (nx23155)
             ) ;
    oai21 ix34725 (.Y (nx34724), .A0 (nx22305), .A1 (nx15523), .B0 (nx15535)) ;
    mux21 ix15524 (.Y (nx15523), .A0 (nx34688), .A1 (nx34716), .S0 (nx22901)) ;
    mux21_ni ix34689 (.Y (nx34688), .A0 (nx34672), .A1 (nx34684), .S0 (nx23633)
             ) ;
    mux21_ni ix34673 (.Y (nx34672), .A0 (inputs_452__8), .A1 (inputs_453__8), .S0 (
             nx24383)) ;
    mux21_ni ix34685 (.Y (nx34684), .A0 (inputs_454__8), .A1 (inputs_455__8), .S0 (
             nx24383)) ;
    mux21_ni ix34717 (.Y (nx34716), .A0 (nx34700), .A1 (nx34712), .S0 (nx23633)
             ) ;
    mux21_ni ix34701 (.Y (nx34700), .A0 (inputs_468__8), .A1 (inputs_469__8), .S0 (
             nx24383)) ;
    mux21_ni ix34713 (.Y (nx34712), .A0 (inputs_470__8), .A1 (inputs_471__8), .S0 (
             nx24383)) ;
    nand04 ix15536 (.Y (nx15535), .A0 (nx22305), .A1 (nx23633), .A2 (nx24383), .A3 (
           nx34660)) ;
    mux21_ni ix34661 (.Y (nx34660), .A0 (inputs_451__8), .A1 (inputs_467__8), .S0 (
             nx22901)) ;
    mux21_ni ix34647 (.Y (nx34646), .A0 (nx34582), .A1 (nx34642), .S0 (nx22901)
             ) ;
    mux21_ni ix34583 (.Y (nx34582), .A0 (nx34550), .A1 (nx34578), .S0 (nx23267)
             ) ;
    mux21_ni ix34551 (.Y (nx34550), .A0 (nx34534), .A1 (nx34546), .S0 (nx23633)
             ) ;
    mux21_ni ix34535 (.Y (nx34534), .A0 (inputs_456__8), .A1 (inputs_457__8), .S0 (
             nx24383)) ;
    mux21_ni ix34547 (.Y (nx34546), .A0 (inputs_458__8), .A1 (inputs_459__8), .S0 (
             nx24383)) ;
    mux21_ni ix34579 (.Y (nx34578), .A0 (nx34562), .A1 (nx34574), .S0 (nx23633)
             ) ;
    mux21_ni ix34563 (.Y (nx34562), .A0 (inputs_460__8), .A1 (inputs_461__8), .S0 (
             nx24385)) ;
    mux21_ni ix34575 (.Y (nx34574), .A0 (inputs_462__8), .A1 (inputs_463__8), .S0 (
             nx24385)) ;
    mux21_ni ix34643 (.Y (nx34642), .A0 (nx34610), .A1 (nx34638), .S0 (nx23267)
             ) ;
    mux21_ni ix34611 (.Y (nx34610), .A0 (nx34594), .A1 (nx34606), .S0 (nx23635)
             ) ;
    mux21_ni ix34595 (.Y (nx34594), .A0 (inputs_472__8), .A1 (inputs_473__8), .S0 (
             nx24385)) ;
    mux21_ni ix34607 (.Y (nx34606), .A0 (inputs_474__8), .A1 (inputs_475__8), .S0 (
             nx24385)) ;
    mux21_ni ix34639 (.Y (nx34638), .A0 (nx34622), .A1 (nx34634), .S0 (nx23635)
             ) ;
    mux21_ni ix34623 (.Y (nx34622), .A0 (inputs_476__8), .A1 (inputs_477__8), .S0 (
             nx24385)) ;
    mux21_ni ix34635 (.Y (nx34634), .A0 (inputs_478__8), .A1 (inputs_479__8), .S0 (
             nx24385)) ;
    mux21_ni ix34939 (.Y (nx34938), .A0 (nx34932), .A1 (nx34854), .S0 (nx23155)
             ) ;
    oai21 ix34933 (.Y (nx34932), .A0 (nx22305), .A1 (nx15567), .B0 (nx15579)) ;
    mux21 ix15568 (.Y (nx15567), .A0 (nx34896), .A1 (nx34924), .S0 (nx22901)) ;
    mux21_ni ix34897 (.Y (nx34896), .A0 (nx34880), .A1 (nx34892), .S0 (nx23635)
             ) ;
    mux21_ni ix34881 (.Y (nx34880), .A0 (inputs_484__8), .A1 (inputs_485__8), .S0 (
             nx24385)) ;
    mux21_ni ix34893 (.Y (nx34892), .A0 (inputs_486__8), .A1 (inputs_487__8), .S0 (
             nx24387)) ;
    mux21_ni ix34925 (.Y (nx34924), .A0 (nx34908), .A1 (nx34920), .S0 (nx23635)
             ) ;
    mux21_ni ix34909 (.Y (nx34908), .A0 (inputs_500__8), .A1 (inputs_501__8), .S0 (
             nx24387)) ;
    mux21_ni ix34921 (.Y (nx34920), .A0 (inputs_502__8), .A1 (inputs_503__8), .S0 (
             nx24387)) ;
    nand04 ix15580 (.Y (nx15579), .A0 (nx22305), .A1 (nx23635), .A2 (nx24387), .A3 (
           nx34868)) ;
    mux21_ni ix34869 (.Y (nx34868), .A0 (inputs_483__8), .A1 (inputs_499__8), .S0 (
             nx22901)) ;
    mux21_ni ix34855 (.Y (nx34854), .A0 (nx34790), .A1 (nx34850), .S0 (nx22903)
             ) ;
    mux21_ni ix34791 (.Y (nx34790), .A0 (nx34758), .A1 (nx34786), .S0 (nx23267)
             ) ;
    mux21_ni ix34759 (.Y (nx34758), .A0 (nx34742), .A1 (nx34754), .S0 (nx23635)
             ) ;
    mux21_ni ix34743 (.Y (nx34742), .A0 (inputs_488__8), .A1 (inputs_489__8), .S0 (
             nx24387)) ;
    mux21_ni ix34755 (.Y (nx34754), .A0 (inputs_490__8), .A1 (inputs_491__8), .S0 (
             nx24387)) ;
    mux21_ni ix34787 (.Y (nx34786), .A0 (nx34770), .A1 (nx34782), .S0 (nx23635)
             ) ;
    mux21_ni ix34771 (.Y (nx34770), .A0 (inputs_492__8), .A1 (inputs_493__8), .S0 (
             nx24387)) ;
    mux21_ni ix34783 (.Y (nx34782), .A0 (inputs_494__8), .A1 (inputs_495__8), .S0 (
             nx24389)) ;
    mux21_ni ix34851 (.Y (nx34850), .A0 (nx34818), .A1 (nx34846), .S0 (nx23267)
             ) ;
    mux21_ni ix34819 (.Y (nx34818), .A0 (nx34802), .A1 (nx34814), .S0 (nx23637)
             ) ;
    mux21_ni ix34803 (.Y (nx34802), .A0 (inputs_504__8), .A1 (inputs_505__8), .S0 (
             nx24389)) ;
    mux21_ni ix34815 (.Y (nx34814), .A0 (inputs_506__8), .A1 (inputs_507__8), .S0 (
             nx24389)) ;
    mux21_ni ix34847 (.Y (nx34846), .A0 (nx34830), .A1 (nx34842), .S0 (nx23637)
             ) ;
    mux21_ni ix34831 (.Y (nx34830), .A0 (inputs_508__8), .A1 (inputs_509__8), .S0 (
             nx24389)) ;
    mux21_ni ix34843 (.Y (nx34842), .A0 (inputs_510__8), .A1 (inputs_511__8), .S0 (
             nx24389)) ;
    aoi32 ix15608 (.Y (nx15607), .A0 (nx35716), .A1 (nx22387), .A2 (nx22307), .B0 (
          nx22221), .B1 (nx37412)) ;
    oai21 ix35717 (.Y (nx35716), .A0 (nx23637), .A1 (nx15611), .B0 (nx15713)) ;
    mux21 ix15612 (.Y (nx15611), .A0 (nx35454), .A1 (nx35706), .S0 (nx24389)) ;
    mux21_ni ix35455 (.Y (nx35454), .A0 (nx35326), .A1 (nx35450), .S0 (nx22399)
             ) ;
    mux21_ni ix35327 (.Y (nx35326), .A0 (nx35262), .A1 (nx35322), .S0 (nx22429)
             ) ;
    mux21_ni ix35263 (.Y (nx35262), .A0 (nx35230), .A1 (nx35258), .S0 (nx22487)
             ) ;
    mux21_ni ix35231 (.Y (nx35230), .A0 (nx35214), .A1 (nx35226), .S0 (nx22601)
             ) ;
    mux21_ni ix35215 (.Y (nx35214), .A0 (inputs_0__8), .A1 (inputs_16__8), .S0 (
             nx22903)) ;
    mux21_ni ix35227 (.Y (nx35226), .A0 (inputs_32__8), .A1 (inputs_48__8), .S0 (
             nx22903)) ;
    mux21_ni ix35259 (.Y (nx35258), .A0 (nx35242), .A1 (nx35254), .S0 (nx22601)
             ) ;
    mux21_ni ix35243 (.Y (nx35242), .A0 (inputs_64__8), .A1 (inputs_80__8), .S0 (
             nx22903)) ;
    mux21_ni ix35255 (.Y (nx35254), .A0 (inputs_96__8), .A1 (inputs_112__8), .S0 (
             nx22903)) ;
    mux21_ni ix35323 (.Y (nx35322), .A0 (nx35290), .A1 (nx35318), .S0 (nx22487)
             ) ;
    mux21_ni ix35291 (.Y (nx35290), .A0 (nx35274), .A1 (nx35286), .S0 (nx22601)
             ) ;
    mux21_ni ix35275 (.Y (nx35274), .A0 (inputs_128__8), .A1 (inputs_144__8), .S0 (
             nx22903)) ;
    mux21_ni ix35287 (.Y (nx35286), .A0 (inputs_160__8), .A1 (inputs_176__8), .S0 (
             nx22903)) ;
    mux21_ni ix35319 (.Y (nx35318), .A0 (nx35302), .A1 (nx35314), .S0 (nx22601)
             ) ;
    mux21_ni ix35303 (.Y (nx35302), .A0 (inputs_192__8), .A1 (inputs_208__8), .S0 (
             nx22905)) ;
    mux21_ni ix35315 (.Y (nx35314), .A0 (inputs_224__8), .A1 (inputs_240__8), .S0 (
             nx22905)) ;
    mux21_ni ix35451 (.Y (nx35450), .A0 (nx35386), .A1 (nx35446), .S0 (nx22429)
             ) ;
    mux21_ni ix35387 (.Y (nx35386), .A0 (nx35354), .A1 (nx35382), .S0 (nx22487)
             ) ;
    mux21_ni ix35355 (.Y (nx35354), .A0 (nx35338), .A1 (nx35350), .S0 (nx22601)
             ) ;
    mux21_ni ix35339 (.Y (nx35338), .A0 (inputs_256__8), .A1 (inputs_272__8), .S0 (
             nx22905)) ;
    mux21_ni ix35351 (.Y (nx35350), .A0 (inputs_288__8), .A1 (inputs_304__8), .S0 (
             nx22905)) ;
    mux21_ni ix35383 (.Y (nx35382), .A0 (nx35366), .A1 (nx35378), .S0 (nx22601)
             ) ;
    mux21_ni ix35367 (.Y (nx35366), .A0 (inputs_320__8), .A1 (inputs_336__8), .S0 (
             nx22905)) ;
    mux21_ni ix35379 (.Y (nx35378), .A0 (inputs_352__8), .A1 (inputs_368__8), .S0 (
             nx22905)) ;
    mux21_ni ix35447 (.Y (nx35446), .A0 (nx35414), .A1 (nx35442), .S0 (nx22489)
             ) ;
    mux21_ni ix35415 (.Y (nx35414), .A0 (nx35398), .A1 (nx35410), .S0 (nx22603)
             ) ;
    mux21_ni ix35399 (.Y (nx35398), .A0 (inputs_384__8), .A1 (inputs_400__8), .S0 (
             nx22905)) ;
    mux21_ni ix35411 (.Y (nx35410), .A0 (inputs_416__8), .A1 (inputs_432__8), .S0 (
             nx22907)) ;
    mux21_ni ix35443 (.Y (nx35442), .A0 (nx35426), .A1 (nx35438), .S0 (nx22603)
             ) ;
    mux21_ni ix35427 (.Y (nx35426), .A0 (inputs_448__8), .A1 (inputs_464__8), .S0 (
             nx22907)) ;
    mux21_ni ix35439 (.Y (nx35438), .A0 (inputs_480__8), .A1 (inputs_496__8), .S0 (
             nx22907)) ;
    mux21_ni ix35707 (.Y (nx35706), .A0 (nx35578), .A1 (nx35702), .S0 (nx22399)
             ) ;
    mux21_ni ix35579 (.Y (nx35578), .A0 (nx35514), .A1 (nx35574), .S0 (nx22429)
             ) ;
    mux21_ni ix35515 (.Y (nx35514), .A0 (nx35482), .A1 (nx35510), .S0 (nx22489)
             ) ;
    mux21_ni ix35483 (.Y (nx35482), .A0 (nx35466), .A1 (nx35478), .S0 (nx22603)
             ) ;
    mux21_ni ix35467 (.Y (nx35466), .A0 (inputs_1__8), .A1 (inputs_17__8), .S0 (
             nx22907)) ;
    mux21_ni ix35479 (.Y (nx35478), .A0 (inputs_33__8), .A1 (inputs_49__8), .S0 (
             nx22907)) ;
    mux21_ni ix35511 (.Y (nx35510), .A0 (nx35494), .A1 (nx35506), .S0 (nx22603)
             ) ;
    mux21_ni ix35495 (.Y (nx35494), .A0 (inputs_65__8), .A1 (inputs_81__8), .S0 (
             nx22907)) ;
    mux21_ni ix35507 (.Y (nx35506), .A0 (inputs_97__8), .A1 (inputs_113__8), .S0 (
             nx22907)) ;
    mux21_ni ix35575 (.Y (nx35574), .A0 (nx35542), .A1 (nx35570), .S0 (nx22489)
             ) ;
    mux21_ni ix35543 (.Y (nx35542), .A0 (nx35526), .A1 (nx35538), .S0 (nx22603)
             ) ;
    mux21_ni ix35527 (.Y (nx35526), .A0 (inputs_129__8), .A1 (inputs_145__8), .S0 (
             nx22909)) ;
    mux21_ni ix35539 (.Y (nx35538), .A0 (inputs_161__8), .A1 (inputs_177__8), .S0 (
             nx22909)) ;
    mux21_ni ix35571 (.Y (nx35570), .A0 (nx35554), .A1 (nx35566), .S0 (nx22603)
             ) ;
    mux21_ni ix35555 (.Y (nx35554), .A0 (inputs_193__8), .A1 (inputs_209__8), .S0 (
             nx22909)) ;
    mux21_ni ix35567 (.Y (nx35566), .A0 (inputs_225__8), .A1 (inputs_241__8), .S0 (
             nx22909)) ;
    mux21_ni ix35703 (.Y (nx35702), .A0 (nx35638), .A1 (nx35698), .S0 (nx22429)
             ) ;
    mux21_ni ix35639 (.Y (nx35638), .A0 (nx35606), .A1 (nx35634), .S0 (nx22489)
             ) ;
    mux21_ni ix35607 (.Y (nx35606), .A0 (nx35590), .A1 (nx35602), .S0 (nx22603)
             ) ;
    mux21_ni ix35591 (.Y (nx35590), .A0 (inputs_257__8), .A1 (inputs_273__8), .S0 (
             nx22909)) ;
    mux21_ni ix35603 (.Y (nx35602), .A0 (inputs_289__8), .A1 (inputs_305__8), .S0 (
             nx22909)) ;
    mux21_ni ix35635 (.Y (nx35634), .A0 (nx35618), .A1 (nx35630), .S0 (nx22605)
             ) ;
    mux21_ni ix35619 (.Y (nx35618), .A0 (inputs_321__8), .A1 (inputs_337__8), .S0 (
             nx22909)) ;
    mux21_ni ix35631 (.Y (nx35630), .A0 (inputs_353__8), .A1 (inputs_369__8), .S0 (
             nx22911)) ;
    mux21_ni ix35699 (.Y (nx35698), .A0 (nx35666), .A1 (nx35694), .S0 (nx22489)
             ) ;
    mux21_ni ix35667 (.Y (nx35666), .A0 (nx35650), .A1 (nx35662), .S0 (nx22605)
             ) ;
    mux21_ni ix35651 (.Y (nx35650), .A0 (inputs_385__8), .A1 (inputs_401__8), .S0 (
             nx22911)) ;
    mux21_ni ix35663 (.Y (nx35662), .A0 (inputs_417__8), .A1 (inputs_433__8), .S0 (
             nx22911)) ;
    mux21_ni ix35695 (.Y (nx35694), .A0 (nx35678), .A1 (nx35690), .S0 (nx22605)
             ) ;
    mux21_ni ix35679 (.Y (nx35678), .A0 (inputs_449__8), .A1 (inputs_465__8), .S0 (
             nx22911)) ;
    mux21_ni ix35691 (.Y (nx35690), .A0 (inputs_481__8), .A1 (inputs_497__8), .S0 (
             nx22911)) ;
    nand03 ix15714 (.Y (nx15713), .A0 (nx35200), .A1 (nx23637), .A2 (nx22381)) ;
    mux21_ni ix35201 (.Y (nx35200), .A0 (nx35072), .A1 (nx35196), .S0 (nx22399)
             ) ;
    mux21_ni ix35073 (.Y (nx35072), .A0 (nx35008), .A1 (nx35068), .S0 (nx22429)
             ) ;
    mux21_ni ix35009 (.Y (nx35008), .A0 (nx34976), .A1 (nx35004), .S0 (nx22489)
             ) ;
    mux21_ni ix34977 (.Y (nx34976), .A0 (nx34960), .A1 (nx34972), .S0 (nx22605)
             ) ;
    mux21_ni ix34961 (.Y (nx34960), .A0 (inputs_2__8), .A1 (inputs_18__8), .S0 (
             nx22911)) ;
    mux21_ni ix34973 (.Y (nx34972), .A0 (inputs_34__8), .A1 (inputs_50__8), .S0 (
             nx22911)) ;
    mux21_ni ix35005 (.Y (nx35004), .A0 (nx34988), .A1 (nx35000), .S0 (nx22605)
             ) ;
    mux21_ni ix34989 (.Y (nx34988), .A0 (inputs_66__8), .A1 (inputs_82__8), .S0 (
             nx22913)) ;
    mux21_ni ix35001 (.Y (nx35000), .A0 (inputs_98__8), .A1 (inputs_114__8), .S0 (
             nx22913)) ;
    mux21_ni ix35069 (.Y (nx35068), .A0 (nx35036), .A1 (nx35064), .S0 (nx22489)
             ) ;
    mux21_ni ix35037 (.Y (nx35036), .A0 (nx35020), .A1 (nx35032), .S0 (nx22605)
             ) ;
    mux21_ni ix35021 (.Y (nx35020), .A0 (inputs_130__8), .A1 (inputs_146__8), .S0 (
             nx22913)) ;
    mux21_ni ix35033 (.Y (nx35032), .A0 (inputs_162__8), .A1 (inputs_178__8), .S0 (
             nx22913)) ;
    mux21_ni ix35065 (.Y (nx35064), .A0 (nx35048), .A1 (nx35060), .S0 (nx22605)
             ) ;
    mux21_ni ix35049 (.Y (nx35048), .A0 (inputs_194__8), .A1 (inputs_210__8), .S0 (
             nx22913)) ;
    mux21_ni ix35061 (.Y (nx35060), .A0 (inputs_226__8), .A1 (inputs_242__8), .S0 (
             nx22913)) ;
    mux21_ni ix35197 (.Y (nx35196), .A0 (nx35132), .A1 (nx35192), .S0 (nx22431)
             ) ;
    mux21_ni ix35133 (.Y (nx35132), .A0 (nx35100), .A1 (nx35128), .S0 (nx22491)
             ) ;
    mux21_ni ix35101 (.Y (nx35100), .A0 (nx35084), .A1 (nx35096), .S0 (nx22607)
             ) ;
    mux21_ni ix35085 (.Y (nx35084), .A0 (inputs_258__8), .A1 (inputs_274__8), .S0 (
             nx22913)) ;
    mux21_ni ix35097 (.Y (nx35096), .A0 (inputs_290__8), .A1 (inputs_306__8), .S0 (
             nx22915)) ;
    mux21_ni ix35129 (.Y (nx35128), .A0 (nx35112), .A1 (nx35124), .S0 (nx22607)
             ) ;
    mux21_ni ix35113 (.Y (nx35112), .A0 (inputs_322__8), .A1 (inputs_338__8), .S0 (
             nx22915)) ;
    mux21_ni ix35125 (.Y (nx35124), .A0 (inputs_354__8), .A1 (inputs_370__8), .S0 (
             nx22915)) ;
    mux21_ni ix35193 (.Y (nx35192), .A0 (nx35160), .A1 (nx35188), .S0 (nx22491)
             ) ;
    mux21_ni ix35161 (.Y (nx35160), .A0 (nx35144), .A1 (nx35156), .S0 (nx22607)
             ) ;
    mux21_ni ix35145 (.Y (nx35144), .A0 (inputs_386__8), .A1 (inputs_402__8), .S0 (
             nx22915)) ;
    mux21_ni ix35157 (.Y (nx35156), .A0 (inputs_418__8), .A1 (inputs_434__8), .S0 (
             nx22915)) ;
    mux21_ni ix35189 (.Y (nx35188), .A0 (nx35172), .A1 (nx35184), .S0 (nx22607)
             ) ;
    mux21_ni ix35173 (.Y (nx35172), .A0 (inputs_450__8), .A1 (inputs_466__8), .S0 (
             nx22915)) ;
    mux21_ni ix35185 (.Y (nx35184), .A0 (inputs_482__8), .A1 (inputs_498__8), .S0 (
             nx22915)) ;
    mux21_ni ix37413 (.Y (nx37412), .A0 (nx36564), .A1 (nx37408), .S0 (nx22431)
             ) ;
    mux21_ni ix36565 (.Y (nx36564), .A0 (nx36140), .A1 (nx36560), .S0 (nx22491)
             ) ;
    mux21_ni ix36141 (.Y (nx36140), .A0 (nx35928), .A1 (nx36136), .S0 (nx22607)
             ) ;
    mux21_ni ix35929 (.Y (nx35928), .A0 (nx35922), .A1 (nx35844), .S0 (nx23155)
             ) ;
    oai21 ix35923 (.Y (nx35922), .A0 (nx22307), .A1 (nx15775), .B0 (nx15785)) ;
    mux21 ix15776 (.Y (nx15775), .A0 (nx35886), .A1 (nx35914), .S0 (nx22917)) ;
    mux21_ni ix35887 (.Y (nx35886), .A0 (nx35870), .A1 (nx35882), .S0 (nx23637)
             ) ;
    mux21_ni ix35871 (.Y (nx35870), .A0 (inputs_4__8), .A1 (inputs_5__8), .S0 (
             nx24389)) ;
    mux21_ni ix35883 (.Y (nx35882), .A0 (inputs_6__8), .A1 (inputs_7__8), .S0 (
             nx24391)) ;
    mux21_ni ix35915 (.Y (nx35914), .A0 (nx35898), .A1 (nx35910), .S0 (nx23637)
             ) ;
    mux21_ni ix35899 (.Y (nx35898), .A0 (inputs_20__8), .A1 (inputs_21__8), .S0 (
             nx24391)) ;
    mux21_ni ix35911 (.Y (nx35910), .A0 (inputs_22__8), .A1 (inputs_23__8), .S0 (
             nx24391)) ;
    nand04 ix15786 (.Y (nx15785), .A0 (nx22307), .A1 (nx23637), .A2 (nx24391), .A3 (
           nx35858)) ;
    mux21_ni ix35859 (.Y (nx35858), .A0 (inputs_3__8), .A1 (inputs_19__8), .S0 (
             nx22917)) ;
    mux21_ni ix35845 (.Y (nx35844), .A0 (nx35780), .A1 (nx35840), .S0 (nx22917)
             ) ;
    mux21_ni ix35781 (.Y (nx35780), .A0 (nx35748), .A1 (nx35776), .S0 (nx23267)
             ) ;
    mux21_ni ix35749 (.Y (nx35748), .A0 (nx35732), .A1 (nx35744), .S0 (nx23639)
             ) ;
    mux21_ni ix35733 (.Y (nx35732), .A0 (inputs_8__8), .A1 (inputs_9__8), .S0 (
             nx24391)) ;
    mux21_ni ix35745 (.Y (nx35744), .A0 (inputs_10__8), .A1 (inputs_11__8), .S0 (
             nx24391)) ;
    mux21_ni ix35777 (.Y (nx35776), .A0 (nx35760), .A1 (nx35772), .S0 (nx23639)
             ) ;
    mux21_ni ix35761 (.Y (nx35760), .A0 (inputs_12__8), .A1 (inputs_13__8), .S0 (
             nx24391)) ;
    mux21_ni ix35773 (.Y (nx35772), .A0 (inputs_14__8), .A1 (inputs_15__8), .S0 (
             nx24393)) ;
    mux21_ni ix35841 (.Y (nx35840), .A0 (nx35808), .A1 (nx35836), .S0 (nx23269)
             ) ;
    mux21_ni ix35809 (.Y (nx35808), .A0 (nx35792), .A1 (nx35804), .S0 (nx23639)
             ) ;
    mux21_ni ix35793 (.Y (nx35792), .A0 (inputs_24__8), .A1 (inputs_25__8), .S0 (
             nx24393)) ;
    mux21_ni ix35805 (.Y (nx35804), .A0 (inputs_26__8), .A1 (inputs_27__8), .S0 (
             nx24393)) ;
    mux21_ni ix35837 (.Y (nx35836), .A0 (nx35820), .A1 (nx35832), .S0 (nx23639)
             ) ;
    mux21_ni ix35821 (.Y (nx35820), .A0 (inputs_28__8), .A1 (inputs_29__8), .S0 (
             nx24393)) ;
    mux21_ni ix35833 (.Y (nx35832), .A0 (inputs_30__8), .A1 (inputs_31__8), .S0 (
             nx24393)) ;
    mux21_ni ix36137 (.Y (nx36136), .A0 (nx36130), .A1 (nx36052), .S0 (nx23155)
             ) ;
    oai21 ix36131 (.Y (nx36130), .A0 (nx22307), .A1 (nx15815), .B0 (nx15825)) ;
    mux21 ix15816 (.Y (nx15815), .A0 (nx36094), .A1 (nx36122), .S0 (nx22917)) ;
    mux21_ni ix36095 (.Y (nx36094), .A0 (nx36078), .A1 (nx36090), .S0 (nx23639)
             ) ;
    mux21_ni ix36079 (.Y (nx36078), .A0 (inputs_36__8), .A1 (inputs_37__8), .S0 (
             nx24393)) ;
    mux21_ni ix36091 (.Y (nx36090), .A0 (inputs_38__8), .A1 (inputs_39__8), .S0 (
             nx24393)) ;
    mux21_ni ix36123 (.Y (nx36122), .A0 (nx36106), .A1 (nx36118), .S0 (nx23639)
             ) ;
    mux21_ni ix36107 (.Y (nx36106), .A0 (inputs_52__8), .A1 (inputs_53__8), .S0 (
             nx24395)) ;
    mux21_ni ix36119 (.Y (nx36118), .A0 (inputs_54__8), .A1 (inputs_55__8), .S0 (
             nx24395)) ;
    nand04 ix15826 (.Y (nx15825), .A0 (nx22307), .A1 (nx23639), .A2 (nx24395), .A3 (
           nx36066)) ;
    mux21_ni ix36067 (.Y (nx36066), .A0 (inputs_35__8), .A1 (inputs_51__8), .S0 (
             nx22917)) ;
    mux21_ni ix36053 (.Y (nx36052), .A0 (nx35988), .A1 (nx36048), .S0 (nx22917)
             ) ;
    mux21_ni ix35989 (.Y (nx35988), .A0 (nx35956), .A1 (nx35984), .S0 (nx23269)
             ) ;
    mux21_ni ix35957 (.Y (nx35956), .A0 (nx35940), .A1 (nx35952), .S0 (nx23641)
             ) ;
    mux21_ni ix35941 (.Y (nx35940), .A0 (inputs_40__8), .A1 (inputs_41__8), .S0 (
             nx24395)) ;
    mux21_ni ix35953 (.Y (nx35952), .A0 (inputs_42__8), .A1 (inputs_43__8), .S0 (
             nx24395)) ;
    mux21_ni ix35985 (.Y (nx35984), .A0 (nx35968), .A1 (nx35980), .S0 (nx23641)
             ) ;
    mux21_ni ix35969 (.Y (nx35968), .A0 (inputs_44__8), .A1 (inputs_45__8), .S0 (
             nx24395)) ;
    mux21_ni ix35981 (.Y (nx35980), .A0 (inputs_46__8), .A1 (inputs_47__8), .S0 (
             nx24395)) ;
    mux21_ni ix36049 (.Y (nx36048), .A0 (nx36016), .A1 (nx36044), .S0 (nx23269)
             ) ;
    mux21_ni ix36017 (.Y (nx36016), .A0 (nx36000), .A1 (nx36012), .S0 (nx23641)
             ) ;
    mux21_ni ix36001 (.Y (nx36000), .A0 (inputs_56__8), .A1 (inputs_57__8), .S0 (
             nx24397)) ;
    mux21_ni ix36013 (.Y (nx36012), .A0 (inputs_58__8), .A1 (inputs_59__8), .S0 (
             nx24397)) ;
    mux21_ni ix36045 (.Y (nx36044), .A0 (nx36028), .A1 (nx36040), .S0 (nx23641)
             ) ;
    mux21_ni ix36029 (.Y (nx36028), .A0 (inputs_60__8), .A1 (inputs_61__8), .S0 (
             nx24397)) ;
    mux21_ni ix36041 (.Y (nx36040), .A0 (inputs_62__8), .A1 (inputs_63__8), .S0 (
             nx24397)) ;
    mux21_ni ix36561 (.Y (nx36560), .A0 (nx36348), .A1 (nx36556), .S0 (nx22607)
             ) ;
    mux21_ni ix36349 (.Y (nx36348), .A0 (nx36342), .A1 (nx36264), .S0 (nx23155)
             ) ;
    oai21 ix36343 (.Y (nx36342), .A0 (nx22307), .A1 (nx15857), .B0 (nx15869)) ;
    mux21 ix15858 (.Y (nx15857), .A0 (nx36306), .A1 (nx36334), .S0 (nx22917)) ;
    mux21_ni ix36307 (.Y (nx36306), .A0 (nx36290), .A1 (nx36302), .S0 (nx23641)
             ) ;
    mux21_ni ix36291 (.Y (nx36290), .A0 (inputs_68__8), .A1 (inputs_69__8), .S0 (
             nx24397)) ;
    mux21_ni ix36303 (.Y (nx36302), .A0 (inputs_70__8), .A1 (inputs_71__8), .S0 (
             nx24397)) ;
    mux21_ni ix36335 (.Y (nx36334), .A0 (nx36318), .A1 (nx36330), .S0 (nx23641)
             ) ;
    mux21_ni ix36319 (.Y (nx36318), .A0 (inputs_84__8), .A1 (inputs_85__8), .S0 (
             nx24397)) ;
    mux21_ni ix36331 (.Y (nx36330), .A0 (inputs_86__8), .A1 (inputs_87__8), .S0 (
             nx24399)) ;
    nand04 ix15870 (.Y (nx15869), .A0 (nx22307), .A1 (nx23641), .A2 (nx24399), .A3 (
           nx36278)) ;
    mux21_ni ix36279 (.Y (nx36278), .A0 (inputs_67__8), .A1 (inputs_83__8), .S0 (
             nx22919)) ;
    mux21_ni ix36265 (.Y (nx36264), .A0 (nx36200), .A1 (nx36260), .S0 (nx22919)
             ) ;
    mux21_ni ix36201 (.Y (nx36200), .A0 (nx36168), .A1 (nx36196), .S0 (nx23269)
             ) ;
    mux21_ni ix36169 (.Y (nx36168), .A0 (nx36152), .A1 (nx36164), .S0 (nx23643)
             ) ;
    mux21_ni ix36153 (.Y (nx36152), .A0 (inputs_72__8), .A1 (inputs_73__8), .S0 (
             nx24399)) ;
    mux21_ni ix36165 (.Y (nx36164), .A0 (inputs_74__8), .A1 (inputs_75__8), .S0 (
             nx24399)) ;
    mux21_ni ix36197 (.Y (nx36196), .A0 (nx36180), .A1 (nx36192), .S0 (nx23643)
             ) ;
    mux21_ni ix36181 (.Y (nx36180), .A0 (inputs_76__8), .A1 (inputs_77__8), .S0 (
             nx24399)) ;
    mux21_ni ix36193 (.Y (nx36192), .A0 (inputs_78__8), .A1 (inputs_79__8), .S0 (
             nx24399)) ;
    mux21_ni ix36261 (.Y (nx36260), .A0 (nx36228), .A1 (nx36256), .S0 (nx23269)
             ) ;
    mux21_ni ix36229 (.Y (nx36228), .A0 (nx36212), .A1 (nx36224), .S0 (nx23643)
             ) ;
    mux21_ni ix36213 (.Y (nx36212), .A0 (inputs_88__8), .A1 (inputs_89__8), .S0 (
             nx24399)) ;
    mux21_ni ix36225 (.Y (nx36224), .A0 (inputs_90__8), .A1 (inputs_91__8), .S0 (
             nx24401)) ;
    mux21_ni ix36257 (.Y (nx36256), .A0 (nx36240), .A1 (nx36252), .S0 (nx23643)
             ) ;
    mux21_ni ix36241 (.Y (nx36240), .A0 (inputs_92__8), .A1 (inputs_93__8), .S0 (
             nx24401)) ;
    mux21_ni ix36253 (.Y (nx36252), .A0 (inputs_94__8), .A1 (inputs_95__8), .S0 (
             nx24401)) ;
    mux21_ni ix36557 (.Y (nx36556), .A0 (nx36550), .A1 (nx36472), .S0 (nx23155)
             ) ;
    oai21 ix36551 (.Y (nx36550), .A0 (nx22309), .A1 (nx15903), .B0 (nx15915)) ;
    mux21 ix15904 (.Y (nx15903), .A0 (nx36514), .A1 (nx36542), .S0 (nx22919)) ;
    mux21_ni ix36515 (.Y (nx36514), .A0 (nx36498), .A1 (nx36510), .S0 (nx23643)
             ) ;
    mux21_ni ix36499 (.Y (nx36498), .A0 (inputs_100__8), .A1 (inputs_101__8), .S0 (
             nx24401)) ;
    mux21_ni ix36511 (.Y (nx36510), .A0 (inputs_102__8), .A1 (inputs_103__8), .S0 (
             nx24401)) ;
    mux21_ni ix36543 (.Y (nx36542), .A0 (nx36526), .A1 (nx36538), .S0 (nx23643)
             ) ;
    mux21_ni ix36527 (.Y (nx36526), .A0 (inputs_116__8), .A1 (inputs_117__8), .S0 (
             nx24401)) ;
    mux21_ni ix36539 (.Y (nx36538), .A0 (inputs_118__8), .A1 (inputs_119__8), .S0 (
             nx24401)) ;
    nand04 ix15916 (.Y (nx15915), .A0 (nx22309), .A1 (nx23643), .A2 (nx24403), .A3 (
           nx36486)) ;
    mux21_ni ix36487 (.Y (nx36486), .A0 (inputs_99__8), .A1 (inputs_115__8), .S0 (
             nx22919)) ;
    mux21_ni ix36473 (.Y (nx36472), .A0 (nx36408), .A1 (nx36468), .S0 (nx22919)
             ) ;
    mux21_ni ix36409 (.Y (nx36408), .A0 (nx36376), .A1 (nx36404), .S0 (nx23269)
             ) ;
    mux21_ni ix36377 (.Y (nx36376), .A0 (nx36360), .A1 (nx36372), .S0 (nx23645)
             ) ;
    mux21_ni ix36361 (.Y (nx36360), .A0 (inputs_104__8), .A1 (inputs_105__8), .S0 (
             nx24403)) ;
    mux21_ni ix36373 (.Y (nx36372), .A0 (inputs_106__8), .A1 (inputs_107__8), .S0 (
             nx24403)) ;
    mux21_ni ix36405 (.Y (nx36404), .A0 (nx36388), .A1 (nx36400), .S0 (nx23645)
             ) ;
    mux21_ni ix36389 (.Y (nx36388), .A0 (inputs_108__8), .A1 (inputs_109__8), .S0 (
             nx24403)) ;
    mux21_ni ix36401 (.Y (nx36400), .A0 (inputs_110__8), .A1 (inputs_111__8), .S0 (
             nx24403)) ;
    mux21_ni ix36469 (.Y (nx36468), .A0 (nx36436), .A1 (nx36464), .S0 (nx23269)
             ) ;
    mux21_ni ix36437 (.Y (nx36436), .A0 (nx36420), .A1 (nx36432), .S0 (nx23645)
             ) ;
    mux21_ni ix36421 (.Y (nx36420), .A0 (inputs_120__8), .A1 (inputs_121__8), .S0 (
             nx24403)) ;
    mux21_ni ix36433 (.Y (nx36432), .A0 (inputs_122__8), .A1 (inputs_123__8), .S0 (
             nx24403)) ;
    mux21_ni ix36465 (.Y (nx36464), .A0 (nx36448), .A1 (nx36460), .S0 (nx23645)
             ) ;
    mux21_ni ix36449 (.Y (nx36448), .A0 (inputs_124__8), .A1 (inputs_125__8), .S0 (
             nx24405)) ;
    mux21_ni ix36461 (.Y (nx36460), .A0 (inputs_126__8), .A1 (inputs_127__8), .S0 (
             nx24405)) ;
    mux21_ni ix37409 (.Y (nx37408), .A0 (nx36984), .A1 (nx37404), .S0 (nx22491)
             ) ;
    mux21_ni ix36985 (.Y (nx36984), .A0 (nx36772), .A1 (nx36980), .S0 (nx22607)
             ) ;
    mux21_ni ix36773 (.Y (nx36772), .A0 (nx36766), .A1 (nx36688), .S0 (nx23157)
             ) ;
    oai21 ix36767 (.Y (nx36766), .A0 (nx22309), .A1 (nx15949), .B0 (nx15961)) ;
    mux21 ix15950 (.Y (nx15949), .A0 (nx36730), .A1 (nx36758), .S0 (nx22919)) ;
    mux21_ni ix36731 (.Y (nx36730), .A0 (nx36714), .A1 (nx36726), .S0 (nx23645)
             ) ;
    mux21_ni ix36715 (.Y (nx36714), .A0 (inputs_132__8), .A1 (inputs_133__8), .S0 (
             nx24405)) ;
    mux21_ni ix36727 (.Y (nx36726), .A0 (inputs_134__8), .A1 (inputs_135__8), .S0 (
             nx24405)) ;
    mux21_ni ix36759 (.Y (nx36758), .A0 (nx36742), .A1 (nx36754), .S0 (nx23645)
             ) ;
    mux21_ni ix36743 (.Y (nx36742), .A0 (inputs_148__8), .A1 (inputs_149__8), .S0 (
             nx24405)) ;
    mux21_ni ix36755 (.Y (nx36754), .A0 (inputs_150__8), .A1 (inputs_151__8), .S0 (
             nx24405)) ;
    nand04 ix15962 (.Y (nx15961), .A0 (nx22309), .A1 (nx23645), .A2 (nx24405), .A3 (
           nx36702)) ;
    mux21_ni ix36703 (.Y (nx36702), .A0 (inputs_131__8), .A1 (inputs_147__8), .S0 (
             nx22919)) ;
    mux21_ni ix36689 (.Y (nx36688), .A0 (nx36624), .A1 (nx36684), .S0 (nx22921)
             ) ;
    mux21_ni ix36625 (.Y (nx36624), .A0 (nx36592), .A1 (nx36620), .S0 (nx23271)
             ) ;
    mux21_ni ix36593 (.Y (nx36592), .A0 (nx36576), .A1 (nx36588), .S0 (nx23647)
             ) ;
    mux21_ni ix36577 (.Y (nx36576), .A0 (inputs_136__8), .A1 (inputs_137__8), .S0 (
             nx24407)) ;
    mux21_ni ix36589 (.Y (nx36588), .A0 (inputs_138__8), .A1 (inputs_139__8), .S0 (
             nx24407)) ;
    mux21_ni ix36621 (.Y (nx36620), .A0 (nx36604), .A1 (nx36616), .S0 (nx23647)
             ) ;
    mux21_ni ix36605 (.Y (nx36604), .A0 (inputs_140__8), .A1 (inputs_141__8), .S0 (
             nx24407)) ;
    mux21_ni ix36617 (.Y (nx36616), .A0 (inputs_142__8), .A1 (inputs_143__8), .S0 (
             nx24407)) ;
    mux21_ni ix36685 (.Y (nx36684), .A0 (nx36652), .A1 (nx36680), .S0 (nx23271)
             ) ;
    mux21_ni ix36653 (.Y (nx36652), .A0 (nx36636), .A1 (nx36648), .S0 (nx23647)
             ) ;
    mux21_ni ix36637 (.Y (nx36636), .A0 (inputs_152__8), .A1 (inputs_153__8), .S0 (
             nx24407)) ;
    mux21_ni ix36649 (.Y (nx36648), .A0 (inputs_154__8), .A1 (inputs_155__8), .S0 (
             nx24407)) ;
    mux21_ni ix36681 (.Y (nx36680), .A0 (nx36664), .A1 (nx36676), .S0 (nx23647)
             ) ;
    mux21_ni ix36665 (.Y (nx36664), .A0 (inputs_156__8), .A1 (inputs_157__8), .S0 (
             nx24407)) ;
    mux21_ni ix36677 (.Y (nx36676), .A0 (inputs_158__8), .A1 (inputs_159__8), .S0 (
             nx24409)) ;
    mux21_ni ix36981 (.Y (nx36980), .A0 (nx36974), .A1 (nx36896), .S0 (nx23157)
             ) ;
    oai21 ix36975 (.Y (nx36974), .A0 (nx22309), .A1 (nx15993), .B0 (nx16003)) ;
    mux21 ix15994 (.Y (nx15993), .A0 (nx36938), .A1 (nx36966), .S0 (nx22921)) ;
    mux21_ni ix36939 (.Y (nx36938), .A0 (nx36922), .A1 (nx36934), .S0 (nx23647)
             ) ;
    mux21_ni ix36923 (.Y (nx36922), .A0 (inputs_164__8), .A1 (inputs_165__8), .S0 (
             nx24409)) ;
    mux21_ni ix36935 (.Y (nx36934), .A0 (inputs_166__8), .A1 (inputs_167__8), .S0 (
             nx24409)) ;
    mux21_ni ix36967 (.Y (nx36966), .A0 (nx36950), .A1 (nx36962), .S0 (nx23647)
             ) ;
    mux21_ni ix36951 (.Y (nx36950), .A0 (inputs_180__8), .A1 (inputs_181__8), .S0 (
             nx24409)) ;
    mux21_ni ix36963 (.Y (nx36962), .A0 (inputs_182__8), .A1 (inputs_183__8), .S0 (
             nx24409)) ;
    nand04 ix16004 (.Y (nx16003), .A0 (nx22309), .A1 (nx23647), .A2 (nx24409), .A3 (
           nx36910)) ;
    mux21_ni ix36911 (.Y (nx36910), .A0 (inputs_163__8), .A1 (inputs_179__8), .S0 (
             nx22921)) ;
    mux21_ni ix36897 (.Y (nx36896), .A0 (nx36832), .A1 (nx36892), .S0 (nx22921)
             ) ;
    mux21_ni ix36833 (.Y (nx36832), .A0 (nx36800), .A1 (nx36828), .S0 (nx23271)
             ) ;
    mux21_ni ix36801 (.Y (nx36800), .A0 (nx36784), .A1 (nx36796), .S0 (nx23649)
             ) ;
    mux21_ni ix36785 (.Y (nx36784), .A0 (inputs_168__8), .A1 (inputs_169__8), .S0 (
             nx24409)) ;
    mux21_ni ix36797 (.Y (nx36796), .A0 (inputs_170__8), .A1 (inputs_171__8), .S0 (
             nx24411)) ;
    mux21_ni ix36829 (.Y (nx36828), .A0 (nx36812), .A1 (nx36824), .S0 (nx23649)
             ) ;
    mux21_ni ix36813 (.Y (nx36812), .A0 (inputs_172__8), .A1 (inputs_173__8), .S0 (
             nx24411)) ;
    mux21_ni ix36825 (.Y (nx36824), .A0 (inputs_174__8), .A1 (inputs_175__8), .S0 (
             nx24411)) ;
    mux21_ni ix36893 (.Y (nx36892), .A0 (nx36860), .A1 (nx36888), .S0 (nx23271)
             ) ;
    mux21_ni ix36861 (.Y (nx36860), .A0 (nx36844), .A1 (nx36856), .S0 (nx23649)
             ) ;
    mux21_ni ix36845 (.Y (nx36844), .A0 (inputs_184__8), .A1 (inputs_185__8), .S0 (
             nx24411)) ;
    mux21_ni ix36857 (.Y (nx36856), .A0 (inputs_186__8), .A1 (inputs_187__8), .S0 (
             nx24411)) ;
    mux21_ni ix36889 (.Y (nx36888), .A0 (nx36872), .A1 (nx36884), .S0 (nx23649)
             ) ;
    mux21_ni ix36873 (.Y (nx36872), .A0 (inputs_188__8), .A1 (inputs_189__8), .S0 (
             nx24411)) ;
    mux21_ni ix36885 (.Y (nx36884), .A0 (inputs_190__8), .A1 (inputs_191__8), .S0 (
             nx24411)) ;
    mux21_ni ix37405 (.Y (nx37404), .A0 (nx37192), .A1 (nx37400), .S0 (nx22609)
             ) ;
    mux21_ni ix37193 (.Y (nx37192), .A0 (nx37186), .A1 (nx37108), .S0 (nx23157)
             ) ;
    oai21 ix37187 (.Y (nx37186), .A0 (nx22309), .A1 (nx16035), .B0 (nx16047)) ;
    mux21 ix16036 (.Y (nx16035), .A0 (nx37150), .A1 (nx37178), .S0 (nx22921)) ;
    mux21_ni ix37151 (.Y (nx37150), .A0 (nx37134), .A1 (nx37146), .S0 (nx23649)
             ) ;
    mux21_ni ix37135 (.Y (nx37134), .A0 (inputs_196__8), .A1 (inputs_197__8), .S0 (
             nx24413)) ;
    mux21_ni ix37147 (.Y (nx37146), .A0 (inputs_198__8), .A1 (inputs_199__8), .S0 (
             nx24413)) ;
    mux21_ni ix37179 (.Y (nx37178), .A0 (nx37162), .A1 (nx37174), .S0 (nx23649)
             ) ;
    mux21_ni ix37163 (.Y (nx37162), .A0 (inputs_212__8), .A1 (inputs_213__8), .S0 (
             nx24413)) ;
    mux21_ni ix37175 (.Y (nx37174), .A0 (inputs_214__8), .A1 (inputs_215__8), .S0 (
             nx24413)) ;
    nand04 ix16048 (.Y (nx16047), .A0 (nx22311), .A1 (nx23649), .A2 (nx24413), .A3 (
           nx37122)) ;
    mux21_ni ix37123 (.Y (nx37122), .A0 (inputs_195__8), .A1 (inputs_211__8), .S0 (
             nx22921)) ;
    mux21_ni ix37109 (.Y (nx37108), .A0 (nx37044), .A1 (nx37104), .S0 (nx22921)
             ) ;
    mux21_ni ix37045 (.Y (nx37044), .A0 (nx37012), .A1 (nx37040), .S0 (nx23271)
             ) ;
    mux21_ni ix37013 (.Y (nx37012), .A0 (nx36996), .A1 (nx37008), .S0 (nx23651)
             ) ;
    mux21_ni ix36997 (.Y (nx36996), .A0 (inputs_200__8), .A1 (inputs_201__8), .S0 (
             nx24413)) ;
    mux21_ni ix37009 (.Y (nx37008), .A0 (inputs_202__8), .A1 (inputs_203__8), .S0 (
             nx24413)) ;
    mux21_ni ix37041 (.Y (nx37040), .A0 (nx37024), .A1 (nx37036), .S0 (nx23651)
             ) ;
    mux21_ni ix37025 (.Y (nx37024), .A0 (inputs_204__8), .A1 (inputs_205__8), .S0 (
             nx24415)) ;
    mux21_ni ix37037 (.Y (nx37036), .A0 (inputs_206__8), .A1 (inputs_207__8), .S0 (
             nx24415)) ;
    mux21_ni ix37105 (.Y (nx37104), .A0 (nx37072), .A1 (nx37100), .S0 (nx23271)
             ) ;
    mux21_ni ix37073 (.Y (nx37072), .A0 (nx37056), .A1 (nx37068), .S0 (nx23651)
             ) ;
    mux21_ni ix37057 (.Y (nx37056), .A0 (inputs_216__8), .A1 (inputs_217__8), .S0 (
             nx24415)) ;
    mux21_ni ix37069 (.Y (nx37068), .A0 (inputs_218__8), .A1 (inputs_219__8), .S0 (
             nx24415)) ;
    mux21_ni ix37101 (.Y (nx37100), .A0 (nx37084), .A1 (nx37096), .S0 (nx23651)
             ) ;
    mux21_ni ix37085 (.Y (nx37084), .A0 (inputs_220__8), .A1 (inputs_221__8), .S0 (
             nx24415)) ;
    mux21_ni ix37097 (.Y (nx37096), .A0 (inputs_222__8), .A1 (inputs_223__8), .S0 (
             nx24415)) ;
    mux21_ni ix37401 (.Y (nx37400), .A0 (nx37394), .A1 (nx37316), .S0 (nx23157)
             ) ;
    oai21 ix37395 (.Y (nx37394), .A0 (nx22311), .A1 (nx16077), .B0 (nx16089)) ;
    mux21 ix16078 (.Y (nx16077), .A0 (nx37358), .A1 (nx37386), .S0 (nx22923)) ;
    mux21_ni ix37359 (.Y (nx37358), .A0 (nx37342), .A1 (nx37354), .S0 (nx23651)
             ) ;
    mux21_ni ix37343 (.Y (nx37342), .A0 (inputs_228__8), .A1 (inputs_229__8), .S0 (
             nx24415)) ;
    mux21_ni ix37355 (.Y (nx37354), .A0 (inputs_230__8), .A1 (inputs_231__8), .S0 (
             nx24417)) ;
    mux21_ni ix37387 (.Y (nx37386), .A0 (nx37370), .A1 (nx37382), .S0 (nx23651)
             ) ;
    mux21_ni ix37371 (.Y (nx37370), .A0 (inputs_244__8), .A1 (inputs_245__8), .S0 (
             nx24417)) ;
    mux21_ni ix37383 (.Y (nx37382), .A0 (inputs_246__8), .A1 (inputs_247__8), .S0 (
             nx24417)) ;
    nand04 ix16090 (.Y (nx16089), .A0 (nx22311), .A1 (nx23651), .A2 (nx24417), .A3 (
           nx37330)) ;
    mux21_ni ix37331 (.Y (nx37330), .A0 (inputs_227__8), .A1 (inputs_243__8), .S0 (
             nx22923)) ;
    mux21_ni ix37317 (.Y (nx37316), .A0 (nx37252), .A1 (nx37312), .S0 (nx22923)
             ) ;
    mux21_ni ix37253 (.Y (nx37252), .A0 (nx37220), .A1 (nx37248), .S0 (nx23271)
             ) ;
    mux21_ni ix37221 (.Y (nx37220), .A0 (nx37204), .A1 (nx37216), .S0 (nx23653)
             ) ;
    mux21_ni ix37205 (.Y (nx37204), .A0 (inputs_232__8), .A1 (inputs_233__8), .S0 (
             nx24417)) ;
    mux21_ni ix37217 (.Y (nx37216), .A0 (inputs_234__8), .A1 (inputs_235__8), .S0 (
             nx24417)) ;
    mux21_ni ix37249 (.Y (nx37248), .A0 (nx37232), .A1 (nx37244), .S0 (nx23653)
             ) ;
    mux21_ni ix37233 (.Y (nx37232), .A0 (inputs_236__8), .A1 (inputs_237__8), .S0 (
             nx24417)) ;
    mux21_ni ix37245 (.Y (nx37244), .A0 (inputs_238__8), .A1 (inputs_239__8), .S0 (
             nx24419)) ;
    mux21_ni ix37313 (.Y (nx37312), .A0 (nx37280), .A1 (nx37308), .S0 (nx23273)
             ) ;
    mux21_ni ix37281 (.Y (nx37280), .A0 (nx37264), .A1 (nx37276), .S0 (nx23653)
             ) ;
    mux21_ni ix37265 (.Y (nx37264), .A0 (inputs_248__8), .A1 (inputs_249__8), .S0 (
             nx24419)) ;
    mux21_ni ix37277 (.Y (nx37276), .A0 (inputs_250__8), .A1 (inputs_251__8), .S0 (
             nx24419)) ;
    mux21_ni ix37309 (.Y (nx37308), .A0 (nx37292), .A1 (nx37304), .S0 (nx23653)
             ) ;
    mux21_ni ix37293 (.Y (nx37292), .A0 (inputs_252__8), .A1 (inputs_253__8), .S0 (
             nx24419)) ;
    mux21_ni ix37305 (.Y (nx37304), .A0 (inputs_254__8), .A1 (inputs_255__8), .S0 (
             nx24419)) ;
    oai21 ix41579 (.Y (\output [9]), .A0 (nx22221), .A1 (nx16121), .B0 (nx16475)
          ) ;
    mux21 ix16122 (.Y (nx16121), .A0 (nx38260), .A1 (nx39104), .S0 (nx22431)) ;
    mux21_ni ix38261 (.Y (nx38260), .A0 (nx37836), .A1 (nx38256), .S0 (nx22491)
             ) ;
    mux21_ni ix37837 (.Y (nx37836), .A0 (nx37624), .A1 (nx37832), .S0 (nx22609)
             ) ;
    mux21_ni ix37625 (.Y (nx37624), .A0 (nx37618), .A1 (nx37540), .S0 (nx23157)
             ) ;
    oai21 ix37619 (.Y (nx37618), .A0 (nx22311), .A1 (nx16129), .B0 (nx16141)) ;
    mux21 ix16130 (.Y (nx16129), .A0 (nx37582), .A1 (nx37610), .S0 (nx22923)) ;
    mux21_ni ix37583 (.Y (nx37582), .A0 (nx37566), .A1 (nx37578), .S0 (nx23653)
             ) ;
    mux21_ni ix37567 (.Y (nx37566), .A0 (inputs_260__9), .A1 (inputs_261__9), .S0 (
             nx24419)) ;
    mux21_ni ix37579 (.Y (nx37578), .A0 (inputs_262__9), .A1 (inputs_263__9), .S0 (
             nx24419)) ;
    mux21_ni ix37611 (.Y (nx37610), .A0 (nx37594), .A1 (nx37606), .S0 (nx23653)
             ) ;
    mux21_ni ix37595 (.Y (nx37594), .A0 (inputs_276__9), .A1 (inputs_277__9), .S0 (
             nx24421)) ;
    mux21_ni ix37607 (.Y (nx37606), .A0 (inputs_278__9), .A1 (inputs_279__9), .S0 (
             nx24421)) ;
    nand04 ix16142 (.Y (nx16141), .A0 (nx22311), .A1 (nx23653), .A2 (nx24421), .A3 (
           nx37554)) ;
    mux21_ni ix37555 (.Y (nx37554), .A0 (inputs_259__9), .A1 (inputs_275__9), .S0 (
             nx22923)) ;
    mux21_ni ix37541 (.Y (nx37540), .A0 (nx37476), .A1 (nx37536), .S0 (nx22923)
             ) ;
    mux21_ni ix37477 (.Y (nx37476), .A0 (nx37444), .A1 (nx37472), .S0 (nx23273)
             ) ;
    mux21_ni ix37445 (.Y (nx37444), .A0 (nx37428), .A1 (nx37440), .S0 (nx23655)
             ) ;
    mux21_ni ix37429 (.Y (nx37428), .A0 (inputs_264__9), .A1 (inputs_265__9), .S0 (
             nx24421)) ;
    mux21_ni ix37441 (.Y (nx37440), .A0 (inputs_266__9), .A1 (inputs_267__9), .S0 (
             nx24421)) ;
    mux21_ni ix37473 (.Y (nx37472), .A0 (nx37456), .A1 (nx37468), .S0 (nx23655)
             ) ;
    mux21_ni ix37457 (.Y (nx37456), .A0 (inputs_268__9), .A1 (inputs_269__9), .S0 (
             nx24421)) ;
    mux21_ni ix37469 (.Y (nx37468), .A0 (inputs_270__9), .A1 (inputs_271__9), .S0 (
             nx24421)) ;
    mux21_ni ix37537 (.Y (nx37536), .A0 (nx37504), .A1 (nx37532), .S0 (nx23273)
             ) ;
    mux21_ni ix37505 (.Y (nx37504), .A0 (nx37488), .A1 (nx37500), .S0 (nx23655)
             ) ;
    mux21_ni ix37489 (.Y (nx37488), .A0 (inputs_280__9), .A1 (inputs_281__9), .S0 (
             nx24423)) ;
    mux21_ni ix37501 (.Y (nx37500), .A0 (inputs_282__9), .A1 (inputs_283__9), .S0 (
             nx24423)) ;
    mux21_ni ix37533 (.Y (nx37532), .A0 (nx37516), .A1 (nx37528), .S0 (nx23655)
             ) ;
    mux21_ni ix37517 (.Y (nx37516), .A0 (inputs_284__9), .A1 (inputs_285__9), .S0 (
             nx24423)) ;
    mux21_ni ix37529 (.Y (nx37528), .A0 (inputs_286__9), .A1 (inputs_287__9), .S0 (
             nx24423)) ;
    mux21_ni ix37833 (.Y (nx37832), .A0 (nx37826), .A1 (nx37748), .S0 (nx23157)
             ) ;
    oai21 ix37827 (.Y (nx37826), .A0 (nx22311), .A1 (nx16171), .B0 (nx16185)) ;
    mux21 ix16172 (.Y (nx16171), .A0 (nx37790), .A1 (nx37818), .S0 (nx22923)) ;
    mux21_ni ix37791 (.Y (nx37790), .A0 (nx37774), .A1 (nx37786), .S0 (nx23655)
             ) ;
    mux21_ni ix37775 (.Y (nx37774), .A0 (inputs_292__9), .A1 (inputs_293__9), .S0 (
             nx24423)) ;
    mux21_ni ix37787 (.Y (nx37786), .A0 (inputs_294__9), .A1 (inputs_295__9), .S0 (
             nx24423)) ;
    mux21_ni ix37819 (.Y (nx37818), .A0 (nx37802), .A1 (nx37814), .S0 (nx23655)
             ) ;
    mux21_ni ix37803 (.Y (nx37802), .A0 (inputs_308__9), .A1 (inputs_309__9), .S0 (
             nx24423)) ;
    mux21_ni ix37815 (.Y (nx37814), .A0 (inputs_310__9), .A1 (inputs_311__9), .S0 (
             nx24425)) ;
    nand04 ix16186 (.Y (nx16185), .A0 (nx22311), .A1 (nx23655), .A2 (nx24425), .A3 (
           nx37762)) ;
    mux21_ni ix37763 (.Y (nx37762), .A0 (inputs_291__9), .A1 (inputs_307__9), .S0 (
             nx22925)) ;
    mux21_ni ix37749 (.Y (nx37748), .A0 (nx37684), .A1 (nx37744), .S0 (nx22925)
             ) ;
    mux21_ni ix37685 (.Y (nx37684), .A0 (nx37652), .A1 (nx37680), .S0 (nx23273)
             ) ;
    mux21_ni ix37653 (.Y (nx37652), .A0 (nx37636), .A1 (nx37648), .S0 (nx23657)
             ) ;
    mux21_ni ix37637 (.Y (nx37636), .A0 (inputs_296__9), .A1 (inputs_297__9), .S0 (
             nx24425)) ;
    mux21_ni ix37649 (.Y (nx37648), .A0 (inputs_298__9), .A1 (inputs_299__9), .S0 (
             nx24425)) ;
    mux21_ni ix37681 (.Y (nx37680), .A0 (nx37664), .A1 (nx37676), .S0 (nx23657)
             ) ;
    mux21_ni ix37665 (.Y (nx37664), .A0 (inputs_300__9), .A1 (inputs_301__9), .S0 (
             nx24425)) ;
    mux21_ni ix37677 (.Y (nx37676), .A0 (inputs_302__9), .A1 (inputs_303__9), .S0 (
             nx24425)) ;
    mux21_ni ix37745 (.Y (nx37744), .A0 (nx37712), .A1 (nx37740), .S0 (nx23273)
             ) ;
    mux21_ni ix37713 (.Y (nx37712), .A0 (nx37696), .A1 (nx37708), .S0 (nx23657)
             ) ;
    mux21_ni ix37697 (.Y (nx37696), .A0 (inputs_312__9), .A1 (inputs_313__9), .S0 (
             nx24425)) ;
    mux21_ni ix37709 (.Y (nx37708), .A0 (inputs_314__9), .A1 (inputs_315__9), .S0 (
             nx24427)) ;
    mux21_ni ix37741 (.Y (nx37740), .A0 (nx37724), .A1 (nx37736), .S0 (nx23657)
             ) ;
    mux21_ni ix37725 (.Y (nx37724), .A0 (inputs_316__9), .A1 (inputs_317__9), .S0 (
             nx24427)) ;
    mux21_ni ix37737 (.Y (nx37736), .A0 (inputs_318__9), .A1 (inputs_319__9), .S0 (
             nx24427)) ;
    mux21_ni ix38257 (.Y (nx38256), .A0 (nx38044), .A1 (nx38252), .S0 (nx22609)
             ) ;
    mux21_ni ix38045 (.Y (nx38044), .A0 (nx38038), .A1 (nx37960), .S0 (nx23157)
             ) ;
    oai21 ix38039 (.Y (nx38038), .A0 (nx22313), .A1 (nx16215), .B0 (nx16227)) ;
    mux21 ix16216 (.Y (nx16215), .A0 (nx38002), .A1 (nx38030), .S0 (nx22925)) ;
    mux21_ni ix38003 (.Y (nx38002), .A0 (nx37986), .A1 (nx37998), .S0 (nx23657)
             ) ;
    mux21_ni ix37987 (.Y (nx37986), .A0 (inputs_324__9), .A1 (inputs_325__9), .S0 (
             nx24427)) ;
    mux21_ni ix37999 (.Y (nx37998), .A0 (inputs_326__9), .A1 (inputs_327__9), .S0 (
             nx24427)) ;
    mux21_ni ix38031 (.Y (nx38030), .A0 (nx38014), .A1 (nx38026), .S0 (nx23657)
             ) ;
    mux21_ni ix38015 (.Y (nx38014), .A0 (inputs_340__9), .A1 (inputs_341__9), .S0 (
             nx24427)) ;
    mux21_ni ix38027 (.Y (nx38026), .A0 (inputs_342__9), .A1 (inputs_343__9), .S0 (
             nx24427)) ;
    nand04 ix16228 (.Y (nx16227), .A0 (nx22313), .A1 (nx23657), .A2 (nx24429), .A3 (
           nx37974)) ;
    mux21_ni ix37975 (.Y (nx37974), .A0 (inputs_323__9), .A1 (inputs_339__9), .S0 (
             nx22925)) ;
    mux21_ni ix37961 (.Y (nx37960), .A0 (nx37896), .A1 (nx37956), .S0 (nx22925)
             ) ;
    mux21_ni ix37897 (.Y (nx37896), .A0 (nx37864), .A1 (nx37892), .S0 (nx23273)
             ) ;
    mux21_ni ix37865 (.Y (nx37864), .A0 (nx37848), .A1 (nx37860), .S0 (nx23659)
             ) ;
    mux21_ni ix37849 (.Y (nx37848), .A0 (inputs_328__9), .A1 (inputs_329__9), .S0 (
             nx24429)) ;
    mux21_ni ix37861 (.Y (nx37860), .A0 (inputs_330__9), .A1 (inputs_331__9), .S0 (
             nx24429)) ;
    mux21_ni ix37893 (.Y (nx37892), .A0 (nx37876), .A1 (nx37888), .S0 (nx23659)
             ) ;
    mux21_ni ix37877 (.Y (nx37876), .A0 (inputs_332__9), .A1 (inputs_333__9), .S0 (
             nx24429)) ;
    mux21_ni ix37889 (.Y (nx37888), .A0 (inputs_334__9), .A1 (inputs_335__9), .S0 (
             nx24429)) ;
    mux21_ni ix37957 (.Y (nx37956), .A0 (nx37924), .A1 (nx37952), .S0 (nx23273)
             ) ;
    mux21_ni ix37925 (.Y (nx37924), .A0 (nx37908), .A1 (nx37920), .S0 (nx23659)
             ) ;
    mux21_ni ix37909 (.Y (nx37908), .A0 (inputs_344__9), .A1 (inputs_345__9), .S0 (
             nx24429)) ;
    mux21_ni ix37921 (.Y (nx37920), .A0 (inputs_346__9), .A1 (inputs_347__9), .S0 (
             nx24429)) ;
    mux21_ni ix37953 (.Y (nx37952), .A0 (nx37936), .A1 (nx37948), .S0 (nx23659)
             ) ;
    mux21_ni ix37937 (.Y (nx37936), .A0 (inputs_348__9), .A1 (inputs_349__9), .S0 (
             nx24431)) ;
    mux21_ni ix37949 (.Y (nx37948), .A0 (inputs_350__9), .A1 (inputs_351__9), .S0 (
             nx24431)) ;
    mux21_ni ix38253 (.Y (nx38252), .A0 (nx38246), .A1 (nx38168), .S0 (nx23159)
             ) ;
    oai21 ix38247 (.Y (nx38246), .A0 (nx22313), .A1 (nx16259), .B0 (nx16271)) ;
    mux21 ix16260 (.Y (nx16259), .A0 (nx38210), .A1 (nx38238), .S0 (nx22925)) ;
    mux21_ni ix38211 (.Y (nx38210), .A0 (nx38194), .A1 (nx38206), .S0 (nx23659)
             ) ;
    mux21_ni ix38195 (.Y (nx38194), .A0 (inputs_356__9), .A1 (inputs_357__9), .S0 (
             nx24431)) ;
    mux21_ni ix38207 (.Y (nx38206), .A0 (inputs_358__9), .A1 (inputs_359__9), .S0 (
             nx24431)) ;
    mux21_ni ix38239 (.Y (nx38238), .A0 (nx38222), .A1 (nx38234), .S0 (nx23659)
             ) ;
    mux21_ni ix38223 (.Y (nx38222), .A0 (inputs_372__9), .A1 (inputs_373__9), .S0 (
             nx24431)) ;
    mux21_ni ix38235 (.Y (nx38234), .A0 (inputs_374__9), .A1 (inputs_375__9), .S0 (
             nx24431)) ;
    nand04 ix16272 (.Y (nx16271), .A0 (nx22313), .A1 (nx23659), .A2 (nx24431), .A3 (
           nx38182)) ;
    mux21_ni ix38183 (.Y (nx38182), .A0 (inputs_355__9), .A1 (inputs_371__9), .S0 (
             nx22925)) ;
    mux21_ni ix38169 (.Y (nx38168), .A0 (nx38104), .A1 (nx38164), .S0 (nx22927)
             ) ;
    mux21_ni ix38105 (.Y (nx38104), .A0 (nx38072), .A1 (nx38100), .S0 (nx23275)
             ) ;
    mux21_ni ix38073 (.Y (nx38072), .A0 (nx38056), .A1 (nx38068), .S0 (nx23661)
             ) ;
    mux21_ni ix38057 (.Y (nx38056), .A0 (inputs_360__9), .A1 (inputs_361__9), .S0 (
             nx24433)) ;
    mux21_ni ix38069 (.Y (nx38068), .A0 (inputs_362__9), .A1 (inputs_363__9), .S0 (
             nx24433)) ;
    mux21_ni ix38101 (.Y (nx38100), .A0 (nx38084), .A1 (nx38096), .S0 (nx23661)
             ) ;
    mux21_ni ix38085 (.Y (nx38084), .A0 (inputs_364__9), .A1 (inputs_365__9), .S0 (
             nx24433)) ;
    mux21_ni ix38097 (.Y (nx38096), .A0 (inputs_366__9), .A1 (inputs_367__9), .S0 (
             nx24433)) ;
    mux21_ni ix38165 (.Y (nx38164), .A0 (nx38132), .A1 (nx38160), .S0 (nx23275)
             ) ;
    mux21_ni ix38133 (.Y (nx38132), .A0 (nx38116), .A1 (nx38128), .S0 (nx23661)
             ) ;
    mux21_ni ix38117 (.Y (nx38116), .A0 (inputs_376__9), .A1 (inputs_377__9), .S0 (
             nx24433)) ;
    mux21_ni ix38129 (.Y (nx38128), .A0 (inputs_378__9), .A1 (inputs_379__9), .S0 (
             nx24433)) ;
    mux21_ni ix38161 (.Y (nx38160), .A0 (nx38144), .A1 (nx38156), .S0 (nx23661)
             ) ;
    mux21_ni ix38145 (.Y (nx38144), .A0 (inputs_380__9), .A1 (inputs_381__9), .S0 (
             nx24433)) ;
    mux21_ni ix38157 (.Y (nx38156), .A0 (inputs_382__9), .A1 (inputs_383__9), .S0 (
             nx24435)) ;
    mux21_ni ix39105 (.Y (nx39104), .A0 (nx38680), .A1 (nx39100), .S0 (nx22491)
             ) ;
    mux21_ni ix38681 (.Y (nx38680), .A0 (nx38468), .A1 (nx38676), .S0 (nx22609)
             ) ;
    mux21_ni ix38469 (.Y (nx38468), .A0 (nx38462), .A1 (nx38384), .S0 (nx23159)
             ) ;
    oai21 ix38463 (.Y (nx38462), .A0 (nx22313), .A1 (nx16303), .B0 (nx16317)) ;
    mux21 ix16304 (.Y (nx16303), .A0 (nx38426), .A1 (nx38454), .S0 (nx22927)) ;
    mux21_ni ix38427 (.Y (nx38426), .A0 (nx38410), .A1 (nx38422), .S0 (nx23661)
             ) ;
    mux21_ni ix38411 (.Y (nx38410), .A0 (inputs_388__9), .A1 (inputs_389__9), .S0 (
             nx24435)) ;
    mux21_ni ix38423 (.Y (nx38422), .A0 (inputs_390__9), .A1 (inputs_391__9), .S0 (
             nx24435)) ;
    mux21_ni ix38455 (.Y (nx38454), .A0 (nx38438), .A1 (nx38450), .S0 (nx23661)
             ) ;
    mux21_ni ix38439 (.Y (nx38438), .A0 (inputs_404__9), .A1 (inputs_405__9), .S0 (
             nx24435)) ;
    mux21_ni ix38451 (.Y (nx38450), .A0 (inputs_406__9), .A1 (inputs_407__9), .S0 (
             nx24435)) ;
    nand04 ix16318 (.Y (nx16317), .A0 (nx22313), .A1 (nx23661), .A2 (nx24435), .A3 (
           nx38398)) ;
    mux21_ni ix38399 (.Y (nx38398), .A0 (inputs_387__9), .A1 (inputs_403__9), .S0 (
             nx22927)) ;
    mux21_ni ix38385 (.Y (nx38384), .A0 (nx38320), .A1 (nx38380), .S0 (nx22927)
             ) ;
    mux21_ni ix38321 (.Y (nx38320), .A0 (nx38288), .A1 (nx38316), .S0 (nx23275)
             ) ;
    mux21_ni ix38289 (.Y (nx38288), .A0 (nx38272), .A1 (nx38284), .S0 (nx23663)
             ) ;
    mux21_ni ix38273 (.Y (nx38272), .A0 (inputs_392__9), .A1 (inputs_393__9), .S0 (
             nx24435)) ;
    mux21_ni ix38285 (.Y (nx38284), .A0 (inputs_394__9), .A1 (inputs_395__9), .S0 (
             nx24437)) ;
    mux21_ni ix38317 (.Y (nx38316), .A0 (nx38300), .A1 (nx38312), .S0 (nx23663)
             ) ;
    mux21_ni ix38301 (.Y (nx38300), .A0 (inputs_396__9), .A1 (inputs_397__9), .S0 (
             nx24437)) ;
    mux21_ni ix38313 (.Y (nx38312), .A0 (inputs_398__9), .A1 (inputs_399__9), .S0 (
             nx24437)) ;
    mux21_ni ix38381 (.Y (nx38380), .A0 (nx38348), .A1 (nx38376), .S0 (nx23275)
             ) ;
    mux21_ni ix38349 (.Y (nx38348), .A0 (nx38332), .A1 (nx38344), .S0 (nx23663)
             ) ;
    mux21_ni ix38333 (.Y (nx38332), .A0 (inputs_408__9), .A1 (inputs_409__9), .S0 (
             nx24437)) ;
    mux21_ni ix38345 (.Y (nx38344), .A0 (inputs_410__9), .A1 (inputs_411__9), .S0 (
             nx24437)) ;
    mux21_ni ix38377 (.Y (nx38376), .A0 (nx38360), .A1 (nx38372), .S0 (nx23663)
             ) ;
    mux21_ni ix38361 (.Y (nx38360), .A0 (inputs_412__9), .A1 (inputs_413__9), .S0 (
             nx24437)) ;
    mux21_ni ix38373 (.Y (nx38372), .A0 (inputs_414__9), .A1 (inputs_415__9), .S0 (
             nx24437)) ;
    mux21_ni ix38677 (.Y (nx38676), .A0 (nx38670), .A1 (nx38592), .S0 (nx23159)
             ) ;
    oai21 ix38671 (.Y (nx38670), .A0 (nx22313), .A1 (nx16349), .B0 (nx16361)) ;
    mux21 ix16350 (.Y (nx16349), .A0 (nx38634), .A1 (nx38662), .S0 (nx22927)) ;
    mux21_ni ix38635 (.Y (nx38634), .A0 (nx38618), .A1 (nx38630), .S0 (nx23663)
             ) ;
    mux21_ni ix38619 (.Y (nx38618), .A0 (inputs_420__9), .A1 (inputs_421__9), .S0 (
             nx24439)) ;
    mux21_ni ix38631 (.Y (nx38630), .A0 (inputs_422__9), .A1 (inputs_423__9), .S0 (
             nx24439)) ;
    mux21_ni ix38663 (.Y (nx38662), .A0 (nx38646), .A1 (nx38658), .S0 (nx23663)
             ) ;
    mux21_ni ix38647 (.Y (nx38646), .A0 (inputs_436__9), .A1 (inputs_437__9), .S0 (
             nx24439)) ;
    mux21_ni ix38659 (.Y (nx38658), .A0 (inputs_438__9), .A1 (inputs_439__9), .S0 (
             nx24439)) ;
    nand04 ix16362 (.Y (nx16361), .A0 (nx22315), .A1 (nx23663), .A2 (nx24439), .A3 (
           nx38606)) ;
    mux21_ni ix38607 (.Y (nx38606), .A0 (inputs_419__9), .A1 (inputs_435__9), .S0 (
             nx22927)) ;
    mux21_ni ix38593 (.Y (nx38592), .A0 (nx38528), .A1 (nx38588), .S0 (nx22927)
             ) ;
    mux21_ni ix38529 (.Y (nx38528), .A0 (nx38496), .A1 (nx38524), .S0 (nx23275)
             ) ;
    mux21_ni ix38497 (.Y (nx38496), .A0 (nx38480), .A1 (nx38492), .S0 (nx23665)
             ) ;
    mux21_ni ix38481 (.Y (nx38480), .A0 (inputs_424__9), .A1 (inputs_425__9), .S0 (
             nx24439)) ;
    mux21_ni ix38493 (.Y (nx38492), .A0 (inputs_426__9), .A1 (inputs_427__9), .S0 (
             nx24439)) ;
    mux21_ni ix38525 (.Y (nx38524), .A0 (nx38508), .A1 (nx38520), .S0 (nx23665)
             ) ;
    mux21_ni ix38509 (.Y (nx38508), .A0 (inputs_428__9), .A1 (inputs_429__9), .S0 (
             nx24441)) ;
    mux21_ni ix38521 (.Y (nx38520), .A0 (inputs_430__9), .A1 (inputs_431__9), .S0 (
             nx24441)) ;
    mux21_ni ix38589 (.Y (nx38588), .A0 (nx38556), .A1 (nx38584), .S0 (nx23275)
             ) ;
    mux21_ni ix38557 (.Y (nx38556), .A0 (nx38540), .A1 (nx38552), .S0 (nx23665)
             ) ;
    mux21_ni ix38541 (.Y (nx38540), .A0 (inputs_440__9), .A1 (inputs_441__9), .S0 (
             nx24441)) ;
    mux21_ni ix38553 (.Y (nx38552), .A0 (inputs_442__9), .A1 (inputs_443__9), .S0 (
             nx24441)) ;
    mux21_ni ix38585 (.Y (nx38584), .A0 (nx38568), .A1 (nx38580), .S0 (nx23665)
             ) ;
    mux21_ni ix38569 (.Y (nx38568), .A0 (inputs_444__9), .A1 (inputs_445__9), .S0 (
             nx24441)) ;
    mux21_ni ix38581 (.Y (nx38580), .A0 (inputs_446__9), .A1 (inputs_447__9), .S0 (
             nx24441)) ;
    mux21_ni ix39101 (.Y (nx39100), .A0 (nx38888), .A1 (nx39096), .S0 (nx22609)
             ) ;
    mux21_ni ix38889 (.Y (nx38888), .A0 (nx38882), .A1 (nx38804), .S0 (nx23159)
             ) ;
    oai21 ix38883 (.Y (nx38882), .A0 (nx22315), .A1 (nx16393), .B0 (nx16405)) ;
    mux21 ix16394 (.Y (nx16393), .A0 (nx38846), .A1 (nx38874), .S0 (nx22929)) ;
    mux21_ni ix38847 (.Y (nx38846), .A0 (nx38830), .A1 (nx38842), .S0 (nx23665)
             ) ;
    mux21_ni ix38831 (.Y (nx38830), .A0 (inputs_452__9), .A1 (inputs_453__9), .S0 (
             nx24441)) ;
    mux21_ni ix38843 (.Y (nx38842), .A0 (inputs_454__9), .A1 (inputs_455__9), .S0 (
             nx24443)) ;
    mux21_ni ix38875 (.Y (nx38874), .A0 (nx38858), .A1 (nx38870), .S0 (nx23665)
             ) ;
    mux21_ni ix38859 (.Y (nx38858), .A0 (inputs_468__9), .A1 (inputs_469__9), .S0 (
             nx24443)) ;
    mux21_ni ix38871 (.Y (nx38870), .A0 (inputs_470__9), .A1 (inputs_471__9), .S0 (
             nx24443)) ;
    nand04 ix16406 (.Y (nx16405), .A0 (nx22315), .A1 (nx23665), .A2 (nx24443), .A3 (
           nx38818)) ;
    mux21_ni ix38819 (.Y (nx38818), .A0 (inputs_451__9), .A1 (inputs_467__9), .S0 (
             nx22929)) ;
    mux21_ni ix38805 (.Y (nx38804), .A0 (nx38740), .A1 (nx38800), .S0 (nx22929)
             ) ;
    mux21_ni ix38741 (.Y (nx38740), .A0 (nx38708), .A1 (nx38736), .S0 (nx23275)
             ) ;
    mux21_ni ix38709 (.Y (nx38708), .A0 (nx38692), .A1 (nx38704), .S0 (nx23667)
             ) ;
    mux21_ni ix38693 (.Y (nx38692), .A0 (inputs_456__9), .A1 (inputs_457__9), .S0 (
             nx24443)) ;
    mux21_ni ix38705 (.Y (nx38704), .A0 (inputs_458__9), .A1 (inputs_459__9), .S0 (
             nx24443)) ;
    mux21_ni ix38737 (.Y (nx38736), .A0 (nx38720), .A1 (nx38732), .S0 (nx23667)
             ) ;
    mux21_ni ix38721 (.Y (nx38720), .A0 (inputs_460__9), .A1 (inputs_461__9), .S0 (
             nx24443)) ;
    mux21_ni ix38733 (.Y (nx38732), .A0 (inputs_462__9), .A1 (inputs_463__9), .S0 (
             nx24445)) ;
    mux21_ni ix38801 (.Y (nx38800), .A0 (nx38768), .A1 (nx38796), .S0 (nx23277)
             ) ;
    mux21_ni ix38769 (.Y (nx38768), .A0 (nx38752), .A1 (nx38764), .S0 (nx23667)
             ) ;
    mux21_ni ix38753 (.Y (nx38752), .A0 (inputs_472__9), .A1 (inputs_473__9), .S0 (
             nx24445)) ;
    mux21_ni ix38765 (.Y (nx38764), .A0 (inputs_474__9), .A1 (inputs_475__9), .S0 (
             nx24445)) ;
    mux21_ni ix38797 (.Y (nx38796), .A0 (nx38780), .A1 (nx38792), .S0 (nx23667)
             ) ;
    mux21_ni ix38781 (.Y (nx38780), .A0 (inputs_476__9), .A1 (inputs_477__9), .S0 (
             nx24445)) ;
    mux21_ni ix38793 (.Y (nx38792), .A0 (inputs_478__9), .A1 (inputs_479__9), .S0 (
             nx24445)) ;
    mux21_ni ix39097 (.Y (nx39096), .A0 (nx39090), .A1 (nx39012), .S0 (nx23159)
             ) ;
    oai21 ix39091 (.Y (nx39090), .A0 (nx22315), .A1 (nx16435), .B0 (nx16447)) ;
    mux21 ix16436 (.Y (nx16435), .A0 (nx39054), .A1 (nx39082), .S0 (nx22929)) ;
    mux21_ni ix39055 (.Y (nx39054), .A0 (nx39038), .A1 (nx39050), .S0 (nx23667)
             ) ;
    mux21_ni ix39039 (.Y (nx39038), .A0 (inputs_484__9), .A1 (inputs_485__9), .S0 (
             nx24445)) ;
    mux21_ni ix39051 (.Y (nx39050), .A0 (inputs_486__9), .A1 (inputs_487__9), .S0 (
             nx24445)) ;
    mux21_ni ix39083 (.Y (nx39082), .A0 (nx39066), .A1 (nx39078), .S0 (nx23667)
             ) ;
    mux21_ni ix39067 (.Y (nx39066), .A0 (inputs_500__9), .A1 (inputs_501__9), .S0 (
             nx24447)) ;
    mux21_ni ix39079 (.Y (nx39078), .A0 (inputs_502__9), .A1 (inputs_503__9), .S0 (
             nx24447)) ;
    nand04 ix16448 (.Y (nx16447), .A0 (nx22315), .A1 (nx23667), .A2 (nx24447), .A3 (
           nx39026)) ;
    mux21_ni ix39027 (.Y (nx39026), .A0 (inputs_483__9), .A1 (inputs_499__9), .S0 (
             nx22929)) ;
    mux21_ni ix39013 (.Y (nx39012), .A0 (nx38948), .A1 (nx39008), .S0 (nx22929)
             ) ;
    mux21_ni ix38949 (.Y (nx38948), .A0 (nx38916), .A1 (nx38944), .S0 (nx23277)
             ) ;
    mux21_ni ix38917 (.Y (nx38916), .A0 (nx38900), .A1 (nx38912), .S0 (nx23669)
             ) ;
    mux21_ni ix38901 (.Y (nx38900), .A0 (inputs_488__9), .A1 (inputs_489__9), .S0 (
             nx24447)) ;
    mux21_ni ix38913 (.Y (nx38912), .A0 (inputs_490__9), .A1 (inputs_491__9), .S0 (
             nx24447)) ;
    mux21_ni ix38945 (.Y (nx38944), .A0 (nx38928), .A1 (nx38940), .S0 (nx23669)
             ) ;
    mux21_ni ix38929 (.Y (nx38928), .A0 (inputs_492__9), .A1 (inputs_493__9), .S0 (
             nx24447)) ;
    mux21_ni ix38941 (.Y (nx38940), .A0 (inputs_494__9), .A1 (inputs_495__9), .S0 (
             nx24447)) ;
    mux21_ni ix39009 (.Y (nx39008), .A0 (nx38976), .A1 (nx39004), .S0 (nx23277)
             ) ;
    mux21_ni ix38977 (.Y (nx38976), .A0 (nx38960), .A1 (nx38972), .S0 (nx23669)
             ) ;
    mux21_ni ix38961 (.Y (nx38960), .A0 (inputs_504__9), .A1 (inputs_505__9), .S0 (
             nx24449)) ;
    mux21_ni ix38973 (.Y (nx38972), .A0 (inputs_506__9), .A1 (inputs_507__9), .S0 (
             nx24449)) ;
    mux21_ni ix39005 (.Y (nx39004), .A0 (nx38988), .A1 (nx39000), .S0 (nx23669)
             ) ;
    mux21_ni ix38989 (.Y (nx38988), .A0 (inputs_508__9), .A1 (inputs_509__9), .S0 (
             nx24449)) ;
    mux21_ni ix39001 (.Y (nx39000), .A0 (inputs_510__9), .A1 (inputs_511__9), .S0 (
             nx24449)) ;
    aoi32 ix16476 (.Y (nx16475), .A0 (nx39874), .A1 (nx22387), .A2 (nx22315), .B0 (
          nx22221), .B1 (nx41570)) ;
    oai21 ix39875 (.Y (nx39874), .A0 (nx23669), .A1 (nx16479), .B0 (nx16581)) ;
    mux21 ix16480 (.Y (nx16479), .A0 (nx39612), .A1 (nx39864), .S0 (nx24449)) ;
    mux21_ni ix39613 (.Y (nx39612), .A0 (nx39484), .A1 (nx39608), .S0 (nx22399)
             ) ;
    mux21_ni ix39485 (.Y (nx39484), .A0 (nx39420), .A1 (nx39480), .S0 (nx22431)
             ) ;
    mux21_ni ix39421 (.Y (nx39420), .A0 (nx39388), .A1 (nx39416), .S0 (nx22491)
             ) ;
    mux21_ni ix39389 (.Y (nx39388), .A0 (nx39372), .A1 (nx39384), .S0 (nx22609)
             ) ;
    mux21_ni ix39373 (.Y (nx39372), .A0 (inputs_0__9), .A1 (inputs_16__9), .S0 (
             nx22929)) ;
    mux21_ni ix39385 (.Y (nx39384), .A0 (inputs_32__9), .A1 (inputs_48__9), .S0 (
             nx22931)) ;
    mux21_ni ix39417 (.Y (nx39416), .A0 (nx39400), .A1 (nx39412), .S0 (nx22609)
             ) ;
    mux21_ni ix39401 (.Y (nx39400), .A0 (inputs_64__9), .A1 (inputs_80__9), .S0 (
             nx22931)) ;
    mux21_ni ix39413 (.Y (nx39412), .A0 (inputs_96__9), .A1 (inputs_112__9), .S0 (
             nx22931)) ;
    mux21_ni ix39481 (.Y (nx39480), .A0 (nx39448), .A1 (nx39476), .S0 (nx22493)
             ) ;
    mux21_ni ix39449 (.Y (nx39448), .A0 (nx39432), .A1 (nx39444), .S0 (nx22611)
             ) ;
    mux21_ni ix39433 (.Y (nx39432), .A0 (inputs_128__9), .A1 (inputs_144__9), .S0 (
             nx22931)) ;
    mux21_ni ix39445 (.Y (nx39444), .A0 (inputs_160__9), .A1 (inputs_176__9), .S0 (
             nx22931)) ;
    mux21_ni ix39477 (.Y (nx39476), .A0 (nx39460), .A1 (nx39472), .S0 (nx22611)
             ) ;
    mux21_ni ix39461 (.Y (nx39460), .A0 (inputs_192__9), .A1 (inputs_208__9), .S0 (
             nx22931)) ;
    mux21_ni ix39473 (.Y (nx39472), .A0 (inputs_224__9), .A1 (inputs_240__9), .S0 (
             nx22931)) ;
    mux21_ni ix39609 (.Y (nx39608), .A0 (nx39544), .A1 (nx39604), .S0 (nx22431)
             ) ;
    mux21_ni ix39545 (.Y (nx39544), .A0 (nx39512), .A1 (nx39540), .S0 (nx22493)
             ) ;
    mux21_ni ix39513 (.Y (nx39512), .A0 (nx39496), .A1 (nx39508), .S0 (nx22611)
             ) ;
    mux21_ni ix39497 (.Y (nx39496), .A0 (inputs_256__9), .A1 (inputs_272__9), .S0 (
             nx22933)) ;
    mux21_ni ix39509 (.Y (nx39508), .A0 (inputs_288__9), .A1 (inputs_304__9), .S0 (
             nx22933)) ;
    mux21_ni ix39541 (.Y (nx39540), .A0 (nx39524), .A1 (nx39536), .S0 (nx22611)
             ) ;
    mux21_ni ix39525 (.Y (nx39524), .A0 (inputs_320__9), .A1 (inputs_336__9), .S0 (
             nx22933)) ;
    mux21_ni ix39537 (.Y (nx39536), .A0 (inputs_352__9), .A1 (inputs_368__9), .S0 (
             nx22933)) ;
    mux21_ni ix39605 (.Y (nx39604), .A0 (nx39572), .A1 (nx39600), .S0 (nx22493)
             ) ;
    mux21_ni ix39573 (.Y (nx39572), .A0 (nx39556), .A1 (nx39568), .S0 (nx22611)
             ) ;
    mux21_ni ix39557 (.Y (nx39556), .A0 (inputs_384__9), .A1 (inputs_400__9), .S0 (
             nx22933)) ;
    mux21_ni ix39569 (.Y (nx39568), .A0 (inputs_416__9), .A1 (inputs_432__9), .S0 (
             nx22933)) ;
    mux21_ni ix39601 (.Y (nx39600), .A0 (nx39584), .A1 (nx39596), .S0 (nx22611)
             ) ;
    mux21_ni ix39585 (.Y (nx39584), .A0 (inputs_448__9), .A1 (inputs_464__9), .S0 (
             nx22933)) ;
    mux21_ni ix39597 (.Y (nx39596), .A0 (inputs_480__9), .A1 (inputs_496__9), .S0 (
             nx22935)) ;
    mux21_ni ix39865 (.Y (nx39864), .A0 (nx39736), .A1 (nx39860), .S0 (nx22401)
             ) ;
    mux21_ni ix39737 (.Y (nx39736), .A0 (nx39672), .A1 (nx39732), .S0 (nx22431)
             ) ;
    mux21_ni ix39673 (.Y (nx39672), .A0 (nx39640), .A1 (nx39668), .S0 (nx22493)
             ) ;
    mux21_ni ix39641 (.Y (nx39640), .A0 (nx39624), .A1 (nx39636), .S0 (nx22611)
             ) ;
    mux21_ni ix39625 (.Y (nx39624), .A0 (inputs_1__9), .A1 (inputs_17__9), .S0 (
             nx22935)) ;
    mux21_ni ix39637 (.Y (nx39636), .A0 (inputs_33__9), .A1 (inputs_49__9), .S0 (
             nx22935)) ;
    mux21_ni ix39669 (.Y (nx39668), .A0 (nx39652), .A1 (nx39664), .S0 (nx22613)
             ) ;
    mux21_ni ix39653 (.Y (nx39652), .A0 (inputs_65__9), .A1 (inputs_81__9), .S0 (
             nx22935)) ;
    mux21_ni ix39665 (.Y (nx39664), .A0 (inputs_97__9), .A1 (inputs_113__9), .S0 (
             nx22935)) ;
    mux21_ni ix39733 (.Y (nx39732), .A0 (nx39700), .A1 (nx39728), .S0 (nx22493)
             ) ;
    mux21_ni ix39701 (.Y (nx39700), .A0 (nx39684), .A1 (nx39696), .S0 (nx22613)
             ) ;
    mux21_ni ix39685 (.Y (nx39684), .A0 (inputs_129__9), .A1 (inputs_145__9), .S0 (
             nx22935)) ;
    mux21_ni ix39697 (.Y (nx39696), .A0 (inputs_161__9), .A1 (inputs_177__9), .S0 (
             nx22935)) ;
    mux21_ni ix39729 (.Y (nx39728), .A0 (nx39712), .A1 (nx39724), .S0 (nx22613)
             ) ;
    mux21_ni ix39713 (.Y (nx39712), .A0 (inputs_193__9), .A1 (inputs_209__9), .S0 (
             nx22937)) ;
    mux21_ni ix39725 (.Y (nx39724), .A0 (inputs_225__9), .A1 (inputs_241__9), .S0 (
             nx22937)) ;
    mux21_ni ix39861 (.Y (nx39860), .A0 (nx39796), .A1 (nx39856), .S0 (nx22431)
             ) ;
    mux21_ni ix39797 (.Y (nx39796), .A0 (nx39764), .A1 (nx39792), .S0 (nx22493)
             ) ;
    mux21_ni ix39765 (.Y (nx39764), .A0 (nx39748), .A1 (nx39760), .S0 (nx22613)
             ) ;
    mux21_ni ix39749 (.Y (nx39748), .A0 (inputs_257__9), .A1 (inputs_273__9), .S0 (
             nx22937)) ;
    mux21_ni ix39761 (.Y (nx39760), .A0 (inputs_289__9), .A1 (inputs_305__9), .S0 (
             nx22937)) ;
    mux21_ni ix39793 (.Y (nx39792), .A0 (nx39776), .A1 (nx39788), .S0 (nx22613)
             ) ;
    mux21_ni ix39777 (.Y (nx39776), .A0 (inputs_321__9), .A1 (inputs_337__9), .S0 (
             nx22937)) ;
    mux21_ni ix39789 (.Y (nx39788), .A0 (inputs_353__9), .A1 (inputs_369__9), .S0 (
             nx22937)) ;
    mux21_ni ix39857 (.Y (nx39856), .A0 (nx39824), .A1 (nx39852), .S0 (nx22493)
             ) ;
    mux21_ni ix39825 (.Y (nx39824), .A0 (nx39808), .A1 (nx39820), .S0 (nx22613)
             ) ;
    mux21_ni ix39809 (.Y (nx39808), .A0 (inputs_385__9), .A1 (inputs_401__9), .S0 (
             nx22937)) ;
    mux21_ni ix39821 (.Y (nx39820), .A0 (inputs_417__9), .A1 (inputs_433__9), .S0 (
             nx22939)) ;
    mux21_ni ix39853 (.Y (nx39852), .A0 (nx39836), .A1 (nx39848), .S0 (nx22613)
             ) ;
    mux21_ni ix39837 (.Y (nx39836), .A0 (inputs_449__9), .A1 (inputs_465__9), .S0 (
             nx22939)) ;
    mux21_ni ix39849 (.Y (nx39848), .A0 (inputs_481__9), .A1 (inputs_497__9), .S0 (
             nx22939)) ;
    nand03 ix16582 (.Y (nx16581), .A0 (nx39358), .A1 (nx23669), .A2 (nx22381)) ;
    mux21_ni ix39359 (.Y (nx39358), .A0 (nx39230), .A1 (nx39354), .S0 (nx22401)
             ) ;
    mux21_ni ix39231 (.Y (nx39230), .A0 (nx39166), .A1 (nx39226), .S0 (nx22433)
             ) ;
    mux21_ni ix39167 (.Y (nx39166), .A0 (nx39134), .A1 (nx39162), .S0 (nx22495)
             ) ;
    mux21_ni ix39135 (.Y (nx39134), .A0 (nx39118), .A1 (nx39130), .S0 (nx22615)
             ) ;
    mux21_ni ix39119 (.Y (nx39118), .A0 (inputs_2__9), .A1 (inputs_18__9), .S0 (
             nx22939)) ;
    mux21_ni ix39131 (.Y (nx39130), .A0 (inputs_34__9), .A1 (inputs_50__9), .S0 (
             nx22939)) ;
    mux21_ni ix39163 (.Y (nx39162), .A0 (nx39146), .A1 (nx39158), .S0 (nx22615)
             ) ;
    mux21_ni ix39147 (.Y (nx39146), .A0 (inputs_66__9), .A1 (inputs_82__9), .S0 (
             nx22939)) ;
    mux21_ni ix39159 (.Y (nx39158), .A0 (inputs_98__9), .A1 (inputs_114__9), .S0 (
             nx22939)) ;
    mux21_ni ix39227 (.Y (nx39226), .A0 (nx39194), .A1 (nx39222), .S0 (nx22495)
             ) ;
    mux21_ni ix39195 (.Y (nx39194), .A0 (nx39178), .A1 (nx39190), .S0 (nx22615)
             ) ;
    mux21_ni ix39179 (.Y (nx39178), .A0 (inputs_130__9), .A1 (inputs_146__9), .S0 (
             nx22941)) ;
    mux21_ni ix39191 (.Y (nx39190), .A0 (inputs_162__9), .A1 (inputs_178__9), .S0 (
             nx22941)) ;
    mux21_ni ix39223 (.Y (nx39222), .A0 (nx39206), .A1 (nx39218), .S0 (nx22615)
             ) ;
    mux21_ni ix39207 (.Y (nx39206), .A0 (inputs_194__9), .A1 (inputs_210__9), .S0 (
             nx22941)) ;
    mux21_ni ix39219 (.Y (nx39218), .A0 (inputs_226__9), .A1 (inputs_242__9), .S0 (
             nx22941)) ;
    mux21_ni ix39355 (.Y (nx39354), .A0 (nx39290), .A1 (nx39350), .S0 (nx22433)
             ) ;
    mux21_ni ix39291 (.Y (nx39290), .A0 (nx39258), .A1 (nx39286), .S0 (nx22495)
             ) ;
    mux21_ni ix39259 (.Y (nx39258), .A0 (nx39242), .A1 (nx39254), .S0 (nx22615)
             ) ;
    mux21_ni ix39243 (.Y (nx39242), .A0 (inputs_258__9), .A1 (inputs_274__9), .S0 (
             nx22941)) ;
    mux21_ni ix39255 (.Y (nx39254), .A0 (inputs_290__9), .A1 (inputs_306__9), .S0 (
             nx22941)) ;
    mux21_ni ix39287 (.Y (nx39286), .A0 (nx39270), .A1 (nx39282), .S0 (nx22615)
             ) ;
    mux21_ni ix39271 (.Y (nx39270), .A0 (inputs_322__9), .A1 (inputs_338__9), .S0 (
             nx22941)) ;
    mux21_ni ix39283 (.Y (nx39282), .A0 (inputs_354__9), .A1 (inputs_370__9), .S0 (
             nx22943)) ;
    mux21_ni ix39351 (.Y (nx39350), .A0 (nx39318), .A1 (nx39346), .S0 (nx22495)
             ) ;
    mux21_ni ix39319 (.Y (nx39318), .A0 (nx39302), .A1 (nx39314), .S0 (nx22615)
             ) ;
    mux21_ni ix39303 (.Y (nx39302), .A0 (inputs_386__9), .A1 (inputs_402__9), .S0 (
             nx22943)) ;
    mux21_ni ix39315 (.Y (nx39314), .A0 (inputs_418__9), .A1 (inputs_434__9), .S0 (
             nx22943)) ;
    mux21_ni ix39347 (.Y (nx39346), .A0 (nx39330), .A1 (nx39342), .S0 (nx22617)
             ) ;
    mux21_ni ix39331 (.Y (nx39330), .A0 (inputs_450__9), .A1 (inputs_466__9), .S0 (
             nx22943)) ;
    mux21_ni ix39343 (.Y (nx39342), .A0 (inputs_482__9), .A1 (inputs_498__9), .S0 (
             nx22943)) ;
    mux21_ni ix41571 (.Y (nx41570), .A0 (nx40722), .A1 (nx41566), .S0 (nx22433)
             ) ;
    mux21_ni ix40723 (.Y (nx40722), .A0 (nx40298), .A1 (nx40718), .S0 (nx22495)
             ) ;
    mux21_ni ix40299 (.Y (nx40298), .A0 (nx40086), .A1 (nx40294), .S0 (nx22617)
             ) ;
    mux21_ni ix40087 (.Y (nx40086), .A0 (nx40080), .A1 (nx40002), .S0 (nx23159)
             ) ;
    oai21 ix40081 (.Y (nx40080), .A0 (nx22315), .A1 (nx16643), .B0 (nx16655)) ;
    mux21 ix16644 (.Y (nx16643), .A0 (nx40044), .A1 (nx40072), .S0 (nx22943)) ;
    mux21_ni ix40045 (.Y (nx40044), .A0 (nx40028), .A1 (nx40040), .S0 (nx23669)
             ) ;
    mux21_ni ix40029 (.Y (nx40028), .A0 (inputs_4__9), .A1 (inputs_5__9), .S0 (
             nx24449)) ;
    mux21_ni ix40041 (.Y (nx40040), .A0 (inputs_6__9), .A1 (inputs_7__9), .S0 (
             nx24449)) ;
    mux21_ni ix40073 (.Y (nx40072), .A0 (nx40056), .A1 (nx40068), .S0 (nx23671)
             ) ;
    mux21_ni ix40057 (.Y (nx40056), .A0 (inputs_20__9), .A1 (inputs_21__9), .S0 (
             nx24451)) ;
    mux21_ni ix40069 (.Y (nx40068), .A0 (inputs_22__9), .A1 (inputs_23__9), .S0 (
             nx24451)) ;
    nand04 ix16656 (.Y (nx16655), .A0 (nx22317), .A1 (nx23671), .A2 (nx24451), .A3 (
           nx40016)) ;
    mux21_ni ix40017 (.Y (nx40016), .A0 (inputs_3__9), .A1 (inputs_19__9), .S0 (
             nx22943)) ;
    mux21_ni ix40003 (.Y (nx40002), .A0 (nx39938), .A1 (nx39998), .S0 (nx22945)
             ) ;
    mux21_ni ix39939 (.Y (nx39938), .A0 (nx39906), .A1 (nx39934), .S0 (nx23277)
             ) ;
    mux21_ni ix39907 (.Y (nx39906), .A0 (nx39890), .A1 (nx39902), .S0 (nx23671)
             ) ;
    mux21_ni ix39891 (.Y (nx39890), .A0 (inputs_8__9), .A1 (inputs_9__9), .S0 (
             nx24451)) ;
    mux21_ni ix39903 (.Y (nx39902), .A0 (inputs_10__9), .A1 (inputs_11__9), .S0 (
             nx24451)) ;
    mux21_ni ix39935 (.Y (nx39934), .A0 (nx39918), .A1 (nx39930), .S0 (nx23671)
             ) ;
    mux21_ni ix39919 (.Y (nx39918), .A0 (inputs_12__9), .A1 (inputs_13__9), .S0 (
             nx24451)) ;
    mux21_ni ix39931 (.Y (nx39930), .A0 (inputs_14__9), .A1 (inputs_15__9), .S0 (
             nx24451)) ;
    mux21_ni ix39999 (.Y (nx39998), .A0 (nx39966), .A1 (nx39994), .S0 (nx23277)
             ) ;
    mux21_ni ix39967 (.Y (nx39966), .A0 (nx39950), .A1 (nx39962), .S0 (nx23671)
             ) ;
    mux21_ni ix39951 (.Y (nx39950), .A0 (inputs_24__9), .A1 (inputs_25__9), .S0 (
             nx24453)) ;
    mux21_ni ix39963 (.Y (nx39962), .A0 (inputs_26__9), .A1 (inputs_27__9), .S0 (
             nx24453)) ;
    mux21_ni ix39995 (.Y (nx39994), .A0 (nx39978), .A1 (nx39990), .S0 (nx23671)
             ) ;
    mux21_ni ix39979 (.Y (nx39978), .A0 (inputs_28__9), .A1 (inputs_29__9), .S0 (
             nx24453)) ;
    mux21_ni ix39991 (.Y (nx39990), .A0 (inputs_30__9), .A1 (inputs_31__9), .S0 (
             nx24453)) ;
    mux21_ni ix40295 (.Y (nx40294), .A0 (nx40288), .A1 (nx40210), .S0 (nx23159)
             ) ;
    oai21 ix40289 (.Y (nx40288), .A0 (nx22317), .A1 (nx16685), .B0 (nx16695)) ;
    mux21 ix16686 (.Y (nx16685), .A0 (nx40252), .A1 (nx40280), .S0 (nx22945)) ;
    mux21_ni ix40253 (.Y (nx40252), .A0 (nx40236), .A1 (nx40248), .S0 (nx23671)
             ) ;
    mux21_ni ix40237 (.Y (nx40236), .A0 (inputs_36__9), .A1 (inputs_37__9), .S0 (
             nx24453)) ;
    mux21_ni ix40249 (.Y (nx40248), .A0 (inputs_38__9), .A1 (inputs_39__9), .S0 (
             nx24453)) ;
    mux21_ni ix40281 (.Y (nx40280), .A0 (nx40264), .A1 (nx40276), .S0 (nx23673)
             ) ;
    mux21_ni ix40265 (.Y (nx40264), .A0 (inputs_52__9), .A1 (inputs_53__9), .S0 (
             nx24453)) ;
    mux21_ni ix40277 (.Y (nx40276), .A0 (inputs_54__9), .A1 (inputs_55__9), .S0 (
             nx24455)) ;
    nand04 ix16696 (.Y (nx16695), .A0 (nx22317), .A1 (nx23673), .A2 (nx24455), .A3 (
           nx40224)) ;
    mux21_ni ix40225 (.Y (nx40224), .A0 (inputs_35__9), .A1 (inputs_51__9), .S0 (
             nx22945)) ;
    mux21_ni ix40211 (.Y (nx40210), .A0 (nx40146), .A1 (nx40206), .S0 (nx22945)
             ) ;
    mux21_ni ix40147 (.Y (nx40146), .A0 (nx40114), .A1 (nx40142), .S0 (nx23277)
             ) ;
    mux21_ni ix40115 (.Y (nx40114), .A0 (nx40098), .A1 (nx40110), .S0 (nx23673)
             ) ;
    mux21_ni ix40099 (.Y (nx40098), .A0 (inputs_40__9), .A1 (inputs_41__9), .S0 (
             nx24455)) ;
    mux21_ni ix40111 (.Y (nx40110), .A0 (inputs_42__9), .A1 (inputs_43__9), .S0 (
             nx24455)) ;
    mux21_ni ix40143 (.Y (nx40142), .A0 (nx40126), .A1 (nx40138), .S0 (nx23673)
             ) ;
    mux21_ni ix40127 (.Y (nx40126), .A0 (inputs_44__9), .A1 (inputs_45__9), .S0 (
             nx24455)) ;
    mux21_ni ix40139 (.Y (nx40138), .A0 (inputs_46__9), .A1 (inputs_47__9), .S0 (
             nx24455)) ;
    mux21_ni ix40207 (.Y (nx40206), .A0 (nx40174), .A1 (nx40202), .S0 (nx23277)
             ) ;
    mux21_ni ix40175 (.Y (nx40174), .A0 (nx40158), .A1 (nx40170), .S0 (nx23673)
             ) ;
    mux21_ni ix40159 (.Y (nx40158), .A0 (inputs_56__9), .A1 (inputs_57__9), .S0 (
             nx24455)) ;
    mux21_ni ix40171 (.Y (nx40170), .A0 (inputs_58__9), .A1 (inputs_59__9), .S0 (
             nx24457)) ;
    mux21_ni ix40203 (.Y (nx40202), .A0 (nx40186), .A1 (nx40198), .S0 (nx23673)
             ) ;
    mux21_ni ix40187 (.Y (nx40186), .A0 (inputs_60__9), .A1 (inputs_61__9), .S0 (
             nx24457)) ;
    mux21_ni ix40199 (.Y (nx40198), .A0 (inputs_62__9), .A1 (inputs_63__9), .S0 (
             nx24457)) ;
    mux21_ni ix40719 (.Y (nx40718), .A0 (nx40506), .A1 (nx40714), .S0 (nx22617)
             ) ;
    mux21_ni ix40507 (.Y (nx40506), .A0 (nx40500), .A1 (nx40422), .S0 (nx23161)
             ) ;
    oai21 ix40501 (.Y (nx40500), .A0 (nx22317), .A1 (nx16727), .B0 (nx16737)) ;
    mux21 ix16728 (.Y (nx16727), .A0 (nx40464), .A1 (nx40492), .S0 (nx22945)) ;
    mux21_ni ix40465 (.Y (nx40464), .A0 (nx40448), .A1 (nx40460), .S0 (nx23673)
             ) ;
    mux21_ni ix40449 (.Y (nx40448), .A0 (inputs_68__9), .A1 (inputs_69__9), .S0 (
             nx24457)) ;
    mux21_ni ix40461 (.Y (nx40460), .A0 (inputs_70__9), .A1 (inputs_71__9), .S0 (
             nx24457)) ;
    mux21_ni ix40493 (.Y (nx40492), .A0 (nx40476), .A1 (nx40488), .S0 (nx23675)
             ) ;
    mux21_ni ix40477 (.Y (nx40476), .A0 (inputs_84__9), .A1 (inputs_85__9), .S0 (
             nx24457)) ;
    mux21_ni ix40489 (.Y (nx40488), .A0 (inputs_86__9), .A1 (inputs_87__9), .S0 (
             nx24457)) ;
    nand04 ix16738 (.Y (nx16737), .A0 (nx22317), .A1 (nx23675), .A2 (nx24459), .A3 (
           nx40436)) ;
    mux21_ni ix40437 (.Y (nx40436), .A0 (inputs_67__9), .A1 (inputs_83__9), .S0 (
             nx22945)) ;
    mux21_ni ix40423 (.Y (nx40422), .A0 (nx40358), .A1 (nx40418), .S0 (nx22945)
             ) ;
    mux21_ni ix40359 (.Y (nx40358), .A0 (nx40326), .A1 (nx40354), .S0 (nx23279)
             ) ;
    mux21_ni ix40327 (.Y (nx40326), .A0 (nx40310), .A1 (nx40322), .S0 (nx23675)
             ) ;
    mux21_ni ix40311 (.Y (nx40310), .A0 (inputs_72__9), .A1 (inputs_73__9), .S0 (
             nx24459)) ;
    mux21_ni ix40323 (.Y (nx40322), .A0 (inputs_74__9), .A1 (inputs_75__9), .S0 (
             nx24459)) ;
    mux21_ni ix40355 (.Y (nx40354), .A0 (nx40338), .A1 (nx40350), .S0 (nx23675)
             ) ;
    mux21_ni ix40339 (.Y (nx40338), .A0 (inputs_76__9), .A1 (inputs_77__9), .S0 (
             nx24459)) ;
    mux21_ni ix40351 (.Y (nx40350), .A0 (inputs_78__9), .A1 (inputs_79__9), .S0 (
             nx24459)) ;
    mux21_ni ix40419 (.Y (nx40418), .A0 (nx40386), .A1 (nx40414), .S0 (nx23279)
             ) ;
    mux21_ni ix40387 (.Y (nx40386), .A0 (nx40370), .A1 (nx40382), .S0 (nx23675)
             ) ;
    mux21_ni ix40371 (.Y (nx40370), .A0 (inputs_88__9), .A1 (inputs_89__9), .S0 (
             nx24459)) ;
    mux21_ni ix40383 (.Y (nx40382), .A0 (inputs_90__9), .A1 (inputs_91__9), .S0 (
             nx24459)) ;
    mux21_ni ix40415 (.Y (nx40414), .A0 (nx40398), .A1 (nx40410), .S0 (nx23675)
             ) ;
    mux21_ni ix40399 (.Y (nx40398), .A0 (inputs_92__9), .A1 (inputs_93__9), .S0 (
             nx24461)) ;
    mux21_ni ix40411 (.Y (nx40410), .A0 (inputs_94__9), .A1 (inputs_95__9), .S0 (
             nx24461)) ;
    mux21_ni ix40715 (.Y (nx40714), .A0 (nx40708), .A1 (nx40630), .S0 (nx23161)
             ) ;
    oai21 ix40709 (.Y (nx40708), .A0 (nx22317), .A1 (nx16771), .B0 (nx16783)) ;
    mux21 ix16772 (.Y (nx16771), .A0 (nx40672), .A1 (nx40700), .S0 (nx22947)) ;
    mux21_ni ix40673 (.Y (nx40672), .A0 (nx40656), .A1 (nx40668), .S0 (nx23675)
             ) ;
    mux21_ni ix40657 (.Y (nx40656), .A0 (inputs_100__9), .A1 (inputs_101__9), .S0 (
             nx24461)) ;
    mux21_ni ix40669 (.Y (nx40668), .A0 (inputs_102__9), .A1 (inputs_103__9), .S0 (
             nx24461)) ;
    mux21_ni ix40701 (.Y (nx40700), .A0 (nx40684), .A1 (nx40696), .S0 (nx23677)
             ) ;
    mux21_ni ix40685 (.Y (nx40684), .A0 (inputs_116__9), .A1 (inputs_117__9), .S0 (
             nx24461)) ;
    mux21_ni ix40697 (.Y (nx40696), .A0 (inputs_118__9), .A1 (inputs_119__9), .S0 (
             nx24461)) ;
    nand04 ix16784 (.Y (nx16783), .A0 (nx22317), .A1 (nx23677), .A2 (nx24461), .A3 (
           nx40644)) ;
    mux21_ni ix40645 (.Y (nx40644), .A0 (inputs_99__9), .A1 (inputs_115__9), .S0 (
             nx22947)) ;
    mux21_ni ix40631 (.Y (nx40630), .A0 (nx40566), .A1 (nx40626), .S0 (nx22947)
             ) ;
    mux21_ni ix40567 (.Y (nx40566), .A0 (nx40534), .A1 (nx40562), .S0 (nx23279)
             ) ;
    mux21_ni ix40535 (.Y (nx40534), .A0 (nx40518), .A1 (nx40530), .S0 (nx23677)
             ) ;
    mux21_ni ix40519 (.Y (nx40518), .A0 (inputs_104__9), .A1 (inputs_105__9), .S0 (
             nx24463)) ;
    mux21_ni ix40531 (.Y (nx40530), .A0 (inputs_106__9), .A1 (inputs_107__9), .S0 (
             nx24463)) ;
    mux21_ni ix40563 (.Y (nx40562), .A0 (nx40546), .A1 (nx40558), .S0 (nx23677)
             ) ;
    mux21_ni ix40547 (.Y (nx40546), .A0 (inputs_108__9), .A1 (inputs_109__9), .S0 (
             nx24463)) ;
    mux21_ni ix40559 (.Y (nx40558), .A0 (inputs_110__9), .A1 (inputs_111__9), .S0 (
             nx24463)) ;
    mux21_ni ix40627 (.Y (nx40626), .A0 (nx40594), .A1 (nx40622), .S0 (nx23279)
             ) ;
    mux21_ni ix40595 (.Y (nx40594), .A0 (nx40578), .A1 (nx40590), .S0 (nx23677)
             ) ;
    mux21_ni ix40579 (.Y (nx40578), .A0 (inputs_120__9), .A1 (inputs_121__9), .S0 (
             nx24463)) ;
    mux21_ni ix40591 (.Y (nx40590), .A0 (inputs_122__9), .A1 (inputs_123__9), .S0 (
             nx24463)) ;
    mux21_ni ix40623 (.Y (nx40622), .A0 (nx40606), .A1 (nx40618), .S0 (nx23677)
             ) ;
    mux21_ni ix40607 (.Y (nx40606), .A0 (inputs_124__9), .A1 (inputs_125__9), .S0 (
             nx24463)) ;
    mux21_ni ix40619 (.Y (nx40618), .A0 (inputs_126__9), .A1 (inputs_127__9), .S0 (
             nx24465)) ;
    mux21_ni ix41567 (.Y (nx41566), .A0 (nx41142), .A1 (nx41562), .S0 (nx22495)
             ) ;
    mux21_ni ix41143 (.Y (nx41142), .A0 (nx40930), .A1 (nx41138), .S0 (nx22617)
             ) ;
    mux21_ni ix40931 (.Y (nx40930), .A0 (nx40924), .A1 (nx40846), .S0 (nx23161)
             ) ;
    oai21 ix40925 (.Y (nx40924), .A0 (nx22319), .A1 (nx16817), .B0 (nx16831)) ;
    mux21 ix16818 (.Y (nx16817), .A0 (nx40888), .A1 (nx40916), .S0 (nx22947)) ;
    mux21_ni ix40889 (.Y (nx40888), .A0 (nx40872), .A1 (nx40884), .S0 (nx23677)
             ) ;
    mux21_ni ix40873 (.Y (nx40872), .A0 (inputs_132__9), .A1 (inputs_133__9), .S0 (
             nx24465)) ;
    mux21_ni ix40885 (.Y (nx40884), .A0 (inputs_134__9), .A1 (inputs_135__9), .S0 (
             nx24465)) ;
    mux21_ni ix40917 (.Y (nx40916), .A0 (nx40900), .A1 (nx40912), .S0 (nx23679)
             ) ;
    mux21_ni ix40901 (.Y (nx40900), .A0 (inputs_148__9), .A1 (inputs_149__9), .S0 (
             nx24465)) ;
    mux21_ni ix40913 (.Y (nx40912), .A0 (inputs_150__9), .A1 (inputs_151__9), .S0 (
             nx24465)) ;
    nand04 ix16832 (.Y (nx16831), .A0 (nx22319), .A1 (nx23679), .A2 (nx24465), .A3 (
           nx40860)) ;
    mux21_ni ix40861 (.Y (nx40860), .A0 (inputs_131__9), .A1 (inputs_147__9), .S0 (
             nx22947)) ;
    mux21_ni ix40847 (.Y (nx40846), .A0 (nx40782), .A1 (nx40842), .S0 (nx22947)
             ) ;
    mux21_ni ix40783 (.Y (nx40782), .A0 (nx40750), .A1 (nx40778), .S0 (nx23279)
             ) ;
    mux21_ni ix40751 (.Y (nx40750), .A0 (nx40734), .A1 (nx40746), .S0 (nx23679)
             ) ;
    mux21_ni ix40735 (.Y (nx40734), .A0 (inputs_136__9), .A1 (inputs_137__9), .S0 (
             nx24465)) ;
    mux21_ni ix40747 (.Y (nx40746), .A0 (inputs_138__9), .A1 (inputs_139__9), .S0 (
             nx24467)) ;
    mux21_ni ix40779 (.Y (nx40778), .A0 (nx40762), .A1 (nx40774), .S0 (nx23679)
             ) ;
    mux21_ni ix40763 (.Y (nx40762), .A0 (inputs_140__9), .A1 (inputs_141__9), .S0 (
             nx24467)) ;
    mux21_ni ix40775 (.Y (nx40774), .A0 (inputs_142__9), .A1 (inputs_143__9), .S0 (
             nx24467)) ;
    mux21_ni ix40843 (.Y (nx40842), .A0 (nx40810), .A1 (nx40838), .S0 (nx23279)
             ) ;
    mux21_ni ix40811 (.Y (nx40810), .A0 (nx40794), .A1 (nx40806), .S0 (nx23679)
             ) ;
    mux21_ni ix40795 (.Y (nx40794), .A0 (inputs_152__9), .A1 (inputs_153__9), .S0 (
             nx24467)) ;
    mux21_ni ix40807 (.Y (nx40806), .A0 (inputs_154__9), .A1 (inputs_155__9), .S0 (
             nx24467)) ;
    mux21_ni ix40839 (.Y (nx40838), .A0 (nx40822), .A1 (nx40834), .S0 (nx23679)
             ) ;
    mux21_ni ix40823 (.Y (nx40822), .A0 (inputs_156__9), .A1 (inputs_157__9), .S0 (
             nx24467)) ;
    mux21_ni ix40835 (.Y (nx40834), .A0 (inputs_158__9), .A1 (inputs_159__9), .S0 (
             nx24467)) ;
    mux21_ni ix41139 (.Y (nx41138), .A0 (nx41132), .A1 (nx41054), .S0 (nx23161)
             ) ;
    oai21 ix41133 (.Y (nx41132), .A0 (nx22319), .A1 (nx16861), .B0 (nx16871)) ;
    mux21 ix16862 (.Y (nx16861), .A0 (nx41096), .A1 (nx41124), .S0 (nx22947)) ;
    mux21_ni ix41097 (.Y (nx41096), .A0 (nx41080), .A1 (nx41092), .S0 (nx23679)
             ) ;
    mux21_ni ix41081 (.Y (nx41080), .A0 (inputs_164__9), .A1 (inputs_165__9), .S0 (
             nx24469)) ;
    mux21_ni ix41093 (.Y (nx41092), .A0 (inputs_166__9), .A1 (inputs_167__9), .S0 (
             nx24469)) ;
    mux21_ni ix41125 (.Y (nx41124), .A0 (nx41108), .A1 (nx41120), .S0 (nx23681)
             ) ;
    mux21_ni ix41109 (.Y (nx41108), .A0 (inputs_180__9), .A1 (inputs_181__9), .S0 (
             nx24469)) ;
    mux21_ni ix41121 (.Y (nx41120), .A0 (inputs_182__9), .A1 (inputs_183__9), .S0 (
             nx24469)) ;
    nand04 ix16872 (.Y (nx16871), .A0 (nx22319), .A1 (nx23681), .A2 (nx24469), .A3 (
           nx41068)) ;
    mux21_ni ix41069 (.Y (nx41068), .A0 (inputs_163__9), .A1 (inputs_179__9), .S0 (
             nx22949)) ;
    mux21_ni ix41055 (.Y (nx41054), .A0 (nx40990), .A1 (nx41050), .S0 (nx22949)
             ) ;
    mux21_ni ix40991 (.Y (nx40990), .A0 (nx40958), .A1 (nx40986), .S0 (nx23279)
             ) ;
    mux21_ni ix40959 (.Y (nx40958), .A0 (nx40942), .A1 (nx40954), .S0 (nx23681)
             ) ;
    mux21_ni ix40943 (.Y (nx40942), .A0 (inputs_168__9), .A1 (inputs_169__9), .S0 (
             nx24469)) ;
    mux21_ni ix40955 (.Y (nx40954), .A0 (inputs_170__9), .A1 (inputs_171__9), .S0 (
             nx24469)) ;
    mux21_ni ix40987 (.Y (nx40986), .A0 (nx40970), .A1 (nx40982), .S0 (nx23681)
             ) ;
    mux21_ni ix40971 (.Y (nx40970), .A0 (inputs_172__9), .A1 (inputs_173__9), .S0 (
             nx24471)) ;
    mux21_ni ix40983 (.Y (nx40982), .A0 (inputs_174__9), .A1 (inputs_175__9), .S0 (
             nx24471)) ;
    mux21_ni ix41051 (.Y (nx41050), .A0 (nx41018), .A1 (nx41046), .S0 (nx23281)
             ) ;
    mux21_ni ix41019 (.Y (nx41018), .A0 (nx41002), .A1 (nx41014), .S0 (nx23681)
             ) ;
    mux21_ni ix41003 (.Y (nx41002), .A0 (inputs_184__9), .A1 (inputs_185__9), .S0 (
             nx24471)) ;
    mux21_ni ix41015 (.Y (nx41014), .A0 (inputs_186__9), .A1 (inputs_187__9), .S0 (
             nx24471)) ;
    mux21_ni ix41047 (.Y (nx41046), .A0 (nx41030), .A1 (nx41042), .S0 (nx23681)
             ) ;
    mux21_ni ix41031 (.Y (nx41030), .A0 (inputs_188__9), .A1 (inputs_189__9), .S0 (
             nx24471)) ;
    mux21_ni ix41043 (.Y (nx41042), .A0 (inputs_190__9), .A1 (inputs_191__9), .S0 (
             nx24471)) ;
    mux21_ni ix41563 (.Y (nx41562), .A0 (nx41350), .A1 (nx41558), .S0 (nx22617)
             ) ;
    mux21_ni ix41351 (.Y (nx41350), .A0 (nx41344), .A1 (nx41266), .S0 (nx23161)
             ) ;
    oai21 ix41345 (.Y (nx41344), .A0 (nx22319), .A1 (nx16903), .B0 (nx16915)) ;
    mux21 ix16904 (.Y (nx16903), .A0 (nx41308), .A1 (nx41336), .S0 (nx22949)) ;
    mux21_ni ix41309 (.Y (nx41308), .A0 (nx41292), .A1 (nx41304), .S0 (nx23681)
             ) ;
    mux21_ni ix41293 (.Y (nx41292), .A0 (inputs_196__9), .A1 (inputs_197__9), .S0 (
             nx24471)) ;
    mux21_ni ix41305 (.Y (nx41304), .A0 (inputs_198__9), .A1 (inputs_199__9), .S0 (
             nx24473)) ;
    mux21_ni ix41337 (.Y (nx41336), .A0 (nx41320), .A1 (nx41332), .S0 (nx23683)
             ) ;
    mux21_ni ix41321 (.Y (nx41320), .A0 (inputs_212__9), .A1 (inputs_213__9), .S0 (
             nx24473)) ;
    mux21_ni ix41333 (.Y (nx41332), .A0 (inputs_214__9), .A1 (inputs_215__9), .S0 (
             nx24473)) ;
    nand04 ix16916 (.Y (nx16915), .A0 (nx22319), .A1 (nx23683), .A2 (nx24473), .A3 (
           nx41280)) ;
    mux21_ni ix41281 (.Y (nx41280), .A0 (inputs_195__9), .A1 (inputs_211__9), .S0 (
             nx22949)) ;
    mux21_ni ix41267 (.Y (nx41266), .A0 (nx41202), .A1 (nx41262), .S0 (nx22949)
             ) ;
    mux21_ni ix41203 (.Y (nx41202), .A0 (nx41170), .A1 (nx41198), .S0 (nx23281)
             ) ;
    mux21_ni ix41171 (.Y (nx41170), .A0 (nx41154), .A1 (nx41166), .S0 (nx23683)
             ) ;
    mux21_ni ix41155 (.Y (nx41154), .A0 (inputs_200__9), .A1 (inputs_201__9), .S0 (
             nx24473)) ;
    mux21_ni ix41167 (.Y (nx41166), .A0 (inputs_202__9), .A1 (inputs_203__9), .S0 (
             nx24473)) ;
    mux21_ni ix41199 (.Y (nx41198), .A0 (nx41182), .A1 (nx41194), .S0 (nx23683)
             ) ;
    mux21_ni ix41183 (.Y (nx41182), .A0 (inputs_204__9), .A1 (inputs_205__9), .S0 (
             nx24473)) ;
    mux21_ni ix41195 (.Y (nx41194), .A0 (inputs_206__9), .A1 (inputs_207__9), .S0 (
             nx24475)) ;
    mux21_ni ix41263 (.Y (nx41262), .A0 (nx41230), .A1 (nx41258), .S0 (nx23281)
             ) ;
    mux21_ni ix41231 (.Y (nx41230), .A0 (nx41214), .A1 (nx41226), .S0 (nx23683)
             ) ;
    mux21_ni ix41215 (.Y (nx41214), .A0 (inputs_216__9), .A1 (inputs_217__9), .S0 (
             nx24475)) ;
    mux21_ni ix41227 (.Y (nx41226), .A0 (inputs_218__9), .A1 (inputs_219__9), .S0 (
             nx24475)) ;
    mux21_ni ix41259 (.Y (nx41258), .A0 (nx41242), .A1 (nx41254), .S0 (nx23683)
             ) ;
    mux21_ni ix41243 (.Y (nx41242), .A0 (inputs_220__9), .A1 (inputs_221__9), .S0 (
             nx24475)) ;
    mux21_ni ix41255 (.Y (nx41254), .A0 (inputs_222__9), .A1 (inputs_223__9), .S0 (
             nx24475)) ;
    mux21_ni ix41559 (.Y (nx41558), .A0 (nx41552), .A1 (nx41474), .S0 (nx23161)
             ) ;
    oai21 ix41553 (.Y (nx41552), .A0 (nx22319), .A1 (nx16945), .B0 (nx16959)) ;
    mux21 ix16946 (.Y (nx16945), .A0 (nx41516), .A1 (nx41544), .S0 (nx22949)) ;
    mux21_ni ix41517 (.Y (nx41516), .A0 (nx41500), .A1 (nx41512), .S0 (nx23683)
             ) ;
    mux21_ni ix41501 (.Y (nx41500), .A0 (inputs_228__9), .A1 (inputs_229__9), .S0 (
             nx24475)) ;
    mux21_ni ix41513 (.Y (nx41512), .A0 (inputs_230__9), .A1 (inputs_231__9), .S0 (
             nx24475)) ;
    mux21_ni ix41545 (.Y (nx41544), .A0 (nx41528), .A1 (nx41540), .S0 (nx23685)
             ) ;
    mux21_ni ix41529 (.Y (nx41528), .A0 (inputs_244__9), .A1 (inputs_245__9), .S0 (
             nx24477)) ;
    mux21_ni ix41541 (.Y (nx41540), .A0 (inputs_246__9), .A1 (inputs_247__9), .S0 (
             nx24477)) ;
    nand04 ix16960 (.Y (nx16959), .A0 (nx22321), .A1 (nx23685), .A2 (nx24477), .A3 (
           nx41488)) ;
    mux21_ni ix41489 (.Y (nx41488), .A0 (inputs_227__9), .A1 (inputs_243__9), .S0 (
             nx22949)) ;
    mux21_ni ix41475 (.Y (nx41474), .A0 (nx41410), .A1 (nx41470), .S0 (nx22951)
             ) ;
    mux21_ni ix41411 (.Y (nx41410), .A0 (nx41378), .A1 (nx41406), .S0 (nx23281)
             ) ;
    mux21_ni ix41379 (.Y (nx41378), .A0 (nx41362), .A1 (nx41374), .S0 (nx23685)
             ) ;
    mux21_ni ix41363 (.Y (nx41362), .A0 (inputs_232__9), .A1 (inputs_233__9), .S0 (
             nx24477)) ;
    mux21_ni ix41375 (.Y (nx41374), .A0 (inputs_234__9), .A1 (inputs_235__9), .S0 (
             nx24477)) ;
    mux21_ni ix41407 (.Y (nx41406), .A0 (nx41390), .A1 (nx41402), .S0 (nx23685)
             ) ;
    mux21_ni ix41391 (.Y (nx41390), .A0 (inputs_236__9), .A1 (inputs_237__9), .S0 (
             nx24477)) ;
    mux21_ni ix41403 (.Y (nx41402), .A0 (inputs_238__9), .A1 (inputs_239__9), .S0 (
             nx24477)) ;
    mux21_ni ix41471 (.Y (nx41470), .A0 (nx41438), .A1 (nx41466), .S0 (nx23281)
             ) ;
    mux21_ni ix41439 (.Y (nx41438), .A0 (nx41422), .A1 (nx41434), .S0 (nx23685)
             ) ;
    mux21_ni ix41423 (.Y (nx41422), .A0 (inputs_248__9), .A1 (inputs_249__9), .S0 (
             nx24479)) ;
    mux21_ni ix41435 (.Y (nx41434), .A0 (inputs_250__9), .A1 (inputs_251__9), .S0 (
             nx24479)) ;
    mux21_ni ix41467 (.Y (nx41466), .A0 (nx41450), .A1 (nx41462), .S0 (nx23685)
             ) ;
    mux21_ni ix41451 (.Y (nx41450), .A0 (inputs_252__9), .A1 (inputs_253__9), .S0 (
             nx24479)) ;
    mux21_ni ix41463 (.Y (nx41462), .A0 (inputs_254__9), .A1 (inputs_255__9), .S0 (
             nx24479)) ;
    oai21 ix45737 (.Y (\output [10]), .A0 (nx22221), .A1 (nx16989), .B0 (nx17347
          )) ;
    mux21 ix16990 (.Y (nx16989), .A0 (nx42418), .A1 (nx43262), .S0 (nx22433)) ;
    mux21_ni ix42419 (.Y (nx42418), .A0 (nx41994), .A1 (nx42414), .S0 (nx22495)
             ) ;
    mux21_ni ix41995 (.Y (nx41994), .A0 (nx41782), .A1 (nx41990), .S0 (nx22617)
             ) ;
    mux21_ni ix41783 (.Y (nx41782), .A0 (nx41776), .A1 (nx41698), .S0 (nx23161)
             ) ;
    oai21 ix41777 (.Y (nx41776), .A0 (nx22321), .A1 (nx16997), .B0 (nx17009)) ;
    mux21 ix16998 (.Y (nx16997), .A0 (nx41740), .A1 (nx41768), .S0 (nx22951)) ;
    mux21_ni ix41741 (.Y (nx41740), .A0 (nx41724), .A1 (nx41736), .S0 (nx23685)
             ) ;
    mux21_ni ix41725 (.Y (nx41724), .A0 (inputs_260__10), .A1 (inputs_261__10), 
             .S0 (nx24479)) ;
    mux21_ni ix41737 (.Y (nx41736), .A0 (inputs_262__10), .A1 (inputs_263__10), 
             .S0 (nx24479)) ;
    mux21_ni ix41769 (.Y (nx41768), .A0 (nx41752), .A1 (nx41764), .S0 (nx23687)
             ) ;
    mux21_ni ix41753 (.Y (nx41752), .A0 (inputs_276__10), .A1 (inputs_277__10), 
             .S0 (nx24479)) ;
    mux21_ni ix41765 (.Y (nx41764), .A0 (inputs_278__10), .A1 (inputs_279__10), 
             .S0 (nx24481)) ;
    nand04 ix17010 (.Y (nx17009), .A0 (nx22321), .A1 (nx23687), .A2 (nx24481), .A3 (
           nx41712)) ;
    mux21_ni ix41713 (.Y (nx41712), .A0 (inputs_259__10), .A1 (inputs_275__10), 
             .S0 (nx22951)) ;
    mux21_ni ix41699 (.Y (nx41698), .A0 (nx41634), .A1 (nx41694), .S0 (nx22951)
             ) ;
    mux21_ni ix41635 (.Y (nx41634), .A0 (nx41602), .A1 (nx41630), .S0 (nx23281)
             ) ;
    mux21_ni ix41603 (.Y (nx41602), .A0 (nx41586), .A1 (nx41598), .S0 (nx23687)
             ) ;
    mux21_ni ix41587 (.Y (nx41586), .A0 (inputs_264__10), .A1 (inputs_265__10), 
             .S0 (nx24481)) ;
    mux21_ni ix41599 (.Y (nx41598), .A0 (inputs_266__10), .A1 (inputs_267__10), 
             .S0 (nx24481)) ;
    mux21_ni ix41631 (.Y (nx41630), .A0 (nx41614), .A1 (nx41626), .S0 (nx23687)
             ) ;
    mux21_ni ix41615 (.Y (nx41614), .A0 (inputs_268__10), .A1 (inputs_269__10), 
             .S0 (nx24481)) ;
    mux21_ni ix41627 (.Y (nx41626), .A0 (inputs_270__10), .A1 (inputs_271__10), 
             .S0 (nx24481)) ;
    mux21_ni ix41695 (.Y (nx41694), .A0 (nx41662), .A1 (nx41690), .S0 (nx23281)
             ) ;
    mux21_ni ix41663 (.Y (nx41662), .A0 (nx41646), .A1 (nx41658), .S0 (nx23687)
             ) ;
    mux21_ni ix41647 (.Y (nx41646), .A0 (inputs_280__10), .A1 (inputs_281__10), 
             .S0 (nx24481)) ;
    mux21_ni ix41659 (.Y (nx41658), .A0 (inputs_282__10), .A1 (inputs_283__10), 
             .S0 (nx24483)) ;
    mux21_ni ix41691 (.Y (nx41690), .A0 (nx41674), .A1 (nx41686), .S0 (nx23687)
             ) ;
    mux21_ni ix41675 (.Y (nx41674), .A0 (inputs_284__10), .A1 (inputs_285__10), 
             .S0 (nx24483)) ;
    mux21_ni ix41687 (.Y (nx41686), .A0 (inputs_286__10), .A1 (inputs_287__10), 
             .S0 (nx24483)) ;
    mux21_ni ix41991 (.Y (nx41990), .A0 (nx41984), .A1 (nx41906), .S0 (nx23163)
             ) ;
    oai21 ix41985 (.Y (nx41984), .A0 (nx22321), .A1 (nx17041), .B0 (nx17053)) ;
    mux21 ix17042 (.Y (nx17041), .A0 (nx41948), .A1 (nx41976), .S0 (nx22951)) ;
    mux21_ni ix41949 (.Y (nx41948), .A0 (nx41932), .A1 (nx41944), .S0 (nx23687)
             ) ;
    mux21_ni ix41933 (.Y (nx41932), .A0 (inputs_292__10), .A1 (inputs_293__10), 
             .S0 (nx24483)) ;
    mux21_ni ix41945 (.Y (nx41944), .A0 (inputs_294__10), .A1 (inputs_295__10), 
             .S0 (nx24483)) ;
    mux21_ni ix41977 (.Y (nx41976), .A0 (nx41960), .A1 (nx41972), .S0 (nx23689)
             ) ;
    mux21_ni ix41961 (.Y (nx41960), .A0 (inputs_308__10), .A1 (inputs_309__10), 
             .S0 (nx24483)) ;
    mux21_ni ix41973 (.Y (nx41972), .A0 (inputs_310__10), .A1 (inputs_311__10), 
             .S0 (nx24483)) ;
    nand04 ix17054 (.Y (nx17053), .A0 (nx22321), .A1 (nx23689), .A2 (nx24485), .A3 (
           nx41920)) ;
    mux21_ni ix41921 (.Y (nx41920), .A0 (inputs_291__10), .A1 (inputs_307__10), 
             .S0 (nx22951)) ;
    mux21_ni ix41907 (.Y (nx41906), .A0 (nx41842), .A1 (nx41902), .S0 (nx22951)
             ) ;
    mux21_ni ix41843 (.Y (nx41842), .A0 (nx41810), .A1 (nx41838), .S0 (nx23283)
             ) ;
    mux21_ni ix41811 (.Y (nx41810), .A0 (nx41794), .A1 (nx41806), .S0 (nx23689)
             ) ;
    mux21_ni ix41795 (.Y (nx41794), .A0 (inputs_296__10), .A1 (inputs_297__10), 
             .S0 (nx24485)) ;
    mux21_ni ix41807 (.Y (nx41806), .A0 (inputs_298__10), .A1 (inputs_299__10), 
             .S0 (nx24485)) ;
    mux21_ni ix41839 (.Y (nx41838), .A0 (nx41822), .A1 (nx41834), .S0 (nx23689)
             ) ;
    mux21_ni ix41823 (.Y (nx41822), .A0 (inputs_300__10), .A1 (inputs_301__10), 
             .S0 (nx24485)) ;
    mux21_ni ix41835 (.Y (nx41834), .A0 (inputs_302__10), .A1 (inputs_303__10), 
             .S0 (nx24485)) ;
    mux21_ni ix41903 (.Y (nx41902), .A0 (nx41870), .A1 (nx41898), .S0 (nx23283)
             ) ;
    mux21_ni ix41871 (.Y (nx41870), .A0 (nx41854), .A1 (nx41866), .S0 (nx23689)
             ) ;
    mux21_ni ix41855 (.Y (nx41854), .A0 (inputs_312__10), .A1 (inputs_313__10), 
             .S0 (nx24485)) ;
    mux21_ni ix41867 (.Y (nx41866), .A0 (inputs_314__10), .A1 (inputs_315__10), 
             .S0 (nx24485)) ;
    mux21_ni ix41899 (.Y (nx41898), .A0 (nx41882), .A1 (nx41894), .S0 (nx23689)
             ) ;
    mux21_ni ix41883 (.Y (nx41882), .A0 (inputs_316__10), .A1 (inputs_317__10), 
             .S0 (nx24487)) ;
    mux21_ni ix41895 (.Y (nx41894), .A0 (inputs_318__10), .A1 (inputs_319__10), 
             .S0 (nx24487)) ;
    mux21_ni ix42415 (.Y (nx42414), .A0 (nx42202), .A1 (nx42410), .S0 (nx22617)
             ) ;
    mux21_ni ix42203 (.Y (nx42202), .A0 (nx42196), .A1 (nx42118), .S0 (nx23163)
             ) ;
    oai21 ix42197 (.Y (nx42196), .A0 (nx22321), .A1 (nx17085), .B0 (nx17095)) ;
    mux21 ix17086 (.Y (nx17085), .A0 (nx42160), .A1 (nx42188), .S0 (nx22953)) ;
    mux21_ni ix42161 (.Y (nx42160), .A0 (nx42144), .A1 (nx42156), .S0 (nx23689)
             ) ;
    mux21_ni ix42145 (.Y (nx42144), .A0 (inputs_324__10), .A1 (inputs_325__10), 
             .S0 (nx24487)) ;
    mux21_ni ix42157 (.Y (nx42156), .A0 (inputs_326__10), .A1 (inputs_327__10), 
             .S0 (nx24487)) ;
    mux21_ni ix42189 (.Y (nx42188), .A0 (nx42172), .A1 (nx42184), .S0 (nx23691)
             ) ;
    mux21_ni ix42173 (.Y (nx42172), .A0 (inputs_340__10), .A1 (inputs_341__10), 
             .S0 (nx24487)) ;
    mux21_ni ix42185 (.Y (nx42184), .A0 (inputs_342__10), .A1 (inputs_343__10), 
             .S0 (nx24487)) ;
    nand04 ix17096 (.Y (nx17095), .A0 (nx22321), .A1 (nx23691), .A2 (nx24487), .A3 (
           nx42132)) ;
    mux21_ni ix42133 (.Y (nx42132), .A0 (inputs_323__10), .A1 (inputs_339__10), 
             .S0 (nx22953)) ;
    mux21_ni ix42119 (.Y (nx42118), .A0 (nx42054), .A1 (nx42114), .S0 (nx22953)
             ) ;
    mux21_ni ix42055 (.Y (nx42054), .A0 (nx42022), .A1 (nx42050), .S0 (nx23283)
             ) ;
    mux21_ni ix42023 (.Y (nx42022), .A0 (nx42006), .A1 (nx42018), .S0 (nx23691)
             ) ;
    mux21_ni ix42007 (.Y (nx42006), .A0 (inputs_328__10), .A1 (inputs_329__10), 
             .S0 (nx24489)) ;
    mux21_ni ix42019 (.Y (nx42018), .A0 (inputs_330__10), .A1 (inputs_331__10), 
             .S0 (nx24489)) ;
    mux21_ni ix42051 (.Y (nx42050), .A0 (nx42034), .A1 (nx42046), .S0 (nx23691)
             ) ;
    mux21_ni ix42035 (.Y (nx42034), .A0 (inputs_332__10), .A1 (inputs_333__10), 
             .S0 (nx24489)) ;
    mux21_ni ix42047 (.Y (nx42046), .A0 (inputs_334__10), .A1 (inputs_335__10), 
             .S0 (nx24489)) ;
    mux21_ni ix42115 (.Y (nx42114), .A0 (nx42082), .A1 (nx42110), .S0 (nx23283)
             ) ;
    mux21_ni ix42083 (.Y (nx42082), .A0 (nx42066), .A1 (nx42078), .S0 (nx23691)
             ) ;
    mux21_ni ix42067 (.Y (nx42066), .A0 (inputs_344__10), .A1 (inputs_345__10), 
             .S0 (nx24489)) ;
    mux21_ni ix42079 (.Y (nx42078), .A0 (inputs_346__10), .A1 (inputs_347__10), 
             .S0 (nx24489)) ;
    mux21_ni ix42111 (.Y (nx42110), .A0 (nx42094), .A1 (nx42106), .S0 (nx23691)
             ) ;
    mux21_ni ix42095 (.Y (nx42094), .A0 (inputs_348__10), .A1 (inputs_349__10), 
             .S0 (nx24489)) ;
    mux21_ni ix42107 (.Y (nx42106), .A0 (inputs_350__10), .A1 (inputs_351__10), 
             .S0 (nx24491)) ;
    mux21_ni ix42411 (.Y (nx42410), .A0 (nx42404), .A1 (nx42326), .S0 (nx23163)
             ) ;
    oai21 ix42405 (.Y (nx42404), .A0 (nx22323), .A1 (nx17127), .B0 (nx17139)) ;
    mux21 ix17128 (.Y (nx17127), .A0 (nx42368), .A1 (nx42396), .S0 (nx22953)) ;
    mux21_ni ix42369 (.Y (nx42368), .A0 (nx42352), .A1 (nx42364), .S0 (nx23691)
             ) ;
    mux21_ni ix42353 (.Y (nx42352), .A0 (inputs_356__10), .A1 (inputs_357__10), 
             .S0 (nx24491)) ;
    mux21_ni ix42365 (.Y (nx42364), .A0 (inputs_358__10), .A1 (inputs_359__10), 
             .S0 (nx24491)) ;
    mux21_ni ix42397 (.Y (nx42396), .A0 (nx42380), .A1 (nx42392), .S0 (nx23693)
             ) ;
    mux21_ni ix42381 (.Y (nx42380), .A0 (inputs_372__10), .A1 (inputs_373__10), 
             .S0 (nx24491)) ;
    mux21_ni ix42393 (.Y (nx42392), .A0 (inputs_374__10), .A1 (inputs_375__10), 
             .S0 (nx24491)) ;
    nand04 ix17140 (.Y (nx17139), .A0 (nx22323), .A1 (nx23693), .A2 (nx24491), .A3 (
           nx42340)) ;
    mux21_ni ix42341 (.Y (nx42340), .A0 (inputs_355__10), .A1 (inputs_371__10), 
             .S0 (nx22953)) ;
    mux21_ni ix42327 (.Y (nx42326), .A0 (nx42262), .A1 (nx42322), .S0 (nx22953)
             ) ;
    mux21_ni ix42263 (.Y (nx42262), .A0 (nx42230), .A1 (nx42258), .S0 (nx23283)
             ) ;
    mux21_ni ix42231 (.Y (nx42230), .A0 (nx42214), .A1 (nx42226), .S0 (nx23693)
             ) ;
    mux21_ni ix42215 (.Y (nx42214), .A0 (inputs_360__10), .A1 (inputs_361__10), 
             .S0 (nx24491)) ;
    mux21_ni ix42227 (.Y (nx42226), .A0 (inputs_362__10), .A1 (inputs_363__10), 
             .S0 (nx24493)) ;
    mux21_ni ix42259 (.Y (nx42258), .A0 (nx42242), .A1 (nx42254), .S0 (nx23693)
             ) ;
    mux21_ni ix42243 (.Y (nx42242), .A0 (inputs_364__10), .A1 (inputs_365__10), 
             .S0 (nx24493)) ;
    mux21_ni ix42255 (.Y (nx42254), .A0 (inputs_366__10), .A1 (inputs_367__10), 
             .S0 (nx24493)) ;
    mux21_ni ix42323 (.Y (nx42322), .A0 (nx42290), .A1 (nx42318), .S0 (nx23283)
             ) ;
    mux21_ni ix42291 (.Y (nx42290), .A0 (nx42274), .A1 (nx42286), .S0 (nx23693)
             ) ;
    mux21_ni ix42275 (.Y (nx42274), .A0 (inputs_376__10), .A1 (inputs_377__10), 
             .S0 (nx24493)) ;
    mux21_ni ix42287 (.Y (nx42286), .A0 (inputs_378__10), .A1 (inputs_379__10), 
             .S0 (nx24493)) ;
    mux21_ni ix42319 (.Y (nx42318), .A0 (nx42302), .A1 (nx42314), .S0 (nx23693)
             ) ;
    mux21_ni ix42303 (.Y (nx42302), .A0 (inputs_380__10), .A1 (inputs_381__10), 
             .S0 (nx24493)) ;
    mux21_ni ix42315 (.Y (nx42314), .A0 (inputs_382__10), .A1 (inputs_383__10), 
             .S0 (nx24493)) ;
    mux21_ni ix43263 (.Y (nx43262), .A0 (nx42838), .A1 (nx43258), .S0 (nx22497)
             ) ;
    mux21_ni ix42839 (.Y (nx42838), .A0 (nx42626), .A1 (nx42834), .S0 (nx22619)
             ) ;
    mux21_ni ix42627 (.Y (nx42626), .A0 (nx42620), .A1 (nx42542), .S0 (nx23163)
             ) ;
    oai21 ix42621 (.Y (nx42620), .A0 (nx22323), .A1 (nx17175), .B0 (nx17187)) ;
    mux21 ix17176 (.Y (nx17175), .A0 (nx42584), .A1 (nx42612), .S0 (nx22953)) ;
    mux21_ni ix42585 (.Y (nx42584), .A0 (nx42568), .A1 (nx42580), .S0 (nx23693)
             ) ;
    mux21_ni ix42569 (.Y (nx42568), .A0 (inputs_388__10), .A1 (inputs_389__10), 
             .S0 (nx24495)) ;
    mux21_ni ix42581 (.Y (nx42580), .A0 (inputs_390__10), .A1 (inputs_391__10), 
             .S0 (nx24495)) ;
    mux21_ni ix42613 (.Y (nx42612), .A0 (nx42596), .A1 (nx42608), .S0 (nx23695)
             ) ;
    mux21_ni ix42597 (.Y (nx42596), .A0 (inputs_404__10), .A1 (inputs_405__10), 
             .S0 (nx24495)) ;
    mux21_ni ix42609 (.Y (nx42608), .A0 (inputs_406__10), .A1 (inputs_407__10), 
             .S0 (nx24495)) ;
    nand04 ix17188 (.Y (nx17187), .A0 (nx22323), .A1 (nx23695), .A2 (nx24495), .A3 (
           nx42556)) ;
    mux21_ni ix42557 (.Y (nx42556), .A0 (inputs_387__10), .A1 (inputs_403__10), 
             .S0 (nx22955)) ;
    mux21_ni ix42543 (.Y (nx42542), .A0 (nx42478), .A1 (nx42538), .S0 (nx22955)
             ) ;
    mux21_ni ix42479 (.Y (nx42478), .A0 (nx42446), .A1 (nx42474), .S0 (nx23283)
             ) ;
    mux21_ni ix42447 (.Y (nx42446), .A0 (nx42430), .A1 (nx42442), .S0 (nx23695)
             ) ;
    mux21_ni ix42431 (.Y (nx42430), .A0 (inputs_392__10), .A1 (inputs_393__10), 
             .S0 (nx24495)) ;
    mux21_ni ix42443 (.Y (nx42442), .A0 (inputs_394__10), .A1 (inputs_395__10), 
             .S0 (nx24495)) ;
    mux21_ni ix42475 (.Y (nx42474), .A0 (nx42458), .A1 (nx42470), .S0 (nx23695)
             ) ;
    mux21_ni ix42459 (.Y (nx42458), .A0 (inputs_396__10), .A1 (inputs_397__10), 
             .S0 (nx24497)) ;
    mux21_ni ix42471 (.Y (nx42470), .A0 (inputs_398__10), .A1 (inputs_399__10), 
             .S0 (nx24497)) ;
    mux21_ni ix42539 (.Y (nx42538), .A0 (nx42506), .A1 (nx42534), .S0 (nx23285)
             ) ;
    mux21_ni ix42507 (.Y (nx42506), .A0 (nx42490), .A1 (nx42502), .S0 (nx23695)
             ) ;
    mux21_ni ix42491 (.Y (nx42490), .A0 (inputs_408__10), .A1 (inputs_409__10), 
             .S0 (nx24497)) ;
    mux21_ni ix42503 (.Y (nx42502), .A0 (inputs_410__10), .A1 (inputs_411__10), 
             .S0 (nx24497)) ;
    mux21_ni ix42535 (.Y (nx42534), .A0 (nx42518), .A1 (nx42530), .S0 (nx23695)
             ) ;
    mux21_ni ix42519 (.Y (nx42518), .A0 (inputs_412__10), .A1 (inputs_413__10), 
             .S0 (nx24497)) ;
    mux21_ni ix42531 (.Y (nx42530), .A0 (inputs_414__10), .A1 (inputs_415__10), 
             .S0 (nx24497)) ;
    mux21_ni ix42835 (.Y (nx42834), .A0 (nx42828), .A1 (nx42750), .S0 (nx23163)
             ) ;
    oai21 ix42829 (.Y (nx42828), .A0 (nx22323), .A1 (nx17217), .B0 (nx17229)) ;
    mux21 ix17218 (.Y (nx17217), .A0 (nx42792), .A1 (nx42820), .S0 (nx22955)) ;
    mux21_ni ix42793 (.Y (nx42792), .A0 (nx42776), .A1 (nx42788), .S0 (nx23695)
             ) ;
    mux21_ni ix42777 (.Y (nx42776), .A0 (inputs_420__10), .A1 (inputs_421__10), 
             .S0 (nx24497)) ;
    mux21_ni ix42789 (.Y (nx42788), .A0 (inputs_422__10), .A1 (inputs_423__10), 
             .S0 (nx24499)) ;
    mux21_ni ix42821 (.Y (nx42820), .A0 (nx42804), .A1 (nx42816), .S0 (nx23697)
             ) ;
    mux21_ni ix42805 (.Y (nx42804), .A0 (inputs_436__10), .A1 (inputs_437__10), 
             .S0 (nx24499)) ;
    mux21_ni ix42817 (.Y (nx42816), .A0 (inputs_438__10), .A1 (inputs_439__10), 
             .S0 (nx24499)) ;
    nand04 ix17230 (.Y (nx17229), .A0 (nx22323), .A1 (nx23697), .A2 (nx24499), .A3 (
           nx42764)) ;
    mux21_ni ix42765 (.Y (nx42764), .A0 (inputs_419__10), .A1 (inputs_435__10), 
             .S0 (nx22955)) ;
    mux21_ni ix42751 (.Y (nx42750), .A0 (nx42686), .A1 (nx42746), .S0 (nx22955)
             ) ;
    mux21_ni ix42687 (.Y (nx42686), .A0 (nx42654), .A1 (nx42682), .S0 (nx23285)
             ) ;
    mux21_ni ix42655 (.Y (nx42654), .A0 (nx42638), .A1 (nx42650), .S0 (nx23697)
             ) ;
    mux21_ni ix42639 (.Y (nx42638), .A0 (inputs_424__10), .A1 (inputs_425__10), 
             .S0 (nx24499)) ;
    mux21_ni ix42651 (.Y (nx42650), .A0 (inputs_426__10), .A1 (inputs_427__10), 
             .S0 (nx24499)) ;
    mux21_ni ix42683 (.Y (nx42682), .A0 (nx42666), .A1 (nx42678), .S0 (nx23697)
             ) ;
    mux21_ni ix42667 (.Y (nx42666), .A0 (inputs_428__10), .A1 (inputs_429__10), 
             .S0 (nx24499)) ;
    mux21_ni ix42679 (.Y (nx42678), .A0 (inputs_430__10), .A1 (inputs_431__10), 
             .S0 (nx24501)) ;
    mux21_ni ix42747 (.Y (nx42746), .A0 (nx42714), .A1 (nx42742), .S0 (nx23285)
             ) ;
    mux21_ni ix42715 (.Y (nx42714), .A0 (nx42698), .A1 (nx42710), .S0 (nx23697)
             ) ;
    mux21_ni ix42699 (.Y (nx42698), .A0 (inputs_440__10), .A1 (inputs_441__10), 
             .S0 (nx24501)) ;
    mux21_ni ix42711 (.Y (nx42710), .A0 (inputs_442__10), .A1 (inputs_443__10), 
             .S0 (nx24501)) ;
    mux21_ni ix42743 (.Y (nx42742), .A0 (nx42726), .A1 (nx42738), .S0 (nx23697)
             ) ;
    mux21_ni ix42727 (.Y (nx42726), .A0 (inputs_444__10), .A1 (inputs_445__10), 
             .S0 (nx24501)) ;
    mux21_ni ix42739 (.Y (nx42738), .A0 (inputs_446__10), .A1 (inputs_447__10), 
             .S0 (nx24501)) ;
    mux21_ni ix43259 (.Y (nx43258), .A0 (nx43046), .A1 (nx43254), .S0 (nx22619)
             ) ;
    mux21_ni ix43047 (.Y (nx43046), .A0 (nx43040), .A1 (nx42962), .S0 (nx23163)
             ) ;
    oai21 ix43041 (.Y (nx43040), .A0 (nx22323), .A1 (nx17263), .B0 (nx17275)) ;
    mux21 ix17264 (.Y (nx17263), .A0 (nx43004), .A1 (nx43032), .S0 (nx22955)) ;
    mux21_ni ix43005 (.Y (nx43004), .A0 (nx42988), .A1 (nx43000), .S0 (nx23697)
             ) ;
    mux21_ni ix42989 (.Y (nx42988), .A0 (inputs_452__10), .A1 (inputs_453__10), 
             .S0 (nx24501)) ;
    mux21_ni ix43001 (.Y (nx43000), .A0 (inputs_454__10), .A1 (inputs_455__10), 
             .S0 (nx24501)) ;
    mux21_ni ix43033 (.Y (nx43032), .A0 (nx43016), .A1 (nx43028), .S0 (nx23699)
             ) ;
    mux21_ni ix43017 (.Y (nx43016), .A0 (inputs_468__10), .A1 (inputs_469__10), 
             .S0 (nx24503)) ;
    mux21_ni ix43029 (.Y (nx43028), .A0 (inputs_470__10), .A1 (inputs_471__10), 
             .S0 (nx24503)) ;
    nand04 ix17276 (.Y (nx17275), .A0 (nx22325), .A1 (nx23699), .A2 (nx24503), .A3 (
           nx42976)) ;
    mux21_ni ix42977 (.Y (nx42976), .A0 (inputs_451__10), .A1 (inputs_467__10), 
             .S0 (nx22955)) ;
    mux21_ni ix42963 (.Y (nx42962), .A0 (nx42898), .A1 (nx42958), .S0 (nx22957)
             ) ;
    mux21_ni ix42899 (.Y (nx42898), .A0 (nx42866), .A1 (nx42894), .S0 (nx23285)
             ) ;
    mux21_ni ix42867 (.Y (nx42866), .A0 (nx42850), .A1 (nx42862), .S0 (nx23699)
             ) ;
    mux21_ni ix42851 (.Y (nx42850), .A0 (inputs_456__10), .A1 (inputs_457__10), 
             .S0 (nx24503)) ;
    mux21_ni ix42863 (.Y (nx42862), .A0 (inputs_458__10), .A1 (inputs_459__10), 
             .S0 (nx24503)) ;
    mux21_ni ix42895 (.Y (nx42894), .A0 (nx42878), .A1 (nx42890), .S0 (nx23699)
             ) ;
    mux21_ni ix42879 (.Y (nx42878), .A0 (inputs_460__10), .A1 (inputs_461__10), 
             .S0 (nx24503)) ;
    mux21_ni ix42891 (.Y (nx42890), .A0 (inputs_462__10), .A1 (inputs_463__10), 
             .S0 (nx24503)) ;
    mux21_ni ix42959 (.Y (nx42958), .A0 (nx42926), .A1 (nx42954), .S0 (nx23285)
             ) ;
    mux21_ni ix42927 (.Y (nx42926), .A0 (nx42910), .A1 (nx42922), .S0 (nx23699)
             ) ;
    mux21_ni ix42911 (.Y (nx42910), .A0 (inputs_472__10), .A1 (inputs_473__10), 
             .S0 (nx24505)) ;
    mux21_ni ix42923 (.Y (nx42922), .A0 (inputs_474__10), .A1 (inputs_475__10), 
             .S0 (nx24505)) ;
    mux21_ni ix42955 (.Y (nx42954), .A0 (nx42938), .A1 (nx42950), .S0 (nx23699)
             ) ;
    mux21_ni ix42939 (.Y (nx42938), .A0 (inputs_476__10), .A1 (inputs_477__10), 
             .S0 (nx24505)) ;
    mux21_ni ix42951 (.Y (nx42950), .A0 (inputs_478__10), .A1 (inputs_479__10), 
             .S0 (nx24505)) ;
    mux21_ni ix43255 (.Y (nx43254), .A0 (nx43248), .A1 (nx43170), .S0 (nx23163)
             ) ;
    oai21 ix43249 (.Y (nx43248), .A0 (nx22325), .A1 (nx17305), .B0 (nx17319)) ;
    mux21 ix17306 (.Y (nx17305), .A0 (nx43212), .A1 (nx43240), .S0 (nx22957)) ;
    mux21_ni ix43213 (.Y (nx43212), .A0 (nx43196), .A1 (nx43208), .S0 (nx23699)
             ) ;
    mux21_ni ix43197 (.Y (nx43196), .A0 (inputs_484__10), .A1 (inputs_485__10), 
             .S0 (nx24505)) ;
    mux21_ni ix43209 (.Y (nx43208), .A0 (inputs_486__10), .A1 (inputs_487__10), 
             .S0 (nx24505)) ;
    mux21_ni ix43241 (.Y (nx43240), .A0 (nx43224), .A1 (nx43236), .S0 (nx23701)
             ) ;
    mux21_ni ix43225 (.Y (nx43224), .A0 (inputs_500__10), .A1 (inputs_501__10), 
             .S0 (nx24505)) ;
    mux21_ni ix43237 (.Y (nx43236), .A0 (inputs_502__10), .A1 (inputs_503__10), 
             .S0 (nx24507)) ;
    nand04 ix17320 (.Y (nx17319), .A0 (nx22325), .A1 (nx23701), .A2 (nx24507), .A3 (
           nx43184)) ;
    mux21_ni ix43185 (.Y (nx43184), .A0 (inputs_483__10), .A1 (inputs_499__10), 
             .S0 (nx22957)) ;
    mux21_ni ix43171 (.Y (nx43170), .A0 (nx43106), .A1 (nx43166), .S0 (nx22957)
             ) ;
    mux21_ni ix43107 (.Y (nx43106), .A0 (nx43074), .A1 (nx43102), .S0 (nx23285)
             ) ;
    mux21_ni ix43075 (.Y (nx43074), .A0 (nx43058), .A1 (nx43070), .S0 (nx23701)
             ) ;
    mux21_ni ix43059 (.Y (nx43058), .A0 (inputs_488__10), .A1 (inputs_489__10), 
             .S0 (nx24507)) ;
    mux21_ni ix43071 (.Y (nx43070), .A0 (inputs_490__10), .A1 (inputs_491__10), 
             .S0 (nx24507)) ;
    mux21_ni ix43103 (.Y (nx43102), .A0 (nx43086), .A1 (nx43098), .S0 (nx23701)
             ) ;
    mux21_ni ix43087 (.Y (nx43086), .A0 (inputs_492__10), .A1 (inputs_493__10), 
             .S0 (nx24507)) ;
    mux21_ni ix43099 (.Y (nx43098), .A0 (inputs_494__10), .A1 (inputs_495__10), 
             .S0 (nx24507)) ;
    mux21_ni ix43167 (.Y (nx43166), .A0 (nx43134), .A1 (nx43162), .S0 (nx23285)
             ) ;
    mux21_ni ix43135 (.Y (nx43134), .A0 (nx43118), .A1 (nx43130), .S0 (nx23701)
             ) ;
    mux21_ni ix43119 (.Y (nx43118), .A0 (inputs_504__10), .A1 (inputs_505__10), 
             .S0 (nx24507)) ;
    mux21_ni ix43131 (.Y (nx43130), .A0 (inputs_506__10), .A1 (inputs_507__10), 
             .S0 (nx24509)) ;
    mux21_ni ix43163 (.Y (nx43162), .A0 (nx43146), .A1 (nx43158), .S0 (nx23701)
             ) ;
    mux21_ni ix43147 (.Y (nx43146), .A0 (inputs_508__10), .A1 (inputs_509__10), 
             .S0 (nx24509)) ;
    mux21_ni ix43159 (.Y (nx43158), .A0 (inputs_510__10), .A1 (inputs_511__10), 
             .S0 (nx24509)) ;
    aoi32 ix17348 (.Y (nx17347), .A0 (nx44032), .A1 (nx22387), .A2 (nx22325), .B0 (
          nx22223), .B1 (nx45728)) ;
    oai21 ix44033 (.Y (nx44032), .A0 (nx23701), .A1 (nx17351), .B0 (nx17455)) ;
    mux21 ix17352 (.Y (nx17351), .A0 (nx43770), .A1 (nx44022), .S0 (nx24509)) ;
    mux21_ni ix43771 (.Y (nx43770), .A0 (nx43642), .A1 (nx43766), .S0 (nx22401)
             ) ;
    mux21_ni ix43643 (.Y (nx43642), .A0 (nx43578), .A1 (nx43638), .S0 (nx22433)
             ) ;
    mux21_ni ix43579 (.Y (nx43578), .A0 (nx43546), .A1 (nx43574), .S0 (nx22497)
             ) ;
    mux21_ni ix43547 (.Y (nx43546), .A0 (nx43530), .A1 (nx43542), .S0 (nx22619)
             ) ;
    mux21_ni ix43531 (.Y (nx43530), .A0 (inputs_0__10), .A1 (inputs_16__10), .S0 (
             nx22957)) ;
    mux21_ni ix43543 (.Y (nx43542), .A0 (inputs_32__10), .A1 (inputs_48__10), .S0 (
             nx22957)) ;
    mux21_ni ix43575 (.Y (nx43574), .A0 (nx43558), .A1 (nx43570), .S0 (nx22619)
             ) ;
    mux21_ni ix43559 (.Y (nx43558), .A0 (inputs_64__10), .A1 (inputs_80__10), .S0 (
             nx22957)) ;
    mux21_ni ix43571 (.Y (nx43570), .A0 (inputs_96__10), .A1 (inputs_112__10), .S0 (
             nx22959)) ;
    mux21_ni ix43639 (.Y (nx43638), .A0 (nx43606), .A1 (nx43634), .S0 (nx22497)
             ) ;
    mux21_ni ix43607 (.Y (nx43606), .A0 (nx43590), .A1 (nx43602), .S0 (nx22619)
             ) ;
    mux21_ni ix43591 (.Y (nx43590), .A0 (inputs_128__10), .A1 (inputs_144__10), 
             .S0 (nx22959)) ;
    mux21_ni ix43603 (.Y (nx43602), .A0 (inputs_160__10), .A1 (inputs_176__10), 
             .S0 (nx22959)) ;
    mux21_ni ix43635 (.Y (nx43634), .A0 (nx43618), .A1 (nx43630), .S0 (nx22619)
             ) ;
    mux21_ni ix43619 (.Y (nx43618), .A0 (inputs_192__10), .A1 (inputs_208__10), 
             .S0 (nx22959)) ;
    mux21_ni ix43631 (.Y (nx43630), .A0 (inputs_224__10), .A1 (inputs_240__10), 
             .S0 (nx22959)) ;
    mux21_ni ix43767 (.Y (nx43766), .A0 (nx43702), .A1 (nx43762), .S0 (nx22433)
             ) ;
    mux21_ni ix43703 (.Y (nx43702), .A0 (nx43670), .A1 (nx43698), .S0 (nx22497)
             ) ;
    mux21_ni ix43671 (.Y (nx43670), .A0 (nx43654), .A1 (nx43666), .S0 (nx22619)
             ) ;
    mux21_ni ix43655 (.Y (nx43654), .A0 (inputs_256__10), .A1 (inputs_272__10), 
             .S0 (nx22959)) ;
    mux21_ni ix43667 (.Y (nx43666), .A0 (inputs_288__10), .A1 (inputs_304__10), 
             .S0 (nx22959)) ;
    mux21_ni ix43699 (.Y (nx43698), .A0 (nx43682), .A1 (nx43694), .S0 (nx22621)
             ) ;
    mux21_ni ix43683 (.Y (nx43682), .A0 (inputs_320__10), .A1 (inputs_336__10), 
             .S0 (nx22961)) ;
    mux21_ni ix43695 (.Y (nx43694), .A0 (inputs_352__10), .A1 (inputs_368__10), 
             .S0 (nx22961)) ;
    mux21_ni ix43763 (.Y (nx43762), .A0 (nx43730), .A1 (nx43758), .S0 (nx22497)
             ) ;
    mux21_ni ix43731 (.Y (nx43730), .A0 (nx43714), .A1 (nx43726), .S0 (nx22621)
             ) ;
    mux21_ni ix43715 (.Y (nx43714), .A0 (inputs_384__10), .A1 (inputs_400__10), 
             .S0 (nx22961)) ;
    mux21_ni ix43727 (.Y (nx43726), .A0 (inputs_416__10), .A1 (inputs_432__10), 
             .S0 (nx22961)) ;
    mux21_ni ix43759 (.Y (nx43758), .A0 (nx43742), .A1 (nx43754), .S0 (nx22621)
             ) ;
    mux21_ni ix43743 (.Y (nx43742), .A0 (inputs_448__10), .A1 (inputs_464__10), 
             .S0 (nx22961)) ;
    mux21_ni ix43755 (.Y (nx43754), .A0 (inputs_480__10), .A1 (inputs_496__10), 
             .S0 (nx22961)) ;
    mux21_ni ix44023 (.Y (nx44022), .A0 (nx43894), .A1 (nx44018), .S0 (nx22401)
             ) ;
    mux21_ni ix43895 (.Y (nx43894), .A0 (nx43830), .A1 (nx43890), .S0 (nx22433)
             ) ;
    mux21_ni ix43831 (.Y (nx43830), .A0 (nx43798), .A1 (nx43826), .S0 (nx22497)
             ) ;
    mux21_ni ix43799 (.Y (nx43798), .A0 (nx43782), .A1 (nx43794), .S0 (nx22621)
             ) ;
    mux21_ni ix43783 (.Y (nx43782), .A0 (inputs_1__10), .A1 (inputs_17__10), .S0 (
             nx22961)) ;
    mux21_ni ix43795 (.Y (nx43794), .A0 (inputs_33__10), .A1 (inputs_49__10), .S0 (
             nx22963)) ;
    mux21_ni ix43827 (.Y (nx43826), .A0 (nx43810), .A1 (nx43822), .S0 (nx22621)
             ) ;
    mux21_ni ix43811 (.Y (nx43810), .A0 (inputs_65__10), .A1 (inputs_81__10), .S0 (
             nx22963)) ;
    mux21_ni ix43823 (.Y (nx43822), .A0 (inputs_97__10), .A1 (inputs_113__10), .S0 (
             nx22963)) ;
    mux21_ni ix43891 (.Y (nx43890), .A0 (nx43858), .A1 (nx43886), .S0 (nx22497)
             ) ;
    mux21_ni ix43859 (.Y (nx43858), .A0 (nx43842), .A1 (nx43854), .S0 (nx22621)
             ) ;
    mux21_ni ix43843 (.Y (nx43842), .A0 (inputs_129__10), .A1 (inputs_145__10), 
             .S0 (nx22963)) ;
    mux21_ni ix43855 (.Y (nx43854), .A0 (inputs_161__10), .A1 (inputs_177__10), 
             .S0 (nx22963)) ;
    mux21_ni ix43887 (.Y (nx43886), .A0 (nx43870), .A1 (nx43882), .S0 (nx22621)
             ) ;
    mux21_ni ix43871 (.Y (nx43870), .A0 (inputs_193__10), .A1 (inputs_209__10), 
             .S0 (nx22963)) ;
    mux21_ni ix43883 (.Y (nx43882), .A0 (inputs_225__10), .A1 (inputs_241__10), 
             .S0 (nx22963)) ;
    mux21_ni ix44019 (.Y (nx44018), .A0 (nx43954), .A1 (nx44014), .S0 (nx22435)
             ) ;
    mux21_ni ix43955 (.Y (nx43954), .A0 (nx43922), .A1 (nx43950), .S0 (nx22499)
             ) ;
    mux21_ni ix43923 (.Y (nx43922), .A0 (nx43906), .A1 (nx43918), .S0 (nx22623)
             ) ;
    mux21_ni ix43907 (.Y (nx43906), .A0 (inputs_257__10), .A1 (inputs_273__10), 
             .S0 (nx22965)) ;
    mux21_ni ix43919 (.Y (nx43918), .A0 (inputs_289__10), .A1 (inputs_305__10), 
             .S0 (nx22965)) ;
    mux21_ni ix43951 (.Y (nx43950), .A0 (nx43934), .A1 (nx43946), .S0 (nx22623)
             ) ;
    mux21_ni ix43935 (.Y (nx43934), .A0 (inputs_321__10), .A1 (inputs_337__10), 
             .S0 (nx22965)) ;
    mux21_ni ix43947 (.Y (nx43946), .A0 (inputs_353__10), .A1 (inputs_369__10), 
             .S0 (nx22965)) ;
    mux21_ni ix44015 (.Y (nx44014), .A0 (nx43982), .A1 (nx44010), .S0 (nx22499)
             ) ;
    mux21_ni ix43983 (.Y (nx43982), .A0 (nx43966), .A1 (nx43978), .S0 (nx22623)
             ) ;
    mux21_ni ix43967 (.Y (nx43966), .A0 (inputs_385__10), .A1 (inputs_401__10), 
             .S0 (nx22965)) ;
    mux21_ni ix43979 (.Y (nx43978), .A0 (inputs_417__10), .A1 (inputs_433__10), 
             .S0 (nx22965)) ;
    mux21_ni ix44011 (.Y (nx44010), .A0 (nx43994), .A1 (nx44006), .S0 (nx22623)
             ) ;
    mux21_ni ix43995 (.Y (nx43994), .A0 (inputs_449__10), .A1 (inputs_465__10), 
             .S0 (nx22965)) ;
    mux21_ni ix44007 (.Y (nx44006), .A0 (inputs_481__10), .A1 (inputs_497__10), 
             .S0 (nx22967)) ;
    nand03 ix17456 (.Y (nx17455), .A0 (nx43516), .A1 (nx23703), .A2 (nx22381)) ;
    mux21_ni ix43517 (.Y (nx43516), .A0 (nx43388), .A1 (nx43512), .S0 (nx22401)
             ) ;
    mux21_ni ix43389 (.Y (nx43388), .A0 (nx43324), .A1 (nx43384), .S0 (nx22435)
             ) ;
    mux21_ni ix43325 (.Y (nx43324), .A0 (nx43292), .A1 (nx43320), .S0 (nx22499)
             ) ;
    mux21_ni ix43293 (.Y (nx43292), .A0 (nx43276), .A1 (nx43288), .S0 (nx22623)
             ) ;
    mux21_ni ix43277 (.Y (nx43276), .A0 (inputs_2__10), .A1 (inputs_18__10), .S0 (
             nx22967)) ;
    mux21_ni ix43289 (.Y (nx43288), .A0 (inputs_34__10), .A1 (inputs_50__10), .S0 (
             nx22967)) ;
    mux21_ni ix43321 (.Y (nx43320), .A0 (nx43304), .A1 (nx43316), .S0 (nx22623)
             ) ;
    mux21_ni ix43305 (.Y (nx43304), .A0 (inputs_66__10), .A1 (inputs_82__10), .S0 (
             nx22967)) ;
    mux21_ni ix43317 (.Y (nx43316), .A0 (inputs_98__10), .A1 (inputs_114__10), .S0 (
             nx22967)) ;
    mux21_ni ix43385 (.Y (nx43384), .A0 (nx43352), .A1 (nx43380), .S0 (nx22499)
             ) ;
    mux21_ni ix43353 (.Y (nx43352), .A0 (nx43336), .A1 (nx43348), .S0 (nx22623)
             ) ;
    mux21_ni ix43337 (.Y (nx43336), .A0 (inputs_130__10), .A1 (inputs_146__10), 
             .S0 (nx22967)) ;
    mux21_ni ix43349 (.Y (nx43348), .A0 (inputs_162__10), .A1 (inputs_178__10), 
             .S0 (nx22967)) ;
    mux21_ni ix43381 (.Y (nx43380), .A0 (nx43364), .A1 (nx43376), .S0 (nx22625)
             ) ;
    mux21_ni ix43365 (.Y (nx43364), .A0 (inputs_194__10), .A1 (inputs_210__10), 
             .S0 (nx22969)) ;
    mux21_ni ix43377 (.Y (nx43376), .A0 (inputs_226__10), .A1 (inputs_242__10), 
             .S0 (nx22969)) ;
    mux21_ni ix43513 (.Y (nx43512), .A0 (nx43448), .A1 (nx43508), .S0 (nx22435)
             ) ;
    mux21_ni ix43449 (.Y (nx43448), .A0 (nx43416), .A1 (nx43444), .S0 (nx22499)
             ) ;
    mux21_ni ix43417 (.Y (nx43416), .A0 (nx43400), .A1 (nx43412), .S0 (nx22625)
             ) ;
    mux21_ni ix43401 (.Y (nx43400), .A0 (inputs_258__10), .A1 (inputs_274__10), 
             .S0 (nx22969)) ;
    mux21_ni ix43413 (.Y (nx43412), .A0 (inputs_290__10), .A1 (inputs_306__10), 
             .S0 (nx22969)) ;
    mux21_ni ix43445 (.Y (nx43444), .A0 (nx43428), .A1 (nx43440), .S0 (nx22625)
             ) ;
    mux21_ni ix43429 (.Y (nx43428), .A0 (inputs_322__10), .A1 (inputs_338__10), 
             .S0 (nx22969)) ;
    mux21_ni ix43441 (.Y (nx43440), .A0 (inputs_354__10), .A1 (inputs_370__10), 
             .S0 (nx22969)) ;
    mux21_ni ix43509 (.Y (nx43508), .A0 (nx43476), .A1 (nx43504), .S0 (nx22499)
             ) ;
    mux21_ni ix43477 (.Y (nx43476), .A0 (nx43460), .A1 (nx43472), .S0 (nx22625)
             ) ;
    mux21_ni ix43461 (.Y (nx43460), .A0 (inputs_386__10), .A1 (inputs_402__10), 
             .S0 (nx22969)) ;
    mux21_ni ix43473 (.Y (nx43472), .A0 (inputs_418__10), .A1 (inputs_434__10), 
             .S0 (nx22971)) ;
    mux21_ni ix43505 (.Y (nx43504), .A0 (nx43488), .A1 (nx43500), .S0 (nx22625)
             ) ;
    mux21_ni ix43489 (.Y (nx43488), .A0 (inputs_450__10), .A1 (inputs_466__10), 
             .S0 (nx22971)) ;
    mux21_ni ix43501 (.Y (nx43500), .A0 (inputs_482__10), .A1 (inputs_498__10), 
             .S0 (nx22971)) ;
    mux21_ni ix45729 (.Y (nx45728), .A0 (nx44880), .A1 (nx45724), .S0 (nx22435)
             ) ;
    mux21_ni ix44881 (.Y (nx44880), .A0 (nx44456), .A1 (nx44876), .S0 (nx22499)
             ) ;
    mux21_ni ix44457 (.Y (nx44456), .A0 (nx44244), .A1 (nx44452), .S0 (nx22625)
             ) ;
    mux21_ni ix44245 (.Y (nx44244), .A0 (nx44238), .A1 (nx44160), .S0 (nx23165)
             ) ;
    oai21 ix44239 (.Y (nx44238), .A0 (nx22325), .A1 (nx17515), .B0 (nx17527)) ;
    mux21 ix17516 (.Y (nx17515), .A0 (nx44202), .A1 (nx44230), .S0 (nx22971)) ;
    mux21_ni ix44203 (.Y (nx44202), .A0 (nx44186), .A1 (nx44198), .S0 (nx23703)
             ) ;
    mux21_ni ix44187 (.Y (nx44186), .A0 (inputs_4__10), .A1 (inputs_5__10), .S0 (
             nx24509)) ;
    mux21_ni ix44199 (.Y (nx44198), .A0 (inputs_6__10), .A1 (inputs_7__10), .S0 (
             nx24509)) ;
    mux21_ni ix44231 (.Y (nx44230), .A0 (nx44214), .A1 (nx44226), .S0 (nx23703)
             ) ;
    mux21_ni ix44215 (.Y (nx44214), .A0 (inputs_20__10), .A1 (inputs_21__10), .S0 (
             nx24509)) ;
    mux21_ni ix44227 (.Y (nx44226), .A0 (inputs_22__10), .A1 (inputs_23__10), .S0 (
             nx24511)) ;
    nand04 ix17528 (.Y (nx17527), .A0 (nx22325), .A1 (nx23703), .A2 (nx24511), .A3 (
           nx44174)) ;
    mux21_ni ix44175 (.Y (nx44174), .A0 (inputs_3__10), .A1 (inputs_19__10), .S0 (
             nx22971)) ;
    mux21_ni ix44161 (.Y (nx44160), .A0 (nx44096), .A1 (nx44156), .S0 (nx22971)
             ) ;
    mux21_ni ix44097 (.Y (nx44096), .A0 (nx44064), .A1 (nx44092), .S0 (nx23287)
             ) ;
    mux21_ni ix44065 (.Y (nx44064), .A0 (nx44048), .A1 (nx44060), .S0 (nx23703)
             ) ;
    mux21_ni ix44049 (.Y (nx44048), .A0 (inputs_8__10), .A1 (inputs_9__10), .S0 (
             nx24511)) ;
    mux21_ni ix44061 (.Y (nx44060), .A0 (inputs_10__10), .A1 (inputs_11__10), .S0 (
             nx24511)) ;
    mux21_ni ix44093 (.Y (nx44092), .A0 (nx44076), .A1 (nx44088), .S0 (nx23703)
             ) ;
    mux21_ni ix44077 (.Y (nx44076), .A0 (inputs_12__10), .A1 (inputs_13__10), .S0 (
             nx24511)) ;
    mux21_ni ix44089 (.Y (nx44088), .A0 (inputs_14__10), .A1 (inputs_15__10), .S0 (
             nx24511)) ;
    mux21_ni ix44157 (.Y (nx44156), .A0 (nx44124), .A1 (nx44152), .S0 (nx23287)
             ) ;
    mux21_ni ix44125 (.Y (nx44124), .A0 (nx44108), .A1 (nx44120), .S0 (nx23703)
             ) ;
    mux21_ni ix44109 (.Y (nx44108), .A0 (inputs_24__10), .A1 (inputs_25__10), .S0 (
             nx24511)) ;
    mux21_ni ix44121 (.Y (nx44120), .A0 (inputs_26__10), .A1 (inputs_27__10), .S0 (
             nx24513)) ;
    mux21_ni ix44153 (.Y (nx44152), .A0 (nx44136), .A1 (nx44148), .S0 (nx23705)
             ) ;
    mux21_ni ix44137 (.Y (nx44136), .A0 (inputs_28__10), .A1 (inputs_29__10), .S0 (
             nx24513)) ;
    mux21_ni ix44149 (.Y (nx44148), .A0 (inputs_30__10), .A1 (inputs_31__10), .S0 (
             nx24513)) ;
    mux21_ni ix44453 (.Y (nx44452), .A0 (nx44446), .A1 (nx44368), .S0 (nx23165)
             ) ;
    oai21 ix44447 (.Y (nx44446), .A0 (nx22325), .A1 (nx17557), .B0 (nx17567)) ;
    mux21 ix17558 (.Y (nx17557), .A0 (nx44410), .A1 (nx44438), .S0 (nx22971)) ;
    mux21_ni ix44411 (.Y (nx44410), .A0 (nx44394), .A1 (nx44406), .S0 (nx23705)
             ) ;
    mux21_ni ix44395 (.Y (nx44394), .A0 (inputs_36__10), .A1 (inputs_37__10), .S0 (
             nx24513)) ;
    mux21_ni ix44407 (.Y (nx44406), .A0 (inputs_38__10), .A1 (inputs_39__10), .S0 (
             nx24513)) ;
    mux21_ni ix44439 (.Y (nx44438), .A0 (nx44422), .A1 (nx44434), .S0 (nx23705)
             ) ;
    mux21_ni ix44423 (.Y (nx44422), .A0 (inputs_52__10), .A1 (inputs_53__10), .S0 (
             nx24513)) ;
    mux21_ni ix44435 (.Y (nx44434), .A0 (inputs_54__10), .A1 (inputs_55__10), .S0 (
             nx24513)) ;
    nand04 ix17568 (.Y (nx17567), .A0 (nx22327), .A1 (nx23705), .A2 (nx24515), .A3 (
           nx44382)) ;
    mux21_ni ix44383 (.Y (nx44382), .A0 (inputs_35__10), .A1 (inputs_51__10), .S0 (
             nx22973)) ;
    mux21_ni ix44369 (.Y (nx44368), .A0 (nx44304), .A1 (nx44364), .S0 (nx22973)
             ) ;
    mux21_ni ix44305 (.Y (nx44304), .A0 (nx44272), .A1 (nx44300), .S0 (nx23287)
             ) ;
    mux21_ni ix44273 (.Y (nx44272), .A0 (nx44256), .A1 (nx44268), .S0 (nx23705)
             ) ;
    mux21_ni ix44257 (.Y (nx44256), .A0 (inputs_40__10), .A1 (inputs_41__10), .S0 (
             nx24515)) ;
    mux21_ni ix44269 (.Y (nx44268), .A0 (inputs_42__10), .A1 (inputs_43__10), .S0 (
             nx24515)) ;
    mux21_ni ix44301 (.Y (nx44300), .A0 (nx44284), .A1 (nx44296), .S0 (nx23705)
             ) ;
    mux21_ni ix44285 (.Y (nx44284), .A0 (inputs_44__10), .A1 (inputs_45__10), .S0 (
             nx24515)) ;
    mux21_ni ix44297 (.Y (nx44296), .A0 (inputs_46__10), .A1 (inputs_47__10), .S0 (
             nx24515)) ;
    mux21_ni ix44365 (.Y (nx44364), .A0 (nx44332), .A1 (nx44360), .S0 (nx23287)
             ) ;
    mux21_ni ix44333 (.Y (nx44332), .A0 (nx44316), .A1 (nx44328), .S0 (nx23705)
             ) ;
    mux21_ni ix44317 (.Y (nx44316), .A0 (inputs_56__10), .A1 (inputs_57__10), .S0 (
             nx24515)) ;
    mux21_ni ix44329 (.Y (nx44328), .A0 (inputs_58__10), .A1 (inputs_59__10), .S0 (
             nx24515)) ;
    mux21_ni ix44361 (.Y (nx44360), .A0 (nx44344), .A1 (nx44356), .S0 (nx23707)
             ) ;
    mux21_ni ix44345 (.Y (nx44344), .A0 (inputs_60__10), .A1 (inputs_61__10), .S0 (
             nx24517)) ;
    mux21_ni ix44357 (.Y (nx44356), .A0 (inputs_62__10), .A1 (inputs_63__10), .S0 (
             nx24517)) ;
    mux21_ni ix44877 (.Y (nx44876), .A0 (nx44664), .A1 (nx44872), .S0 (nx22625)
             ) ;
    mux21_ni ix44665 (.Y (nx44664), .A0 (nx44658), .A1 (nx44580), .S0 (nx23165)
             ) ;
    oai21 ix44659 (.Y (nx44658), .A0 (nx22327), .A1 (nx17601), .B0 (nx17613)) ;
    mux21 ix17602 (.Y (nx17601), .A0 (nx44622), .A1 (nx44650), .S0 (nx22973)) ;
    mux21_ni ix44623 (.Y (nx44622), .A0 (nx44606), .A1 (nx44618), .S0 (nx23707)
             ) ;
    mux21_ni ix44607 (.Y (nx44606), .A0 (inputs_68__10), .A1 (inputs_69__10), .S0 (
             nx24517)) ;
    mux21_ni ix44619 (.Y (nx44618), .A0 (inputs_70__10), .A1 (inputs_71__10), .S0 (
             nx24517)) ;
    mux21_ni ix44651 (.Y (nx44650), .A0 (nx44634), .A1 (nx44646), .S0 (nx23707)
             ) ;
    mux21_ni ix44635 (.Y (nx44634), .A0 (inputs_84__10), .A1 (inputs_85__10), .S0 (
             nx24517)) ;
    mux21_ni ix44647 (.Y (nx44646), .A0 (inputs_86__10), .A1 (inputs_87__10), .S0 (
             nx24517)) ;
    nand04 ix17614 (.Y (nx17613), .A0 (nx22327), .A1 (nx23707), .A2 (nx24517), .A3 (
           nx44594)) ;
    mux21_ni ix44595 (.Y (nx44594), .A0 (inputs_67__10), .A1 (inputs_83__10), .S0 (
             nx22973)) ;
    mux21_ni ix44581 (.Y (nx44580), .A0 (nx44516), .A1 (nx44576), .S0 (nx22973)
             ) ;
    mux21_ni ix44517 (.Y (nx44516), .A0 (nx44484), .A1 (nx44512), .S0 (nx23287)
             ) ;
    mux21_ni ix44485 (.Y (nx44484), .A0 (nx44468), .A1 (nx44480), .S0 (nx23707)
             ) ;
    mux21_ni ix44469 (.Y (nx44468), .A0 (inputs_72__10), .A1 (inputs_73__10), .S0 (
             nx24519)) ;
    mux21_ni ix44481 (.Y (nx44480), .A0 (inputs_74__10), .A1 (inputs_75__10), .S0 (
             nx24519)) ;
    mux21_ni ix44513 (.Y (nx44512), .A0 (nx44496), .A1 (nx44508), .S0 (nx23707)
             ) ;
    mux21_ni ix44497 (.Y (nx44496), .A0 (inputs_76__10), .A1 (inputs_77__10), .S0 (
             nx24519)) ;
    mux21_ni ix44509 (.Y (nx44508), .A0 (inputs_78__10), .A1 (inputs_79__10), .S0 (
             nx24519)) ;
    mux21_ni ix44577 (.Y (nx44576), .A0 (nx44544), .A1 (nx44572), .S0 (nx23287)
             ) ;
    mux21_ni ix44545 (.Y (nx44544), .A0 (nx44528), .A1 (nx44540), .S0 (nx23707)
             ) ;
    mux21_ni ix44529 (.Y (nx44528), .A0 (inputs_88__10), .A1 (inputs_89__10), .S0 (
             nx24519)) ;
    mux21_ni ix44541 (.Y (nx44540), .A0 (inputs_90__10), .A1 (inputs_91__10), .S0 (
             nx24519)) ;
    mux21_ni ix44573 (.Y (nx44572), .A0 (nx44556), .A1 (nx44568), .S0 (nx23709)
             ) ;
    mux21_ni ix44557 (.Y (nx44556), .A0 (inputs_92__10), .A1 (inputs_93__10), .S0 (
             nx24519)) ;
    mux21_ni ix44569 (.Y (nx44568), .A0 (inputs_94__10), .A1 (inputs_95__10), .S0 (
             nx24521)) ;
    mux21_ni ix44873 (.Y (nx44872), .A0 (nx44866), .A1 (nx44788), .S0 (nx23165)
             ) ;
    oai21 ix44867 (.Y (nx44866), .A0 (nx22327), .A1 (nx17643), .B0 (nx17655)) ;
    mux21 ix17644 (.Y (nx17643), .A0 (nx44830), .A1 (nx44858), .S0 (nx22973)) ;
    mux21_ni ix44831 (.Y (nx44830), .A0 (nx44814), .A1 (nx44826), .S0 (nx23709)
             ) ;
    mux21_ni ix44815 (.Y (nx44814), .A0 (inputs_100__10), .A1 (inputs_101__10), 
             .S0 (nx24521)) ;
    mux21_ni ix44827 (.Y (nx44826), .A0 (inputs_102__10), .A1 (inputs_103__10), 
             .S0 (nx24521)) ;
    mux21_ni ix44859 (.Y (nx44858), .A0 (nx44842), .A1 (nx44854), .S0 (nx23709)
             ) ;
    mux21_ni ix44843 (.Y (nx44842), .A0 (inputs_116__10), .A1 (inputs_117__10), 
             .S0 (nx24521)) ;
    mux21_ni ix44855 (.Y (nx44854), .A0 (inputs_118__10), .A1 (inputs_119__10), 
             .S0 (nx24521)) ;
    nand04 ix17656 (.Y (nx17655), .A0 (nx22327), .A1 (nx23709), .A2 (nx24521), .A3 (
           nx44802)) ;
    mux21_ni ix44803 (.Y (nx44802), .A0 (inputs_99__10), .A1 (inputs_115__10), .S0 (
             nx22973)) ;
    mux21_ni ix44789 (.Y (nx44788), .A0 (nx44724), .A1 (nx44784), .S0 (nx22975)
             ) ;
    mux21_ni ix44725 (.Y (nx44724), .A0 (nx44692), .A1 (nx44720), .S0 (nx23287)
             ) ;
    mux21_ni ix44693 (.Y (nx44692), .A0 (nx44676), .A1 (nx44688), .S0 (nx23709)
             ) ;
    mux21_ni ix44677 (.Y (nx44676), .A0 (inputs_104__10), .A1 (inputs_105__10), 
             .S0 (nx24521)) ;
    mux21_ni ix44689 (.Y (nx44688), .A0 (inputs_106__10), .A1 (inputs_107__10), 
             .S0 (nx24523)) ;
    mux21_ni ix44721 (.Y (nx44720), .A0 (nx44704), .A1 (nx44716), .S0 (nx23709)
             ) ;
    mux21_ni ix44705 (.Y (nx44704), .A0 (inputs_108__10), .A1 (inputs_109__10), 
             .S0 (nx24523)) ;
    mux21_ni ix44717 (.Y (nx44716), .A0 (inputs_110__10), .A1 (inputs_111__10), 
             .S0 (nx24523)) ;
    mux21_ni ix44785 (.Y (nx44784), .A0 (nx44752), .A1 (nx44780), .S0 (nx23289)
             ) ;
    mux21_ni ix44753 (.Y (nx44752), .A0 (nx44736), .A1 (nx44748), .S0 (nx23709)
             ) ;
    mux21_ni ix44737 (.Y (nx44736), .A0 (inputs_120__10), .A1 (inputs_121__10), 
             .S0 (nx24523)) ;
    mux21_ni ix44749 (.Y (nx44748), .A0 (inputs_122__10), .A1 (inputs_123__10), 
             .S0 (nx24523)) ;
    mux21_ni ix44781 (.Y (nx44780), .A0 (nx44764), .A1 (nx44776), .S0 (nx23711)
             ) ;
    mux21_ni ix44765 (.Y (nx44764), .A0 (inputs_124__10), .A1 (inputs_125__10), 
             .S0 (nx24523)) ;
    mux21_ni ix44777 (.Y (nx44776), .A0 (inputs_126__10), .A1 (inputs_127__10), 
             .S0 (nx24523)) ;
    mux21_ni ix45725 (.Y (nx45724), .A0 (nx45300), .A1 (nx45720), .S0 (nx22501)
             ) ;
    mux21_ni ix45301 (.Y (nx45300), .A0 (nx45088), .A1 (nx45296), .S0 (nx22627)
             ) ;
    mux21_ni ix45089 (.Y (nx45088), .A0 (nx45082), .A1 (nx45004), .S0 (nx23165)
             ) ;
    oai21 ix45083 (.Y (nx45082), .A0 (nx22327), .A1 (nx17691), .B0 (nx17701)) ;
    mux21 ix17692 (.Y (nx17691), .A0 (nx45046), .A1 (nx45074), .S0 (nx22975)) ;
    mux21_ni ix45047 (.Y (nx45046), .A0 (nx45030), .A1 (nx45042), .S0 (nx23711)
             ) ;
    mux21_ni ix45031 (.Y (nx45030), .A0 (inputs_132__10), .A1 (inputs_133__10), 
             .S0 (nx24525)) ;
    mux21_ni ix45043 (.Y (nx45042), .A0 (inputs_134__10), .A1 (inputs_135__10), 
             .S0 (nx24525)) ;
    mux21_ni ix45075 (.Y (nx45074), .A0 (nx45058), .A1 (nx45070), .S0 (nx23711)
             ) ;
    mux21_ni ix45059 (.Y (nx45058), .A0 (inputs_148__10), .A1 (inputs_149__10), 
             .S0 (nx24525)) ;
    mux21_ni ix45071 (.Y (nx45070), .A0 (inputs_150__10), .A1 (inputs_151__10), 
             .S0 (nx24525)) ;
    nand04 ix17702 (.Y (nx17701), .A0 (nx22327), .A1 (nx23711), .A2 (nx24525), .A3 (
           nx45018)) ;
    mux21_ni ix45019 (.Y (nx45018), .A0 (inputs_131__10), .A1 (inputs_147__10), 
             .S0 (nx22975)) ;
    mux21_ni ix45005 (.Y (nx45004), .A0 (nx44940), .A1 (nx45000), .S0 (nx22975)
             ) ;
    mux21_ni ix44941 (.Y (nx44940), .A0 (nx44908), .A1 (nx44936), .S0 (nx23289)
             ) ;
    mux21_ni ix44909 (.Y (nx44908), .A0 (nx44892), .A1 (nx44904), .S0 (nx23711)
             ) ;
    mux21_ni ix44893 (.Y (nx44892), .A0 (inputs_136__10), .A1 (inputs_137__10), 
             .S0 (nx24525)) ;
    mux21_ni ix44905 (.Y (nx44904), .A0 (inputs_138__10), .A1 (inputs_139__10), 
             .S0 (nx24525)) ;
    mux21_ni ix44937 (.Y (nx44936), .A0 (nx44920), .A1 (nx44932), .S0 (nx23711)
             ) ;
    mux21_ni ix44921 (.Y (nx44920), .A0 (inputs_140__10), .A1 (inputs_141__10), 
             .S0 (nx24527)) ;
    mux21_ni ix44933 (.Y (nx44932), .A0 (inputs_142__10), .A1 (inputs_143__10), 
             .S0 (nx24527)) ;
    mux21_ni ix45001 (.Y (nx45000), .A0 (nx44968), .A1 (nx44996), .S0 (nx23289)
             ) ;
    mux21_ni ix44969 (.Y (nx44968), .A0 (nx44952), .A1 (nx44964), .S0 (nx23711)
             ) ;
    mux21_ni ix44953 (.Y (nx44952), .A0 (inputs_152__10), .A1 (inputs_153__10), 
             .S0 (nx24527)) ;
    mux21_ni ix44965 (.Y (nx44964), .A0 (inputs_154__10), .A1 (inputs_155__10), 
             .S0 (nx24527)) ;
    mux21_ni ix44997 (.Y (nx44996), .A0 (nx44980), .A1 (nx44992), .S0 (nx23713)
             ) ;
    mux21_ni ix44981 (.Y (nx44980), .A0 (inputs_156__10), .A1 (inputs_157__10), 
             .S0 (nx24527)) ;
    mux21_ni ix44993 (.Y (nx44992), .A0 (inputs_158__10), .A1 (inputs_159__10), 
             .S0 (nx24527)) ;
    mux21_ni ix45297 (.Y (nx45296), .A0 (nx45290), .A1 (nx45212), .S0 (nx23165)
             ) ;
    oai21 ix45291 (.Y (nx45290), .A0 (nx22329), .A1 (nx17731), .B0 (nx17743)) ;
    mux21 ix17732 (.Y (nx17731), .A0 (nx45254), .A1 (nx45282), .S0 (nx22975)) ;
    mux21_ni ix45255 (.Y (nx45254), .A0 (nx45238), .A1 (nx45250), .S0 (nx23713)
             ) ;
    mux21_ni ix45239 (.Y (nx45238), .A0 (inputs_164__10), .A1 (inputs_165__10), 
             .S0 (nx24527)) ;
    mux21_ni ix45251 (.Y (nx45250), .A0 (inputs_166__10), .A1 (inputs_167__10), 
             .S0 (nx24529)) ;
    mux21_ni ix45283 (.Y (nx45282), .A0 (nx45266), .A1 (nx45278), .S0 (nx23713)
             ) ;
    mux21_ni ix45267 (.Y (nx45266), .A0 (inputs_180__10), .A1 (inputs_181__10), 
             .S0 (nx24529)) ;
    mux21_ni ix45279 (.Y (nx45278), .A0 (inputs_182__10), .A1 (inputs_183__10), 
             .S0 (nx24529)) ;
    nand04 ix17744 (.Y (nx17743), .A0 (nx22329), .A1 (nx23713), .A2 (nx24529), .A3 (
           nx45226)) ;
    mux21_ni ix45227 (.Y (nx45226), .A0 (inputs_163__10), .A1 (inputs_179__10), 
             .S0 (nx22975)) ;
    mux21_ni ix45213 (.Y (nx45212), .A0 (nx45148), .A1 (nx45208), .S0 (nx22975)
             ) ;
    mux21_ni ix45149 (.Y (nx45148), .A0 (nx45116), .A1 (nx45144), .S0 (nx23289)
             ) ;
    mux21_ni ix45117 (.Y (nx45116), .A0 (nx45100), .A1 (nx45112), .S0 (nx23713)
             ) ;
    mux21_ni ix45101 (.Y (nx45100), .A0 (inputs_168__10), .A1 (inputs_169__10), 
             .S0 (nx24529)) ;
    mux21_ni ix45113 (.Y (nx45112), .A0 (inputs_170__10), .A1 (inputs_171__10), 
             .S0 (nx24529)) ;
    mux21_ni ix45145 (.Y (nx45144), .A0 (nx45128), .A1 (nx45140), .S0 (nx23713)
             ) ;
    mux21_ni ix45129 (.Y (nx45128), .A0 (inputs_172__10), .A1 (inputs_173__10), 
             .S0 (nx24529)) ;
    mux21_ni ix45141 (.Y (nx45140), .A0 (inputs_174__10), .A1 (inputs_175__10), 
             .S0 (nx24531)) ;
    mux21_ni ix45209 (.Y (nx45208), .A0 (nx45176), .A1 (nx45204), .S0 (nx23289)
             ) ;
    mux21_ni ix45177 (.Y (nx45176), .A0 (nx45160), .A1 (nx45172), .S0 (nx23713)
             ) ;
    mux21_ni ix45161 (.Y (nx45160), .A0 (inputs_184__10), .A1 (inputs_185__10), 
             .S0 (nx24531)) ;
    mux21_ni ix45173 (.Y (nx45172), .A0 (inputs_186__10), .A1 (inputs_187__10), 
             .S0 (nx24531)) ;
    mux21_ni ix45205 (.Y (nx45204), .A0 (nx45188), .A1 (nx45200), .S0 (nx23715)
             ) ;
    mux21_ni ix45189 (.Y (nx45188), .A0 (inputs_188__10), .A1 (inputs_189__10), 
             .S0 (nx24531)) ;
    mux21_ni ix45201 (.Y (nx45200), .A0 (inputs_190__10), .A1 (inputs_191__10), 
             .S0 (nx24531)) ;
    mux21_ni ix45721 (.Y (nx45720), .A0 (nx45508), .A1 (nx45716), .S0 (nx22627)
             ) ;
    mux21_ni ix45509 (.Y (nx45508), .A0 (nx45502), .A1 (nx45424), .S0 (nx23165)
             ) ;
    oai21 ix45503 (.Y (nx45502), .A0 (nx22329), .A1 (nx17775), .B0 (nx17787)) ;
    mux21 ix17776 (.Y (nx17775), .A0 (nx45466), .A1 (nx45494), .S0 (nx22977)) ;
    mux21_ni ix45467 (.Y (nx45466), .A0 (nx45450), .A1 (nx45462), .S0 (nx23715)
             ) ;
    mux21_ni ix45451 (.Y (nx45450), .A0 (inputs_196__10), .A1 (inputs_197__10), 
             .S0 (nx24531)) ;
    mux21_ni ix45463 (.Y (nx45462), .A0 (inputs_198__10), .A1 (inputs_199__10), 
             .S0 (nx24531)) ;
    mux21_ni ix45495 (.Y (nx45494), .A0 (nx45478), .A1 (nx45490), .S0 (nx23715)
             ) ;
    mux21_ni ix45479 (.Y (nx45478), .A0 (inputs_212__10), .A1 (inputs_213__10), 
             .S0 (nx24533)) ;
    mux21_ni ix45491 (.Y (nx45490), .A0 (inputs_214__10), .A1 (inputs_215__10), 
             .S0 (nx24533)) ;
    nand04 ix17788 (.Y (nx17787), .A0 (nx22329), .A1 (nx23715), .A2 (nx24533), .A3 (
           nx45438)) ;
    mux21_ni ix45439 (.Y (nx45438), .A0 (inputs_195__10), .A1 (inputs_211__10), 
             .S0 (nx22977)) ;
    mux21_ni ix45425 (.Y (nx45424), .A0 (nx45360), .A1 (nx45420), .S0 (nx22977)
             ) ;
    mux21_ni ix45361 (.Y (nx45360), .A0 (nx45328), .A1 (nx45356), .S0 (nx23289)
             ) ;
    mux21_ni ix45329 (.Y (nx45328), .A0 (nx45312), .A1 (nx45324), .S0 (nx23715)
             ) ;
    mux21_ni ix45313 (.Y (nx45312), .A0 (inputs_200__10), .A1 (inputs_201__10), 
             .S0 (nx24533)) ;
    mux21_ni ix45325 (.Y (nx45324), .A0 (inputs_202__10), .A1 (inputs_203__10), 
             .S0 (nx24533)) ;
    mux21_ni ix45357 (.Y (nx45356), .A0 (nx45340), .A1 (nx45352), .S0 (nx23715)
             ) ;
    mux21_ni ix45341 (.Y (nx45340), .A0 (inputs_204__10), .A1 (inputs_205__10), 
             .S0 (nx24533)) ;
    mux21_ni ix45353 (.Y (nx45352), .A0 (inputs_206__10), .A1 (inputs_207__10), 
             .S0 (nx24533)) ;
    mux21_ni ix45421 (.Y (nx45420), .A0 (nx45388), .A1 (nx45416), .S0 (nx23289)
             ) ;
    mux21_ni ix45389 (.Y (nx45388), .A0 (nx45372), .A1 (nx45384), .S0 (nx23715)
             ) ;
    mux21_ni ix45373 (.Y (nx45372), .A0 (inputs_216__10), .A1 (inputs_217__10), 
             .S0 (nx24535)) ;
    mux21_ni ix45385 (.Y (nx45384), .A0 (inputs_218__10), .A1 (inputs_219__10), 
             .S0 (nx24535)) ;
    mux21_ni ix45417 (.Y (nx45416), .A0 (nx45400), .A1 (nx45412), .S0 (nx23717)
             ) ;
    mux21_ni ix45401 (.Y (nx45400), .A0 (inputs_220__10), .A1 (inputs_221__10), 
             .S0 (nx24535)) ;
    mux21_ni ix45413 (.Y (nx45412), .A0 (inputs_222__10), .A1 (inputs_223__10), 
             .S0 (nx24535)) ;
    mux21_ni ix45717 (.Y (nx45716), .A0 (nx45710), .A1 (nx45632), .S0 (nx23167)
             ) ;
    oai21 ix45711 (.Y (nx45710), .A0 (nx22329), .A1 (nx17821), .B0 (nx17833)) ;
    mux21 ix17822 (.Y (nx17821), .A0 (nx45674), .A1 (nx45702), .S0 (nx22977)) ;
    mux21_ni ix45675 (.Y (nx45674), .A0 (nx45658), .A1 (nx45670), .S0 (nx23717)
             ) ;
    mux21_ni ix45659 (.Y (nx45658), .A0 (inputs_228__10), .A1 (inputs_229__10), 
             .S0 (nx24535)) ;
    mux21_ni ix45671 (.Y (nx45670), .A0 (inputs_230__10), .A1 (inputs_231__10), 
             .S0 (nx24535)) ;
    mux21_ni ix45703 (.Y (nx45702), .A0 (nx45686), .A1 (nx45698), .S0 (nx23717)
             ) ;
    mux21_ni ix45687 (.Y (nx45686), .A0 (inputs_244__10), .A1 (inputs_245__10), 
             .S0 (nx24535)) ;
    mux21_ni ix45699 (.Y (nx45698), .A0 (inputs_246__10), .A1 (inputs_247__10), 
             .S0 (nx24537)) ;
    nand04 ix17834 (.Y (nx17833), .A0 (nx22329), .A1 (nx23717), .A2 (nx24537), .A3 (
           nx45646)) ;
    mux21_ni ix45647 (.Y (nx45646), .A0 (inputs_227__10), .A1 (inputs_243__10), 
             .S0 (nx22977)) ;
    mux21_ni ix45633 (.Y (nx45632), .A0 (nx45568), .A1 (nx45628), .S0 (nx22977)
             ) ;
    mux21_ni ix45569 (.Y (nx45568), .A0 (nx45536), .A1 (nx45564), .S0 (nx23291)
             ) ;
    mux21_ni ix45537 (.Y (nx45536), .A0 (nx45520), .A1 (nx45532), .S0 (nx23717)
             ) ;
    mux21_ni ix45521 (.Y (nx45520), .A0 (inputs_232__10), .A1 (inputs_233__10), 
             .S0 (nx24537)) ;
    mux21_ni ix45533 (.Y (nx45532), .A0 (inputs_234__10), .A1 (inputs_235__10), 
             .S0 (nx24537)) ;
    mux21_ni ix45565 (.Y (nx45564), .A0 (nx45548), .A1 (nx45560), .S0 (nx23717)
             ) ;
    mux21_ni ix45549 (.Y (nx45548), .A0 (inputs_236__10), .A1 (inputs_237__10), 
             .S0 (nx24537)) ;
    mux21_ni ix45561 (.Y (nx45560), .A0 (inputs_238__10), .A1 (inputs_239__10), 
             .S0 (nx24537)) ;
    mux21_ni ix45629 (.Y (nx45628), .A0 (nx45596), .A1 (nx45624), .S0 (nx23291)
             ) ;
    mux21_ni ix45597 (.Y (nx45596), .A0 (nx45580), .A1 (nx45592), .S0 (nx23717)
             ) ;
    mux21_ni ix45581 (.Y (nx45580), .A0 (inputs_248__10), .A1 (inputs_249__10), 
             .S0 (nx24537)) ;
    mux21_ni ix45593 (.Y (nx45592), .A0 (inputs_250__10), .A1 (inputs_251__10), 
             .S0 (nx24539)) ;
    mux21_ni ix45625 (.Y (nx45624), .A0 (nx45608), .A1 (nx45620), .S0 (nx23719)
             ) ;
    mux21_ni ix45609 (.Y (nx45608), .A0 (inputs_252__10), .A1 (inputs_253__10), 
             .S0 (nx24539)) ;
    mux21_ni ix45621 (.Y (nx45620), .A0 (inputs_254__10), .A1 (inputs_255__10), 
             .S0 (nx24539)) ;
    oai21 ix49895 (.Y (\output [11]), .A0 (nx22223), .A1 (nx17861), .B0 (nx18219
          )) ;
    mux21 ix17862 (.Y (nx17861), .A0 (nx46576), .A1 (nx47420), .S0 (nx22435)) ;
    mux21_ni ix46577 (.Y (nx46576), .A0 (nx46152), .A1 (nx46572), .S0 (nx22501)
             ) ;
    mux21_ni ix46153 (.Y (nx46152), .A0 (nx45940), .A1 (nx46148), .S0 (nx22627)
             ) ;
    mux21_ni ix45941 (.Y (nx45940), .A0 (nx45934), .A1 (nx45856), .S0 (nx23167)
             ) ;
    oai21 ix45935 (.Y (nx45934), .A0 (nx22329), .A1 (nx17869), .B0 (nx17883)) ;
    mux21 ix17870 (.Y (nx17869), .A0 (nx45898), .A1 (nx45926), .S0 (nx22977)) ;
    mux21_ni ix45899 (.Y (nx45898), .A0 (nx45882), .A1 (nx45894), .S0 (nx23719)
             ) ;
    mux21_ni ix45883 (.Y (nx45882), .A0 (inputs_260__11), .A1 (inputs_261__11), 
             .S0 (nx24539)) ;
    mux21_ni ix45895 (.Y (nx45894), .A0 (inputs_262__11), .A1 (inputs_263__11), 
             .S0 (nx24539)) ;
    mux21_ni ix45927 (.Y (nx45926), .A0 (nx45910), .A1 (nx45922), .S0 (nx23719)
             ) ;
    mux21_ni ix45911 (.Y (nx45910), .A0 (inputs_276__11), .A1 (inputs_277__11), 
             .S0 (nx24539)) ;
    mux21_ni ix45923 (.Y (nx45922), .A0 (inputs_278__11), .A1 (inputs_279__11), 
             .S0 (nx24539)) ;
    nand04 ix17884 (.Y (nx17883), .A0 (nx22331), .A1 (nx23719), .A2 (nx24541), .A3 (
           nx45870)) ;
    mux21_ni ix45871 (.Y (nx45870), .A0 (inputs_259__11), .A1 (inputs_275__11), 
             .S0 (nx22979)) ;
    mux21_ni ix45857 (.Y (nx45856), .A0 (nx45792), .A1 (nx45852), .S0 (nx22979)
             ) ;
    mux21_ni ix45793 (.Y (nx45792), .A0 (nx45760), .A1 (nx45788), .S0 (nx23291)
             ) ;
    mux21_ni ix45761 (.Y (nx45760), .A0 (nx45744), .A1 (nx45756), .S0 (nx23719)
             ) ;
    mux21_ni ix45745 (.Y (nx45744), .A0 (inputs_264__11), .A1 (inputs_265__11), 
             .S0 (nx24541)) ;
    mux21_ni ix45757 (.Y (nx45756), .A0 (inputs_266__11), .A1 (inputs_267__11), 
             .S0 (nx24541)) ;
    mux21_ni ix45789 (.Y (nx45788), .A0 (nx45772), .A1 (nx45784), .S0 (nx23719)
             ) ;
    mux21_ni ix45773 (.Y (nx45772), .A0 (inputs_268__11), .A1 (inputs_269__11), 
             .S0 (nx24541)) ;
    mux21_ni ix45785 (.Y (nx45784), .A0 (inputs_270__11), .A1 (inputs_271__11), 
             .S0 (nx24541)) ;
    mux21_ni ix45853 (.Y (nx45852), .A0 (nx45820), .A1 (nx45848), .S0 (nx23291)
             ) ;
    mux21_ni ix45821 (.Y (nx45820), .A0 (nx45804), .A1 (nx45816), .S0 (nx23719)
             ) ;
    mux21_ni ix45805 (.Y (nx45804), .A0 (inputs_280__11), .A1 (inputs_281__11), 
             .S0 (nx24541)) ;
    mux21_ni ix45817 (.Y (nx45816), .A0 (inputs_282__11), .A1 (inputs_283__11), 
             .S0 (nx24541)) ;
    mux21_ni ix45849 (.Y (nx45848), .A0 (nx45832), .A1 (nx45844), .S0 (nx23721)
             ) ;
    mux21_ni ix45833 (.Y (nx45832), .A0 (inputs_284__11), .A1 (inputs_285__11), 
             .S0 (nx24543)) ;
    mux21_ni ix45845 (.Y (nx45844), .A0 (inputs_286__11), .A1 (inputs_287__11), 
             .S0 (nx24543)) ;
    mux21_ni ix46149 (.Y (nx46148), .A0 (nx46142), .A1 (nx46064), .S0 (nx23167)
             ) ;
    oai21 ix46143 (.Y (nx46142), .A0 (nx22331), .A1 (nx17913), .B0 (nx17925)) ;
    mux21 ix17914 (.Y (nx17913), .A0 (nx46106), .A1 (nx46134), .S0 (nx22979)) ;
    mux21_ni ix46107 (.Y (nx46106), .A0 (nx46090), .A1 (nx46102), .S0 (nx23721)
             ) ;
    mux21_ni ix46091 (.Y (nx46090), .A0 (inputs_292__11), .A1 (inputs_293__11), 
             .S0 (nx24543)) ;
    mux21_ni ix46103 (.Y (nx46102), .A0 (inputs_294__11), .A1 (inputs_295__11), 
             .S0 (nx24543)) ;
    mux21_ni ix46135 (.Y (nx46134), .A0 (nx46118), .A1 (nx46130), .S0 (nx23721)
             ) ;
    mux21_ni ix46119 (.Y (nx46118), .A0 (inputs_308__11), .A1 (inputs_309__11), 
             .S0 (nx24543)) ;
    mux21_ni ix46131 (.Y (nx46130), .A0 (inputs_310__11), .A1 (inputs_311__11), 
             .S0 (nx24543)) ;
    nand04 ix17926 (.Y (nx17925), .A0 (nx22331), .A1 (nx23721), .A2 (nx24543), .A3 (
           nx46078)) ;
    mux21_ni ix46079 (.Y (nx46078), .A0 (inputs_291__11), .A1 (inputs_307__11), 
             .S0 (nx22979)) ;
    mux21_ni ix46065 (.Y (nx46064), .A0 (nx46000), .A1 (nx46060), .S0 (nx22979)
             ) ;
    mux21_ni ix46001 (.Y (nx46000), .A0 (nx45968), .A1 (nx45996), .S0 (nx23291)
             ) ;
    mux21_ni ix45969 (.Y (nx45968), .A0 (nx45952), .A1 (nx45964), .S0 (nx23721)
             ) ;
    mux21_ni ix45953 (.Y (nx45952), .A0 (inputs_296__11), .A1 (inputs_297__11), 
             .S0 (nx24545)) ;
    mux21_ni ix45965 (.Y (nx45964), .A0 (inputs_298__11), .A1 (inputs_299__11), 
             .S0 (nx24545)) ;
    mux21_ni ix45997 (.Y (nx45996), .A0 (nx45980), .A1 (nx45992), .S0 (nx23721)
             ) ;
    mux21_ni ix45981 (.Y (nx45980), .A0 (inputs_300__11), .A1 (inputs_301__11), 
             .S0 (nx24545)) ;
    mux21_ni ix45993 (.Y (nx45992), .A0 (inputs_302__11), .A1 (inputs_303__11), 
             .S0 (nx24545)) ;
    mux21_ni ix46061 (.Y (nx46060), .A0 (nx46028), .A1 (nx46056), .S0 (nx23291)
             ) ;
    mux21_ni ix46029 (.Y (nx46028), .A0 (nx46012), .A1 (nx46024), .S0 (nx23721)
             ) ;
    mux21_ni ix46013 (.Y (nx46012), .A0 (inputs_312__11), .A1 (inputs_313__11), 
             .S0 (nx24545)) ;
    mux21_ni ix46025 (.Y (nx46024), .A0 (inputs_314__11), .A1 (inputs_315__11), 
             .S0 (nx24545)) ;
    mux21_ni ix46057 (.Y (nx46056), .A0 (nx46040), .A1 (nx46052), .S0 (nx23723)
             ) ;
    mux21_ni ix46041 (.Y (nx46040), .A0 (inputs_316__11), .A1 (inputs_317__11), 
             .S0 (nx24545)) ;
    mux21_ni ix46053 (.Y (nx46052), .A0 (inputs_318__11), .A1 (inputs_319__11), 
             .S0 (nx24547)) ;
    mux21_ni ix46573 (.Y (nx46572), .A0 (nx46360), .A1 (nx46568), .S0 (nx22627)
             ) ;
    mux21_ni ix46361 (.Y (nx46360), .A0 (nx46354), .A1 (nx46276), .S0 (nx23167)
             ) ;
    oai21 ix46355 (.Y (nx46354), .A0 (nx22331), .A1 (nx17959), .B0 (nx17971)) ;
    mux21 ix17960 (.Y (nx17959), .A0 (nx46318), .A1 (nx46346), .S0 (nx22979)) ;
    mux21_ni ix46319 (.Y (nx46318), .A0 (nx46302), .A1 (nx46314), .S0 (nx23723)
             ) ;
    mux21_ni ix46303 (.Y (nx46302), .A0 (inputs_324__11), .A1 (inputs_325__11), 
             .S0 (nx24547)) ;
    mux21_ni ix46315 (.Y (nx46314), .A0 (inputs_326__11), .A1 (inputs_327__11), 
             .S0 (nx24547)) ;
    mux21_ni ix46347 (.Y (nx46346), .A0 (nx46330), .A1 (nx46342), .S0 (nx23723)
             ) ;
    mux21_ni ix46331 (.Y (nx46330), .A0 (inputs_340__11), .A1 (inputs_341__11), 
             .S0 (nx24547)) ;
    mux21_ni ix46343 (.Y (nx46342), .A0 (inputs_342__11), .A1 (inputs_343__11), 
             .S0 (nx24547)) ;
    nand04 ix17972 (.Y (nx17971), .A0 (nx22331), .A1 (nx23723), .A2 (nx24547), .A3 (
           nx46290)) ;
    mux21_ni ix46291 (.Y (nx46290), .A0 (inputs_323__11), .A1 (inputs_339__11), 
             .S0 (nx22979)) ;
    mux21_ni ix46277 (.Y (nx46276), .A0 (nx46212), .A1 (nx46272), .S0 (nx22981)
             ) ;
    mux21_ni ix46213 (.Y (nx46212), .A0 (nx46180), .A1 (nx46208), .S0 (nx23291)
             ) ;
    mux21_ni ix46181 (.Y (nx46180), .A0 (nx46164), .A1 (nx46176), .S0 (nx23723)
             ) ;
    mux21_ni ix46165 (.Y (nx46164), .A0 (inputs_328__11), .A1 (inputs_329__11), 
             .S0 (nx24547)) ;
    mux21_ni ix46177 (.Y (nx46176), .A0 (inputs_330__11), .A1 (inputs_331__11), 
             .S0 (nx24549)) ;
    mux21_ni ix46209 (.Y (nx46208), .A0 (nx46192), .A1 (nx46204), .S0 (nx23723)
             ) ;
    mux21_ni ix46193 (.Y (nx46192), .A0 (inputs_332__11), .A1 (inputs_333__11), 
             .S0 (nx24549)) ;
    mux21_ni ix46205 (.Y (nx46204), .A0 (inputs_334__11), .A1 (inputs_335__11), 
             .S0 (nx24549)) ;
    mux21_ni ix46273 (.Y (nx46272), .A0 (nx46240), .A1 (nx46268), .S0 (nx23293)
             ) ;
    mux21_ni ix46241 (.Y (nx46240), .A0 (nx46224), .A1 (nx46236), .S0 (nx23723)
             ) ;
    mux21_ni ix46225 (.Y (nx46224), .A0 (inputs_344__11), .A1 (inputs_345__11), 
             .S0 (nx24549)) ;
    mux21_ni ix46237 (.Y (nx46236), .A0 (inputs_346__11), .A1 (inputs_347__11), 
             .S0 (nx24549)) ;
    mux21_ni ix46269 (.Y (nx46268), .A0 (nx46252), .A1 (nx46264), .S0 (nx23725)
             ) ;
    mux21_ni ix46253 (.Y (nx46252), .A0 (inputs_348__11), .A1 (inputs_349__11), 
             .S0 (nx24549)) ;
    mux21_ni ix46265 (.Y (nx46264), .A0 (inputs_350__11), .A1 (inputs_351__11), 
             .S0 (nx24549)) ;
    mux21_ni ix46569 (.Y (nx46568), .A0 (nx46562), .A1 (nx46484), .S0 (nx23167)
             ) ;
    oai21 ix46563 (.Y (nx46562), .A0 (nx22331), .A1 (nx18001), .B0 (nx18015)) ;
    mux21 ix18002 (.Y (nx18001), .A0 (nx46526), .A1 (nx46554), .S0 (nx22981)) ;
    mux21_ni ix46527 (.Y (nx46526), .A0 (nx46510), .A1 (nx46522), .S0 (nx23725)
             ) ;
    mux21_ni ix46511 (.Y (nx46510), .A0 (inputs_356__11), .A1 (inputs_357__11), 
             .S0 (nx24551)) ;
    mux21_ni ix46523 (.Y (nx46522), .A0 (inputs_358__11), .A1 (inputs_359__11), 
             .S0 (nx24551)) ;
    mux21_ni ix46555 (.Y (nx46554), .A0 (nx46538), .A1 (nx46550), .S0 (nx23725)
             ) ;
    mux21_ni ix46539 (.Y (nx46538), .A0 (inputs_372__11), .A1 (inputs_373__11), 
             .S0 (nx24551)) ;
    mux21_ni ix46551 (.Y (nx46550), .A0 (inputs_374__11), .A1 (inputs_375__11), 
             .S0 (nx24551)) ;
    nand04 ix18016 (.Y (nx18015), .A0 (nx22331), .A1 (nx23725), .A2 (nx24551), .A3 (
           nx46498)) ;
    mux21_ni ix46499 (.Y (nx46498), .A0 (inputs_355__11), .A1 (inputs_371__11), 
             .S0 (nx22981)) ;
    mux21_ni ix46485 (.Y (nx46484), .A0 (nx46420), .A1 (nx46480), .S0 (nx22981)
             ) ;
    mux21_ni ix46421 (.Y (nx46420), .A0 (nx46388), .A1 (nx46416), .S0 (nx23293)
             ) ;
    mux21_ni ix46389 (.Y (nx46388), .A0 (nx46372), .A1 (nx46384), .S0 (nx23725)
             ) ;
    mux21_ni ix46373 (.Y (nx46372), .A0 (inputs_360__11), .A1 (inputs_361__11), 
             .S0 (nx24551)) ;
    mux21_ni ix46385 (.Y (nx46384), .A0 (inputs_362__11), .A1 (inputs_363__11), 
             .S0 (nx24551)) ;
    mux21_ni ix46417 (.Y (nx46416), .A0 (nx46400), .A1 (nx46412), .S0 (nx23725)
             ) ;
    mux21_ni ix46401 (.Y (nx46400), .A0 (inputs_364__11), .A1 (inputs_365__11), 
             .S0 (nx24553)) ;
    mux21_ni ix46413 (.Y (nx46412), .A0 (inputs_366__11), .A1 (inputs_367__11), 
             .S0 (nx24553)) ;
    mux21_ni ix46481 (.Y (nx46480), .A0 (nx46448), .A1 (nx46476), .S0 (nx23293)
             ) ;
    mux21_ni ix46449 (.Y (nx46448), .A0 (nx46432), .A1 (nx46444), .S0 (nx23725)
             ) ;
    mux21_ni ix46433 (.Y (nx46432), .A0 (inputs_376__11), .A1 (inputs_377__11), 
             .S0 (nx24553)) ;
    mux21_ni ix46445 (.Y (nx46444), .A0 (inputs_378__11), .A1 (inputs_379__11), 
             .S0 (nx24553)) ;
    mux21_ni ix46477 (.Y (nx46476), .A0 (nx46460), .A1 (nx46472), .S0 (nx23727)
             ) ;
    mux21_ni ix46461 (.Y (nx46460), .A0 (inputs_380__11), .A1 (inputs_381__11), 
             .S0 (nx24553)) ;
    mux21_ni ix46473 (.Y (nx46472), .A0 (inputs_382__11), .A1 (inputs_383__11), 
             .S0 (nx24553)) ;
    mux21_ni ix47421 (.Y (nx47420), .A0 (nx46996), .A1 (nx47416), .S0 (nx22501)
             ) ;
    mux21_ni ix46997 (.Y (nx46996), .A0 (nx46784), .A1 (nx46992), .S0 (nx22627)
             ) ;
    mux21_ni ix46785 (.Y (nx46784), .A0 (nx46778), .A1 (nx46700), .S0 (nx23167)
             ) ;
    oai21 ix46779 (.Y (nx46778), .A0 (nx22333), .A1 (nx18049), .B0 (nx18061)) ;
    mux21 ix18050 (.Y (nx18049), .A0 (nx46742), .A1 (nx46770), .S0 (nx22981)) ;
    mux21_ni ix46743 (.Y (nx46742), .A0 (nx46726), .A1 (nx46738), .S0 (nx23727)
             ) ;
    mux21_ni ix46727 (.Y (nx46726), .A0 (inputs_388__11), .A1 (inputs_389__11), 
             .S0 (nx24553)) ;
    mux21_ni ix46739 (.Y (nx46738), .A0 (inputs_390__11), .A1 (inputs_391__11), 
             .S0 (nx24555)) ;
    mux21_ni ix46771 (.Y (nx46770), .A0 (nx46754), .A1 (nx46766), .S0 (nx23727)
             ) ;
    mux21_ni ix46755 (.Y (nx46754), .A0 (inputs_404__11), .A1 (inputs_405__11), 
             .S0 (nx24555)) ;
    mux21_ni ix46767 (.Y (nx46766), .A0 (inputs_406__11), .A1 (inputs_407__11), 
             .S0 (nx24555)) ;
    nand04 ix18062 (.Y (nx18061), .A0 (nx22333), .A1 (nx23727), .A2 (nx24555), .A3 (
           nx46714)) ;
    mux21_ni ix46715 (.Y (nx46714), .A0 (inputs_387__11), .A1 (inputs_403__11), 
             .S0 (nx22981)) ;
    mux21_ni ix46701 (.Y (nx46700), .A0 (nx46636), .A1 (nx46696), .S0 (nx22981)
             ) ;
    mux21_ni ix46637 (.Y (nx46636), .A0 (nx46604), .A1 (nx46632), .S0 (nx23293)
             ) ;
    mux21_ni ix46605 (.Y (nx46604), .A0 (nx46588), .A1 (nx46600), .S0 (nx23727)
             ) ;
    mux21_ni ix46589 (.Y (nx46588), .A0 (inputs_392__11), .A1 (inputs_393__11), 
             .S0 (nx24555)) ;
    mux21_ni ix46601 (.Y (nx46600), .A0 (inputs_394__11), .A1 (inputs_395__11), 
             .S0 (nx24555)) ;
    mux21_ni ix46633 (.Y (nx46632), .A0 (nx46616), .A1 (nx46628), .S0 (nx23727)
             ) ;
    mux21_ni ix46617 (.Y (nx46616), .A0 (inputs_396__11), .A1 (inputs_397__11), 
             .S0 (nx24555)) ;
    mux21_ni ix46629 (.Y (nx46628), .A0 (inputs_398__11), .A1 (inputs_399__11), 
             .S0 (nx24557)) ;
    mux21_ni ix46697 (.Y (nx46696), .A0 (nx46664), .A1 (nx46692), .S0 (nx23293)
             ) ;
    mux21_ni ix46665 (.Y (nx46664), .A0 (nx46648), .A1 (nx46660), .S0 (nx23727)
             ) ;
    mux21_ni ix46649 (.Y (nx46648), .A0 (inputs_408__11), .A1 (inputs_409__11), 
             .S0 (nx24557)) ;
    mux21_ni ix46661 (.Y (nx46660), .A0 (inputs_410__11), .A1 (inputs_411__11), 
             .S0 (nx24557)) ;
    mux21_ni ix46693 (.Y (nx46692), .A0 (nx46676), .A1 (nx46688), .S0 (nx23729)
             ) ;
    mux21_ni ix46677 (.Y (nx46676), .A0 (inputs_412__11), .A1 (inputs_413__11), 
             .S0 (nx24557)) ;
    mux21_ni ix46689 (.Y (nx46688), .A0 (inputs_414__11), .A1 (inputs_415__11), 
             .S0 (nx24557)) ;
    mux21_ni ix46993 (.Y (nx46992), .A0 (nx46986), .A1 (nx46908), .S0 (nx23167)
             ) ;
    oai21 ix46987 (.Y (nx46986), .A0 (nx22333), .A1 (nx18093), .B0 (nx18103)) ;
    mux21 ix18094 (.Y (nx18093), .A0 (nx46950), .A1 (nx46978), .S0 (nx22983)) ;
    mux21_ni ix46951 (.Y (nx46950), .A0 (nx46934), .A1 (nx46946), .S0 (nx23729)
             ) ;
    mux21_ni ix46935 (.Y (nx46934), .A0 (inputs_420__11), .A1 (inputs_421__11), 
             .S0 (nx24557)) ;
    mux21_ni ix46947 (.Y (nx46946), .A0 (inputs_422__11), .A1 (inputs_423__11), 
             .S0 (nx24557)) ;
    mux21_ni ix46979 (.Y (nx46978), .A0 (nx46962), .A1 (nx46974), .S0 (nx23729)
             ) ;
    mux21_ni ix46963 (.Y (nx46962), .A0 (inputs_436__11), .A1 (inputs_437__11), 
             .S0 (nx24559)) ;
    mux21_ni ix46975 (.Y (nx46974), .A0 (inputs_438__11), .A1 (inputs_439__11), 
             .S0 (nx24559)) ;
    nand04 ix18104 (.Y (nx18103), .A0 (nx22333), .A1 (nx23729), .A2 (nx24559), .A3 (
           nx46922)) ;
    mux21_ni ix46923 (.Y (nx46922), .A0 (inputs_419__11), .A1 (inputs_435__11), 
             .S0 (nx22983)) ;
    mux21_ni ix46909 (.Y (nx46908), .A0 (nx46844), .A1 (nx46904), .S0 (nx22983)
             ) ;
    mux21_ni ix46845 (.Y (nx46844), .A0 (nx46812), .A1 (nx46840), .S0 (nx23293)
             ) ;
    mux21_ni ix46813 (.Y (nx46812), .A0 (nx46796), .A1 (nx46808), .S0 (nx23729)
             ) ;
    mux21_ni ix46797 (.Y (nx46796), .A0 (inputs_424__11), .A1 (inputs_425__11), 
             .S0 (nx24559)) ;
    mux21_ni ix46809 (.Y (nx46808), .A0 (inputs_426__11), .A1 (inputs_427__11), 
             .S0 (nx24559)) ;
    mux21_ni ix46841 (.Y (nx46840), .A0 (nx46824), .A1 (nx46836), .S0 (nx23729)
             ) ;
    mux21_ni ix46825 (.Y (nx46824), .A0 (inputs_428__11), .A1 (inputs_429__11), 
             .S0 (nx24559)) ;
    mux21_ni ix46837 (.Y (nx46836), .A0 (inputs_430__11), .A1 (inputs_431__11), 
             .S0 (nx24559)) ;
    mux21_ni ix46905 (.Y (nx46904), .A0 (nx46872), .A1 (nx46900), .S0 (nx23293)
             ) ;
    mux21_ni ix46873 (.Y (nx46872), .A0 (nx46856), .A1 (nx46868), .S0 (nx23729)
             ) ;
    mux21_ni ix46857 (.Y (nx46856), .A0 (inputs_440__11), .A1 (inputs_441__11), 
             .S0 (nx24561)) ;
    mux21_ni ix46869 (.Y (nx46868), .A0 (inputs_442__11), .A1 (inputs_443__11), 
             .S0 (nx24561)) ;
    mux21_ni ix46901 (.Y (nx46900), .A0 (nx46884), .A1 (nx46896), .S0 (nx23731)
             ) ;
    mux21_ni ix46885 (.Y (nx46884), .A0 (inputs_444__11), .A1 (inputs_445__11), 
             .S0 (nx24561)) ;
    mux21_ni ix46897 (.Y (nx46896), .A0 (inputs_446__11), .A1 (inputs_447__11), 
             .S0 (nx24561)) ;
    mux21_ni ix47417 (.Y (nx47416), .A0 (nx47204), .A1 (nx47412), .S0 (nx22627)
             ) ;
    mux21_ni ix47205 (.Y (nx47204), .A0 (nx47198), .A1 (nx47120), .S0 (nx23169)
             ) ;
    oai21 ix47199 (.Y (nx47198), .A0 (nx22333), .A1 (nx18135), .B0 (nx18147)) ;
    mux21 ix18136 (.Y (nx18135), .A0 (nx47162), .A1 (nx47190), .S0 (nx22983)) ;
    mux21_ni ix47163 (.Y (nx47162), .A0 (nx47146), .A1 (nx47158), .S0 (nx23731)
             ) ;
    mux21_ni ix47147 (.Y (nx47146), .A0 (inputs_452__11), .A1 (inputs_453__11), 
             .S0 (nx24561)) ;
    mux21_ni ix47159 (.Y (nx47158), .A0 (inputs_454__11), .A1 (inputs_455__11), 
             .S0 (nx24561)) ;
    mux21_ni ix47191 (.Y (nx47190), .A0 (nx47174), .A1 (nx47186), .S0 (nx23731)
             ) ;
    mux21_ni ix47175 (.Y (nx47174), .A0 (inputs_468__11), .A1 (inputs_469__11), 
             .S0 (nx24561)) ;
    mux21_ni ix47187 (.Y (nx47186), .A0 (inputs_470__11), .A1 (inputs_471__11), 
             .S0 (nx24563)) ;
    nand04 ix18148 (.Y (nx18147), .A0 (nx22333), .A1 (nx23731), .A2 (nx24563), .A3 (
           nx47134)) ;
    mux21_ni ix47135 (.Y (nx47134), .A0 (inputs_451__11), .A1 (inputs_467__11), 
             .S0 (nx22983)) ;
    mux21_ni ix47121 (.Y (nx47120), .A0 (nx47056), .A1 (nx47116), .S0 (nx22983)
             ) ;
    mux21_ni ix47057 (.Y (nx47056), .A0 (nx47024), .A1 (nx47052), .S0 (nx23295)
             ) ;
    mux21_ni ix47025 (.Y (nx47024), .A0 (nx47008), .A1 (nx47020), .S0 (nx23731)
             ) ;
    mux21_ni ix47009 (.Y (nx47008), .A0 (inputs_456__11), .A1 (inputs_457__11), 
             .S0 (nx24563)) ;
    mux21_ni ix47021 (.Y (nx47020), .A0 (inputs_458__11), .A1 (inputs_459__11), 
             .S0 (nx24563)) ;
    mux21_ni ix47053 (.Y (nx47052), .A0 (nx47036), .A1 (nx47048), .S0 (nx23731)
             ) ;
    mux21_ni ix47037 (.Y (nx47036), .A0 (inputs_460__11), .A1 (inputs_461__11), 
             .S0 (nx24563)) ;
    mux21_ni ix47049 (.Y (nx47048), .A0 (inputs_462__11), .A1 (inputs_463__11), 
             .S0 (nx24563)) ;
    mux21_ni ix47117 (.Y (nx47116), .A0 (nx47084), .A1 (nx47112), .S0 (nx23295)
             ) ;
    mux21_ni ix47085 (.Y (nx47084), .A0 (nx47068), .A1 (nx47080), .S0 (nx23731)
             ) ;
    mux21_ni ix47069 (.Y (nx47068), .A0 (inputs_472__11), .A1 (inputs_473__11), 
             .S0 (nx24563)) ;
    mux21_ni ix47081 (.Y (nx47080), .A0 (inputs_474__11), .A1 (inputs_475__11), 
             .S0 (nx24565)) ;
    mux21_ni ix47113 (.Y (nx47112), .A0 (nx47096), .A1 (nx47108), .S0 (nx23733)
             ) ;
    mux21_ni ix47097 (.Y (nx47096), .A0 (inputs_476__11), .A1 (inputs_477__11), 
             .S0 (nx24565)) ;
    mux21_ni ix47109 (.Y (nx47108), .A0 (inputs_478__11), .A1 (inputs_479__11), 
             .S0 (nx24565)) ;
    mux21_ni ix47413 (.Y (nx47412), .A0 (nx47406), .A1 (nx47328), .S0 (nx23169)
             ) ;
    oai21 ix47407 (.Y (nx47406), .A0 (nx22333), .A1 (nx18179), .B0 (nx18191)) ;
    mux21 ix18180 (.Y (nx18179), .A0 (nx47370), .A1 (nx47398), .S0 (nx22983)) ;
    mux21_ni ix47371 (.Y (nx47370), .A0 (nx47354), .A1 (nx47366), .S0 (nx23733)
             ) ;
    mux21_ni ix47355 (.Y (nx47354), .A0 (inputs_484__11), .A1 (inputs_485__11), 
             .S0 (nx24565)) ;
    mux21_ni ix47367 (.Y (nx47366), .A0 (inputs_486__11), .A1 (inputs_487__11), 
             .S0 (nx24565)) ;
    mux21_ni ix47399 (.Y (nx47398), .A0 (nx47382), .A1 (nx47394), .S0 (nx23733)
             ) ;
    mux21_ni ix47383 (.Y (nx47382), .A0 (inputs_500__11), .A1 (inputs_501__11), 
             .S0 (nx24565)) ;
    mux21_ni ix47395 (.Y (nx47394), .A0 (inputs_502__11), .A1 (inputs_503__11), 
             .S0 (nx24565)) ;
    nand04 ix18192 (.Y (nx18191), .A0 (nx22335), .A1 (nx23733), .A2 (nx24567), .A3 (
           nx47342)) ;
    mux21_ni ix47343 (.Y (nx47342), .A0 (inputs_483__11), .A1 (inputs_499__11), 
             .S0 (nx22985)) ;
    mux21_ni ix47329 (.Y (nx47328), .A0 (nx47264), .A1 (nx47324), .S0 (nx22985)
             ) ;
    mux21_ni ix47265 (.Y (nx47264), .A0 (nx47232), .A1 (nx47260), .S0 (nx23295)
             ) ;
    mux21_ni ix47233 (.Y (nx47232), .A0 (nx47216), .A1 (nx47228), .S0 (nx23733)
             ) ;
    mux21_ni ix47217 (.Y (nx47216), .A0 (inputs_488__11), .A1 (inputs_489__11), 
             .S0 (nx24567)) ;
    mux21_ni ix47229 (.Y (nx47228), .A0 (inputs_490__11), .A1 (inputs_491__11), 
             .S0 (nx24567)) ;
    mux21_ni ix47261 (.Y (nx47260), .A0 (nx47244), .A1 (nx47256), .S0 (nx23733)
             ) ;
    mux21_ni ix47245 (.Y (nx47244), .A0 (inputs_492__11), .A1 (inputs_493__11), 
             .S0 (nx24567)) ;
    mux21_ni ix47257 (.Y (nx47256), .A0 (inputs_494__11), .A1 (inputs_495__11), 
             .S0 (nx24567)) ;
    mux21_ni ix47325 (.Y (nx47324), .A0 (nx47292), .A1 (nx47320), .S0 (nx23295)
             ) ;
    mux21_ni ix47293 (.Y (nx47292), .A0 (nx47276), .A1 (nx47288), .S0 (nx23733)
             ) ;
    mux21_ni ix47277 (.Y (nx47276), .A0 (inputs_504__11), .A1 (inputs_505__11), 
             .S0 (nx24567)) ;
    mux21_ni ix47289 (.Y (nx47288), .A0 (inputs_506__11), .A1 (inputs_507__11), 
             .S0 (nx24567)) ;
    mux21_ni ix47321 (.Y (nx47320), .A0 (nx47304), .A1 (nx47316), .S0 (nx23735)
             ) ;
    mux21_ni ix47305 (.Y (nx47304), .A0 (inputs_508__11), .A1 (inputs_509__11), 
             .S0 (nx24569)) ;
    mux21_ni ix47317 (.Y (nx47316), .A0 (inputs_510__11), .A1 (inputs_511__11), 
             .S0 (nx24569)) ;
    aoi32 ix18220 (.Y (nx18219), .A0 (nx48190), .A1 (nx22387), .A2 (nx22335), .B0 (
          nx22223), .B1 (nx49886)) ;
    oai21 ix48191 (.Y (nx48190), .A0 (nx23735), .A1 (nx18223), .B0 (nx18327)) ;
    mux21 ix18224 (.Y (nx18223), .A0 (nx47928), .A1 (nx48180), .S0 (nx24569)) ;
    mux21_ni ix47929 (.Y (nx47928), .A0 (nx47800), .A1 (nx47924), .S0 (nx22401)
             ) ;
    mux21_ni ix47801 (.Y (nx47800), .A0 (nx47736), .A1 (nx47796), .S0 (nx22435)
             ) ;
    mux21_ni ix47737 (.Y (nx47736), .A0 (nx47704), .A1 (nx47732), .S0 (nx22501)
             ) ;
    mux21_ni ix47705 (.Y (nx47704), .A0 (nx47688), .A1 (nx47700), .S0 (nx22627)
             ) ;
    mux21_ni ix47689 (.Y (nx47688), .A0 (inputs_0__11), .A1 (inputs_16__11), .S0 (
             nx22985)) ;
    mux21_ni ix47701 (.Y (nx47700), .A0 (inputs_32__11), .A1 (inputs_48__11), .S0 (
             nx22985)) ;
    mux21_ni ix47733 (.Y (nx47732), .A0 (nx47716), .A1 (nx47728), .S0 (nx22629)
             ) ;
    mux21_ni ix47717 (.Y (nx47716), .A0 (inputs_64__11), .A1 (inputs_80__11), .S0 (
             nx22985)) ;
    mux21_ni ix47729 (.Y (nx47728), .A0 (inputs_96__11), .A1 (inputs_112__11), .S0 (
             nx22985)) ;
    mux21_ni ix47797 (.Y (nx47796), .A0 (nx47764), .A1 (nx47792), .S0 (nx22501)
             ) ;
    mux21_ni ix47765 (.Y (nx47764), .A0 (nx47748), .A1 (nx47760), .S0 (nx22629)
             ) ;
    mux21_ni ix47749 (.Y (nx47748), .A0 (inputs_128__11), .A1 (inputs_144__11), 
             .S0 (nx22985)) ;
    mux21_ni ix47761 (.Y (nx47760), .A0 (inputs_160__11), .A1 (inputs_176__11), 
             .S0 (nx22987)) ;
    mux21_ni ix47793 (.Y (nx47792), .A0 (nx47776), .A1 (nx47788), .S0 (nx22629)
             ) ;
    mux21_ni ix47777 (.Y (nx47776), .A0 (inputs_192__11), .A1 (inputs_208__11), 
             .S0 (nx22987)) ;
    mux21_ni ix47789 (.Y (nx47788), .A0 (inputs_224__11), .A1 (inputs_240__11), 
             .S0 (nx22987)) ;
    mux21_ni ix47925 (.Y (nx47924), .A0 (nx47860), .A1 (nx47920), .S0 (nx22435)
             ) ;
    mux21_ni ix47861 (.Y (nx47860), .A0 (nx47828), .A1 (nx47856), .S0 (nx22501)
             ) ;
    mux21_ni ix47829 (.Y (nx47828), .A0 (nx47812), .A1 (nx47824), .S0 (nx22629)
             ) ;
    mux21_ni ix47813 (.Y (nx47812), .A0 (inputs_256__11), .A1 (inputs_272__11), 
             .S0 (nx22987)) ;
    mux21_ni ix47825 (.Y (nx47824), .A0 (inputs_288__11), .A1 (inputs_304__11), 
             .S0 (nx22987)) ;
    mux21_ni ix47857 (.Y (nx47856), .A0 (nx47840), .A1 (nx47852), .S0 (nx22629)
             ) ;
    mux21_ni ix47841 (.Y (nx47840), .A0 (inputs_320__11), .A1 (inputs_336__11), 
             .S0 (nx22987)) ;
    mux21_ni ix47853 (.Y (nx47852), .A0 (inputs_352__11), .A1 (inputs_368__11), 
             .S0 (nx22987)) ;
    mux21_ni ix47921 (.Y (nx47920), .A0 (nx47888), .A1 (nx47916), .S0 (nx22501)
             ) ;
    mux21_ni ix47889 (.Y (nx47888), .A0 (nx47872), .A1 (nx47884), .S0 (nx22629)
             ) ;
    mux21_ni ix47873 (.Y (nx47872), .A0 (inputs_384__11), .A1 (inputs_400__11), 
             .S0 (nx22989)) ;
    mux21_ni ix47885 (.Y (nx47884), .A0 (inputs_416__11), .A1 (inputs_432__11), 
             .S0 (nx22989)) ;
    mux21_ni ix47917 (.Y (nx47916), .A0 (nx47900), .A1 (nx47912), .S0 (nx22629)
             ) ;
    mux21_ni ix47901 (.Y (nx47900), .A0 (inputs_448__11), .A1 (inputs_464__11), 
             .S0 (nx22989)) ;
    mux21_ni ix47913 (.Y (nx47912), .A0 (inputs_480__11), .A1 (inputs_496__11), 
             .S0 (nx22989)) ;
    mux21_ni ix48181 (.Y (nx48180), .A0 (nx48052), .A1 (nx48176), .S0 (nx22401)
             ) ;
    mux21_ni ix48053 (.Y (nx48052), .A0 (nx47988), .A1 (nx48048), .S0 (nx22437)
             ) ;
    mux21_ni ix47989 (.Y (nx47988), .A0 (nx47956), .A1 (nx47984), .S0 (nx22503)
             ) ;
    mux21_ni ix47957 (.Y (nx47956), .A0 (nx47940), .A1 (nx47952), .S0 (nx22631)
             ) ;
    mux21_ni ix47941 (.Y (nx47940), .A0 (inputs_1__11), .A1 (inputs_17__11), .S0 (
             nx22989)) ;
    mux21_ni ix47953 (.Y (nx47952), .A0 (inputs_33__11), .A1 (inputs_49__11), .S0 (
             nx22989)) ;
    mux21_ni ix47985 (.Y (nx47984), .A0 (nx47968), .A1 (nx47980), .S0 (nx22631)
             ) ;
    mux21_ni ix47969 (.Y (nx47968), .A0 (inputs_65__11), .A1 (inputs_81__11), .S0 (
             nx22989)) ;
    mux21_ni ix47981 (.Y (nx47980), .A0 (inputs_97__11), .A1 (inputs_113__11), .S0 (
             nx22991)) ;
    mux21_ni ix48049 (.Y (nx48048), .A0 (nx48016), .A1 (nx48044), .S0 (nx22503)
             ) ;
    mux21_ni ix48017 (.Y (nx48016), .A0 (nx48000), .A1 (nx48012), .S0 (nx22631)
             ) ;
    mux21_ni ix48001 (.Y (nx48000), .A0 (inputs_129__11), .A1 (inputs_145__11), 
             .S0 (nx22991)) ;
    mux21_ni ix48013 (.Y (nx48012), .A0 (inputs_161__11), .A1 (inputs_177__11), 
             .S0 (nx22991)) ;
    mux21_ni ix48045 (.Y (nx48044), .A0 (nx48028), .A1 (nx48040), .S0 (nx22631)
             ) ;
    mux21_ni ix48029 (.Y (nx48028), .A0 (inputs_193__11), .A1 (inputs_209__11), 
             .S0 (nx22991)) ;
    mux21_ni ix48041 (.Y (nx48040), .A0 (inputs_225__11), .A1 (inputs_241__11), 
             .S0 (nx22991)) ;
    mux21_ni ix48177 (.Y (nx48176), .A0 (nx48112), .A1 (nx48172), .S0 (nx22437)
             ) ;
    mux21_ni ix48113 (.Y (nx48112), .A0 (nx48080), .A1 (nx48108), .S0 (nx22503)
             ) ;
    mux21_ni ix48081 (.Y (nx48080), .A0 (nx48064), .A1 (nx48076), .S0 (nx22631)
             ) ;
    mux21_ni ix48065 (.Y (nx48064), .A0 (inputs_257__11), .A1 (inputs_273__11), 
             .S0 (nx22991)) ;
    mux21_ni ix48077 (.Y (nx48076), .A0 (inputs_289__11), .A1 (inputs_305__11), 
             .S0 (nx22991)) ;
    mux21_ni ix48109 (.Y (nx48108), .A0 (nx48092), .A1 (nx48104), .S0 (nx22631)
             ) ;
    mux21_ni ix48093 (.Y (nx48092), .A0 (inputs_321__11), .A1 (inputs_337__11), 
             .S0 (nx22993)) ;
    mux21_ni ix48105 (.Y (nx48104), .A0 (inputs_353__11), .A1 (inputs_369__11), 
             .S0 (nx22993)) ;
    mux21_ni ix48173 (.Y (nx48172), .A0 (nx48140), .A1 (nx48168), .S0 (nx22503)
             ) ;
    mux21_ni ix48141 (.Y (nx48140), .A0 (nx48124), .A1 (nx48136), .S0 (nx22631)
             ) ;
    mux21_ni ix48125 (.Y (nx48124), .A0 (inputs_385__11), .A1 (inputs_401__11), 
             .S0 (nx22993)) ;
    mux21_ni ix48137 (.Y (nx48136), .A0 (inputs_417__11), .A1 (inputs_433__11), 
             .S0 (nx22993)) ;
    mux21_ni ix48169 (.Y (nx48168), .A0 (nx48152), .A1 (nx48164), .S0 (nx22633)
             ) ;
    mux21_ni ix48153 (.Y (nx48152), .A0 (inputs_449__11), .A1 (inputs_465__11), 
             .S0 (nx22993)) ;
    mux21_ni ix48165 (.Y (nx48164), .A0 (inputs_481__11), .A1 (inputs_497__11), 
             .S0 (nx22993)) ;
    nand03 ix18328 (.Y (nx18327), .A0 (nx47674), .A1 (nx23735), .A2 (nx22381)) ;
    mux21_ni ix47675 (.Y (nx47674), .A0 (nx47546), .A1 (nx47670), .S0 (nx22403)
             ) ;
    mux21_ni ix47547 (.Y (nx47546), .A0 (nx47482), .A1 (nx47542), .S0 (nx22437)
             ) ;
    mux21_ni ix47483 (.Y (nx47482), .A0 (nx47450), .A1 (nx47478), .S0 (nx22503)
             ) ;
    mux21_ni ix47451 (.Y (nx47450), .A0 (nx47434), .A1 (nx47446), .S0 (nx22633)
             ) ;
    mux21_ni ix47435 (.Y (nx47434), .A0 (inputs_2__11), .A1 (inputs_18__11), .S0 (
             nx22993)) ;
    mux21_ni ix47447 (.Y (nx47446), .A0 (inputs_34__11), .A1 (inputs_50__11), .S0 (
             nx22995)) ;
    mux21_ni ix47479 (.Y (nx47478), .A0 (nx47462), .A1 (nx47474), .S0 (nx22633)
             ) ;
    mux21_ni ix47463 (.Y (nx47462), .A0 (inputs_66__11), .A1 (inputs_82__11), .S0 (
             nx22995)) ;
    mux21_ni ix47475 (.Y (nx47474), .A0 (inputs_98__11), .A1 (inputs_114__11), .S0 (
             nx22995)) ;
    mux21_ni ix47543 (.Y (nx47542), .A0 (nx47510), .A1 (nx47538), .S0 (nx22503)
             ) ;
    mux21_ni ix47511 (.Y (nx47510), .A0 (nx47494), .A1 (nx47506), .S0 (nx22633)
             ) ;
    mux21_ni ix47495 (.Y (nx47494), .A0 (inputs_130__11), .A1 (inputs_146__11), 
             .S0 (nx22995)) ;
    mux21_ni ix47507 (.Y (nx47506), .A0 (inputs_162__11), .A1 (inputs_178__11), 
             .S0 (nx22995)) ;
    mux21_ni ix47539 (.Y (nx47538), .A0 (nx47522), .A1 (nx47534), .S0 (nx22633)
             ) ;
    mux21_ni ix47523 (.Y (nx47522), .A0 (inputs_194__11), .A1 (inputs_210__11), 
             .S0 (nx22995)) ;
    mux21_ni ix47535 (.Y (nx47534), .A0 (inputs_226__11), .A1 (inputs_242__11), 
             .S0 (nx22995)) ;
    mux21_ni ix47671 (.Y (nx47670), .A0 (nx47606), .A1 (nx47666), .S0 (nx22437)
             ) ;
    mux21_ni ix47607 (.Y (nx47606), .A0 (nx47574), .A1 (nx47602), .S0 (nx22503)
             ) ;
    mux21_ni ix47575 (.Y (nx47574), .A0 (nx47558), .A1 (nx47570), .S0 (nx22633)
             ) ;
    mux21_ni ix47559 (.Y (nx47558), .A0 (inputs_258__11), .A1 (inputs_274__11), 
             .S0 (nx22997)) ;
    mux21_ni ix47571 (.Y (nx47570), .A0 (inputs_290__11), .A1 (inputs_306__11), 
             .S0 (nx22997)) ;
    mux21_ni ix47603 (.Y (nx47602), .A0 (nx47586), .A1 (nx47598), .S0 (nx22633)
             ) ;
    mux21_ni ix47587 (.Y (nx47586), .A0 (inputs_322__11), .A1 (inputs_338__11), 
             .S0 (nx22997)) ;
    mux21_ni ix47599 (.Y (nx47598), .A0 (inputs_354__11), .A1 (inputs_370__11), 
             .S0 (nx22997)) ;
    mux21_ni ix47667 (.Y (nx47666), .A0 (nx47634), .A1 (nx47662), .S0 (nx22505)
             ) ;
    mux21_ni ix47635 (.Y (nx47634), .A0 (nx47618), .A1 (nx47630), .S0 (nx22635)
             ) ;
    mux21_ni ix47619 (.Y (nx47618), .A0 (inputs_386__11), .A1 (inputs_402__11), 
             .S0 (nx22997)) ;
    mux21_ni ix47631 (.Y (nx47630), .A0 (inputs_418__11), .A1 (inputs_434__11), 
             .S0 (nx22997)) ;
    mux21_ni ix47663 (.Y (nx47662), .A0 (nx47646), .A1 (nx47658), .S0 (nx22635)
             ) ;
    mux21_ni ix47647 (.Y (nx47646), .A0 (inputs_450__11), .A1 (inputs_466__11), 
             .S0 (nx22997)) ;
    mux21_ni ix47659 (.Y (nx47658), .A0 (inputs_482__11), .A1 (inputs_498__11), 
             .S0 (nx22999)) ;
    mux21_ni ix49887 (.Y (nx49886), .A0 (nx49038), .A1 (nx49882), .S0 (nx22437)
             ) ;
    mux21_ni ix49039 (.Y (nx49038), .A0 (nx48614), .A1 (nx49034), .S0 (nx22505)
             ) ;
    mux21_ni ix48615 (.Y (nx48614), .A0 (nx48402), .A1 (nx48610), .S0 (nx22635)
             ) ;
    mux21_ni ix48403 (.Y (nx48402), .A0 (nx48396), .A1 (nx48318), .S0 (nx23169)
             ) ;
    oai21 ix48397 (.Y (nx48396), .A0 (nx22335), .A1 (nx18385), .B0 (nx18397)) ;
    mux21 ix18386 (.Y (nx18385), .A0 (nx48360), .A1 (nx48388), .S0 (nx22999)) ;
    mux21_ni ix48361 (.Y (nx48360), .A0 (nx48344), .A1 (nx48356), .S0 (nx23735)
             ) ;
    mux21_ni ix48345 (.Y (nx48344), .A0 (inputs_4__11), .A1 (inputs_5__11), .S0 (
             nx24569)) ;
    mux21_ni ix48357 (.Y (nx48356), .A0 (inputs_6__11), .A1 (inputs_7__11), .S0 (
             nx24569)) ;
    mux21_ni ix48389 (.Y (nx48388), .A0 (nx48372), .A1 (nx48384), .S0 (nx23735)
             ) ;
    mux21_ni ix48373 (.Y (nx48372), .A0 (inputs_20__11), .A1 (inputs_21__11), .S0 (
             nx24569)) ;
    mux21_ni ix48385 (.Y (nx48384), .A0 (inputs_22__11), .A1 (inputs_23__11), .S0 (
             nx24569)) ;
    nand04 ix18398 (.Y (nx18397), .A0 (nx22335), .A1 (nx23735), .A2 (nx24571), .A3 (
           nx48332)) ;
    mux21_ni ix48333 (.Y (nx48332), .A0 (inputs_3__11), .A1 (inputs_19__11), .S0 (
             nx22999)) ;
    mux21_ni ix48319 (.Y (nx48318), .A0 (nx48254), .A1 (nx48314), .S0 (nx22999)
             ) ;
    mux21_ni ix48255 (.Y (nx48254), .A0 (nx48222), .A1 (nx48250), .S0 (nx23295)
             ) ;
    mux21_ni ix48223 (.Y (nx48222), .A0 (nx48206), .A1 (nx48218), .S0 (nx23735)
             ) ;
    mux21_ni ix48207 (.Y (nx48206), .A0 (inputs_8__11), .A1 (inputs_9__11), .S0 (
             nx24571)) ;
    mux21_ni ix48219 (.Y (nx48218), .A0 (inputs_10__11), .A1 (inputs_11__11), .S0 (
             nx24571)) ;
    mux21_ni ix48251 (.Y (nx48250), .A0 (nx48234), .A1 (nx48246), .S0 (nx23737)
             ) ;
    mux21_ni ix48235 (.Y (nx48234), .A0 (inputs_12__11), .A1 (inputs_13__11), .S0 (
             nx24571)) ;
    mux21_ni ix48247 (.Y (nx48246), .A0 (inputs_14__11), .A1 (inputs_15__11), .S0 (
             nx24571)) ;
    mux21_ni ix48315 (.Y (nx48314), .A0 (nx48282), .A1 (nx48310), .S0 (nx23295)
             ) ;
    mux21_ni ix48283 (.Y (nx48282), .A0 (nx48266), .A1 (nx48278), .S0 (nx23737)
             ) ;
    mux21_ni ix48267 (.Y (nx48266), .A0 (inputs_24__11), .A1 (inputs_25__11), .S0 (
             nx24571)) ;
    mux21_ni ix48279 (.Y (nx48278), .A0 (inputs_26__11), .A1 (inputs_27__11), .S0 (
             nx24571)) ;
    mux21_ni ix48311 (.Y (nx48310), .A0 (nx48294), .A1 (nx48306), .S0 (nx23737)
             ) ;
    mux21_ni ix48295 (.Y (nx48294), .A0 (inputs_28__11), .A1 (inputs_29__11), .S0 (
             nx24573)) ;
    mux21_ni ix48307 (.Y (nx48306), .A0 (inputs_30__11), .A1 (inputs_31__11), .S0 (
             nx24573)) ;
    mux21_ni ix48611 (.Y (nx48610), .A0 (nx48604), .A1 (nx48526), .S0 (nx23169)
             ) ;
    oai21 ix48605 (.Y (nx48604), .A0 (nx22335), .A1 (nx18427), .B0 (nx18441)) ;
    mux21 ix18428 (.Y (nx18427), .A0 (nx48568), .A1 (nx48596), .S0 (nx22999)) ;
    mux21_ni ix48569 (.Y (nx48568), .A0 (nx48552), .A1 (nx48564), .S0 (nx23737)
             ) ;
    mux21_ni ix48553 (.Y (nx48552), .A0 (inputs_36__11), .A1 (inputs_37__11), .S0 (
             nx24573)) ;
    mux21_ni ix48565 (.Y (nx48564), .A0 (inputs_38__11), .A1 (inputs_39__11), .S0 (
             nx24573)) ;
    mux21_ni ix48597 (.Y (nx48596), .A0 (nx48580), .A1 (nx48592), .S0 (nx23737)
             ) ;
    mux21_ni ix48581 (.Y (nx48580), .A0 (inputs_52__11), .A1 (inputs_53__11), .S0 (
             nx24573)) ;
    mux21_ni ix48593 (.Y (nx48592), .A0 (inputs_54__11), .A1 (inputs_55__11), .S0 (
             nx24573)) ;
    nand04 ix18442 (.Y (nx18441), .A0 (nx22335), .A1 (nx23737), .A2 (nx24573), .A3 (
           nx48540)) ;
    mux21_ni ix48541 (.Y (nx48540), .A0 (inputs_35__11), .A1 (inputs_51__11), .S0 (
             nx22999)) ;
    mux21_ni ix48527 (.Y (nx48526), .A0 (nx48462), .A1 (nx48522), .S0 (nx22999)
             ) ;
    mux21_ni ix48463 (.Y (nx48462), .A0 (nx48430), .A1 (nx48458), .S0 (nx23295)
             ) ;
    mux21_ni ix48431 (.Y (nx48430), .A0 (nx48414), .A1 (nx48426), .S0 (nx23737)
             ) ;
    mux21_ni ix48415 (.Y (nx48414), .A0 (inputs_40__11), .A1 (inputs_41__11), .S0 (
             nx24575)) ;
    mux21_ni ix48427 (.Y (nx48426), .A0 (inputs_42__11), .A1 (inputs_43__11), .S0 (
             nx24575)) ;
    mux21_ni ix48459 (.Y (nx48458), .A0 (nx48442), .A1 (nx48454), .S0 (nx23739)
             ) ;
    mux21_ni ix48443 (.Y (nx48442), .A0 (inputs_44__11), .A1 (inputs_45__11), .S0 (
             nx24575)) ;
    mux21_ni ix48455 (.Y (nx48454), .A0 (inputs_46__11), .A1 (inputs_47__11), .S0 (
             nx24575)) ;
    mux21_ni ix48523 (.Y (nx48522), .A0 (nx48490), .A1 (nx48518), .S0 (nx23297)
             ) ;
    mux21_ni ix48491 (.Y (nx48490), .A0 (nx48474), .A1 (nx48486), .S0 (nx23739)
             ) ;
    mux21_ni ix48475 (.Y (nx48474), .A0 (inputs_56__11), .A1 (inputs_57__11), .S0 (
             nx24575)) ;
    mux21_ni ix48487 (.Y (nx48486), .A0 (inputs_58__11), .A1 (inputs_59__11), .S0 (
             nx24575)) ;
    mux21_ni ix48519 (.Y (nx48518), .A0 (nx48502), .A1 (nx48514), .S0 (nx23739)
             ) ;
    mux21_ni ix48503 (.Y (nx48502), .A0 (inputs_60__11), .A1 (inputs_61__11), .S0 (
             nx24575)) ;
    mux21_ni ix48515 (.Y (nx48514), .A0 (inputs_62__11), .A1 (inputs_63__11), .S0 (
             nx24577)) ;
    mux21_ni ix49035 (.Y (nx49034), .A0 (nx48822), .A1 (nx49030), .S0 (nx22635)
             ) ;
    mux21_ni ix48823 (.Y (nx48822), .A0 (nx48816), .A1 (nx48738), .S0 (nx23169)
             ) ;
    oai21 ix48817 (.Y (nx48816), .A0 (nx22335), .A1 (nx18473), .B0 (nx18485)) ;
    mux21 ix18474 (.Y (nx18473), .A0 (nx48780), .A1 (nx48808), .S0 (nx23001)) ;
    mux21_ni ix48781 (.Y (nx48780), .A0 (nx48764), .A1 (nx48776), .S0 (nx23739)
             ) ;
    mux21_ni ix48765 (.Y (nx48764), .A0 (inputs_68__11), .A1 (inputs_69__11), .S0 (
             nx24577)) ;
    mux21_ni ix48777 (.Y (nx48776), .A0 (inputs_70__11), .A1 (inputs_71__11), .S0 (
             nx24577)) ;
    mux21_ni ix48809 (.Y (nx48808), .A0 (nx48792), .A1 (nx48804), .S0 (nx23739)
             ) ;
    mux21_ni ix48793 (.Y (nx48792), .A0 (inputs_84__11), .A1 (inputs_85__11), .S0 (
             nx24577)) ;
    mux21_ni ix48805 (.Y (nx48804), .A0 (inputs_86__11), .A1 (inputs_87__11), .S0 (
             nx24577)) ;
    nand04 ix18486 (.Y (nx18485), .A0 (nx22337), .A1 (nx23739), .A2 (nx24577), .A3 (
           nx48752)) ;
    mux21_ni ix48753 (.Y (nx48752), .A0 (inputs_67__11), .A1 (inputs_83__11), .S0 (
             nx23001)) ;
    mux21_ni ix48739 (.Y (nx48738), .A0 (nx48674), .A1 (nx48734), .S0 (nx23001)
             ) ;
    mux21_ni ix48675 (.Y (nx48674), .A0 (nx48642), .A1 (nx48670), .S0 (nx23297)
             ) ;
    mux21_ni ix48643 (.Y (nx48642), .A0 (nx48626), .A1 (nx48638), .S0 (nx23739)
             ) ;
    mux21_ni ix48627 (.Y (nx48626), .A0 (inputs_72__11), .A1 (inputs_73__11), .S0 (
             nx24577)) ;
    mux21_ni ix48639 (.Y (nx48638), .A0 (inputs_74__11), .A1 (inputs_75__11), .S0 (
             nx24579)) ;
    mux21_ni ix48671 (.Y (nx48670), .A0 (nx48654), .A1 (nx48666), .S0 (nx23741)
             ) ;
    mux21_ni ix48655 (.Y (nx48654), .A0 (inputs_76__11), .A1 (inputs_77__11), .S0 (
             nx24579)) ;
    mux21_ni ix48667 (.Y (nx48666), .A0 (inputs_78__11), .A1 (inputs_79__11), .S0 (
             nx24579)) ;
    mux21_ni ix48735 (.Y (nx48734), .A0 (nx48702), .A1 (nx48730), .S0 (nx23297)
             ) ;
    mux21_ni ix48703 (.Y (nx48702), .A0 (nx48686), .A1 (nx48698), .S0 (nx23741)
             ) ;
    mux21_ni ix48687 (.Y (nx48686), .A0 (inputs_88__11), .A1 (inputs_89__11), .S0 (
             nx24579)) ;
    mux21_ni ix48699 (.Y (nx48698), .A0 (inputs_90__11), .A1 (inputs_91__11), .S0 (
             nx24579)) ;
    mux21_ni ix48731 (.Y (nx48730), .A0 (nx48714), .A1 (nx48726), .S0 (nx23741)
             ) ;
    mux21_ni ix48715 (.Y (nx48714), .A0 (inputs_92__11), .A1 (inputs_93__11), .S0 (
             nx24579)) ;
    mux21_ni ix48727 (.Y (nx48726), .A0 (inputs_94__11), .A1 (inputs_95__11), .S0 (
             nx24579)) ;
    mux21_ni ix49031 (.Y (nx49030), .A0 (nx49024), .A1 (nx48946), .S0 (nx23169)
             ) ;
    oai21 ix49025 (.Y (nx49024), .A0 (nx22337), .A1 (nx18517), .B0 (nx18529)) ;
    mux21 ix18518 (.Y (nx18517), .A0 (nx48988), .A1 (nx49016), .S0 (nx23001)) ;
    mux21_ni ix48989 (.Y (nx48988), .A0 (nx48972), .A1 (nx48984), .S0 (nx23741)
             ) ;
    mux21_ni ix48973 (.Y (nx48972), .A0 (inputs_100__11), .A1 (inputs_101__11), 
             .S0 (nx24581)) ;
    mux21_ni ix48985 (.Y (nx48984), .A0 (inputs_102__11), .A1 (inputs_103__11), 
             .S0 (nx24581)) ;
    mux21_ni ix49017 (.Y (nx49016), .A0 (nx49000), .A1 (nx49012), .S0 (nx23741)
             ) ;
    mux21_ni ix49001 (.Y (nx49000), .A0 (inputs_116__11), .A1 (inputs_117__11), 
             .S0 (nx24581)) ;
    mux21_ni ix49013 (.Y (nx49012), .A0 (inputs_118__11), .A1 (inputs_119__11), 
             .S0 (nx24581)) ;
    nand04 ix18530 (.Y (nx18529), .A0 (nx22337), .A1 (nx23741), .A2 (nx24581), .A3 (
           nx48960)) ;
    mux21_ni ix48961 (.Y (nx48960), .A0 (inputs_99__11), .A1 (inputs_115__11), .S0 (
             nx23001)) ;
    mux21_ni ix48947 (.Y (nx48946), .A0 (nx48882), .A1 (nx48942), .S0 (nx23001)
             ) ;
    mux21_ni ix48883 (.Y (nx48882), .A0 (nx48850), .A1 (nx48878), .S0 (nx23297)
             ) ;
    mux21_ni ix48851 (.Y (nx48850), .A0 (nx48834), .A1 (nx48846), .S0 (nx23741)
             ) ;
    mux21_ni ix48835 (.Y (nx48834), .A0 (inputs_104__11), .A1 (inputs_105__11), 
             .S0 (nx24581)) ;
    mux21_ni ix48847 (.Y (nx48846), .A0 (inputs_106__11), .A1 (inputs_107__11), 
             .S0 (nx24581)) ;
    mux21_ni ix48879 (.Y (nx48878), .A0 (nx48862), .A1 (nx48874), .S0 (nx23743)
             ) ;
    mux21_ni ix48863 (.Y (nx48862), .A0 (inputs_108__11), .A1 (inputs_109__11), 
             .S0 (nx24583)) ;
    mux21_ni ix48875 (.Y (nx48874), .A0 (inputs_110__11), .A1 (inputs_111__11), 
             .S0 (nx24583)) ;
    mux21_ni ix48943 (.Y (nx48942), .A0 (nx48910), .A1 (nx48938), .S0 (nx23297)
             ) ;
    mux21_ni ix48911 (.Y (nx48910), .A0 (nx48894), .A1 (nx48906), .S0 (nx23743)
             ) ;
    mux21_ni ix48895 (.Y (nx48894), .A0 (inputs_120__11), .A1 (inputs_121__11), 
             .S0 (nx24583)) ;
    mux21_ni ix48907 (.Y (nx48906), .A0 (inputs_122__11), .A1 (inputs_123__11), 
             .S0 (nx24583)) ;
    mux21_ni ix48939 (.Y (nx48938), .A0 (nx48922), .A1 (nx48934), .S0 (nx23743)
             ) ;
    mux21_ni ix48923 (.Y (nx48922), .A0 (inputs_124__11), .A1 (inputs_125__11), 
             .S0 (nx24583)) ;
    mux21_ni ix48935 (.Y (nx48934), .A0 (inputs_126__11), .A1 (inputs_127__11), 
             .S0 (nx24583)) ;
    mux21_ni ix49883 (.Y (nx49882), .A0 (nx49458), .A1 (nx49878), .S0 (nx22505)
             ) ;
    mux21_ni ix49459 (.Y (nx49458), .A0 (nx49246), .A1 (nx49454), .S0 (nx22635)
             ) ;
    mux21_ni ix49247 (.Y (nx49246), .A0 (nx49240), .A1 (nx49162), .S0 (nx23169)
             ) ;
    oai21 ix49241 (.Y (nx49240), .A0 (nx22337), .A1 (nx18563), .B0 (nx18575)) ;
    mux21 ix18564 (.Y (nx18563), .A0 (nx49204), .A1 (nx49232), .S0 (nx23001)) ;
    mux21_ni ix49205 (.Y (nx49204), .A0 (nx49188), .A1 (nx49200), .S0 (nx23743)
             ) ;
    mux21_ni ix49189 (.Y (nx49188), .A0 (inputs_132__11), .A1 (inputs_133__11), 
             .S0 (nx24583)) ;
    mux21_ni ix49201 (.Y (nx49200), .A0 (inputs_134__11), .A1 (inputs_135__11), 
             .S0 (nx24585)) ;
    mux21_ni ix49233 (.Y (nx49232), .A0 (nx49216), .A1 (nx49228), .S0 (nx23743)
             ) ;
    mux21_ni ix49217 (.Y (nx49216), .A0 (inputs_148__11), .A1 (inputs_149__11), 
             .S0 (nx24585)) ;
    mux21_ni ix49229 (.Y (nx49228), .A0 (inputs_150__11), .A1 (inputs_151__11), 
             .S0 (nx24585)) ;
    nand04 ix18576 (.Y (nx18575), .A0 (nx22337), .A1 (nx23743), .A2 (nx24585), .A3 (
           nx49176)) ;
    mux21_ni ix49177 (.Y (nx49176), .A0 (inputs_131__11), .A1 (inputs_147__11), 
             .S0 (nx23003)) ;
    mux21_ni ix49163 (.Y (nx49162), .A0 (nx49098), .A1 (nx49158), .S0 (nx23003)
             ) ;
    mux21_ni ix49099 (.Y (nx49098), .A0 (nx49066), .A1 (nx49094), .S0 (nx23297)
             ) ;
    mux21_ni ix49067 (.Y (nx49066), .A0 (nx49050), .A1 (nx49062), .S0 (nx23743)
             ) ;
    mux21_ni ix49051 (.Y (nx49050), .A0 (inputs_136__11), .A1 (inputs_137__11), 
             .S0 (nx24585)) ;
    mux21_ni ix49063 (.Y (nx49062), .A0 (inputs_138__11), .A1 (inputs_139__11), 
             .S0 (nx24585)) ;
    mux21_ni ix49095 (.Y (nx49094), .A0 (nx49078), .A1 (nx49090), .S0 (nx23745)
             ) ;
    mux21_ni ix49079 (.Y (nx49078), .A0 (inputs_140__11), .A1 (inputs_141__11), 
             .S0 (nx24585)) ;
    mux21_ni ix49091 (.Y (nx49090), .A0 (inputs_142__11), .A1 (inputs_143__11), 
             .S0 (nx24587)) ;
    mux21_ni ix49159 (.Y (nx49158), .A0 (nx49126), .A1 (nx49154), .S0 (nx23297)
             ) ;
    mux21_ni ix49127 (.Y (nx49126), .A0 (nx49110), .A1 (nx49122), .S0 (nx23745)
             ) ;
    mux21_ni ix49111 (.Y (nx49110), .A0 (inputs_152__11), .A1 (inputs_153__11), 
             .S0 (nx24587)) ;
    mux21_ni ix49123 (.Y (nx49122), .A0 (inputs_154__11), .A1 (inputs_155__11), 
             .S0 (nx24587)) ;
    mux21_ni ix49155 (.Y (nx49154), .A0 (nx49138), .A1 (nx49150), .S0 (nx23745)
             ) ;
    mux21_ni ix49139 (.Y (nx49138), .A0 (inputs_156__11), .A1 (inputs_157__11), 
             .S0 (nx24587)) ;
    mux21_ni ix49151 (.Y (nx49150), .A0 (inputs_158__11), .A1 (inputs_159__11), 
             .S0 (nx24587)) ;
    mux21_ni ix49455 (.Y (nx49454), .A0 (nx49448), .A1 (nx49370), .S0 (nx23171)
             ) ;
    oai21 ix49449 (.Y (nx49448), .A0 (nx22337), .A1 (nx18605), .B0 (nx18617)) ;
    mux21 ix18606 (.Y (nx18605), .A0 (nx49412), .A1 (nx49440), .S0 (nx23003)) ;
    mux21_ni ix49413 (.Y (nx49412), .A0 (nx49396), .A1 (nx49408), .S0 (nx23745)
             ) ;
    mux21_ni ix49397 (.Y (nx49396), .A0 (inputs_164__11), .A1 (inputs_165__11), 
             .S0 (nx24587)) ;
    mux21_ni ix49409 (.Y (nx49408), .A0 (inputs_166__11), .A1 (inputs_167__11), 
             .S0 (nx24587)) ;
    mux21_ni ix49441 (.Y (nx49440), .A0 (nx49424), .A1 (nx49436), .S0 (nx23745)
             ) ;
    mux21_ni ix49425 (.Y (nx49424), .A0 (inputs_180__11), .A1 (inputs_181__11), 
             .S0 (nx24589)) ;
    mux21_ni ix49437 (.Y (nx49436), .A0 (inputs_182__11), .A1 (inputs_183__11), 
             .S0 (nx24589)) ;
    nand04 ix18618 (.Y (nx18617), .A0 (nx22337), .A1 (nx23745), .A2 (nx24589), .A3 (
           nx49384)) ;
    mux21_ni ix49385 (.Y (nx49384), .A0 (inputs_163__11), .A1 (inputs_179__11), 
             .S0 (nx23003)) ;
    mux21_ni ix49371 (.Y (nx49370), .A0 (nx49306), .A1 (nx49366), .S0 (nx23003)
             ) ;
    mux21_ni ix49307 (.Y (nx49306), .A0 (nx49274), .A1 (nx49302), .S0 (nx23299)
             ) ;
    mux21_ni ix49275 (.Y (nx49274), .A0 (nx49258), .A1 (nx49270), .S0 (nx23745)
             ) ;
    mux21_ni ix49259 (.Y (nx49258), .A0 (inputs_168__11), .A1 (inputs_169__11), 
             .S0 (nx24589)) ;
    mux21_ni ix49271 (.Y (nx49270), .A0 (inputs_170__11), .A1 (inputs_171__11), 
             .S0 (nx24589)) ;
    mux21_ni ix49303 (.Y (nx49302), .A0 (nx49286), .A1 (nx49298), .S0 (nx23747)
             ) ;
    mux21_ni ix49287 (.Y (nx49286), .A0 (inputs_172__11), .A1 (inputs_173__11), 
             .S0 (nx24589)) ;
    mux21_ni ix49299 (.Y (nx49298), .A0 (inputs_174__11), .A1 (inputs_175__11), 
             .S0 (nx24589)) ;
    mux21_ni ix49367 (.Y (nx49366), .A0 (nx49334), .A1 (nx49362), .S0 (nx23299)
             ) ;
    mux21_ni ix49335 (.Y (nx49334), .A0 (nx49318), .A1 (nx49330), .S0 (nx23747)
             ) ;
    mux21_ni ix49319 (.Y (nx49318), .A0 (inputs_184__11), .A1 (inputs_185__11), 
             .S0 (nx24591)) ;
    mux21_ni ix49331 (.Y (nx49330), .A0 (inputs_186__11), .A1 (inputs_187__11), 
             .S0 (nx24591)) ;
    mux21_ni ix49363 (.Y (nx49362), .A0 (nx49346), .A1 (nx49358), .S0 (nx23747)
             ) ;
    mux21_ni ix49347 (.Y (nx49346), .A0 (inputs_188__11), .A1 (inputs_189__11), 
             .S0 (nx24591)) ;
    mux21_ni ix49359 (.Y (nx49358), .A0 (inputs_190__11), .A1 (inputs_191__11), 
             .S0 (nx24591)) ;
    mux21_ni ix49879 (.Y (nx49878), .A0 (nx49666), .A1 (nx49874), .S0 (nx22635)
             ) ;
    mux21_ni ix49667 (.Y (nx49666), .A0 (nx49660), .A1 (nx49582), .S0 (nx23171)
             ) ;
    oai21 ix49661 (.Y (nx49660), .A0 (nx22339), .A1 (nx18651), .B0 (nx18663)) ;
    mux21 ix18652 (.Y (nx18651), .A0 (nx49624), .A1 (nx49652), .S0 (nx23003)) ;
    mux21_ni ix49625 (.Y (nx49624), .A0 (nx49608), .A1 (nx49620), .S0 (nx23747)
             ) ;
    mux21_ni ix49609 (.Y (nx49608), .A0 (inputs_196__11), .A1 (inputs_197__11), 
             .S0 (nx24591)) ;
    mux21_ni ix49621 (.Y (nx49620), .A0 (inputs_198__11), .A1 (inputs_199__11), 
             .S0 (nx24591)) ;
    mux21_ni ix49653 (.Y (nx49652), .A0 (nx49636), .A1 (nx49648), .S0 (nx23747)
             ) ;
    mux21_ni ix49637 (.Y (nx49636), .A0 (inputs_212__11), .A1 (inputs_213__11), 
             .S0 (nx24591)) ;
    mux21_ni ix49649 (.Y (nx49648), .A0 (inputs_214__11), .A1 (inputs_215__11), 
             .S0 (nx24593)) ;
    nand04 ix18664 (.Y (nx18663), .A0 (nx22339), .A1 (nx23747), .A2 (nx24593), .A3 (
           nx49596)) ;
    mux21_ni ix49597 (.Y (nx49596), .A0 (inputs_195__11), .A1 (inputs_211__11), 
             .S0 (nx23003)) ;
    mux21_ni ix49583 (.Y (nx49582), .A0 (nx49518), .A1 (nx49578), .S0 (nx23005)
             ) ;
    mux21_ni ix49519 (.Y (nx49518), .A0 (nx49486), .A1 (nx49514), .S0 (nx23299)
             ) ;
    mux21_ni ix49487 (.Y (nx49486), .A0 (nx49470), .A1 (nx49482), .S0 (nx23747)
             ) ;
    mux21_ni ix49471 (.Y (nx49470), .A0 (inputs_200__11), .A1 (inputs_201__11), 
             .S0 (nx24593)) ;
    mux21_ni ix49483 (.Y (nx49482), .A0 (inputs_202__11), .A1 (inputs_203__11), 
             .S0 (nx24593)) ;
    mux21_ni ix49515 (.Y (nx49514), .A0 (nx49498), .A1 (nx49510), .S0 (nx23749)
             ) ;
    mux21_ni ix49499 (.Y (nx49498), .A0 (inputs_204__11), .A1 (inputs_205__11), 
             .S0 (nx24593)) ;
    mux21_ni ix49511 (.Y (nx49510), .A0 (inputs_206__11), .A1 (inputs_207__11), 
             .S0 (nx24593)) ;
    mux21_ni ix49579 (.Y (nx49578), .A0 (nx49546), .A1 (nx49574), .S0 (nx23299)
             ) ;
    mux21_ni ix49547 (.Y (nx49546), .A0 (nx49530), .A1 (nx49542), .S0 (nx23749)
             ) ;
    mux21_ni ix49531 (.Y (nx49530), .A0 (inputs_216__11), .A1 (inputs_217__11), 
             .S0 (nx24593)) ;
    mux21_ni ix49543 (.Y (nx49542), .A0 (inputs_218__11), .A1 (inputs_219__11), 
             .S0 (nx24595)) ;
    mux21_ni ix49575 (.Y (nx49574), .A0 (nx49558), .A1 (nx49570), .S0 (nx23749)
             ) ;
    mux21_ni ix49559 (.Y (nx49558), .A0 (inputs_220__11), .A1 (inputs_221__11), 
             .S0 (nx24595)) ;
    mux21_ni ix49571 (.Y (nx49570), .A0 (inputs_222__11), .A1 (inputs_223__11), 
             .S0 (nx24595)) ;
    mux21_ni ix49875 (.Y (nx49874), .A0 (nx49868), .A1 (nx49790), .S0 (nx23171)
             ) ;
    oai21 ix49869 (.Y (nx49868), .A0 (nx22339), .A1 (nx18695), .B0 (nx18705)) ;
    mux21 ix18696 (.Y (nx18695), .A0 (nx49832), .A1 (nx49860), .S0 (nx23005)) ;
    mux21_ni ix49833 (.Y (nx49832), .A0 (nx49816), .A1 (nx49828), .S0 (nx23749)
             ) ;
    mux21_ni ix49817 (.Y (nx49816), .A0 (inputs_228__11), .A1 (inputs_229__11), 
             .S0 (nx24595)) ;
    mux21_ni ix49829 (.Y (nx49828), .A0 (inputs_230__11), .A1 (inputs_231__11), 
             .S0 (nx24595)) ;
    mux21_ni ix49861 (.Y (nx49860), .A0 (nx49844), .A1 (nx49856), .S0 (nx23749)
             ) ;
    mux21_ni ix49845 (.Y (nx49844), .A0 (inputs_244__11), .A1 (inputs_245__11), 
             .S0 (nx24595)) ;
    mux21_ni ix49857 (.Y (nx49856), .A0 (inputs_246__11), .A1 (inputs_247__11), 
             .S0 (nx24595)) ;
    nand04 ix18706 (.Y (nx18705), .A0 (nx22339), .A1 (nx23749), .A2 (nx24597), .A3 (
           nx49804)) ;
    mux21_ni ix49805 (.Y (nx49804), .A0 (inputs_227__11), .A1 (inputs_243__11), 
             .S0 (nx23005)) ;
    mux21_ni ix49791 (.Y (nx49790), .A0 (nx49726), .A1 (nx49786), .S0 (nx23005)
             ) ;
    mux21_ni ix49727 (.Y (nx49726), .A0 (nx49694), .A1 (nx49722), .S0 (nx23299)
             ) ;
    mux21_ni ix49695 (.Y (nx49694), .A0 (nx49678), .A1 (nx49690), .S0 (nx23749)
             ) ;
    mux21_ni ix49679 (.Y (nx49678), .A0 (inputs_232__11), .A1 (inputs_233__11), 
             .S0 (nx24597)) ;
    mux21_ni ix49691 (.Y (nx49690), .A0 (inputs_234__11), .A1 (inputs_235__11), 
             .S0 (nx24597)) ;
    mux21_ni ix49723 (.Y (nx49722), .A0 (nx49706), .A1 (nx49718), .S0 (nx23751)
             ) ;
    mux21_ni ix49707 (.Y (nx49706), .A0 (inputs_236__11), .A1 (inputs_237__11), 
             .S0 (nx24597)) ;
    mux21_ni ix49719 (.Y (nx49718), .A0 (inputs_238__11), .A1 (inputs_239__11), 
             .S0 (nx24597)) ;
    mux21_ni ix49787 (.Y (nx49786), .A0 (nx49754), .A1 (nx49782), .S0 (nx23299)
             ) ;
    mux21_ni ix49755 (.Y (nx49754), .A0 (nx49738), .A1 (nx49750), .S0 (nx23751)
             ) ;
    mux21_ni ix49739 (.Y (nx49738), .A0 (inputs_248__11), .A1 (inputs_249__11), 
             .S0 (nx24597)) ;
    mux21_ni ix49751 (.Y (nx49750), .A0 (inputs_250__11), .A1 (inputs_251__11), 
             .S0 (nx24597)) ;
    mux21_ni ix49783 (.Y (nx49782), .A0 (nx49766), .A1 (nx49778), .S0 (nx23751)
             ) ;
    mux21_ni ix49767 (.Y (nx49766), .A0 (inputs_252__11), .A1 (inputs_253__11), 
             .S0 (nx24599)) ;
    mux21_ni ix49779 (.Y (nx49778), .A0 (inputs_254__11), .A1 (inputs_255__11), 
             .S0 (nx24599)) ;
    oai21 ix54053 (.Y (\output [12]), .A0 (nx22223), .A1 (nx18733), .B0 (nx19088
          )) ;
    mux21 ix18734 (.Y (nx18733), .A0 (nx50734), .A1 (nx51578), .S0 (nx22437)) ;
    mux21_ni ix50735 (.Y (nx50734), .A0 (nx50310), .A1 (nx50730), .S0 (nx22505)
             ) ;
    mux21_ni ix50311 (.Y (nx50310), .A0 (nx50098), .A1 (nx50306), .S0 (nx22635)
             ) ;
    mux21_ni ix50099 (.Y (nx50098), .A0 (nx50092), .A1 (nx50014), .S0 (nx23171)
             ) ;
    oai21 ix50093 (.Y (nx50092), .A0 (nx22339), .A1 (nx18741), .B0 (nx18755)) ;
    mux21 ix18742 (.Y (nx18741), .A0 (nx50056), .A1 (nx50084), .S0 (nx23005)) ;
    mux21_ni ix50057 (.Y (nx50056), .A0 (nx50040), .A1 (nx50052), .S0 (nx23751)
             ) ;
    mux21_ni ix50041 (.Y (nx50040), .A0 (inputs_260__12), .A1 (inputs_261__12), 
             .S0 (nx24599)) ;
    mux21_ni ix50053 (.Y (nx50052), .A0 (inputs_262__12), .A1 (inputs_263__12), 
             .S0 (nx24599)) ;
    mux21_ni ix50085 (.Y (nx50084), .A0 (nx50068), .A1 (nx50080), .S0 (nx23751)
             ) ;
    mux21_ni ix50069 (.Y (nx50068), .A0 (inputs_276__12), .A1 (inputs_277__12), 
             .S0 (nx24599)) ;
    mux21_ni ix50081 (.Y (nx50080), .A0 (inputs_278__12), .A1 (inputs_279__12), 
             .S0 (nx24599)) ;
    nand04 ix18756 (.Y (nx18755), .A0 (nx22339), .A1 (nx23751), .A2 (nx24599), .A3 (
           nx50028)) ;
    mux21_ni ix50029 (.Y (nx50028), .A0 (inputs_259__12), .A1 (inputs_275__12), 
             .S0 (nx23005)) ;
    mux21_ni ix50015 (.Y (nx50014), .A0 (nx49950), .A1 (nx50010), .S0 (nx23005)
             ) ;
    mux21_ni ix49951 (.Y (nx49950), .A0 (nx49918), .A1 (nx49946), .S0 (nx23299)
             ) ;
    mux21_ni ix49919 (.Y (nx49918), .A0 (nx49902), .A1 (nx49914), .S0 (nx23751)
             ) ;
    mux21_ni ix49903 (.Y (nx49902), .A0 (inputs_264__12), .A1 (inputs_265__12), 
             .S0 (nx24601)) ;
    mux21_ni ix49915 (.Y (nx49914), .A0 (inputs_266__12), .A1 (inputs_267__12), 
             .S0 (nx24601)) ;
    mux21_ni ix49947 (.Y (nx49946), .A0 (nx49930), .A1 (nx49942), .S0 (nx23753)
             ) ;
    mux21_ni ix49931 (.Y (nx49930), .A0 (inputs_268__12), .A1 (inputs_269__12), 
             .S0 (nx24601)) ;
    mux21_ni ix49943 (.Y (nx49942), .A0 (inputs_270__12), .A1 (inputs_271__12), 
             .S0 (nx24601)) ;
    mux21_ni ix50011 (.Y (nx50010), .A0 (nx49978), .A1 (nx50006), .S0 (nx23301)
             ) ;
    mux21_ni ix49979 (.Y (nx49978), .A0 (nx49962), .A1 (nx49974), .S0 (nx23753)
             ) ;
    mux21_ni ix49963 (.Y (nx49962), .A0 (inputs_280__12), .A1 (inputs_281__12), 
             .S0 (nx24601)) ;
    mux21_ni ix49975 (.Y (nx49974), .A0 (inputs_282__12), .A1 (inputs_283__12), 
             .S0 (nx24601)) ;
    mux21_ni ix50007 (.Y (nx50006), .A0 (nx49990), .A1 (nx50002), .S0 (nx23753)
             ) ;
    mux21_ni ix49991 (.Y (nx49990), .A0 (inputs_284__12), .A1 (inputs_285__12), 
             .S0 (nx24601)) ;
    mux21_ni ix50003 (.Y (nx50002), .A0 (inputs_286__12), .A1 (inputs_287__12), 
             .S0 (nx24603)) ;
    mux21_ni ix50307 (.Y (nx50306), .A0 (nx50300), .A1 (nx50222), .S0 (nx23171)
             ) ;
    oai21 ix50301 (.Y (nx50300), .A0 (nx22339), .A1 (nx18785), .B0 (nx18797)) ;
    mux21 ix18786 (.Y (nx18785), .A0 (nx50264), .A1 (nx50292), .S0 (nx23007)) ;
    mux21_ni ix50265 (.Y (nx50264), .A0 (nx50248), .A1 (nx50260), .S0 (nx23753)
             ) ;
    mux21_ni ix50249 (.Y (nx50248), .A0 (inputs_292__12), .A1 (inputs_293__12), 
             .S0 (nx24603)) ;
    mux21_ni ix50261 (.Y (nx50260), .A0 (inputs_294__12), .A1 (inputs_295__12), 
             .S0 (nx24603)) ;
    mux21_ni ix50293 (.Y (nx50292), .A0 (nx50276), .A1 (nx50288), .S0 (nx23753)
             ) ;
    mux21_ni ix50277 (.Y (nx50276), .A0 (inputs_308__12), .A1 (inputs_309__12), 
             .S0 (nx24603)) ;
    mux21_ni ix50289 (.Y (nx50288), .A0 (inputs_310__12), .A1 (inputs_311__12), 
             .S0 (nx24603)) ;
    nand04 ix18798 (.Y (nx18797), .A0 (nx22341), .A1 (nx23753), .A2 (nx24603), .A3 (
           nx50236)) ;
    mux21_ni ix50237 (.Y (nx50236), .A0 (inputs_291__12), .A1 (inputs_307__12), 
             .S0 (nx23007)) ;
    mux21_ni ix50223 (.Y (nx50222), .A0 (nx50158), .A1 (nx50218), .S0 (nx23007)
             ) ;
    mux21_ni ix50159 (.Y (nx50158), .A0 (nx50126), .A1 (nx50154), .S0 (nx23301)
             ) ;
    mux21_ni ix50127 (.Y (nx50126), .A0 (nx50110), .A1 (nx50122), .S0 (nx23753)
             ) ;
    mux21_ni ix50111 (.Y (nx50110), .A0 (inputs_296__12), .A1 (inputs_297__12), 
             .S0 (nx24603)) ;
    mux21_ni ix50123 (.Y (nx50122), .A0 (inputs_298__12), .A1 (inputs_299__12), 
             .S0 (nx24605)) ;
    mux21_ni ix50155 (.Y (nx50154), .A0 (nx50138), .A1 (nx50150), .S0 (nx23755)
             ) ;
    mux21_ni ix50139 (.Y (nx50138), .A0 (inputs_300__12), .A1 (inputs_301__12), 
             .S0 (nx24605)) ;
    mux21_ni ix50151 (.Y (nx50150), .A0 (inputs_302__12), .A1 (inputs_303__12), 
             .S0 (nx24605)) ;
    mux21_ni ix50219 (.Y (nx50218), .A0 (nx50186), .A1 (nx50214), .S0 (nx23301)
             ) ;
    mux21_ni ix50187 (.Y (nx50186), .A0 (nx50170), .A1 (nx50182), .S0 (nx23755)
             ) ;
    mux21_ni ix50171 (.Y (nx50170), .A0 (inputs_312__12), .A1 (inputs_313__12), 
             .S0 (nx24605)) ;
    mux21_ni ix50183 (.Y (nx50182), .A0 (inputs_314__12), .A1 (inputs_315__12), 
             .S0 (nx24605)) ;
    mux21_ni ix50215 (.Y (nx50214), .A0 (nx50198), .A1 (nx50210), .S0 (nx23755)
             ) ;
    mux21_ni ix50199 (.Y (nx50198), .A0 (inputs_316__12), .A1 (inputs_317__12), 
             .S0 (nx24605)) ;
    mux21_ni ix50211 (.Y (nx50210), .A0 (inputs_318__12), .A1 (inputs_319__12), 
             .S0 (nx24605)) ;
    mux21_ni ix50731 (.Y (nx50730), .A0 (nx50518), .A1 (nx50726), .S0 (nx22637)
             ) ;
    mux21_ni ix50519 (.Y (nx50518), .A0 (nx50512), .A1 (nx50434), .S0 (nx23171)
             ) ;
    oai21 ix50513 (.Y (nx50512), .A0 (nx22341), .A1 (nx18831), .B0 (nx18843)) ;
    mux21 ix18832 (.Y (nx18831), .A0 (nx50476), .A1 (nx50504), .S0 (nx23007)) ;
    mux21_ni ix50477 (.Y (nx50476), .A0 (nx50460), .A1 (nx50472), .S0 (nx23755)
             ) ;
    mux21_ni ix50461 (.Y (nx50460), .A0 (inputs_324__12), .A1 (inputs_325__12), 
             .S0 (nx24607)) ;
    mux21_ni ix50473 (.Y (nx50472), .A0 (inputs_326__12), .A1 (inputs_327__12), 
             .S0 (nx24607)) ;
    mux21_ni ix50505 (.Y (nx50504), .A0 (nx50488), .A1 (nx50500), .S0 (nx23755)
             ) ;
    mux21_ni ix50489 (.Y (nx50488), .A0 (inputs_340__12), .A1 (inputs_341__12), 
             .S0 (nx24607)) ;
    mux21_ni ix50501 (.Y (nx50500), .A0 (inputs_342__12), .A1 (inputs_343__12), 
             .S0 (nx24607)) ;
    nand04 ix18844 (.Y (nx18843), .A0 (nx22341), .A1 (nx23755), .A2 (nx24607), .A3 (
           nx50448)) ;
    mux21_ni ix50449 (.Y (nx50448), .A0 (inputs_323__12), .A1 (inputs_339__12), 
             .S0 (nx23007)) ;
    mux21_ni ix50435 (.Y (nx50434), .A0 (nx50370), .A1 (nx50430), .S0 (nx23007)
             ) ;
    mux21_ni ix50371 (.Y (nx50370), .A0 (nx50338), .A1 (nx50366), .S0 (nx23301)
             ) ;
    mux21_ni ix50339 (.Y (nx50338), .A0 (nx50322), .A1 (nx50334), .S0 (nx23755)
             ) ;
    mux21_ni ix50323 (.Y (nx50322), .A0 (inputs_328__12), .A1 (inputs_329__12), 
             .S0 (nx24607)) ;
    mux21_ni ix50335 (.Y (nx50334), .A0 (inputs_330__12), .A1 (inputs_331__12), 
             .S0 (nx24607)) ;
    mux21_ni ix50367 (.Y (nx50366), .A0 (nx50350), .A1 (nx50362), .S0 (nx23757)
             ) ;
    mux21_ni ix50351 (.Y (nx50350), .A0 (inputs_332__12), .A1 (inputs_333__12), 
             .S0 (nx24609)) ;
    mux21_ni ix50363 (.Y (nx50362), .A0 (inputs_334__12), .A1 (inputs_335__12), 
             .S0 (nx24609)) ;
    mux21_ni ix50431 (.Y (nx50430), .A0 (nx50398), .A1 (nx50426), .S0 (nx23301)
             ) ;
    mux21_ni ix50399 (.Y (nx50398), .A0 (nx50382), .A1 (nx50394), .S0 (nx23757)
             ) ;
    mux21_ni ix50383 (.Y (nx50382), .A0 (inputs_344__12), .A1 (inputs_345__12), 
             .S0 (nx24609)) ;
    mux21_ni ix50395 (.Y (nx50394), .A0 (inputs_346__12), .A1 (inputs_347__12), 
             .S0 (nx24609)) ;
    mux21_ni ix50427 (.Y (nx50426), .A0 (nx50410), .A1 (nx50422), .S0 (nx23757)
             ) ;
    mux21_ni ix50411 (.Y (nx50410), .A0 (inputs_348__12), .A1 (inputs_349__12), 
             .S0 (nx24609)) ;
    mux21_ni ix50423 (.Y (nx50422), .A0 (inputs_350__12), .A1 (inputs_351__12), 
             .S0 (nx24609)) ;
    mux21_ni ix50727 (.Y (nx50726), .A0 (nx50720), .A1 (nx50642), .S0 (nx23171)
             ) ;
    oai21 ix50721 (.Y (nx50720), .A0 (nx22341), .A1 (nx18873), .B0 (nx18887)) ;
    mux21 ix18874 (.Y (nx18873), .A0 (nx50684), .A1 (nx50712), .S0 (nx23007)) ;
    mux21_ni ix50685 (.Y (nx50684), .A0 (nx50668), .A1 (nx50680), .S0 (nx23757)
             ) ;
    mux21_ni ix50669 (.Y (nx50668), .A0 (inputs_356__12), .A1 (inputs_357__12), 
             .S0 (nx24609)) ;
    mux21_ni ix50681 (.Y (nx50680), .A0 (inputs_358__12), .A1 (inputs_359__12), 
             .S0 (nx24611)) ;
    mux21_ni ix50713 (.Y (nx50712), .A0 (nx50696), .A1 (nx50708), .S0 (nx23757)
             ) ;
    mux21_ni ix50697 (.Y (nx50696), .A0 (inputs_372__12), .A1 (inputs_373__12), 
             .S0 (nx24611)) ;
    mux21_ni ix50709 (.Y (nx50708), .A0 (inputs_374__12), .A1 (inputs_375__12), 
             .S0 (nx24611)) ;
    nand04 ix18888 (.Y (nx18887), .A0 (nx22341), .A1 (nx23757), .A2 (nx24611), .A3 (
           nx50656)) ;
    mux21_ni ix50657 (.Y (nx50656), .A0 (inputs_355__12), .A1 (inputs_371__12), 
             .S0 (nx23009)) ;
    mux21_ni ix50643 (.Y (nx50642), .A0 (nx50578), .A1 (nx50638), .S0 (nx23009)
             ) ;
    mux21_ni ix50579 (.Y (nx50578), .A0 (nx50546), .A1 (nx50574), .S0 (nx23301)
             ) ;
    mux21_ni ix50547 (.Y (nx50546), .A0 (nx50530), .A1 (nx50542), .S0 (nx23757)
             ) ;
    mux21_ni ix50531 (.Y (nx50530), .A0 (inputs_360__12), .A1 (inputs_361__12), 
             .S0 (nx24611)) ;
    mux21_ni ix50543 (.Y (nx50542), .A0 (inputs_362__12), .A1 (inputs_363__12), 
             .S0 (nx24611)) ;
    mux21_ni ix50575 (.Y (nx50574), .A0 (nx50558), .A1 (nx50570), .S0 (nx23759)
             ) ;
    mux21_ni ix50559 (.Y (nx50558), .A0 (inputs_364__12), .A1 (inputs_365__12), 
             .S0 (nx24611)) ;
    mux21_ni ix50571 (.Y (nx50570), .A0 (inputs_366__12), .A1 (inputs_367__12), 
             .S0 (nx24613)) ;
    mux21_ni ix50639 (.Y (nx50638), .A0 (nx50606), .A1 (nx50634), .S0 (nx23301)
             ) ;
    mux21_ni ix50607 (.Y (nx50606), .A0 (nx50590), .A1 (nx50602), .S0 (nx23759)
             ) ;
    mux21_ni ix50591 (.Y (nx50590), .A0 (inputs_376__12), .A1 (inputs_377__12), 
             .S0 (nx24613)) ;
    mux21_ni ix50603 (.Y (nx50602), .A0 (inputs_378__12), .A1 (inputs_379__12), 
             .S0 (nx24613)) ;
    mux21_ni ix50635 (.Y (nx50634), .A0 (nx50618), .A1 (nx50630), .S0 (nx23759)
             ) ;
    mux21_ni ix50619 (.Y (nx50618), .A0 (inputs_380__12), .A1 (inputs_381__12), 
             .S0 (nx24613)) ;
    mux21_ni ix50631 (.Y (nx50630), .A0 (inputs_382__12), .A1 (inputs_383__12), 
             .S0 (nx24613)) ;
    mux21_ni ix51579 (.Y (nx51578), .A0 (nx51154), .A1 (nx51574), .S0 (nx22505)
             ) ;
    mux21_ni ix51155 (.Y (nx51154), .A0 (nx50942), .A1 (nx51150), .S0 (nx22637)
             ) ;
    mux21_ni ix50943 (.Y (nx50942), .A0 (nx50936), .A1 (nx50858), .S0 (nx23173)
             ) ;
    oai21 ix50937 (.Y (nx50936), .A0 (nx22341), .A1 (nx18919), .B0 (nx18931)) ;
    mux21 ix18920 (.Y (nx18919), .A0 (nx50900), .A1 (nx50928), .S0 (nx23009)) ;
    mux21_ni ix50901 (.Y (nx50900), .A0 (nx50884), .A1 (nx50896), .S0 (nx23759)
             ) ;
    mux21_ni ix50885 (.Y (nx50884), .A0 (inputs_388__12), .A1 (inputs_389__12), 
             .S0 (nx24613)) ;
    mux21_ni ix50897 (.Y (nx50896), .A0 (inputs_390__12), .A1 (inputs_391__12), 
             .S0 (nx24613)) ;
    mux21_ni ix50929 (.Y (nx50928), .A0 (nx50912), .A1 (nx50924), .S0 (nx23759)
             ) ;
    mux21_ni ix50913 (.Y (nx50912), .A0 (inputs_404__12), .A1 (inputs_405__12), 
             .S0 (nx24615)) ;
    mux21_ni ix50925 (.Y (nx50924), .A0 (inputs_406__12), .A1 (inputs_407__12), 
             .S0 (nx24615)) ;
    nand04 ix18932 (.Y (nx18931), .A0 (nx22341), .A1 (nx23759), .A2 (nx24615), .A3 (
           nx50872)) ;
    mux21_ni ix50873 (.Y (nx50872), .A0 (inputs_387__12), .A1 (inputs_403__12), 
             .S0 (nx23009)) ;
    mux21_ni ix50859 (.Y (nx50858), .A0 (nx50794), .A1 (nx50854), .S0 (nx23009)
             ) ;
    mux21_ni ix50795 (.Y (nx50794), .A0 (nx50762), .A1 (nx50790), .S0 (nx23303)
             ) ;
    mux21_ni ix50763 (.Y (nx50762), .A0 (nx50746), .A1 (nx50758), .S0 (nx23759)
             ) ;
    mux21_ni ix50747 (.Y (nx50746), .A0 (inputs_392__12), .A1 (inputs_393__12), 
             .S0 (nx24615)) ;
    mux21_ni ix50759 (.Y (nx50758), .A0 (inputs_394__12), .A1 (inputs_395__12), 
             .S0 (nx24615)) ;
    mux21_ni ix50791 (.Y (nx50790), .A0 (nx50774), .A1 (nx50786), .S0 (nx23761)
             ) ;
    mux21_ni ix50775 (.Y (nx50774), .A0 (inputs_396__12), .A1 (inputs_397__12), 
             .S0 (nx24615)) ;
    mux21_ni ix50787 (.Y (nx50786), .A0 (inputs_398__12), .A1 (inputs_399__12), 
             .S0 (nx24615)) ;
    mux21_ni ix50855 (.Y (nx50854), .A0 (nx50822), .A1 (nx50850), .S0 (nx23303)
             ) ;
    mux21_ni ix50823 (.Y (nx50822), .A0 (nx50806), .A1 (nx50818), .S0 (nx23761)
             ) ;
    mux21_ni ix50807 (.Y (nx50806), .A0 (inputs_408__12), .A1 (inputs_409__12), 
             .S0 (nx24617)) ;
    mux21_ni ix50819 (.Y (nx50818), .A0 (inputs_410__12), .A1 (inputs_411__12), 
             .S0 (nx24617)) ;
    mux21_ni ix50851 (.Y (nx50850), .A0 (nx50834), .A1 (nx50846), .S0 (nx23761)
             ) ;
    mux21_ni ix50835 (.Y (nx50834), .A0 (inputs_412__12), .A1 (inputs_413__12), 
             .S0 (nx24617)) ;
    mux21_ni ix50847 (.Y (nx50846), .A0 (inputs_414__12), .A1 (inputs_415__12), 
             .S0 (nx24617)) ;
    mux21_ni ix51151 (.Y (nx51150), .A0 (nx51144), .A1 (nx51066), .S0 (nx23173)
             ) ;
    oai21 ix51145 (.Y (nx51144), .A0 (nx22343), .A1 (nx18963), .B0 (nx18975)) ;
    mux21 ix18964 (.Y (nx18963), .A0 (nx51108), .A1 (nx51136), .S0 (nx23009)) ;
    mux21_ni ix51109 (.Y (nx51108), .A0 (nx51092), .A1 (nx51104), .S0 (nx23761)
             ) ;
    mux21_ni ix51093 (.Y (nx51092), .A0 (inputs_420__12), .A1 (inputs_421__12), 
             .S0 (nx24617)) ;
    mux21_ni ix51105 (.Y (nx51104), .A0 (inputs_422__12), .A1 (inputs_423__12), 
             .S0 (nx24617)) ;
    mux21_ni ix51137 (.Y (nx51136), .A0 (nx51120), .A1 (nx51132), .S0 (nx23761)
             ) ;
    mux21_ni ix51121 (.Y (nx51120), .A0 (inputs_436__12), .A1 (inputs_437__12), 
             .S0 (nx24617)) ;
    mux21_ni ix51133 (.Y (nx51132), .A0 (inputs_438__12), .A1 (inputs_439__12), 
             .S0 (nx24619)) ;
    nand04 ix18976 (.Y (nx18975), .A0 (nx22343), .A1 (nx23761), .A2 (nx24619), .A3 (
           nx51080)) ;
    mux21_ni ix51081 (.Y (nx51080), .A0 (inputs_419__12), .A1 (inputs_435__12), 
             .S0 (nx23009)) ;
    mux21_ni ix51067 (.Y (nx51066), .A0 (nx51002), .A1 (nx51062), .S0 (nx23011)
             ) ;
    mux21_ni ix51003 (.Y (nx51002), .A0 (nx50970), .A1 (nx50998), .S0 (nx23303)
             ) ;
    mux21_ni ix50971 (.Y (nx50970), .A0 (nx50954), .A1 (nx50966), .S0 (nx23761)
             ) ;
    mux21_ni ix50955 (.Y (nx50954), .A0 (inputs_424__12), .A1 (inputs_425__12), 
             .S0 (nx24619)) ;
    mux21_ni ix50967 (.Y (nx50966), .A0 (inputs_426__12), .A1 (inputs_427__12), 
             .S0 (nx24619)) ;
    mux21_ni ix50999 (.Y (nx50998), .A0 (nx50982), .A1 (nx50994), .S0 (nx23763)
             ) ;
    mux21_ni ix50983 (.Y (nx50982), .A0 (inputs_428__12), .A1 (inputs_429__12), 
             .S0 (nx24619)) ;
    mux21_ni ix50995 (.Y (nx50994), .A0 (inputs_430__12), .A1 (inputs_431__12), 
             .S0 (nx24619)) ;
    mux21_ni ix51063 (.Y (nx51062), .A0 (nx51030), .A1 (nx51058), .S0 (nx23303)
             ) ;
    mux21_ni ix51031 (.Y (nx51030), .A0 (nx51014), .A1 (nx51026), .S0 (nx23763)
             ) ;
    mux21_ni ix51015 (.Y (nx51014), .A0 (inputs_440__12), .A1 (inputs_441__12), 
             .S0 (nx24619)) ;
    mux21_ni ix51027 (.Y (nx51026), .A0 (inputs_442__12), .A1 (inputs_443__12), 
             .S0 (nx24621)) ;
    mux21_ni ix51059 (.Y (nx51058), .A0 (nx51042), .A1 (nx51054), .S0 (nx23763)
             ) ;
    mux21_ni ix51043 (.Y (nx51042), .A0 (inputs_444__12), .A1 (inputs_445__12), 
             .S0 (nx24621)) ;
    mux21_ni ix51055 (.Y (nx51054), .A0 (inputs_446__12), .A1 (inputs_447__12), 
             .S0 (nx24621)) ;
    mux21_ni ix51575 (.Y (nx51574), .A0 (nx51362), .A1 (nx51570), .S0 (nx22637)
             ) ;
    mux21_ni ix51363 (.Y (nx51362), .A0 (nx51356), .A1 (nx51278), .S0 (nx23173)
             ) ;
    oai21 ix51357 (.Y (nx51356), .A0 (nx22343), .A1 (nx19007), .B0 (nx19017)) ;
    mux21 ix19008 (.Y (nx19007), .A0 (nx51320), .A1 (nx51348), .S0 (nx23011)) ;
    mux21_ni ix51321 (.Y (nx51320), .A0 (nx51304), .A1 (nx51316), .S0 (nx23763)
             ) ;
    mux21_ni ix51305 (.Y (nx51304), .A0 (inputs_452__12), .A1 (inputs_453__12), 
             .S0 (nx24621)) ;
    mux21_ni ix51317 (.Y (nx51316), .A0 (inputs_454__12), .A1 (inputs_455__12), 
             .S0 (nx24621)) ;
    mux21_ni ix51349 (.Y (nx51348), .A0 (nx51332), .A1 (nx51344), .S0 (nx23763)
             ) ;
    mux21_ni ix51333 (.Y (nx51332), .A0 (inputs_468__12), .A1 (inputs_469__12), 
             .S0 (nx24621)) ;
    mux21_ni ix51345 (.Y (nx51344), .A0 (inputs_470__12), .A1 (inputs_471__12), 
             .S0 (nx24621)) ;
    nand04 ix19018 (.Y (nx19017), .A0 (nx22343), .A1 (nx23763), .A2 (nx24623), .A3 (
           nx51292)) ;
    mux21_ni ix51293 (.Y (nx51292), .A0 (inputs_451__12), .A1 (inputs_467__12), 
             .S0 (nx23011)) ;
    mux21_ni ix51279 (.Y (nx51278), .A0 (nx51214), .A1 (nx51274), .S0 (nx23011)
             ) ;
    mux21_ni ix51215 (.Y (nx51214), .A0 (nx51182), .A1 (nx51210), .S0 (nx23303)
             ) ;
    mux21_ni ix51183 (.Y (nx51182), .A0 (nx51166), .A1 (nx51178), .S0 (nx23763)
             ) ;
    mux21_ni ix51167 (.Y (nx51166), .A0 (inputs_456__12), .A1 (inputs_457__12), 
             .S0 (nx24623)) ;
    mux21_ni ix51179 (.Y (nx51178), .A0 (inputs_458__12), .A1 (inputs_459__12), 
             .S0 (nx24623)) ;
    mux21_ni ix51211 (.Y (nx51210), .A0 (nx51194), .A1 (nx51206), .S0 (nx23765)
             ) ;
    mux21_ni ix51195 (.Y (nx51194), .A0 (inputs_460__12), .A1 (inputs_461__12), 
             .S0 (nx24623)) ;
    mux21_ni ix51207 (.Y (nx51206), .A0 (inputs_462__12), .A1 (inputs_463__12), 
             .S0 (nx24623)) ;
    mux21_ni ix51275 (.Y (nx51274), .A0 (nx51242), .A1 (nx51270), .S0 (nx23303)
             ) ;
    mux21_ni ix51243 (.Y (nx51242), .A0 (nx51226), .A1 (nx51238), .S0 (nx23765)
             ) ;
    mux21_ni ix51227 (.Y (nx51226), .A0 (inputs_472__12), .A1 (inputs_473__12), 
             .S0 (nx24623)) ;
    mux21_ni ix51239 (.Y (nx51238), .A0 (inputs_474__12), .A1 (inputs_475__12), 
             .S0 (nx24623)) ;
    mux21_ni ix51271 (.Y (nx51270), .A0 (nx51254), .A1 (nx51266), .S0 (nx23765)
             ) ;
    mux21_ni ix51255 (.Y (nx51254), .A0 (inputs_476__12), .A1 (inputs_477__12), 
             .S0 (nx24625)) ;
    mux21_ni ix51267 (.Y (nx51266), .A0 (inputs_478__12), .A1 (inputs_479__12), 
             .S0 (nx24625)) ;
    mux21_ni ix51571 (.Y (nx51570), .A0 (nx51564), .A1 (nx51486), .S0 (nx23173)
             ) ;
    oai21 ix51565 (.Y (nx51564), .A0 (nx22343), .A1 (nx19047), .B0 (nx19057)) ;
    mux21 ix19048 (.Y (nx19047), .A0 (nx51528), .A1 (nx51556), .S0 (nx23011)) ;
    mux21_ni ix51529 (.Y (nx51528), .A0 (nx51512), .A1 (nx51524), .S0 (nx23765)
             ) ;
    mux21_ni ix51513 (.Y (nx51512), .A0 (inputs_484__12), .A1 (inputs_485__12), 
             .S0 (nx24625)) ;
    mux21_ni ix51525 (.Y (nx51524), .A0 (inputs_486__12), .A1 (inputs_487__12), 
             .S0 (nx24625)) ;
    mux21_ni ix51557 (.Y (nx51556), .A0 (nx51540), .A1 (nx51552), .S0 (nx23765)
             ) ;
    mux21_ni ix51541 (.Y (nx51540), .A0 (inputs_500__12), .A1 (inputs_501__12), 
             .S0 (nx24625)) ;
    mux21_ni ix51553 (.Y (nx51552), .A0 (inputs_502__12), .A1 (inputs_503__12), 
             .S0 (nx24625)) ;
    nand04 ix19058 (.Y (nx19057), .A0 (nx22343), .A1 (nx23765), .A2 (nx24625), .A3 (
           nx51500)) ;
    mux21_ni ix51501 (.Y (nx51500), .A0 (inputs_483__12), .A1 (inputs_499__12), 
             .S0 (nx23011)) ;
    mux21_ni ix51487 (.Y (nx51486), .A0 (nx51422), .A1 (nx51482), .S0 (nx23011)
             ) ;
    mux21_ni ix51423 (.Y (nx51422), .A0 (nx51390), .A1 (nx51418), .S0 (nx23303)
             ) ;
    mux21_ni ix51391 (.Y (nx51390), .A0 (nx51374), .A1 (nx51386), .S0 (nx23765)
             ) ;
    mux21_ni ix51375 (.Y (nx51374), .A0 (inputs_488__12), .A1 (inputs_489__12), 
             .S0 (nx24627)) ;
    mux21_ni ix51387 (.Y (nx51386), .A0 (inputs_490__12), .A1 (inputs_491__12), 
             .S0 (nx24627)) ;
    mux21_ni ix51419 (.Y (nx51418), .A0 (nx51402), .A1 (nx51414), .S0 (nx23767)
             ) ;
    mux21_ni ix51403 (.Y (nx51402), .A0 (inputs_492__12), .A1 (inputs_493__12), 
             .S0 (nx24627)) ;
    mux21_ni ix51415 (.Y (nx51414), .A0 (inputs_494__12), .A1 (inputs_495__12), 
             .S0 (nx24627)) ;
    mux21_ni ix51483 (.Y (nx51482), .A0 (nx51450), .A1 (nx51478), .S0 (nx23305)
             ) ;
    mux21_ni ix51451 (.Y (nx51450), .A0 (nx51434), .A1 (nx51446), .S0 (nx23767)
             ) ;
    mux21_ni ix51435 (.Y (nx51434), .A0 (inputs_504__12), .A1 (inputs_505__12), 
             .S0 (nx24627)) ;
    mux21_ni ix51447 (.Y (nx51446), .A0 (inputs_506__12), .A1 (inputs_507__12), 
             .S0 (nx24627)) ;
    mux21_ni ix51479 (.Y (nx51478), .A0 (nx51462), .A1 (nx51474), .S0 (nx23767)
             ) ;
    mux21_ni ix51463 (.Y (nx51462), .A0 (inputs_508__12), .A1 (inputs_509__12), 
             .S0 (nx24627)) ;
    mux21_ni ix51475 (.Y (nx51474), .A0 (inputs_510__12), .A1 (inputs_511__12), 
             .S0 (nx24629)) ;
    aoi32 ix19089 (.Y (nx19088), .A0 (nx52348), .A1 (nx24839), .A2 (nx22343), .B0 (
          nx22223), .B1 (nx54044)) ;
    oai21 ix52349 (.Y (nx52348), .A0 (nx23767), .A1 (nx19091), .B0 (nx19191)) ;
    mux21 ix19092 (.Y (nx19091), .A0 (nx52086), .A1 (nx52338), .S0 (nx24629)) ;
    mux21_ni ix52087 (.Y (nx52086), .A0 (nx51958), .A1 (nx52082), .S0 (nx22403)
             ) ;
    mux21_ni ix51959 (.Y (nx51958), .A0 (nx51894), .A1 (nx51954), .S0 (nx22437)
             ) ;
    mux21_ni ix51895 (.Y (nx51894), .A0 (nx51862), .A1 (nx51890), .S0 (nx22505)
             ) ;
    mux21_ni ix51863 (.Y (nx51862), .A0 (nx51846), .A1 (nx51858), .S0 (nx22637)
             ) ;
    mux21_ni ix51847 (.Y (nx51846), .A0 (inputs_0__12), .A1 (inputs_16__12), .S0 (
             nx23013)) ;
    mux21_ni ix51859 (.Y (nx51858), .A0 (inputs_32__12), .A1 (inputs_48__12), .S0 (
             nx23013)) ;
    mux21_ni ix51891 (.Y (nx51890), .A0 (nx51874), .A1 (nx51886), .S0 (nx22637)
             ) ;
    mux21_ni ix51875 (.Y (nx51874), .A0 (inputs_64__12), .A1 (inputs_80__12), .S0 (
             nx23013)) ;
    mux21_ni ix51887 (.Y (nx51886), .A0 (inputs_96__12), .A1 (inputs_112__12), .S0 (
             nx23013)) ;
    mux21_ni ix51955 (.Y (nx51954), .A0 (nx51922), .A1 (nx51950), .S0 (nx22505)
             ) ;
    mux21_ni ix51923 (.Y (nx51922), .A0 (nx51906), .A1 (nx51918), .S0 (nx22637)
             ) ;
    mux21_ni ix51907 (.Y (nx51906), .A0 (inputs_128__12), .A1 (inputs_144__12), 
             .S0 (nx23013)) ;
    mux21_ni ix51919 (.Y (nx51918), .A0 (inputs_160__12), .A1 (inputs_176__12), 
             .S0 (nx23013)) ;
    mux21_ni ix51951 (.Y (nx51950), .A0 (nx51934), .A1 (nx51946), .S0 (nx22637)
             ) ;
    mux21_ni ix51935 (.Y (nx51934), .A0 (inputs_192__12), .A1 (inputs_208__12), 
             .S0 (nx23013)) ;
    mux21_ni ix51947 (.Y (nx51946), .A0 (inputs_224__12), .A1 (inputs_240__12), 
             .S0 (nx23015)) ;
    mux21_ni ix52083 (.Y (nx52082), .A0 (nx52018), .A1 (nx52078), .S0 (nx22439)
             ) ;
    mux21_ni ix52019 (.Y (nx52018), .A0 (nx51986), .A1 (nx52014), .S0 (nx22507)
             ) ;
    mux21_ni ix51987 (.Y (nx51986), .A0 (nx51970), .A1 (nx51982), .S0 (nx22639)
             ) ;
    mux21_ni ix51971 (.Y (nx51970), .A0 (inputs_256__12), .A1 (inputs_272__12), 
             .S0 (nx23015)) ;
    mux21_ni ix51983 (.Y (nx51982), .A0 (inputs_288__12), .A1 (inputs_304__12), 
             .S0 (nx23015)) ;
    mux21_ni ix52015 (.Y (nx52014), .A0 (nx51998), .A1 (nx52010), .S0 (nx22639)
             ) ;
    mux21_ni ix51999 (.Y (nx51998), .A0 (inputs_320__12), .A1 (inputs_336__12), 
             .S0 (nx23015)) ;
    mux21_ni ix52011 (.Y (nx52010), .A0 (inputs_352__12), .A1 (inputs_368__12), 
             .S0 (nx23015)) ;
    mux21_ni ix52079 (.Y (nx52078), .A0 (nx52046), .A1 (nx52074), .S0 (nx22507)
             ) ;
    mux21_ni ix52047 (.Y (nx52046), .A0 (nx52030), .A1 (nx52042), .S0 (nx22639)
             ) ;
    mux21_ni ix52031 (.Y (nx52030), .A0 (inputs_384__12), .A1 (inputs_400__12), 
             .S0 (nx23015)) ;
    mux21_ni ix52043 (.Y (nx52042), .A0 (inputs_416__12), .A1 (inputs_432__12), 
             .S0 (nx23015)) ;
    mux21_ni ix52075 (.Y (nx52074), .A0 (nx52058), .A1 (nx52070), .S0 (nx22639)
             ) ;
    mux21_ni ix52059 (.Y (nx52058), .A0 (inputs_448__12), .A1 (inputs_464__12), 
             .S0 (nx23017)) ;
    mux21_ni ix52071 (.Y (nx52070), .A0 (inputs_480__12), .A1 (inputs_496__12), 
             .S0 (nx23017)) ;
    mux21_ni ix52339 (.Y (nx52338), .A0 (nx52210), .A1 (nx52334), .S0 (nx22403)
             ) ;
    mux21_ni ix52211 (.Y (nx52210), .A0 (nx52146), .A1 (nx52206), .S0 (nx22439)
             ) ;
    mux21_ni ix52147 (.Y (nx52146), .A0 (nx52114), .A1 (nx52142), .S0 (nx22507)
             ) ;
    mux21_ni ix52115 (.Y (nx52114), .A0 (nx52098), .A1 (nx52110), .S0 (nx22639)
             ) ;
    mux21_ni ix52099 (.Y (nx52098), .A0 (inputs_1__12), .A1 (inputs_17__12), .S0 (
             nx23017)) ;
    mux21_ni ix52111 (.Y (nx52110), .A0 (inputs_33__12), .A1 (inputs_49__12), .S0 (
             nx23017)) ;
    mux21_ni ix52143 (.Y (nx52142), .A0 (nx52126), .A1 (nx52138), .S0 (nx22639)
             ) ;
    mux21_ni ix52127 (.Y (nx52126), .A0 (inputs_65__12), .A1 (inputs_81__12), .S0 (
             nx23017)) ;
    mux21_ni ix52139 (.Y (nx52138), .A0 (inputs_97__12), .A1 (inputs_113__12), .S0 (
             nx23017)) ;
    mux21_ni ix52207 (.Y (nx52206), .A0 (nx52174), .A1 (nx52202), .S0 (nx22507)
             ) ;
    mux21_ni ix52175 (.Y (nx52174), .A0 (nx52158), .A1 (nx52170), .S0 (nx22639)
             ) ;
    mux21_ni ix52159 (.Y (nx52158), .A0 (inputs_129__12), .A1 (inputs_145__12), 
             .S0 (nx23017)) ;
    mux21_ni ix52171 (.Y (nx52170), .A0 (inputs_161__12), .A1 (inputs_177__12), 
             .S0 (nx23019)) ;
    mux21_ni ix52203 (.Y (nx52202), .A0 (nx52186), .A1 (nx52198), .S0 (nx22641)
             ) ;
    mux21_ni ix52187 (.Y (nx52186), .A0 (inputs_193__12), .A1 (inputs_209__12), 
             .S0 (nx23019)) ;
    mux21_ni ix52199 (.Y (nx52198), .A0 (inputs_225__12), .A1 (inputs_241__12), 
             .S0 (nx23019)) ;
    mux21_ni ix52335 (.Y (nx52334), .A0 (nx52270), .A1 (nx52330), .S0 (nx22439)
             ) ;
    mux21_ni ix52271 (.Y (nx52270), .A0 (nx52238), .A1 (nx52266), .S0 (nx22507)
             ) ;
    mux21_ni ix52239 (.Y (nx52238), .A0 (nx52222), .A1 (nx52234), .S0 (nx22641)
             ) ;
    mux21_ni ix52223 (.Y (nx52222), .A0 (inputs_257__12), .A1 (inputs_273__12), 
             .S0 (nx23019)) ;
    mux21_ni ix52235 (.Y (nx52234), .A0 (inputs_289__12), .A1 (inputs_305__12), 
             .S0 (nx23019)) ;
    mux21_ni ix52267 (.Y (nx52266), .A0 (nx52250), .A1 (nx52262), .S0 (nx22641)
             ) ;
    mux21_ni ix52251 (.Y (nx52250), .A0 (inputs_321__12), .A1 (inputs_337__12), 
             .S0 (nx23019)) ;
    mux21_ni ix52263 (.Y (nx52262), .A0 (inputs_353__12), .A1 (inputs_369__12), 
             .S0 (nx23019)) ;
    mux21_ni ix52331 (.Y (nx52330), .A0 (nx52298), .A1 (nx52326), .S0 (nx22507)
             ) ;
    mux21_ni ix52299 (.Y (nx52298), .A0 (nx52282), .A1 (nx52294), .S0 (nx22641)
             ) ;
    mux21_ni ix52283 (.Y (nx52282), .A0 (inputs_385__12), .A1 (inputs_401__12), 
             .S0 (nx23021)) ;
    mux21_ni ix52295 (.Y (nx52294), .A0 (inputs_417__12), .A1 (inputs_433__12), 
             .S0 (nx23021)) ;
    mux21_ni ix52327 (.Y (nx52326), .A0 (nx52310), .A1 (nx52322), .S0 (nx22641)
             ) ;
    mux21_ni ix52311 (.Y (nx52310), .A0 (inputs_449__12), .A1 (inputs_465__12), 
             .S0 (nx23021)) ;
    mux21_ni ix52323 (.Y (nx52322), .A0 (inputs_481__12), .A1 (inputs_497__12), 
             .S0 (nx23021)) ;
    nand03 ix19192 (.Y (nx19191), .A0 (nx51832), .A1 (nx23767), .A2 (nx22381)) ;
    mux21_ni ix51833 (.Y (nx51832), .A0 (nx51704), .A1 (nx51828), .S0 (nx22403)
             ) ;
    mux21_ni ix51705 (.Y (nx51704), .A0 (nx51640), .A1 (nx51700), .S0 (nx22439)
             ) ;
    mux21_ni ix51641 (.Y (nx51640), .A0 (nx51608), .A1 (nx51636), .S0 (nx22507)
             ) ;
    mux21_ni ix51609 (.Y (nx51608), .A0 (nx51592), .A1 (nx51604), .S0 (nx22641)
             ) ;
    mux21_ni ix51593 (.Y (nx51592), .A0 (inputs_2__12), .A1 (inputs_18__12), .S0 (
             nx23021)) ;
    mux21_ni ix51605 (.Y (nx51604), .A0 (inputs_34__12), .A1 (inputs_50__12), .S0 (
             nx23021)) ;
    mux21_ni ix51637 (.Y (nx51636), .A0 (nx51620), .A1 (nx51632), .S0 (nx22641)
             ) ;
    mux21_ni ix51621 (.Y (nx51620), .A0 (inputs_66__12), .A1 (inputs_82__12), .S0 (
             nx23021)) ;
    mux21_ni ix51633 (.Y (nx51632), .A0 (inputs_98__12), .A1 (inputs_114__12), .S0 (
             nx23023)) ;
    mux21_ni ix51701 (.Y (nx51700), .A0 (nx51668), .A1 (nx51696), .S0 (nx22509)
             ) ;
    mux21_ni ix51669 (.Y (nx51668), .A0 (nx51652), .A1 (nx51664), .S0 (nx22643)
             ) ;
    mux21_ni ix51653 (.Y (nx51652), .A0 (inputs_130__12), .A1 (inputs_146__12), 
             .S0 (nx23023)) ;
    mux21_ni ix51665 (.Y (nx51664), .A0 (inputs_162__12), .A1 (inputs_178__12), 
             .S0 (nx23023)) ;
    mux21_ni ix51697 (.Y (nx51696), .A0 (nx51680), .A1 (nx51692), .S0 (nx22643)
             ) ;
    mux21_ni ix51681 (.Y (nx51680), .A0 (inputs_194__12), .A1 (inputs_210__12), 
             .S0 (nx23023)) ;
    mux21_ni ix51693 (.Y (nx51692), .A0 (inputs_226__12), .A1 (inputs_242__12), 
             .S0 (nx23023)) ;
    mux21_ni ix51829 (.Y (nx51828), .A0 (nx51764), .A1 (nx51824), .S0 (nx22439)
             ) ;
    mux21_ni ix51765 (.Y (nx51764), .A0 (nx51732), .A1 (nx51760), .S0 (nx22509)
             ) ;
    mux21_ni ix51733 (.Y (nx51732), .A0 (nx51716), .A1 (nx51728), .S0 (nx22643)
             ) ;
    mux21_ni ix51717 (.Y (nx51716), .A0 (inputs_258__12), .A1 (inputs_274__12), 
             .S0 (nx23023)) ;
    mux21_ni ix51729 (.Y (nx51728), .A0 (inputs_290__12), .A1 (inputs_306__12), 
             .S0 (nx23023)) ;
    mux21_ni ix51761 (.Y (nx51760), .A0 (nx51744), .A1 (nx51756), .S0 (nx22643)
             ) ;
    mux21_ni ix51745 (.Y (nx51744), .A0 (inputs_322__12), .A1 (inputs_338__12), 
             .S0 (nx23025)) ;
    mux21_ni ix51757 (.Y (nx51756), .A0 (inputs_354__12), .A1 (inputs_370__12), 
             .S0 (nx23025)) ;
    mux21_ni ix51825 (.Y (nx51824), .A0 (nx51792), .A1 (nx51820), .S0 (nx22509)
             ) ;
    mux21_ni ix51793 (.Y (nx51792), .A0 (nx51776), .A1 (nx51788), .S0 (nx22643)
             ) ;
    mux21_ni ix51777 (.Y (nx51776), .A0 (inputs_386__12), .A1 (inputs_402__12), 
             .S0 (nx23025)) ;
    mux21_ni ix51789 (.Y (nx51788), .A0 (inputs_418__12), .A1 (inputs_434__12), 
             .S0 (nx23025)) ;
    mux21_ni ix51821 (.Y (nx51820), .A0 (nx51804), .A1 (nx51816), .S0 (nx22643)
             ) ;
    mux21_ni ix51805 (.Y (nx51804), .A0 (inputs_450__12), .A1 (inputs_466__12), 
             .S0 (nx23025)) ;
    mux21_ni ix51817 (.Y (nx51816), .A0 (inputs_482__12), .A1 (inputs_498__12), 
             .S0 (nx23025)) ;
    mux21_ni ix54045 (.Y (nx54044), .A0 (nx53196), .A1 (nx54040), .S0 (nx22439)
             ) ;
    mux21_ni ix53197 (.Y (nx53196), .A0 (nx52772), .A1 (nx53192), .S0 (nx22509)
             ) ;
    mux21_ni ix52773 (.Y (nx52772), .A0 (nx52560), .A1 (nx52768), .S0 (nx22643)
             ) ;
    mux21_ni ix52561 (.Y (nx52560), .A0 (nx52554), .A1 (nx52476), .S0 (nx23173)
             ) ;
    oai21 ix52555 (.Y (nx52554), .A0 (nx22345), .A1 (nx19253), .B0 (nx19263)) ;
    mux21 ix19254 (.Y (nx19253), .A0 (nx52518), .A1 (nx52546), .S0 (nx23025)) ;
    mux21_ni ix52519 (.Y (nx52518), .A0 (nx52502), .A1 (nx52514), .S0 (nx23767)
             ) ;
    mux21_ni ix52503 (.Y (nx52502), .A0 (inputs_4__12), .A1 (inputs_5__12), .S0 (
             nx24629)) ;
    mux21_ni ix52515 (.Y (nx52514), .A0 (inputs_6__12), .A1 (inputs_7__12), .S0 (
             nx24629)) ;
    mux21_ni ix52547 (.Y (nx52546), .A0 (nx52530), .A1 (nx52542), .S0 (nx23767)
             ) ;
    mux21_ni ix52531 (.Y (nx52530), .A0 (inputs_20__12), .A1 (inputs_21__12), .S0 (
             nx24629)) ;
    mux21_ni ix52543 (.Y (nx52542), .A0 (inputs_22__12), .A1 (inputs_23__12), .S0 (
             nx24629)) ;
    nand04 ix19264 (.Y (nx19263), .A0 (nx22345), .A1 (nx23769), .A2 (nx24629), .A3 (
           nx52490)) ;
    mux21_ni ix52491 (.Y (nx52490), .A0 (inputs_3__12), .A1 (inputs_19__12), .S0 (
             nx23027)) ;
    mux21_ni ix52477 (.Y (nx52476), .A0 (nx52412), .A1 (nx52472), .S0 (nx23027)
             ) ;
    mux21_ni ix52413 (.Y (nx52412), .A0 (nx52380), .A1 (nx52408), .S0 (nx23305)
             ) ;
    mux21_ni ix52381 (.Y (nx52380), .A0 (nx52364), .A1 (nx52376), .S0 (nx23769)
             ) ;
    mux21_ni ix52365 (.Y (nx52364), .A0 (inputs_8__12), .A1 (inputs_9__12), .S0 (
             nx24631)) ;
    mux21_ni ix52377 (.Y (nx52376), .A0 (inputs_10__12), .A1 (inputs_11__12), .S0 (
             nx24631)) ;
    mux21_ni ix52409 (.Y (nx52408), .A0 (nx52392), .A1 (nx52404), .S0 (nx23769)
             ) ;
    mux21_ni ix52393 (.Y (nx52392), .A0 (inputs_12__12), .A1 (inputs_13__12), .S0 (
             nx24631)) ;
    mux21_ni ix52405 (.Y (nx52404), .A0 (inputs_14__12), .A1 (inputs_15__12), .S0 (
             nx24631)) ;
    mux21_ni ix52473 (.Y (nx52472), .A0 (nx52440), .A1 (nx52468), .S0 (nx23305)
             ) ;
    mux21_ni ix52441 (.Y (nx52440), .A0 (nx52424), .A1 (nx52436), .S0 (nx23769)
             ) ;
    mux21_ni ix52425 (.Y (nx52424), .A0 (inputs_24__12), .A1 (inputs_25__12), .S0 (
             nx24631)) ;
    mux21_ni ix52437 (.Y (nx52436), .A0 (inputs_26__12), .A1 (inputs_27__12), .S0 (
             nx24631)) ;
    mux21_ni ix52469 (.Y (nx52468), .A0 (nx52452), .A1 (nx52464), .S0 (nx23769)
             ) ;
    mux21_ni ix52453 (.Y (nx52452), .A0 (inputs_28__12), .A1 (inputs_29__12), .S0 (
             nx24631)) ;
    mux21_ni ix52465 (.Y (nx52464), .A0 (inputs_30__12), .A1 (inputs_31__12), .S0 (
             nx24633)) ;
    mux21_ni ix52769 (.Y (nx52768), .A0 (nx52762), .A1 (nx52684), .S0 (nx23173)
             ) ;
    oai21 ix52763 (.Y (nx52762), .A0 (nx22345), .A1 (nx19295), .B0 (nx19305)) ;
    mux21 ix19296 (.Y (nx19295), .A0 (nx52726), .A1 (nx52754), .S0 (nx23027)) ;
    mux21_ni ix52727 (.Y (nx52726), .A0 (nx52710), .A1 (nx52722), .S0 (nx23769)
             ) ;
    mux21_ni ix52711 (.Y (nx52710), .A0 (inputs_36__12), .A1 (inputs_37__12), .S0 (
             nx24633)) ;
    mux21_ni ix52723 (.Y (nx52722), .A0 (inputs_38__12), .A1 (inputs_39__12), .S0 (
             nx24633)) ;
    mux21_ni ix52755 (.Y (nx52754), .A0 (nx52738), .A1 (nx52750), .S0 (nx23769)
             ) ;
    mux21_ni ix52739 (.Y (nx52738), .A0 (inputs_52__12), .A1 (inputs_53__12), .S0 (
             nx24633)) ;
    mux21_ni ix52751 (.Y (nx52750), .A0 (inputs_54__12), .A1 (inputs_55__12), .S0 (
             nx24633)) ;
    nand04 ix19306 (.Y (nx19305), .A0 (nx22345), .A1 (nx23771), .A2 (nx24633), .A3 (
           nx52698)) ;
    mux21_ni ix52699 (.Y (nx52698), .A0 (inputs_35__12), .A1 (inputs_51__12), .S0 (
             nx23027)) ;
    mux21_ni ix52685 (.Y (nx52684), .A0 (nx52620), .A1 (nx52680), .S0 (nx23027)
             ) ;
    mux21_ni ix52621 (.Y (nx52620), .A0 (nx52588), .A1 (nx52616), .S0 (nx23305)
             ) ;
    mux21_ni ix52589 (.Y (nx52588), .A0 (nx52572), .A1 (nx52584), .S0 (nx23771)
             ) ;
    mux21_ni ix52573 (.Y (nx52572), .A0 (inputs_40__12), .A1 (inputs_41__12), .S0 (
             nx24633)) ;
    mux21_ni ix52585 (.Y (nx52584), .A0 (inputs_42__12), .A1 (inputs_43__12), .S0 (
             nx24635)) ;
    mux21_ni ix52617 (.Y (nx52616), .A0 (nx52600), .A1 (nx52612), .S0 (nx23771)
             ) ;
    mux21_ni ix52601 (.Y (nx52600), .A0 (inputs_44__12), .A1 (inputs_45__12), .S0 (
             nx24635)) ;
    mux21_ni ix52613 (.Y (nx52612), .A0 (inputs_46__12), .A1 (inputs_47__12), .S0 (
             nx24635)) ;
    mux21_ni ix52681 (.Y (nx52680), .A0 (nx52648), .A1 (nx52676), .S0 (nx23305)
             ) ;
    mux21_ni ix52649 (.Y (nx52648), .A0 (nx52632), .A1 (nx52644), .S0 (nx23771)
             ) ;
    mux21_ni ix52633 (.Y (nx52632), .A0 (inputs_56__12), .A1 (inputs_57__12), .S0 (
             nx24635)) ;
    mux21_ni ix52645 (.Y (nx52644), .A0 (inputs_58__12), .A1 (inputs_59__12), .S0 (
             nx24635)) ;
    mux21_ni ix52677 (.Y (nx52676), .A0 (nx52660), .A1 (nx52672), .S0 (nx23771)
             ) ;
    mux21_ni ix52661 (.Y (nx52660), .A0 (inputs_60__12), .A1 (inputs_61__12), .S0 (
             nx24635)) ;
    mux21_ni ix52673 (.Y (nx52672), .A0 (inputs_62__12), .A1 (inputs_63__12), .S0 (
             nx24635)) ;
    mux21_ni ix53193 (.Y (nx53192), .A0 (nx52980), .A1 (nx53188), .S0 (nx22645)
             ) ;
    mux21_ni ix52981 (.Y (nx52980), .A0 (nx52974), .A1 (nx52896), .S0 (nx23173)
             ) ;
    oai21 ix52975 (.Y (nx52974), .A0 (nx22345), .A1 (nx19337), .B0 (nx19347)) ;
    mux21 ix19338 (.Y (nx19337), .A0 (nx52938), .A1 (nx52966), .S0 (nx23027)) ;
    mux21_ni ix52939 (.Y (nx52938), .A0 (nx52922), .A1 (nx52934), .S0 (nx23771)
             ) ;
    mux21_ni ix52923 (.Y (nx52922), .A0 (inputs_68__12), .A1 (inputs_69__12), .S0 (
             nx24637)) ;
    mux21_ni ix52935 (.Y (nx52934), .A0 (inputs_70__12), .A1 (inputs_71__12), .S0 (
             nx24637)) ;
    mux21_ni ix52967 (.Y (nx52966), .A0 (nx52950), .A1 (nx52962), .S0 (nx23771)
             ) ;
    mux21_ni ix52951 (.Y (nx52950), .A0 (inputs_84__12), .A1 (inputs_85__12), .S0 (
             nx24637)) ;
    mux21_ni ix52963 (.Y (nx52962), .A0 (inputs_86__12), .A1 (inputs_87__12), .S0 (
             nx24637)) ;
    nand04 ix19348 (.Y (nx19347), .A0 (nx22345), .A1 (nx23773), .A2 (nx24637), .A3 (
           nx52910)) ;
    mux21_ni ix52911 (.Y (nx52910), .A0 (inputs_67__12), .A1 (inputs_83__12), .S0 (
             nx23027)) ;
    mux21_ni ix52897 (.Y (nx52896), .A0 (nx52832), .A1 (nx52892), .S0 (nx23029)
             ) ;
    mux21_ni ix52833 (.Y (nx52832), .A0 (nx52800), .A1 (nx52828), .S0 (nx23305)
             ) ;
    mux21_ni ix52801 (.Y (nx52800), .A0 (nx52784), .A1 (nx52796), .S0 (nx23773)
             ) ;
    mux21_ni ix52785 (.Y (nx52784), .A0 (inputs_72__12), .A1 (inputs_73__12), .S0 (
             nx24637)) ;
    mux21_ni ix52797 (.Y (nx52796), .A0 (inputs_74__12), .A1 (inputs_75__12), .S0 (
             nx24637)) ;
    mux21_ni ix52829 (.Y (nx52828), .A0 (nx52812), .A1 (nx52824), .S0 (nx23773)
             ) ;
    mux21_ni ix52813 (.Y (nx52812), .A0 (inputs_76__12), .A1 (inputs_77__12), .S0 (
             nx24639)) ;
    mux21_ni ix52825 (.Y (nx52824), .A0 (inputs_78__12), .A1 (inputs_79__12), .S0 (
             nx24639)) ;
    mux21_ni ix52893 (.Y (nx52892), .A0 (nx52860), .A1 (nx52888), .S0 (nx23305)
             ) ;
    mux21_ni ix52861 (.Y (nx52860), .A0 (nx52844), .A1 (nx52856), .S0 (nx23773)
             ) ;
    mux21_ni ix52845 (.Y (nx52844), .A0 (inputs_88__12), .A1 (inputs_89__12), .S0 (
             nx24639)) ;
    mux21_ni ix52857 (.Y (nx52856), .A0 (inputs_90__12), .A1 (inputs_91__12), .S0 (
             nx24639)) ;
    mux21_ni ix52889 (.Y (nx52888), .A0 (nx52872), .A1 (nx52884), .S0 (nx23773)
             ) ;
    mux21_ni ix52873 (.Y (nx52872), .A0 (inputs_92__12), .A1 (inputs_93__12), .S0 (
             nx24639)) ;
    mux21_ni ix52885 (.Y (nx52884), .A0 (inputs_94__12), .A1 (inputs_95__12), .S0 (
             nx24639)) ;
    mux21_ni ix53189 (.Y (nx53188), .A0 (nx53182), .A1 (nx53104), .S0 (nx23175)
             ) ;
    oai21 ix53183 (.Y (nx53182), .A0 (nx22345), .A1 (nx19377), .B0 (nx19389)) ;
    mux21 ix19378 (.Y (nx19377), .A0 (nx53146), .A1 (nx53174), .S0 (nx23029)) ;
    mux21_ni ix53147 (.Y (nx53146), .A0 (nx53130), .A1 (nx53142), .S0 (nx23773)
             ) ;
    mux21_ni ix53131 (.Y (nx53130), .A0 (inputs_100__12), .A1 (inputs_101__12), 
             .S0 (nx24639)) ;
    mux21_ni ix53143 (.Y (nx53142), .A0 (inputs_102__12), .A1 (inputs_103__12), 
             .S0 (nx24641)) ;
    mux21_ni ix53175 (.Y (nx53174), .A0 (nx53158), .A1 (nx53170), .S0 (nx23773)
             ) ;
    mux21_ni ix53159 (.Y (nx53158), .A0 (inputs_116__12), .A1 (inputs_117__12), 
             .S0 (nx24641)) ;
    mux21_ni ix53171 (.Y (nx53170), .A0 (inputs_118__12), .A1 (inputs_119__12), 
             .S0 (nx24641)) ;
    nand04 ix19390 (.Y (nx19389), .A0 (nx22347), .A1 (nx23775), .A2 (nx24641), .A3 (
           nx53118)) ;
    mux21_ni ix53119 (.Y (nx53118), .A0 (inputs_99__12), .A1 (inputs_115__12), .S0 (
             nx23029)) ;
    mux21_ni ix53105 (.Y (nx53104), .A0 (nx53040), .A1 (nx53100), .S0 (nx23029)
             ) ;
    mux21_ni ix53041 (.Y (nx53040), .A0 (nx53008), .A1 (nx53036), .S0 (nx23307)
             ) ;
    mux21_ni ix53009 (.Y (nx53008), .A0 (nx52992), .A1 (nx53004), .S0 (nx23775)
             ) ;
    mux21_ni ix52993 (.Y (nx52992), .A0 (inputs_104__12), .A1 (inputs_105__12), 
             .S0 (nx24641)) ;
    mux21_ni ix53005 (.Y (nx53004), .A0 (inputs_106__12), .A1 (inputs_107__12), 
             .S0 (nx24641)) ;
    mux21_ni ix53037 (.Y (nx53036), .A0 (nx53020), .A1 (nx53032), .S0 (nx23775)
             ) ;
    mux21_ni ix53021 (.Y (nx53020), .A0 (inputs_108__12), .A1 (inputs_109__12), 
             .S0 (nx24641)) ;
    mux21_ni ix53033 (.Y (nx53032), .A0 (inputs_110__12), .A1 (inputs_111__12), 
             .S0 (nx24643)) ;
    mux21_ni ix53101 (.Y (nx53100), .A0 (nx53068), .A1 (nx53096), .S0 (nx23307)
             ) ;
    mux21_ni ix53069 (.Y (nx53068), .A0 (nx53052), .A1 (nx53064), .S0 (nx23775)
             ) ;
    mux21_ni ix53053 (.Y (nx53052), .A0 (inputs_120__12), .A1 (inputs_121__12), 
             .S0 (nx24643)) ;
    mux21_ni ix53065 (.Y (nx53064), .A0 (inputs_122__12), .A1 (inputs_123__12), 
             .S0 (nx24643)) ;
    mux21_ni ix53097 (.Y (nx53096), .A0 (nx53080), .A1 (nx53092), .S0 (nx23775)
             ) ;
    mux21_ni ix53081 (.Y (nx53080), .A0 (inputs_124__12), .A1 (inputs_125__12), 
             .S0 (nx24643)) ;
    mux21_ni ix53093 (.Y (nx53092), .A0 (inputs_126__12), .A1 (inputs_127__12), 
             .S0 (nx24643)) ;
    mux21_ni ix54041 (.Y (nx54040), .A0 (nx53616), .A1 (nx54036), .S0 (nx22509)
             ) ;
    mux21_ni ix53617 (.Y (nx53616), .A0 (nx53404), .A1 (nx53612), .S0 (nx22645)
             ) ;
    mux21_ni ix53405 (.Y (nx53404), .A0 (nx53398), .A1 (nx53320), .S0 (nx23175)
             ) ;
    oai21 ix53399 (.Y (nx53398), .A0 (nx22347), .A1 (nx19425), .B0 (nx19437)) ;
    mux21 ix19426 (.Y (nx19425), .A0 (nx53362), .A1 (nx53390), .S0 (nx23029)) ;
    mux21_ni ix53363 (.Y (nx53362), .A0 (nx53346), .A1 (nx53358), .S0 (nx23775)
             ) ;
    mux21_ni ix53347 (.Y (nx53346), .A0 (inputs_132__12), .A1 (inputs_133__12), 
             .S0 (nx24643)) ;
    mux21_ni ix53359 (.Y (nx53358), .A0 (inputs_134__12), .A1 (inputs_135__12), 
             .S0 (nx24643)) ;
    mux21_ni ix53391 (.Y (nx53390), .A0 (nx53374), .A1 (nx53386), .S0 (nx23775)
             ) ;
    mux21_ni ix53375 (.Y (nx53374), .A0 (inputs_148__12), .A1 (inputs_149__12), 
             .S0 (nx24645)) ;
    mux21_ni ix53387 (.Y (nx53386), .A0 (inputs_150__12), .A1 (inputs_151__12), 
             .S0 (nx24645)) ;
    nand04 ix19438 (.Y (nx19437), .A0 (nx22347), .A1 (nx23777), .A2 (nx24645), .A3 (
           nx53334)) ;
    mux21_ni ix53335 (.Y (nx53334), .A0 (inputs_131__12), .A1 (inputs_147__12), 
             .S0 (nx23029)) ;
    mux21_ni ix53321 (.Y (nx53320), .A0 (nx53256), .A1 (nx53316), .S0 (nx23029)
             ) ;
    mux21_ni ix53257 (.Y (nx53256), .A0 (nx53224), .A1 (nx53252), .S0 (nx23307)
             ) ;
    mux21_ni ix53225 (.Y (nx53224), .A0 (nx53208), .A1 (nx53220), .S0 (nx23777)
             ) ;
    mux21_ni ix53209 (.Y (nx53208), .A0 (inputs_136__12), .A1 (inputs_137__12), 
             .S0 (nx24645)) ;
    mux21_ni ix53221 (.Y (nx53220), .A0 (inputs_138__12), .A1 (inputs_139__12), 
             .S0 (nx24645)) ;
    mux21_ni ix53253 (.Y (nx53252), .A0 (nx53236), .A1 (nx53248), .S0 (nx23777)
             ) ;
    mux21_ni ix53237 (.Y (nx53236), .A0 (inputs_140__12), .A1 (inputs_141__12), 
             .S0 (nx24645)) ;
    mux21_ni ix53249 (.Y (nx53248), .A0 (inputs_142__12), .A1 (inputs_143__12), 
             .S0 (nx24645)) ;
    mux21_ni ix53317 (.Y (nx53316), .A0 (nx53284), .A1 (nx53312), .S0 (nx23307)
             ) ;
    mux21_ni ix53285 (.Y (nx53284), .A0 (nx53268), .A1 (nx53280), .S0 (nx23777)
             ) ;
    mux21_ni ix53269 (.Y (nx53268), .A0 (inputs_152__12), .A1 (inputs_153__12), 
             .S0 (nx24647)) ;
    mux21_ni ix53281 (.Y (nx53280), .A0 (inputs_154__12), .A1 (inputs_155__12), 
             .S0 (nx24647)) ;
    mux21_ni ix53313 (.Y (nx53312), .A0 (nx53296), .A1 (nx53308), .S0 (nx23777)
             ) ;
    mux21_ni ix53297 (.Y (nx53296), .A0 (inputs_156__12), .A1 (inputs_157__12), 
             .S0 (nx24647)) ;
    mux21_ni ix53309 (.Y (nx53308), .A0 (inputs_158__12), .A1 (inputs_159__12), 
             .S0 (nx24647)) ;
    mux21_ni ix53613 (.Y (nx53612), .A0 (nx53606), .A1 (nx53528), .S0 (nx23175)
             ) ;
    oai21 ix53607 (.Y (nx53606), .A0 (nx22347), .A1 (nx19467), .B0 (nx19479)) ;
    mux21 ix19468 (.Y (nx19467), .A0 (nx53570), .A1 (nx53598), .S0 (nx23031)) ;
    mux21_ni ix53571 (.Y (nx53570), .A0 (nx53554), .A1 (nx53566), .S0 (nx23777)
             ) ;
    mux21_ni ix53555 (.Y (nx53554), .A0 (inputs_164__12), .A1 (inputs_165__12), 
             .S0 (nx24647)) ;
    mux21_ni ix53567 (.Y (nx53566), .A0 (inputs_166__12), .A1 (inputs_167__12), 
             .S0 (nx24647)) ;
    mux21_ni ix53599 (.Y (nx53598), .A0 (nx53582), .A1 (nx53594), .S0 (nx23777)
             ) ;
    mux21_ni ix53583 (.Y (nx53582), .A0 (inputs_180__12), .A1 (inputs_181__12), 
             .S0 (nx24647)) ;
    mux21_ni ix53595 (.Y (nx53594), .A0 (inputs_182__12), .A1 (inputs_183__12), 
             .S0 (nx24649)) ;
    nand04 ix19480 (.Y (nx19479), .A0 (nx22347), .A1 (nx23779), .A2 (nx24649), .A3 (
           nx53542)) ;
    mux21_ni ix53543 (.Y (nx53542), .A0 (inputs_163__12), .A1 (inputs_179__12), 
             .S0 (nx23031)) ;
    mux21_ni ix53529 (.Y (nx53528), .A0 (nx53464), .A1 (nx53524), .S0 (nx23031)
             ) ;
    mux21_ni ix53465 (.Y (nx53464), .A0 (nx53432), .A1 (nx53460), .S0 (nx23307)
             ) ;
    mux21_ni ix53433 (.Y (nx53432), .A0 (nx53416), .A1 (nx53428), .S0 (nx23779)
             ) ;
    mux21_ni ix53417 (.Y (nx53416), .A0 (inputs_168__12), .A1 (inputs_169__12), 
             .S0 (nx24649)) ;
    mux21_ni ix53429 (.Y (nx53428), .A0 (inputs_170__12), .A1 (inputs_171__12), 
             .S0 (nx24649)) ;
    mux21_ni ix53461 (.Y (nx53460), .A0 (nx53444), .A1 (nx53456), .S0 (nx23779)
             ) ;
    mux21_ni ix53445 (.Y (nx53444), .A0 (inputs_172__12), .A1 (inputs_173__12), 
             .S0 (nx24649)) ;
    mux21_ni ix53457 (.Y (nx53456), .A0 (inputs_174__12), .A1 (inputs_175__12), 
             .S0 (nx24649)) ;
    mux21_ni ix53525 (.Y (nx53524), .A0 (nx53492), .A1 (nx53520), .S0 (nx23307)
             ) ;
    mux21_ni ix53493 (.Y (nx53492), .A0 (nx53476), .A1 (nx53488), .S0 (nx23779)
             ) ;
    mux21_ni ix53477 (.Y (nx53476), .A0 (inputs_184__12), .A1 (inputs_185__12), 
             .S0 (nx24649)) ;
    mux21_ni ix53489 (.Y (nx53488), .A0 (inputs_186__12), .A1 (inputs_187__12), 
             .S0 (nx24651)) ;
    mux21_ni ix53521 (.Y (nx53520), .A0 (nx53504), .A1 (nx53516), .S0 (nx23779)
             ) ;
    mux21_ni ix53505 (.Y (nx53504), .A0 (inputs_188__12), .A1 (inputs_189__12), 
             .S0 (nx24651)) ;
    mux21_ni ix53517 (.Y (nx53516), .A0 (inputs_190__12), .A1 (inputs_191__12), 
             .S0 (nx24651)) ;
    mux21_ni ix54037 (.Y (nx54036), .A0 (nx53824), .A1 (nx54032), .S0 (nx22645)
             ) ;
    mux21_ni ix53825 (.Y (nx53824), .A0 (nx53818), .A1 (nx53740), .S0 (nx23175)
             ) ;
    oai21 ix53819 (.Y (nx53818), .A0 (nx22347), .A1 (nx19513), .B0 (nx19525)) ;
    mux21 ix19514 (.Y (nx19513), .A0 (nx53782), .A1 (nx53810), .S0 (nx23031)) ;
    mux21_ni ix53783 (.Y (nx53782), .A0 (nx53766), .A1 (nx53778), .S0 (nx23779)
             ) ;
    mux21_ni ix53767 (.Y (nx53766), .A0 (inputs_196__12), .A1 (inputs_197__12), 
             .S0 (nx24651)) ;
    mux21_ni ix53779 (.Y (nx53778), .A0 (inputs_198__12), .A1 (inputs_199__12), 
             .S0 (nx24651)) ;
    mux21_ni ix53811 (.Y (nx53810), .A0 (nx53794), .A1 (nx53806), .S0 (nx23779)
             ) ;
    mux21_ni ix53795 (.Y (nx53794), .A0 (inputs_212__12), .A1 (inputs_213__12), 
             .S0 (nx24651)) ;
    mux21_ni ix53807 (.Y (nx53806), .A0 (inputs_214__12), .A1 (inputs_215__12), 
             .S0 (nx24651)) ;
    nand04 ix19526 (.Y (nx19525), .A0 (nx22347), .A1 (nx23781), .A2 (nx24653), .A3 (
           nx53754)) ;
    mux21_ni ix53755 (.Y (nx53754), .A0 (inputs_195__12), .A1 (inputs_211__12), 
             .S0 (nx23031)) ;
    mux21_ni ix53741 (.Y (nx53740), .A0 (nx53676), .A1 (nx53736), .S0 (nx23031)
             ) ;
    mux21_ni ix53677 (.Y (nx53676), .A0 (nx53644), .A1 (nx53672), .S0 (nx23307)
             ) ;
    mux21_ni ix53645 (.Y (nx53644), .A0 (nx53628), .A1 (nx53640), .S0 (nx23781)
             ) ;
    mux21_ni ix53629 (.Y (nx53628), .A0 (inputs_200__12), .A1 (inputs_201__12), 
             .S0 (nx24653)) ;
    mux21_ni ix53641 (.Y (nx53640), .A0 (inputs_202__12), .A1 (inputs_203__12), 
             .S0 (nx24653)) ;
    mux21_ni ix53673 (.Y (nx53672), .A0 (nx53656), .A1 (nx53668), .S0 (nx23781)
             ) ;
    mux21_ni ix53657 (.Y (nx53656), .A0 (inputs_204__12), .A1 (inputs_205__12), 
             .S0 (nx24653)) ;
    mux21_ni ix53669 (.Y (nx53668), .A0 (inputs_206__12), .A1 (inputs_207__12), 
             .S0 (nx24653)) ;
    mux21_ni ix53737 (.Y (nx53736), .A0 (nx53704), .A1 (nx53732), .S0 (nx23309)
             ) ;
    mux21_ni ix53705 (.Y (nx53704), .A0 (nx53688), .A1 (nx53700), .S0 (nx23781)
             ) ;
    mux21_ni ix53689 (.Y (nx53688), .A0 (inputs_216__12), .A1 (inputs_217__12), 
             .S0 (nx24653)) ;
    mux21_ni ix53701 (.Y (nx53700), .A0 (inputs_218__12), .A1 (inputs_219__12), 
             .S0 (nx24653)) ;
    mux21_ni ix53733 (.Y (nx53732), .A0 (nx53716), .A1 (nx53728), .S0 (nx23781)
             ) ;
    mux21_ni ix53717 (.Y (nx53716), .A0 (inputs_220__12), .A1 (inputs_221__12), 
             .S0 (nx24655)) ;
    mux21_ni ix53729 (.Y (nx53728), .A0 (inputs_222__12), .A1 (inputs_223__12), 
             .S0 (nx24655)) ;
    mux21_ni ix54033 (.Y (nx54032), .A0 (nx54026), .A1 (nx53948), .S0 (nx23175)
             ) ;
    oai21 ix54027 (.Y (nx54026), .A0 (nx22349), .A1 (nx19555), .B0 (nx19569)) ;
    mux21 ix19556 (.Y (nx19555), .A0 (nx53990), .A1 (nx54018), .S0 (nx23031)) ;
    mux21_ni ix53991 (.Y (nx53990), .A0 (nx53974), .A1 (nx53986), .S0 (nx23781)
             ) ;
    mux21_ni ix53975 (.Y (nx53974), .A0 (inputs_228__12), .A1 (inputs_229__12), 
             .S0 (nx24655)) ;
    mux21_ni ix53987 (.Y (nx53986), .A0 (inputs_230__12), .A1 (inputs_231__12), 
             .S0 (nx24655)) ;
    mux21_ni ix54019 (.Y (nx54018), .A0 (nx54002), .A1 (nx54014), .S0 (nx23781)
             ) ;
    mux21_ni ix54003 (.Y (nx54002), .A0 (inputs_244__12), .A1 (inputs_245__12), 
             .S0 (nx24655)) ;
    mux21_ni ix54015 (.Y (nx54014), .A0 (inputs_246__12), .A1 (inputs_247__12), 
             .S0 (nx24655)) ;
    nand04 ix19570 (.Y (nx19569), .A0 (nx22349), .A1 (nx23783), .A2 (nx24655), .A3 (
           nx53962)) ;
    mux21_ni ix53963 (.Y (nx53962), .A0 (inputs_227__12), .A1 (inputs_243__12), 
             .S0 (nx23033)) ;
    mux21_ni ix53949 (.Y (nx53948), .A0 (nx53884), .A1 (nx53944), .S0 (nx23033)
             ) ;
    mux21_ni ix53885 (.Y (nx53884), .A0 (nx53852), .A1 (nx53880), .S0 (nx23309)
             ) ;
    mux21_ni ix53853 (.Y (nx53852), .A0 (nx53836), .A1 (nx53848), .S0 (nx23783)
             ) ;
    mux21_ni ix53837 (.Y (nx53836), .A0 (inputs_232__12), .A1 (inputs_233__12), 
             .S0 (nx24657)) ;
    mux21_ni ix53849 (.Y (nx53848), .A0 (inputs_234__12), .A1 (inputs_235__12), 
             .S0 (nx24657)) ;
    mux21_ni ix53881 (.Y (nx53880), .A0 (nx53864), .A1 (nx53876), .S0 (nx23783)
             ) ;
    mux21_ni ix53865 (.Y (nx53864), .A0 (inputs_236__12), .A1 (inputs_237__12), 
             .S0 (nx24657)) ;
    mux21_ni ix53877 (.Y (nx53876), .A0 (inputs_238__12), .A1 (inputs_239__12), 
             .S0 (nx24657)) ;
    mux21_ni ix53945 (.Y (nx53944), .A0 (nx53912), .A1 (nx53940), .S0 (nx23309)
             ) ;
    mux21_ni ix53913 (.Y (nx53912), .A0 (nx53896), .A1 (nx53908), .S0 (nx23783)
             ) ;
    mux21_ni ix53897 (.Y (nx53896), .A0 (inputs_248__12), .A1 (inputs_249__12), 
             .S0 (nx24657)) ;
    mux21_ni ix53909 (.Y (nx53908), .A0 (inputs_250__12), .A1 (inputs_251__12), 
             .S0 (nx24657)) ;
    mux21_ni ix53941 (.Y (nx53940), .A0 (nx53924), .A1 (nx53936), .S0 (nx23783)
             ) ;
    mux21_ni ix53925 (.Y (nx53924), .A0 (inputs_252__12), .A1 (inputs_253__12), 
             .S0 (nx24657)) ;
    mux21_ni ix53937 (.Y (nx53936), .A0 (inputs_254__12), .A1 (inputs_255__12), 
             .S0 (nx24659)) ;
    oai21 ix58211 (.Y (\output [13]), .A0 (nx22223), .A1 (nx19597), .B0 (nx19953
          )) ;
    mux21 ix19598 (.Y (nx19597), .A0 (nx54892), .A1 (nx55736), .S0 (nx22439)) ;
    mux21_ni ix54893 (.Y (nx54892), .A0 (nx54468), .A1 (nx54888), .S0 (nx22509)
             ) ;
    mux21_ni ix54469 (.Y (nx54468), .A0 (nx54256), .A1 (nx54464), .S0 (nx22645)
             ) ;
    mux21_ni ix54257 (.Y (nx54256), .A0 (nx54250), .A1 (nx54172), .S0 (nx23175)
             ) ;
    oai21 ix54251 (.Y (nx54250), .A0 (nx22349), .A1 (nx19605), .B0 (nx19617)) ;
    mux21 ix19606 (.Y (nx19605), .A0 (nx54214), .A1 (nx54242), .S0 (nx23033)) ;
    mux21_ni ix54215 (.Y (nx54214), .A0 (nx54198), .A1 (nx54210), .S0 (nx23783)
             ) ;
    mux21_ni ix54199 (.Y (nx54198), .A0 (inputs_260__13), .A1 (inputs_261__13), 
             .S0 (nx24659)) ;
    mux21_ni ix54211 (.Y (nx54210), .A0 (inputs_262__13), .A1 (inputs_263__13), 
             .S0 (nx24659)) ;
    mux21_ni ix54243 (.Y (nx54242), .A0 (nx54226), .A1 (nx54238), .S0 (nx23783)
             ) ;
    mux21_ni ix54227 (.Y (nx54226), .A0 (inputs_276__13), .A1 (inputs_277__13), 
             .S0 (nx24659)) ;
    mux21_ni ix54239 (.Y (nx54238), .A0 (inputs_278__13), .A1 (inputs_279__13), 
             .S0 (nx24659)) ;
    nand04 ix19618 (.Y (nx19617), .A0 (nx22349), .A1 (nx23785), .A2 (nx24659), .A3 (
           nx54186)) ;
    mux21_ni ix54187 (.Y (nx54186), .A0 (inputs_259__13), .A1 (inputs_275__13), 
             .S0 (nx23033)) ;
    mux21_ni ix54173 (.Y (nx54172), .A0 (nx54108), .A1 (nx54168), .S0 (nx23033)
             ) ;
    mux21_ni ix54109 (.Y (nx54108), .A0 (nx54076), .A1 (nx54104), .S0 (nx23309)
             ) ;
    mux21_ni ix54077 (.Y (nx54076), .A0 (nx54060), .A1 (nx54072), .S0 (nx23785)
             ) ;
    mux21_ni ix54061 (.Y (nx54060), .A0 (inputs_264__13), .A1 (inputs_265__13), 
             .S0 (nx24659)) ;
    mux21_ni ix54073 (.Y (nx54072), .A0 (inputs_266__13), .A1 (inputs_267__13), 
             .S0 (nx24661)) ;
    mux21_ni ix54105 (.Y (nx54104), .A0 (nx54088), .A1 (nx54100), .S0 (nx23785)
             ) ;
    mux21_ni ix54089 (.Y (nx54088), .A0 (inputs_268__13), .A1 (inputs_269__13), 
             .S0 (nx24661)) ;
    mux21_ni ix54101 (.Y (nx54100), .A0 (inputs_270__13), .A1 (inputs_271__13), 
             .S0 (nx24661)) ;
    mux21_ni ix54169 (.Y (nx54168), .A0 (nx54136), .A1 (nx54164), .S0 (nx23309)
             ) ;
    mux21_ni ix54137 (.Y (nx54136), .A0 (nx54120), .A1 (nx54132), .S0 (nx23785)
             ) ;
    mux21_ni ix54121 (.Y (nx54120), .A0 (inputs_280__13), .A1 (inputs_281__13), 
             .S0 (nx24661)) ;
    mux21_ni ix54133 (.Y (nx54132), .A0 (inputs_282__13), .A1 (inputs_283__13), 
             .S0 (nx24661)) ;
    mux21_ni ix54165 (.Y (nx54164), .A0 (nx54148), .A1 (nx54160), .S0 (nx23785)
             ) ;
    mux21_ni ix54149 (.Y (nx54148), .A0 (inputs_284__13), .A1 (inputs_285__13), 
             .S0 (nx24661)) ;
    mux21_ni ix54161 (.Y (nx54160), .A0 (inputs_286__13), .A1 (inputs_287__13), 
             .S0 (nx24661)) ;
    mux21_ni ix54465 (.Y (nx54464), .A0 (nx54458), .A1 (nx54380), .S0 (nx23175)
             ) ;
    oai21 ix54459 (.Y (nx54458), .A0 (nx22349), .A1 (nx19651), .B0 (nx19663)) ;
    mux21 ix19652 (.Y (nx19651), .A0 (nx54422), .A1 (nx54450), .S0 (nx23033)) ;
    mux21_ni ix54423 (.Y (nx54422), .A0 (nx54406), .A1 (nx54418), .S0 (nx23785)
             ) ;
    mux21_ni ix54407 (.Y (nx54406), .A0 (inputs_292__13), .A1 (inputs_293__13), 
             .S0 (nx24663)) ;
    mux21_ni ix54419 (.Y (nx54418), .A0 (inputs_294__13), .A1 (inputs_295__13), 
             .S0 (nx24663)) ;
    mux21_ni ix54451 (.Y (nx54450), .A0 (nx54434), .A1 (nx54446), .S0 (nx23785)
             ) ;
    mux21_ni ix54435 (.Y (nx54434), .A0 (inputs_308__13), .A1 (inputs_309__13), 
             .S0 (nx24663)) ;
    mux21_ni ix54447 (.Y (nx54446), .A0 (inputs_310__13), .A1 (inputs_311__13), 
             .S0 (nx24663)) ;
    nand04 ix19664 (.Y (nx19663), .A0 (nx22349), .A1 (nx23787), .A2 (nx24663), .A3 (
           nx54394)) ;
    mux21_ni ix54395 (.Y (nx54394), .A0 (inputs_291__13), .A1 (inputs_307__13), 
             .S0 (nx23033)) ;
    mux21_ni ix54381 (.Y (nx54380), .A0 (nx54316), .A1 (nx54376), .S0 (nx23035)
             ) ;
    mux21_ni ix54317 (.Y (nx54316), .A0 (nx54284), .A1 (nx54312), .S0 (nx23309)
             ) ;
    mux21_ni ix54285 (.Y (nx54284), .A0 (nx54268), .A1 (nx54280), .S0 (nx23787)
             ) ;
    mux21_ni ix54269 (.Y (nx54268), .A0 (inputs_296__13), .A1 (inputs_297__13), 
             .S0 (nx24663)) ;
    mux21_ni ix54281 (.Y (nx54280), .A0 (inputs_298__13), .A1 (inputs_299__13), 
             .S0 (nx24663)) ;
    mux21_ni ix54313 (.Y (nx54312), .A0 (nx54296), .A1 (nx54308), .S0 (nx23787)
             ) ;
    mux21_ni ix54297 (.Y (nx54296), .A0 (inputs_300__13), .A1 (inputs_301__13), 
             .S0 (nx24665)) ;
    mux21_ni ix54309 (.Y (nx54308), .A0 (inputs_302__13), .A1 (inputs_303__13), 
             .S0 (nx24665)) ;
    mux21_ni ix54377 (.Y (nx54376), .A0 (nx54344), .A1 (nx54372), .S0 (nx23309)
             ) ;
    mux21_ni ix54345 (.Y (nx54344), .A0 (nx54328), .A1 (nx54340), .S0 (nx23787)
             ) ;
    mux21_ni ix54329 (.Y (nx54328), .A0 (inputs_312__13), .A1 (inputs_313__13), 
             .S0 (nx24665)) ;
    mux21_ni ix54341 (.Y (nx54340), .A0 (inputs_314__13), .A1 (inputs_315__13), 
             .S0 (nx24665)) ;
    mux21_ni ix54373 (.Y (nx54372), .A0 (nx54356), .A1 (nx54368), .S0 (nx23787)
             ) ;
    mux21_ni ix54357 (.Y (nx54356), .A0 (inputs_316__13), .A1 (inputs_317__13), 
             .S0 (nx24665)) ;
    mux21_ni ix54369 (.Y (nx54368), .A0 (inputs_318__13), .A1 (inputs_319__13), 
             .S0 (nx24665)) ;
    mux21_ni ix54889 (.Y (nx54888), .A0 (nx54676), .A1 (nx54884), .S0 (nx22645)
             ) ;
    mux21_ni ix54677 (.Y (nx54676), .A0 (nx54670), .A1 (nx54592), .S0 (nx23177)
             ) ;
    oai21 ix54671 (.Y (nx54670), .A0 (nx22349), .A1 (nx19695), .B0 (nx19709)) ;
    mux21 ix19696 (.Y (nx19695), .A0 (nx54634), .A1 (nx54662), .S0 (nx23035)) ;
    mux21_ni ix54635 (.Y (nx54634), .A0 (nx54618), .A1 (nx54630), .S0 (nx23787)
             ) ;
    mux21_ni ix54619 (.Y (nx54618), .A0 (inputs_324__13), .A1 (inputs_325__13), 
             .S0 (nx24665)) ;
    mux21_ni ix54631 (.Y (nx54630), .A0 (inputs_326__13), .A1 (inputs_327__13), 
             .S0 (nx24667)) ;
    mux21_ni ix54663 (.Y (nx54662), .A0 (nx54646), .A1 (nx54658), .S0 (nx23787)
             ) ;
    mux21_ni ix54647 (.Y (nx54646), .A0 (inputs_340__13), .A1 (inputs_341__13), 
             .S0 (nx24667)) ;
    mux21_ni ix54659 (.Y (nx54658), .A0 (inputs_342__13), .A1 (inputs_343__13), 
             .S0 (nx24667)) ;
    nand04 ix19710 (.Y (nx19709), .A0 (nx22351), .A1 (nx23789), .A2 (nx24667), .A3 (
           nx54606)) ;
    mux21_ni ix54607 (.Y (nx54606), .A0 (inputs_323__13), .A1 (inputs_339__13), 
             .S0 (nx23035)) ;
    mux21_ni ix54593 (.Y (nx54592), .A0 (nx54528), .A1 (nx54588), .S0 (nx23035)
             ) ;
    mux21_ni ix54529 (.Y (nx54528), .A0 (nx54496), .A1 (nx54524), .S0 (nx23311)
             ) ;
    mux21_ni ix54497 (.Y (nx54496), .A0 (nx54480), .A1 (nx54492), .S0 (nx23789)
             ) ;
    mux21_ni ix54481 (.Y (nx54480), .A0 (inputs_328__13), .A1 (inputs_329__13), 
             .S0 (nx24667)) ;
    mux21_ni ix54493 (.Y (nx54492), .A0 (inputs_330__13), .A1 (inputs_331__13), 
             .S0 (nx24667)) ;
    mux21_ni ix54525 (.Y (nx54524), .A0 (nx54508), .A1 (nx54520), .S0 (nx23789)
             ) ;
    mux21_ni ix54509 (.Y (nx54508), .A0 (inputs_332__13), .A1 (inputs_333__13), 
             .S0 (nx24667)) ;
    mux21_ni ix54521 (.Y (nx54520), .A0 (inputs_334__13), .A1 (inputs_335__13), 
             .S0 (nx24669)) ;
    mux21_ni ix54589 (.Y (nx54588), .A0 (nx54556), .A1 (nx54584), .S0 (nx23311)
             ) ;
    mux21_ni ix54557 (.Y (nx54556), .A0 (nx54540), .A1 (nx54552), .S0 (nx23789)
             ) ;
    mux21_ni ix54541 (.Y (nx54540), .A0 (inputs_344__13), .A1 (inputs_345__13), 
             .S0 (nx24669)) ;
    mux21_ni ix54553 (.Y (nx54552), .A0 (inputs_346__13), .A1 (inputs_347__13), 
             .S0 (nx24669)) ;
    mux21_ni ix54585 (.Y (nx54584), .A0 (nx54568), .A1 (nx54580), .S0 (nx23789)
             ) ;
    mux21_ni ix54569 (.Y (nx54568), .A0 (inputs_348__13), .A1 (inputs_349__13), 
             .S0 (nx24669)) ;
    mux21_ni ix54581 (.Y (nx54580), .A0 (inputs_350__13), .A1 (inputs_351__13), 
             .S0 (nx24669)) ;
    mux21_ni ix54885 (.Y (nx54884), .A0 (nx54878), .A1 (nx54800), .S0 (nx23177)
             ) ;
    oai21 ix54879 (.Y (nx54878), .A0 (nx22351), .A1 (nx19737), .B0 (nx19749)) ;
    mux21 ix19738 (.Y (nx19737), .A0 (nx54842), .A1 (nx54870), .S0 (nx23035)) ;
    mux21_ni ix54843 (.Y (nx54842), .A0 (nx54826), .A1 (nx54838), .S0 (nx23789)
             ) ;
    mux21_ni ix54827 (.Y (nx54826), .A0 (inputs_356__13), .A1 (inputs_357__13), 
             .S0 (nx24669)) ;
    mux21_ni ix54839 (.Y (nx54838), .A0 (inputs_358__13), .A1 (inputs_359__13), 
             .S0 (nx24669)) ;
    mux21_ni ix54871 (.Y (nx54870), .A0 (nx54854), .A1 (nx54866), .S0 (nx23789)
             ) ;
    mux21_ni ix54855 (.Y (nx54854), .A0 (inputs_372__13), .A1 (inputs_373__13), 
             .S0 (nx24671)) ;
    mux21_ni ix54867 (.Y (nx54866), .A0 (inputs_374__13), .A1 (inputs_375__13), 
             .S0 (nx24671)) ;
    nand04 ix19750 (.Y (nx19749), .A0 (nx22351), .A1 (nx23791), .A2 (nx24671), .A3 (
           nx54814)) ;
    mux21_ni ix54815 (.Y (nx54814), .A0 (inputs_355__13), .A1 (inputs_371__13), 
             .S0 (nx23035)) ;
    mux21_ni ix54801 (.Y (nx54800), .A0 (nx54736), .A1 (nx54796), .S0 (nx23035)
             ) ;
    mux21_ni ix54737 (.Y (nx54736), .A0 (nx54704), .A1 (nx54732), .S0 (nx23311)
             ) ;
    mux21_ni ix54705 (.Y (nx54704), .A0 (nx54688), .A1 (nx54700), .S0 (nx23791)
             ) ;
    mux21_ni ix54689 (.Y (nx54688), .A0 (inputs_360__13), .A1 (inputs_361__13), 
             .S0 (nx24671)) ;
    mux21_ni ix54701 (.Y (nx54700), .A0 (inputs_362__13), .A1 (inputs_363__13), 
             .S0 (nx24671)) ;
    mux21_ni ix54733 (.Y (nx54732), .A0 (nx54716), .A1 (nx54728), .S0 (nx23791)
             ) ;
    mux21_ni ix54717 (.Y (nx54716), .A0 (inputs_364__13), .A1 (inputs_365__13), 
             .S0 (nx24671)) ;
    mux21_ni ix54729 (.Y (nx54728), .A0 (inputs_366__13), .A1 (inputs_367__13), 
             .S0 (nx24671)) ;
    mux21_ni ix54797 (.Y (nx54796), .A0 (nx54764), .A1 (nx54792), .S0 (nx23311)
             ) ;
    mux21_ni ix54765 (.Y (nx54764), .A0 (nx54748), .A1 (nx54760), .S0 (nx23791)
             ) ;
    mux21_ni ix54749 (.Y (nx54748), .A0 (inputs_376__13), .A1 (inputs_377__13), 
             .S0 (nx24673)) ;
    mux21_ni ix54761 (.Y (nx54760), .A0 (inputs_378__13), .A1 (inputs_379__13), 
             .S0 (nx24673)) ;
    mux21_ni ix54793 (.Y (nx54792), .A0 (nx54776), .A1 (nx54788), .S0 (nx23791)
             ) ;
    mux21_ni ix54777 (.Y (nx54776), .A0 (inputs_380__13), .A1 (inputs_381__13), 
             .S0 (nx24673)) ;
    mux21_ni ix54789 (.Y (nx54788), .A0 (inputs_382__13), .A1 (inputs_383__13), 
             .S0 (nx24673)) ;
    mux21_ni ix55737 (.Y (nx55736), .A0 (nx55312), .A1 (nx55732), .S0 (nx22509)
             ) ;
    mux21_ni ix55313 (.Y (nx55312), .A0 (nx55100), .A1 (nx55308), .S0 (nx22645)
             ) ;
    mux21_ni ix55101 (.Y (nx55100), .A0 (nx55094), .A1 (nx55016), .S0 (nx23177)
             ) ;
    oai21 ix55095 (.Y (nx55094), .A0 (nx22351), .A1 (nx19783), .B0 (nx19795)) ;
    mux21 ix19784 (.Y (nx19783), .A0 (nx55058), .A1 (nx55086), .S0 (nx23037)) ;
    mux21_ni ix55059 (.Y (nx55058), .A0 (nx55042), .A1 (nx55054), .S0 (nx23791)
             ) ;
    mux21_ni ix55043 (.Y (nx55042), .A0 (inputs_388__13), .A1 (inputs_389__13), 
             .S0 (nx24673)) ;
    mux21_ni ix55055 (.Y (nx55054), .A0 (inputs_390__13), .A1 (inputs_391__13), 
             .S0 (nx24673)) ;
    mux21_ni ix55087 (.Y (nx55086), .A0 (nx55070), .A1 (nx55082), .S0 (nx23791)
             ) ;
    mux21_ni ix55071 (.Y (nx55070), .A0 (inputs_404__13), .A1 (inputs_405__13), 
             .S0 (nx24673)) ;
    mux21_ni ix55083 (.Y (nx55082), .A0 (inputs_406__13), .A1 (inputs_407__13), 
             .S0 (nx24675)) ;
    nand04 ix19796 (.Y (nx19795), .A0 (nx22351), .A1 (nx23793), .A2 (nx24675), .A3 (
           nx55030)) ;
    mux21_ni ix55031 (.Y (nx55030), .A0 (inputs_387__13), .A1 (inputs_403__13), 
             .S0 (nx23037)) ;
    mux21_ni ix55017 (.Y (nx55016), .A0 (nx54952), .A1 (nx55012), .S0 (nx23037)
             ) ;
    mux21_ni ix54953 (.Y (nx54952), .A0 (nx54920), .A1 (nx54948), .S0 (nx23311)
             ) ;
    mux21_ni ix54921 (.Y (nx54920), .A0 (nx54904), .A1 (nx54916), .S0 (nx23793)
             ) ;
    mux21_ni ix54905 (.Y (nx54904), .A0 (inputs_392__13), .A1 (inputs_393__13), 
             .S0 (nx24675)) ;
    mux21_ni ix54917 (.Y (nx54916), .A0 (inputs_394__13), .A1 (inputs_395__13), 
             .S0 (nx24675)) ;
    mux21_ni ix54949 (.Y (nx54948), .A0 (nx54932), .A1 (nx54944), .S0 (nx23793)
             ) ;
    mux21_ni ix54933 (.Y (nx54932), .A0 (inputs_396__13), .A1 (inputs_397__13), 
             .S0 (nx24675)) ;
    mux21_ni ix54945 (.Y (nx54944), .A0 (inputs_398__13), .A1 (inputs_399__13), 
             .S0 (nx24675)) ;
    mux21_ni ix55013 (.Y (nx55012), .A0 (nx54980), .A1 (nx55008), .S0 (nx23311)
             ) ;
    mux21_ni ix54981 (.Y (nx54980), .A0 (nx54964), .A1 (nx54976), .S0 (nx23793)
             ) ;
    mux21_ni ix54965 (.Y (nx54964), .A0 (inputs_408__13), .A1 (inputs_409__13), 
             .S0 (nx24675)) ;
    mux21_ni ix54977 (.Y (nx54976), .A0 (inputs_410__13), .A1 (inputs_411__13), 
             .S0 (nx24677)) ;
    mux21_ni ix55009 (.Y (nx55008), .A0 (nx54992), .A1 (nx55004), .S0 (nx23793)
             ) ;
    mux21_ni ix54993 (.Y (nx54992), .A0 (inputs_412__13), .A1 (inputs_413__13), 
             .S0 (nx24677)) ;
    mux21_ni ix55005 (.Y (nx55004), .A0 (inputs_414__13), .A1 (inputs_415__13), 
             .S0 (nx24677)) ;
    mux21_ni ix55309 (.Y (nx55308), .A0 (nx55302), .A1 (nx55224), .S0 (nx23177)
             ) ;
    oai21 ix55303 (.Y (nx55302), .A0 (nx22351), .A1 (nx19825), .B0 (nx19839)) ;
    mux21 ix19826 (.Y (nx19825), .A0 (nx55266), .A1 (nx55294), .S0 (nx23037)) ;
    mux21_ni ix55267 (.Y (nx55266), .A0 (nx55250), .A1 (nx55262), .S0 (nx23793)
             ) ;
    mux21_ni ix55251 (.Y (nx55250), .A0 (inputs_420__13), .A1 (inputs_421__13), 
             .S0 (nx24677)) ;
    mux21_ni ix55263 (.Y (nx55262), .A0 (inputs_422__13), .A1 (inputs_423__13), 
             .S0 (nx24677)) ;
    mux21_ni ix55295 (.Y (nx55294), .A0 (nx55278), .A1 (nx55290), .S0 (nx23793)
             ) ;
    mux21_ni ix55279 (.Y (nx55278), .A0 (inputs_436__13), .A1 (inputs_437__13), 
             .S0 (nx24677)) ;
    mux21_ni ix55291 (.Y (nx55290), .A0 (inputs_438__13), .A1 (inputs_439__13), 
             .S0 (nx24677)) ;
    nand04 ix19840 (.Y (nx19839), .A0 (nx22351), .A1 (nx23795), .A2 (nx24679), .A3 (
           nx55238)) ;
    mux21_ni ix55239 (.Y (nx55238), .A0 (inputs_419__13), .A1 (inputs_435__13), 
             .S0 (nx23037)) ;
    mux21_ni ix55225 (.Y (nx55224), .A0 (nx55160), .A1 (nx55220), .S0 (nx23037)
             ) ;
    mux21_ni ix55161 (.Y (nx55160), .A0 (nx55128), .A1 (nx55156), .S0 (nx23311)
             ) ;
    mux21_ni ix55129 (.Y (nx55128), .A0 (nx55112), .A1 (nx55124), .S0 (nx23795)
             ) ;
    mux21_ni ix55113 (.Y (nx55112), .A0 (inputs_424__13), .A1 (inputs_425__13), 
             .S0 (nx24679)) ;
    mux21_ni ix55125 (.Y (nx55124), .A0 (inputs_426__13), .A1 (inputs_427__13), 
             .S0 (nx24679)) ;
    mux21_ni ix55157 (.Y (nx55156), .A0 (nx55140), .A1 (nx55152), .S0 (nx23795)
             ) ;
    mux21_ni ix55141 (.Y (nx55140), .A0 (inputs_428__13), .A1 (inputs_429__13), 
             .S0 (nx24679)) ;
    mux21_ni ix55153 (.Y (nx55152), .A0 (inputs_430__13), .A1 (inputs_431__13), 
             .S0 (nx24679)) ;
    mux21_ni ix55221 (.Y (nx55220), .A0 (nx55188), .A1 (nx55216), .S0 (nx23313)
             ) ;
    mux21_ni ix55189 (.Y (nx55188), .A0 (nx55172), .A1 (nx55184), .S0 (nx23795)
             ) ;
    mux21_ni ix55173 (.Y (nx55172), .A0 (inputs_440__13), .A1 (inputs_441__13), 
             .S0 (nx24679)) ;
    mux21_ni ix55185 (.Y (nx55184), .A0 (inputs_442__13), .A1 (inputs_443__13), 
             .S0 (nx24679)) ;
    mux21_ni ix55217 (.Y (nx55216), .A0 (nx55200), .A1 (nx55212), .S0 (nx23795)
             ) ;
    mux21_ni ix55201 (.Y (nx55200), .A0 (inputs_444__13), .A1 (inputs_445__13), 
             .S0 (nx24681)) ;
    mux21_ni ix55213 (.Y (nx55212), .A0 (inputs_446__13), .A1 (inputs_447__13), 
             .S0 (nx24681)) ;
    mux21_ni ix55733 (.Y (nx55732), .A0 (nx55520), .A1 (nx55728), .S0 (nx22645)
             ) ;
    mux21_ni ix55521 (.Y (nx55520), .A0 (nx55514), .A1 (nx55436), .S0 (nx23177)
             ) ;
    oai21 ix55515 (.Y (nx55514), .A0 (nx22353), .A1 (nx19871), .B0 (nx19883)) ;
    mux21 ix19872 (.Y (nx19871), .A0 (nx55478), .A1 (nx55506), .S0 (nx23037)) ;
    mux21_ni ix55479 (.Y (nx55478), .A0 (nx55462), .A1 (nx55474), .S0 (nx23795)
             ) ;
    mux21_ni ix55463 (.Y (nx55462), .A0 (inputs_452__13), .A1 (inputs_453__13), 
             .S0 (nx24681)) ;
    mux21_ni ix55475 (.Y (nx55474), .A0 (inputs_454__13), .A1 (inputs_455__13), 
             .S0 (nx24681)) ;
    mux21_ni ix55507 (.Y (nx55506), .A0 (nx55490), .A1 (nx55502), .S0 (nx23795)
             ) ;
    mux21_ni ix55491 (.Y (nx55490), .A0 (inputs_468__13), .A1 (inputs_469__13), 
             .S0 (nx24681)) ;
    mux21_ni ix55503 (.Y (nx55502), .A0 (inputs_470__13), .A1 (inputs_471__13), 
             .S0 (nx24681)) ;
    nand04 ix19884 (.Y (nx19883), .A0 (nx22353), .A1 (nx23797), .A2 (nx24681), .A3 (
           nx55450)) ;
    mux21_ni ix55451 (.Y (nx55450), .A0 (inputs_451__13), .A1 (inputs_467__13), 
             .S0 (nx23039)) ;
    mux21_ni ix55437 (.Y (nx55436), .A0 (nx55372), .A1 (nx55432), .S0 (nx23039)
             ) ;
    mux21_ni ix55373 (.Y (nx55372), .A0 (nx55340), .A1 (nx55368), .S0 (nx23313)
             ) ;
    mux21_ni ix55341 (.Y (nx55340), .A0 (nx55324), .A1 (nx55336), .S0 (nx23797)
             ) ;
    mux21_ni ix55325 (.Y (nx55324), .A0 (inputs_456__13), .A1 (inputs_457__13), 
             .S0 (nx24683)) ;
    mux21_ni ix55337 (.Y (nx55336), .A0 (inputs_458__13), .A1 (inputs_459__13), 
             .S0 (nx24683)) ;
    mux21_ni ix55369 (.Y (nx55368), .A0 (nx55352), .A1 (nx55364), .S0 (nx23797)
             ) ;
    mux21_ni ix55353 (.Y (nx55352), .A0 (inputs_460__13), .A1 (inputs_461__13), 
             .S0 (nx24683)) ;
    mux21_ni ix55365 (.Y (nx55364), .A0 (inputs_462__13), .A1 (inputs_463__13), 
             .S0 (nx24683)) ;
    mux21_ni ix55433 (.Y (nx55432), .A0 (nx55400), .A1 (nx55428), .S0 (nx23313)
             ) ;
    mux21_ni ix55401 (.Y (nx55400), .A0 (nx55384), .A1 (nx55396), .S0 (nx23797)
             ) ;
    mux21_ni ix55385 (.Y (nx55384), .A0 (inputs_472__13), .A1 (inputs_473__13), 
             .S0 (nx24683)) ;
    mux21_ni ix55397 (.Y (nx55396), .A0 (inputs_474__13), .A1 (inputs_475__13), 
             .S0 (nx24683)) ;
    mux21_ni ix55429 (.Y (nx55428), .A0 (nx55412), .A1 (nx55424), .S0 (nx23797)
             ) ;
    mux21_ni ix55413 (.Y (nx55412), .A0 (inputs_476__13), .A1 (inputs_477__13), 
             .S0 (nx24683)) ;
    mux21_ni ix55425 (.Y (nx55424), .A0 (inputs_478__13), .A1 (inputs_479__13), 
             .S0 (nx24685)) ;
    mux21_ni ix55729 (.Y (nx55728), .A0 (nx55722), .A1 (nx55644), .S0 (nx23177)
             ) ;
    oai21 ix55723 (.Y (nx55722), .A0 (nx22353), .A1 (nx19913), .B0 (nx19925)) ;
    mux21 ix19914 (.Y (nx19913), .A0 (nx55686), .A1 (nx55714), .S0 (nx23039)) ;
    mux21_ni ix55687 (.Y (nx55686), .A0 (nx55670), .A1 (nx55682), .S0 (nx23797)
             ) ;
    mux21_ni ix55671 (.Y (nx55670), .A0 (inputs_484__13), .A1 (inputs_485__13), 
             .S0 (nx24685)) ;
    mux21_ni ix55683 (.Y (nx55682), .A0 (inputs_486__13), .A1 (inputs_487__13), 
             .S0 (nx24685)) ;
    mux21_ni ix55715 (.Y (nx55714), .A0 (nx55698), .A1 (nx55710), .S0 (nx23797)
             ) ;
    mux21_ni ix55699 (.Y (nx55698), .A0 (inputs_500__13), .A1 (inputs_501__13), 
             .S0 (nx24685)) ;
    mux21_ni ix55711 (.Y (nx55710), .A0 (inputs_502__13), .A1 (inputs_503__13), 
             .S0 (nx24685)) ;
    nand04 ix19926 (.Y (nx19925), .A0 (nx22353), .A1 (nx23799), .A2 (nx24685), .A3 (
           nx55658)) ;
    mux21_ni ix55659 (.Y (nx55658), .A0 (inputs_483__13), .A1 (inputs_499__13), 
             .S0 (nx23039)) ;
    mux21_ni ix55645 (.Y (nx55644), .A0 (nx55580), .A1 (nx55640), .S0 (nx23039)
             ) ;
    mux21_ni ix55581 (.Y (nx55580), .A0 (nx55548), .A1 (nx55576), .S0 (nx23313)
             ) ;
    mux21_ni ix55549 (.Y (nx55548), .A0 (nx55532), .A1 (nx55544), .S0 (nx23799)
             ) ;
    mux21_ni ix55533 (.Y (nx55532), .A0 (inputs_488__13), .A1 (inputs_489__13), 
             .S0 (nx24685)) ;
    mux21_ni ix55545 (.Y (nx55544), .A0 (inputs_490__13), .A1 (inputs_491__13), 
             .S0 (nx24687)) ;
    mux21_ni ix55577 (.Y (nx55576), .A0 (nx55560), .A1 (nx55572), .S0 (nx23799)
             ) ;
    mux21_ni ix55561 (.Y (nx55560), .A0 (inputs_492__13), .A1 (inputs_493__13), 
             .S0 (nx24687)) ;
    mux21_ni ix55573 (.Y (nx55572), .A0 (inputs_494__13), .A1 (inputs_495__13), 
             .S0 (nx24687)) ;
    mux21_ni ix55641 (.Y (nx55640), .A0 (nx55608), .A1 (nx55636), .S0 (nx23313)
             ) ;
    mux21_ni ix55609 (.Y (nx55608), .A0 (nx55592), .A1 (nx55604), .S0 (nx23799)
             ) ;
    mux21_ni ix55593 (.Y (nx55592), .A0 (inputs_504__13), .A1 (inputs_505__13), 
             .S0 (nx24687)) ;
    mux21_ni ix55605 (.Y (nx55604), .A0 (inputs_506__13), .A1 (inputs_507__13), 
             .S0 (nx24687)) ;
    mux21_ni ix55637 (.Y (nx55636), .A0 (nx55620), .A1 (nx55632), .S0 (nx23799)
             ) ;
    mux21_ni ix55621 (.Y (nx55620), .A0 (inputs_508__13), .A1 (inputs_509__13), 
             .S0 (nx24687)) ;
    mux21_ni ix55633 (.Y (nx55632), .A0 (inputs_510__13), .A1 (inputs_511__13), 
             .S0 (nx24687)) ;
    aoi32 ix19954 (.Y (nx19953), .A0 (nx56506), .A1 (nx24839), .A2 (nx22353), .B0 (
          nx22223), .B1 (nx58202)) ;
    oai21 ix56507 (.Y (nx56506), .A0 (nx23799), .A1 (nx19957), .B0 (nx20059)) ;
    mux21 ix19958 (.Y (nx19957), .A0 (nx56244), .A1 (nx56496), .S0 (nx24689)) ;
    mux21_ni ix56245 (.Y (nx56244), .A0 (nx56116), .A1 (nx56240), .S0 (nx22403)
             ) ;
    mux21_ni ix56117 (.Y (nx56116), .A0 (nx56052), .A1 (nx56112), .S0 (nx22441)
             ) ;
    mux21_ni ix56053 (.Y (nx56052), .A0 (nx56020), .A1 (nx56048), .S0 (nx22511)
             ) ;
    mux21_ni ix56021 (.Y (nx56020), .A0 (nx56004), .A1 (nx56016), .S0 (nx22647)
             ) ;
    mux21_ni ix56005 (.Y (nx56004), .A0 (inputs_0__13), .A1 (inputs_16__13), .S0 (
             nx23039)) ;
    mux21_ni ix56017 (.Y (nx56016), .A0 (inputs_32__13), .A1 (inputs_48__13), .S0 (
             nx23039)) ;
    mux21_ni ix56049 (.Y (nx56048), .A0 (nx56032), .A1 (nx56044), .S0 (nx22647)
             ) ;
    mux21_ni ix56033 (.Y (nx56032), .A0 (inputs_64__13), .A1 (inputs_80__13), .S0 (
             nx23041)) ;
    mux21_ni ix56045 (.Y (nx56044), .A0 (inputs_96__13), .A1 (inputs_112__13), .S0 (
             nx23041)) ;
    mux21_ni ix56113 (.Y (nx56112), .A0 (nx56080), .A1 (nx56108), .S0 (nx22511)
             ) ;
    mux21_ni ix56081 (.Y (nx56080), .A0 (nx56064), .A1 (nx56076), .S0 (nx22647)
             ) ;
    mux21_ni ix56065 (.Y (nx56064), .A0 (inputs_128__13), .A1 (inputs_144__13), 
             .S0 (nx23041)) ;
    mux21_ni ix56077 (.Y (nx56076), .A0 (inputs_160__13), .A1 (inputs_176__13), 
             .S0 (nx23041)) ;
    mux21_ni ix56109 (.Y (nx56108), .A0 (nx56092), .A1 (nx56104), .S0 (nx22647)
             ) ;
    mux21_ni ix56093 (.Y (nx56092), .A0 (inputs_192__13), .A1 (inputs_208__13), 
             .S0 (nx23041)) ;
    mux21_ni ix56105 (.Y (nx56104), .A0 (inputs_224__13), .A1 (inputs_240__13), 
             .S0 (nx23041)) ;
    mux21_ni ix56241 (.Y (nx56240), .A0 (nx56176), .A1 (nx56236), .S0 (nx22441)
             ) ;
    mux21_ni ix56177 (.Y (nx56176), .A0 (nx56144), .A1 (nx56172), .S0 (nx22511)
             ) ;
    mux21_ni ix56145 (.Y (nx56144), .A0 (nx56128), .A1 (nx56140), .S0 (nx22647)
             ) ;
    mux21_ni ix56129 (.Y (nx56128), .A0 (inputs_256__13), .A1 (inputs_272__13), 
             .S0 (nx23041)) ;
    mux21_ni ix56141 (.Y (nx56140), .A0 (inputs_288__13), .A1 (inputs_304__13), 
             .S0 (nx23043)) ;
    mux21_ni ix56173 (.Y (nx56172), .A0 (nx56156), .A1 (nx56168), .S0 (nx22647)
             ) ;
    mux21_ni ix56157 (.Y (nx56156), .A0 (inputs_320__13), .A1 (inputs_336__13), 
             .S0 (nx23043)) ;
    mux21_ni ix56169 (.Y (nx56168), .A0 (inputs_352__13), .A1 (inputs_368__13), 
             .S0 (nx23043)) ;
    mux21_ni ix56237 (.Y (nx56236), .A0 (nx56204), .A1 (nx56232), .S0 (nx22511)
             ) ;
    mux21_ni ix56205 (.Y (nx56204), .A0 (nx56188), .A1 (nx56200), .S0 (nx22647)
             ) ;
    mux21_ni ix56189 (.Y (nx56188), .A0 (inputs_384__13), .A1 (inputs_400__13), 
             .S0 (nx23043)) ;
    mux21_ni ix56201 (.Y (nx56200), .A0 (inputs_416__13), .A1 (inputs_432__13), 
             .S0 (nx23043)) ;
    mux21_ni ix56233 (.Y (nx56232), .A0 (nx56216), .A1 (nx56228), .S0 (nx22649)
             ) ;
    mux21_ni ix56217 (.Y (nx56216), .A0 (inputs_448__13), .A1 (inputs_464__13), 
             .S0 (nx23043)) ;
    mux21_ni ix56229 (.Y (nx56228), .A0 (inputs_480__13), .A1 (inputs_496__13), 
             .S0 (nx23043)) ;
    mux21_ni ix56497 (.Y (nx56496), .A0 (nx56368), .A1 (nx56492), .S0 (nx22403)
             ) ;
    mux21_ni ix56369 (.Y (nx56368), .A0 (nx56304), .A1 (nx56364), .S0 (nx22441)
             ) ;
    mux21_ni ix56305 (.Y (nx56304), .A0 (nx56272), .A1 (nx56300), .S0 (nx22511)
             ) ;
    mux21_ni ix56273 (.Y (nx56272), .A0 (nx56256), .A1 (nx56268), .S0 (nx22649)
             ) ;
    mux21_ni ix56257 (.Y (nx56256), .A0 (inputs_1__13), .A1 (inputs_17__13), .S0 (
             nx23045)) ;
    mux21_ni ix56269 (.Y (nx56268), .A0 (inputs_33__13), .A1 (inputs_49__13), .S0 (
             nx23045)) ;
    mux21_ni ix56301 (.Y (nx56300), .A0 (nx56284), .A1 (nx56296), .S0 (nx22649)
             ) ;
    mux21_ni ix56285 (.Y (nx56284), .A0 (inputs_65__13), .A1 (inputs_81__13), .S0 (
             nx23045)) ;
    mux21_ni ix56297 (.Y (nx56296), .A0 (inputs_97__13), .A1 (inputs_113__13), .S0 (
             nx23045)) ;
    mux21_ni ix56365 (.Y (nx56364), .A0 (nx56332), .A1 (nx56360), .S0 (nx22511)
             ) ;
    mux21_ni ix56333 (.Y (nx56332), .A0 (nx56316), .A1 (nx56328), .S0 (nx22649)
             ) ;
    mux21_ni ix56317 (.Y (nx56316), .A0 (inputs_129__13), .A1 (inputs_145__13), 
             .S0 (nx23045)) ;
    mux21_ni ix56329 (.Y (nx56328), .A0 (inputs_161__13), .A1 (inputs_177__13), 
             .S0 (nx23045)) ;
    mux21_ni ix56361 (.Y (nx56360), .A0 (nx56344), .A1 (nx56356), .S0 (nx22649)
             ) ;
    mux21_ni ix56345 (.Y (nx56344), .A0 (inputs_193__13), .A1 (inputs_209__13), 
             .S0 (nx23045)) ;
    mux21_ni ix56357 (.Y (nx56356), .A0 (inputs_225__13), .A1 (inputs_241__13), 
             .S0 (nx23047)) ;
    mux21_ni ix56493 (.Y (nx56492), .A0 (nx56428), .A1 (nx56488), .S0 (nx22441)
             ) ;
    mux21_ni ix56429 (.Y (nx56428), .A0 (nx56396), .A1 (nx56424), .S0 (nx22511)
             ) ;
    mux21_ni ix56397 (.Y (nx56396), .A0 (nx56380), .A1 (nx56392), .S0 (nx22649)
             ) ;
    mux21_ni ix56381 (.Y (nx56380), .A0 (inputs_257__13), .A1 (inputs_273__13), 
             .S0 (nx23047)) ;
    mux21_ni ix56393 (.Y (nx56392), .A0 (inputs_289__13), .A1 (inputs_305__13), 
             .S0 (nx23047)) ;
    mux21_ni ix56425 (.Y (nx56424), .A0 (nx56408), .A1 (nx56420), .S0 (nx22649)
             ) ;
    mux21_ni ix56409 (.Y (nx56408), .A0 (inputs_321__13), .A1 (inputs_337__13), 
             .S0 (nx23047)) ;
    mux21_ni ix56421 (.Y (nx56420), .A0 (inputs_353__13), .A1 (inputs_369__13), 
             .S0 (nx23047)) ;
    mux21_ni ix56489 (.Y (nx56488), .A0 (nx56456), .A1 (nx56484), .S0 (nx22513)
             ) ;
    mux21_ni ix56457 (.Y (nx56456), .A0 (nx56440), .A1 (nx56452), .S0 (nx22651)
             ) ;
    mux21_ni ix56441 (.Y (nx56440), .A0 (inputs_385__13), .A1 (inputs_401__13), 
             .S0 (nx23047)) ;
    mux21_ni ix56453 (.Y (nx56452), .A0 (inputs_417__13), .A1 (inputs_433__13), 
             .S0 (nx23047)) ;
    mux21_ni ix56485 (.Y (nx56484), .A0 (nx56468), .A1 (nx56480), .S0 (nx22651)
             ) ;
    mux21_ni ix56469 (.Y (nx56468), .A0 (inputs_449__13), .A1 (inputs_465__13), 
             .S0 (nx23049)) ;
    mux21_ni ix56481 (.Y (nx56480), .A0 (inputs_481__13), .A1 (inputs_497__13), 
             .S0 (nx23049)) ;
    nand03 ix20060 (.Y (nx20059), .A0 (nx55990), .A1 (nx23799), .A2 (nx22381)) ;
    mux21_ni ix55991 (.Y (nx55990), .A0 (nx55862), .A1 (nx55986), .S0 (nx22403)
             ) ;
    mux21_ni ix55863 (.Y (nx55862), .A0 (nx55798), .A1 (nx55858), .S0 (nx22441)
             ) ;
    mux21_ni ix55799 (.Y (nx55798), .A0 (nx55766), .A1 (nx55794), .S0 (nx22513)
             ) ;
    mux21_ni ix55767 (.Y (nx55766), .A0 (nx55750), .A1 (nx55762), .S0 (nx22651)
             ) ;
    mux21_ni ix55751 (.Y (nx55750), .A0 (inputs_2__13), .A1 (inputs_18__13), .S0 (
             nx23049)) ;
    mux21_ni ix55763 (.Y (nx55762), .A0 (inputs_34__13), .A1 (inputs_50__13), .S0 (
             nx23049)) ;
    mux21_ni ix55795 (.Y (nx55794), .A0 (nx55778), .A1 (nx55790), .S0 (nx22651)
             ) ;
    mux21_ni ix55779 (.Y (nx55778), .A0 (inputs_66__13), .A1 (inputs_82__13), .S0 (
             nx23049)) ;
    mux21_ni ix55791 (.Y (nx55790), .A0 (inputs_98__13), .A1 (inputs_114__13), .S0 (
             nx23049)) ;
    mux21_ni ix55859 (.Y (nx55858), .A0 (nx55826), .A1 (nx55854), .S0 (nx22513)
             ) ;
    mux21_ni ix55827 (.Y (nx55826), .A0 (nx55810), .A1 (nx55822), .S0 (nx22651)
             ) ;
    mux21_ni ix55811 (.Y (nx55810), .A0 (inputs_130__13), .A1 (inputs_146__13), 
             .S0 (nx23049)) ;
    mux21_ni ix55823 (.Y (nx55822), .A0 (inputs_162__13), .A1 (inputs_178__13), 
             .S0 (nx23051)) ;
    mux21_ni ix55855 (.Y (nx55854), .A0 (nx55838), .A1 (nx55850), .S0 (nx22651)
             ) ;
    mux21_ni ix55839 (.Y (nx55838), .A0 (inputs_194__13), .A1 (inputs_210__13), 
             .S0 (nx23051)) ;
    mux21_ni ix55851 (.Y (nx55850), .A0 (inputs_226__13), .A1 (inputs_242__13), 
             .S0 (nx23051)) ;
    mux21_ni ix55987 (.Y (nx55986), .A0 (nx55922), .A1 (nx55982), .S0 (nx22441)
             ) ;
    mux21_ni ix55923 (.Y (nx55922), .A0 (nx55890), .A1 (nx55918), .S0 (nx22513)
             ) ;
    mux21_ni ix55891 (.Y (nx55890), .A0 (nx55874), .A1 (nx55886), .S0 (nx22651)
             ) ;
    mux21_ni ix55875 (.Y (nx55874), .A0 (inputs_258__13), .A1 (inputs_274__13), 
             .S0 (nx23051)) ;
    mux21_ni ix55887 (.Y (nx55886), .A0 (inputs_290__13), .A1 (inputs_306__13), 
             .S0 (nx23051)) ;
    mux21_ni ix55919 (.Y (nx55918), .A0 (nx55902), .A1 (nx55914), .S0 (nx22653)
             ) ;
    mux21_ni ix55903 (.Y (nx55902), .A0 (inputs_322__13), .A1 (inputs_338__13), 
             .S0 (nx23051)) ;
    mux21_ni ix55915 (.Y (nx55914), .A0 (inputs_354__13), .A1 (inputs_370__13), 
             .S0 (nx23051)) ;
    mux21_ni ix55983 (.Y (nx55982), .A0 (nx55950), .A1 (nx55978), .S0 (nx22513)
             ) ;
    mux21_ni ix55951 (.Y (nx55950), .A0 (nx55934), .A1 (nx55946), .S0 (nx22653)
             ) ;
    mux21_ni ix55935 (.Y (nx55934), .A0 (inputs_386__13), .A1 (inputs_402__13), 
             .S0 (nx23053)) ;
    mux21_ni ix55947 (.Y (nx55946), .A0 (inputs_418__13), .A1 (inputs_434__13), 
             .S0 (nx23053)) ;
    mux21_ni ix55979 (.Y (nx55978), .A0 (nx55962), .A1 (nx55974), .S0 (nx22653)
             ) ;
    mux21_ni ix55963 (.Y (nx55962), .A0 (inputs_450__13), .A1 (inputs_466__13), 
             .S0 (nx23053)) ;
    mux21_ni ix55975 (.Y (nx55974), .A0 (inputs_482__13), .A1 (inputs_498__13), 
             .S0 (nx23053)) ;
    mux21_ni ix58203 (.Y (nx58202), .A0 (nx57354), .A1 (nx58198), .S0 (nx22441)
             ) ;
    mux21_ni ix57355 (.Y (nx57354), .A0 (nx56930), .A1 (nx57350), .S0 (nx22513)
             ) ;
    mux21_ni ix56931 (.Y (nx56930), .A0 (nx56718), .A1 (nx56926), .S0 (nx22653)
             ) ;
    mux21_ni ix56719 (.Y (nx56718), .A0 (nx56712), .A1 (nx56634), .S0 (nx23177)
             ) ;
    oai21 ix56713 (.Y (nx56712), .A0 (nx22353), .A1 (nx20117), .B0 (nx20131)) ;
    mux21 ix20118 (.Y (nx20117), .A0 (nx56676), .A1 (nx56704), .S0 (nx23053)) ;
    mux21_ni ix56677 (.Y (nx56676), .A0 (nx56660), .A1 (nx56672), .S0 (nx23801)
             ) ;
    mux21_ni ix56661 (.Y (nx56660), .A0 (inputs_4__13), .A1 (inputs_5__13), .S0 (
             nx24689)) ;
    mux21_ni ix56673 (.Y (nx56672), .A0 (inputs_6__13), .A1 (inputs_7__13), .S0 (
             nx24689)) ;
    mux21_ni ix56705 (.Y (nx56704), .A0 (nx56688), .A1 (nx56700), .S0 (nx23801)
             ) ;
    mux21_ni ix56689 (.Y (nx56688), .A0 (inputs_20__13), .A1 (inputs_21__13), .S0 (
             nx24689)) ;
    mux21_ni ix56701 (.Y (nx56700), .A0 (inputs_22__13), .A1 (inputs_23__13), .S0 (
             nx24689)) ;
    nand04 ix20132 (.Y (nx20131), .A0 (nx22353), .A1 (nx23801), .A2 (nx24689), .A3 (
           nx56648)) ;
    mux21_ni ix56649 (.Y (nx56648), .A0 (inputs_3__13), .A1 (inputs_19__13), .S0 (
             nx23053)) ;
    mux21_ni ix56635 (.Y (nx56634), .A0 (nx56570), .A1 (nx56630), .S0 (nx23053)
             ) ;
    mux21_ni ix56571 (.Y (nx56570), .A0 (nx56538), .A1 (nx56566), .S0 (nx23313)
             ) ;
    mux21_ni ix56539 (.Y (nx56538), .A0 (nx56522), .A1 (nx56534), .S0 (nx23801)
             ) ;
    mux21_ni ix56523 (.Y (nx56522), .A0 (inputs_8__13), .A1 (inputs_9__13), .S0 (
             nx24689)) ;
    mux21_ni ix56535 (.Y (nx56534), .A0 (inputs_10__13), .A1 (inputs_11__13), .S0 (
             nx24691)) ;
    mux21_ni ix56567 (.Y (nx56566), .A0 (nx56550), .A1 (nx56562), .S0 (nx23801)
             ) ;
    mux21_ni ix56551 (.Y (nx56550), .A0 (inputs_12__13), .A1 (inputs_13__13), .S0 (
             nx24691)) ;
    mux21_ni ix56563 (.Y (nx56562), .A0 (inputs_14__13), .A1 (inputs_15__13), .S0 (
             nx24691)) ;
    mux21_ni ix56631 (.Y (nx56630), .A0 (nx56598), .A1 (nx56626), .S0 (nx23313)
             ) ;
    mux21_ni ix56599 (.Y (nx56598), .A0 (nx56582), .A1 (nx56594), .S0 (nx23801)
             ) ;
    mux21_ni ix56583 (.Y (nx56582), .A0 (inputs_24__13), .A1 (inputs_25__13), .S0 (
             nx24691)) ;
    mux21_ni ix56595 (.Y (nx56594), .A0 (inputs_26__13), .A1 (inputs_27__13), .S0 (
             nx24691)) ;
    mux21_ni ix56627 (.Y (nx56626), .A0 (nx56610), .A1 (nx56622), .S0 (nx23801)
             ) ;
    mux21_ni ix56611 (.Y (nx56610), .A0 (inputs_28__13), .A1 (inputs_29__13), .S0 (
             nx24691)) ;
    mux21_ni ix56623 (.Y (nx56622), .A0 (inputs_30__13), .A1 (inputs_31__13), .S0 (
             nx24691)) ;
    mux21_ni ix56927 (.Y (nx56926), .A0 (nx56920), .A1 (nx56842), .S0 (nx23179)
             ) ;
    oai21 ix56921 (.Y (nx56920), .A0 (nx22355), .A1 (nx20161), .B0 (nx20173)) ;
    mux21 ix20162 (.Y (nx20161), .A0 (nx56884), .A1 (nx56912), .S0 (nx23055)) ;
    mux21_ni ix56885 (.Y (nx56884), .A0 (nx56868), .A1 (nx56880), .S0 (nx23803)
             ) ;
    mux21_ni ix56869 (.Y (nx56868), .A0 (inputs_36__13), .A1 (inputs_37__13), .S0 (
             nx24693)) ;
    mux21_ni ix56881 (.Y (nx56880), .A0 (inputs_38__13), .A1 (inputs_39__13), .S0 (
             nx24693)) ;
    mux21_ni ix56913 (.Y (nx56912), .A0 (nx56896), .A1 (nx56908), .S0 (nx23803)
             ) ;
    mux21_ni ix56897 (.Y (nx56896), .A0 (inputs_52__13), .A1 (inputs_53__13), .S0 (
             nx24693)) ;
    mux21_ni ix56909 (.Y (nx56908), .A0 (inputs_54__13), .A1 (inputs_55__13), .S0 (
             nx24693)) ;
    nand04 ix20174 (.Y (nx20173), .A0 (nx22355), .A1 (nx23803), .A2 (nx24693), .A3 (
           nx56856)) ;
    mux21_ni ix56857 (.Y (nx56856), .A0 (inputs_35__13), .A1 (inputs_51__13), .S0 (
             nx23055)) ;
    mux21_ni ix56843 (.Y (nx56842), .A0 (nx56778), .A1 (nx56838), .S0 (nx23055)
             ) ;
    mux21_ni ix56779 (.Y (nx56778), .A0 (nx56746), .A1 (nx56774), .S0 (nx23315)
             ) ;
    mux21_ni ix56747 (.Y (nx56746), .A0 (nx56730), .A1 (nx56742), .S0 (nx23803)
             ) ;
    mux21_ni ix56731 (.Y (nx56730), .A0 (inputs_40__13), .A1 (inputs_41__13), .S0 (
             nx24693)) ;
    mux21_ni ix56743 (.Y (nx56742), .A0 (inputs_42__13), .A1 (inputs_43__13), .S0 (
             nx24693)) ;
    mux21_ni ix56775 (.Y (nx56774), .A0 (nx56758), .A1 (nx56770), .S0 (nx23803)
             ) ;
    mux21_ni ix56759 (.Y (nx56758), .A0 (inputs_44__13), .A1 (inputs_45__13), .S0 (
             nx24695)) ;
    mux21_ni ix56771 (.Y (nx56770), .A0 (inputs_46__13), .A1 (inputs_47__13), .S0 (
             nx24695)) ;
    mux21_ni ix56839 (.Y (nx56838), .A0 (nx56806), .A1 (nx56834), .S0 (nx23315)
             ) ;
    mux21_ni ix56807 (.Y (nx56806), .A0 (nx56790), .A1 (nx56802), .S0 (nx23803)
             ) ;
    mux21_ni ix56791 (.Y (nx56790), .A0 (inputs_56__13), .A1 (inputs_57__13), .S0 (
             nx24695)) ;
    mux21_ni ix56803 (.Y (nx56802), .A0 (inputs_58__13), .A1 (inputs_59__13), .S0 (
             nx24695)) ;
    mux21_ni ix56835 (.Y (nx56834), .A0 (nx56818), .A1 (nx56830), .S0 (nx23803)
             ) ;
    mux21_ni ix56819 (.Y (nx56818), .A0 (inputs_60__13), .A1 (inputs_61__13), .S0 (
             nx24695)) ;
    mux21_ni ix56831 (.Y (nx56830), .A0 (inputs_62__13), .A1 (inputs_63__13), .S0 (
             nx24695)) ;
    mux21_ni ix57351 (.Y (nx57350), .A0 (nx57138), .A1 (nx57346), .S0 (nx22653)
             ) ;
    mux21_ni ix57139 (.Y (nx57138), .A0 (nx57132), .A1 (nx57054), .S0 (nx23179)
             ) ;
    oai21 ix57133 (.Y (nx57132), .A0 (nx22355), .A1 (nx20205), .B0 (nx20217)) ;
    mux21 ix20206 (.Y (nx20205), .A0 (nx57096), .A1 (nx57124), .S0 (nx23055)) ;
    mux21_ni ix57097 (.Y (nx57096), .A0 (nx57080), .A1 (nx57092), .S0 (nx23805)
             ) ;
    mux21_ni ix57081 (.Y (nx57080), .A0 (inputs_68__13), .A1 (inputs_69__13), .S0 (
             nx24695)) ;
    mux21_ni ix57093 (.Y (nx57092), .A0 (inputs_70__13), .A1 (inputs_71__13), .S0 (
             nx24697)) ;
    mux21_ni ix57125 (.Y (nx57124), .A0 (nx57108), .A1 (nx57120), .S0 (nx23805)
             ) ;
    mux21_ni ix57109 (.Y (nx57108), .A0 (inputs_84__13), .A1 (inputs_85__13), .S0 (
             nx24697)) ;
    mux21_ni ix57121 (.Y (nx57120), .A0 (inputs_86__13), .A1 (inputs_87__13), .S0 (
             nx24697)) ;
    nand04 ix20218 (.Y (nx20217), .A0 (nx22355), .A1 (nx23805), .A2 (nx24697), .A3 (
           nx57068)) ;
    mux21_ni ix57069 (.Y (nx57068), .A0 (inputs_67__13), .A1 (inputs_83__13), .S0 (
             nx23055)) ;
    mux21_ni ix57055 (.Y (nx57054), .A0 (nx56990), .A1 (nx57050), .S0 (nx23055)
             ) ;
    mux21_ni ix56991 (.Y (nx56990), .A0 (nx56958), .A1 (nx56986), .S0 (nx23315)
             ) ;
    mux21_ni ix56959 (.Y (nx56958), .A0 (nx56942), .A1 (nx56954), .S0 (nx23805)
             ) ;
    mux21_ni ix56943 (.Y (nx56942), .A0 (inputs_72__13), .A1 (inputs_73__13), .S0 (
             nx24697)) ;
    mux21_ni ix56955 (.Y (nx56954), .A0 (inputs_74__13), .A1 (inputs_75__13), .S0 (
             nx24697)) ;
    mux21_ni ix56987 (.Y (nx56986), .A0 (nx56970), .A1 (nx56982), .S0 (nx23805)
             ) ;
    mux21_ni ix56971 (.Y (nx56970), .A0 (inputs_76__13), .A1 (inputs_77__13), .S0 (
             nx24697)) ;
    mux21_ni ix56983 (.Y (nx56982), .A0 (inputs_78__13), .A1 (inputs_79__13), .S0 (
             nx24699)) ;
    mux21_ni ix57051 (.Y (nx57050), .A0 (nx57018), .A1 (nx57046), .S0 (nx23315)
             ) ;
    mux21_ni ix57019 (.Y (nx57018), .A0 (nx57002), .A1 (nx57014), .S0 (nx23805)
             ) ;
    mux21_ni ix57003 (.Y (nx57002), .A0 (inputs_88__13), .A1 (inputs_89__13), .S0 (
             nx24699)) ;
    mux21_ni ix57015 (.Y (nx57014), .A0 (inputs_90__13), .A1 (inputs_91__13), .S0 (
             nx24699)) ;
    mux21_ni ix57047 (.Y (nx57046), .A0 (nx57030), .A1 (nx57042), .S0 (nx23805)
             ) ;
    mux21_ni ix57031 (.Y (nx57030), .A0 (inputs_92__13), .A1 (inputs_93__13), .S0 (
             nx24699)) ;
    mux21_ni ix57043 (.Y (nx57042), .A0 (inputs_94__13), .A1 (inputs_95__13), .S0 (
             nx24699)) ;
    mux21_ni ix57347 (.Y (nx57346), .A0 (nx57340), .A1 (nx57262), .S0 (nx23179)
             ) ;
    oai21 ix57341 (.Y (nx57340), .A0 (nx22355), .A1 (nx20247), .B0 (nx20261)) ;
    mux21 ix20248 (.Y (nx20247), .A0 (nx57304), .A1 (nx57332), .S0 (nx23055)) ;
    mux21_ni ix57305 (.Y (nx57304), .A0 (nx57288), .A1 (nx57300), .S0 (nx23807)
             ) ;
    mux21_ni ix57289 (.Y (nx57288), .A0 (inputs_100__13), .A1 (inputs_101__13), 
             .S0 (nx24699)) ;
    mux21_ni ix57301 (.Y (nx57300), .A0 (inputs_102__13), .A1 (inputs_103__13), 
             .S0 (nx24699)) ;
    mux21_ni ix57333 (.Y (nx57332), .A0 (nx57316), .A1 (nx57328), .S0 (nx23807)
             ) ;
    mux21_ni ix57317 (.Y (nx57316), .A0 (inputs_116__13), .A1 (inputs_117__13), 
             .S0 (nx24701)) ;
    mux21_ni ix57329 (.Y (nx57328), .A0 (inputs_118__13), .A1 (inputs_119__13), 
             .S0 (nx24701)) ;
    nand04 ix20262 (.Y (nx20261), .A0 (nx22355), .A1 (nx23807), .A2 (nx24701), .A3 (
           nx57276)) ;
    mux21_ni ix57277 (.Y (nx57276), .A0 (inputs_99__13), .A1 (inputs_115__13), .S0 (
             nx23057)) ;
    mux21_ni ix57263 (.Y (nx57262), .A0 (nx57198), .A1 (nx57258), .S0 (nx23057)
             ) ;
    mux21_ni ix57199 (.Y (nx57198), .A0 (nx57166), .A1 (nx57194), .S0 (nx23315)
             ) ;
    mux21_ni ix57167 (.Y (nx57166), .A0 (nx57150), .A1 (nx57162), .S0 (nx23807)
             ) ;
    mux21_ni ix57151 (.Y (nx57150), .A0 (inputs_104__13), .A1 (inputs_105__13), 
             .S0 (nx24701)) ;
    mux21_ni ix57163 (.Y (nx57162), .A0 (inputs_106__13), .A1 (inputs_107__13), 
             .S0 (nx24701)) ;
    mux21_ni ix57195 (.Y (nx57194), .A0 (nx57178), .A1 (nx57190), .S0 (nx23807)
             ) ;
    mux21_ni ix57179 (.Y (nx57178), .A0 (inputs_108__13), .A1 (inputs_109__13), 
             .S0 (nx24701)) ;
    mux21_ni ix57191 (.Y (nx57190), .A0 (inputs_110__13), .A1 (inputs_111__13), 
             .S0 (nx24701)) ;
    mux21_ni ix57259 (.Y (nx57258), .A0 (nx57226), .A1 (nx57254), .S0 (nx23315)
             ) ;
    mux21_ni ix57227 (.Y (nx57226), .A0 (nx57210), .A1 (nx57222), .S0 (nx23807)
             ) ;
    mux21_ni ix57211 (.Y (nx57210), .A0 (inputs_120__13), .A1 (inputs_121__13), 
             .S0 (nx24703)) ;
    mux21_ni ix57223 (.Y (nx57222), .A0 (inputs_122__13), .A1 (inputs_123__13), 
             .S0 (nx24703)) ;
    mux21_ni ix57255 (.Y (nx57254), .A0 (nx57238), .A1 (nx57250), .S0 (nx23807)
             ) ;
    mux21_ni ix57239 (.Y (nx57238), .A0 (inputs_124__13), .A1 (inputs_125__13), 
             .S0 (nx24703)) ;
    mux21_ni ix57251 (.Y (nx57250), .A0 (inputs_126__13), .A1 (inputs_127__13), 
             .S0 (nx24703)) ;
    mux21_ni ix58199 (.Y (nx58198), .A0 (nx57774), .A1 (nx58194), .S0 (nx22513)
             ) ;
    mux21_ni ix57775 (.Y (nx57774), .A0 (nx57562), .A1 (nx57770), .S0 (nx22653)
             ) ;
    mux21_ni ix57563 (.Y (nx57562), .A0 (nx57556), .A1 (nx57478), .S0 (nx23179)
             ) ;
    oai21 ix57557 (.Y (nx57556), .A0 (nx22355), .A1 (nx20295), .B0 (nx20307)) ;
    mux21 ix20296 (.Y (nx20295), .A0 (nx57520), .A1 (nx57548), .S0 (nx23057)) ;
    mux21_ni ix57521 (.Y (nx57520), .A0 (nx57504), .A1 (nx57516), .S0 (nx23809)
             ) ;
    mux21_ni ix57505 (.Y (nx57504), .A0 (inputs_132__13), .A1 (inputs_133__13), 
             .S0 (nx24703)) ;
    mux21_ni ix57517 (.Y (nx57516), .A0 (inputs_134__13), .A1 (inputs_135__13), 
             .S0 (nx24703)) ;
    mux21_ni ix57549 (.Y (nx57548), .A0 (nx57532), .A1 (nx57544), .S0 (nx23809)
             ) ;
    mux21_ni ix57533 (.Y (nx57532), .A0 (inputs_148__13), .A1 (inputs_149__13), 
             .S0 (nx24703)) ;
    mux21_ni ix57545 (.Y (nx57544), .A0 (inputs_150__13), .A1 (inputs_151__13), 
             .S0 (nx24705)) ;
    nand04 ix20308 (.Y (nx20307), .A0 (nx22357), .A1 (nx23809), .A2 (nx24705), .A3 (
           nx57492)) ;
    mux21_ni ix57493 (.Y (nx57492), .A0 (inputs_131__13), .A1 (inputs_147__13), 
             .S0 (nx23057)) ;
    mux21_ni ix57479 (.Y (nx57478), .A0 (nx57414), .A1 (nx57474), .S0 (nx23057)
             ) ;
    mux21_ni ix57415 (.Y (nx57414), .A0 (nx57382), .A1 (nx57410), .S0 (nx23315)
             ) ;
    mux21_ni ix57383 (.Y (nx57382), .A0 (nx57366), .A1 (nx57378), .S0 (nx23809)
             ) ;
    mux21_ni ix57367 (.Y (nx57366), .A0 (inputs_136__13), .A1 (inputs_137__13), 
             .S0 (nx24705)) ;
    mux21_ni ix57379 (.Y (nx57378), .A0 (inputs_138__13), .A1 (inputs_139__13), 
             .S0 (nx24705)) ;
    mux21_ni ix57411 (.Y (nx57410), .A0 (nx57394), .A1 (nx57406), .S0 (nx23809)
             ) ;
    mux21_ni ix57395 (.Y (nx57394), .A0 (inputs_140__13), .A1 (inputs_141__13), 
             .S0 (nx24705)) ;
    mux21_ni ix57407 (.Y (nx57406), .A0 (inputs_142__13), .A1 (inputs_143__13), 
             .S0 (nx24705)) ;
    mux21_ni ix57475 (.Y (nx57474), .A0 (nx57442), .A1 (nx57470), .S0 (nx23317)
             ) ;
    mux21_ni ix57443 (.Y (nx57442), .A0 (nx57426), .A1 (nx57438), .S0 (nx23809)
             ) ;
    mux21_ni ix57427 (.Y (nx57426), .A0 (inputs_152__13), .A1 (inputs_153__13), 
             .S0 (nx24705)) ;
    mux21_ni ix57439 (.Y (nx57438), .A0 (inputs_154__13), .A1 (inputs_155__13), 
             .S0 (nx24707)) ;
    mux21_ni ix57471 (.Y (nx57470), .A0 (nx57454), .A1 (nx57466), .S0 (nx23809)
             ) ;
    mux21_ni ix57455 (.Y (nx57454), .A0 (inputs_156__13), .A1 (inputs_157__13), 
             .S0 (nx24707)) ;
    mux21_ni ix57467 (.Y (nx57466), .A0 (inputs_158__13), .A1 (inputs_159__13), 
             .S0 (nx24707)) ;
    mux21_ni ix57771 (.Y (nx57770), .A0 (nx57764), .A1 (nx57686), .S0 (nx23179)
             ) ;
    oai21 ix57765 (.Y (nx57764), .A0 (nx22357), .A1 (nx20337), .B0 (nx20349)) ;
    mux21 ix20338 (.Y (nx20337), .A0 (nx57728), .A1 (nx57756), .S0 (nx23057)) ;
    mux21_ni ix57729 (.Y (nx57728), .A0 (nx57712), .A1 (nx57724), .S0 (nx23811)
             ) ;
    mux21_ni ix57713 (.Y (nx57712), .A0 (inputs_164__13), .A1 (inputs_165__13), 
             .S0 (nx24707)) ;
    mux21_ni ix57725 (.Y (nx57724), .A0 (inputs_166__13), .A1 (inputs_167__13), 
             .S0 (nx24707)) ;
    mux21_ni ix57757 (.Y (nx57756), .A0 (nx57740), .A1 (nx57752), .S0 (nx23811)
             ) ;
    mux21_ni ix57741 (.Y (nx57740), .A0 (inputs_180__13), .A1 (inputs_181__13), 
             .S0 (nx24707)) ;
    mux21_ni ix57753 (.Y (nx57752), .A0 (inputs_182__13), .A1 (inputs_183__13), 
             .S0 (nx24707)) ;
    nand04 ix20350 (.Y (nx20349), .A0 (nx22357), .A1 (nx23811), .A2 (nx24709), .A3 (
           nx57700)) ;
    mux21_ni ix57701 (.Y (nx57700), .A0 (inputs_163__13), .A1 (inputs_179__13), 
             .S0 (nx23057)) ;
    mux21_ni ix57687 (.Y (nx57686), .A0 (nx57622), .A1 (nx57682), .S0 (nx23059)
             ) ;
    mux21_ni ix57623 (.Y (nx57622), .A0 (nx57590), .A1 (nx57618), .S0 (nx23317)
             ) ;
    mux21_ni ix57591 (.Y (nx57590), .A0 (nx57574), .A1 (nx57586), .S0 (nx23811)
             ) ;
    mux21_ni ix57575 (.Y (nx57574), .A0 (inputs_168__13), .A1 (inputs_169__13), 
             .S0 (nx24709)) ;
    mux21_ni ix57587 (.Y (nx57586), .A0 (inputs_170__13), .A1 (inputs_171__13), 
             .S0 (nx24709)) ;
    mux21_ni ix57619 (.Y (nx57618), .A0 (nx57602), .A1 (nx57614), .S0 (nx23811)
             ) ;
    mux21_ni ix57603 (.Y (nx57602), .A0 (inputs_172__13), .A1 (inputs_173__13), 
             .S0 (nx24709)) ;
    mux21_ni ix57615 (.Y (nx57614), .A0 (inputs_174__13), .A1 (inputs_175__13), 
             .S0 (nx24709)) ;
    mux21_ni ix57683 (.Y (nx57682), .A0 (nx57650), .A1 (nx57678), .S0 (nx23317)
             ) ;
    mux21_ni ix57651 (.Y (nx57650), .A0 (nx57634), .A1 (nx57646), .S0 (nx23811)
             ) ;
    mux21_ni ix57635 (.Y (nx57634), .A0 (inputs_184__13), .A1 (inputs_185__13), 
             .S0 (nx24709)) ;
    mux21_ni ix57647 (.Y (nx57646), .A0 (inputs_186__13), .A1 (inputs_187__13), 
             .S0 (nx24709)) ;
    mux21_ni ix57679 (.Y (nx57678), .A0 (nx57662), .A1 (nx57674), .S0 (nx23811)
             ) ;
    mux21_ni ix57663 (.Y (nx57662), .A0 (inputs_188__13), .A1 (inputs_189__13), 
             .S0 (nx24711)) ;
    mux21_ni ix57675 (.Y (nx57674), .A0 (inputs_190__13), .A1 (inputs_191__13), 
             .S0 (nx24711)) ;
    mux21_ni ix58195 (.Y (nx58194), .A0 (nx57982), .A1 (nx58190), .S0 (nx22653)
             ) ;
    mux21_ni ix57983 (.Y (nx57982), .A0 (nx57976), .A1 (nx57898), .S0 (nx23179)
             ) ;
    oai21 ix57977 (.Y (nx57976), .A0 (nx22357), .A1 (nx20381), .B0 (nx20391)) ;
    mux21 ix20382 (.Y (nx20381), .A0 (nx57940), .A1 (nx57968), .S0 (nx23059)) ;
    mux21_ni ix57941 (.Y (nx57940), .A0 (nx57924), .A1 (nx57936), .S0 (nx23813)
             ) ;
    mux21_ni ix57925 (.Y (nx57924), .A0 (inputs_196__13), .A1 (inputs_197__13), 
             .S0 (nx24711)) ;
    mux21_ni ix57937 (.Y (nx57936), .A0 (inputs_198__13), .A1 (inputs_199__13), 
             .S0 (nx24711)) ;
    mux21_ni ix57969 (.Y (nx57968), .A0 (nx57952), .A1 (nx57964), .S0 (nx23813)
             ) ;
    mux21_ni ix57953 (.Y (nx57952), .A0 (inputs_212__13), .A1 (inputs_213__13), 
             .S0 (nx24711)) ;
    mux21_ni ix57965 (.Y (nx57964), .A0 (inputs_214__13), .A1 (inputs_215__13), 
             .S0 (nx24711)) ;
    nand04 ix20392 (.Y (nx20391), .A0 (nx22357), .A1 (nx23813), .A2 (nx24711), .A3 (
           nx57912)) ;
    mux21_ni ix57913 (.Y (nx57912), .A0 (inputs_195__13), .A1 (inputs_211__13), 
             .S0 (nx23059)) ;
    mux21_ni ix57899 (.Y (nx57898), .A0 (nx57834), .A1 (nx57894), .S0 (nx23059)
             ) ;
    mux21_ni ix57835 (.Y (nx57834), .A0 (nx57802), .A1 (nx57830), .S0 (nx23317)
             ) ;
    mux21_ni ix57803 (.Y (nx57802), .A0 (nx57786), .A1 (nx57798), .S0 (nx23813)
             ) ;
    mux21_ni ix57787 (.Y (nx57786), .A0 (inputs_200__13), .A1 (inputs_201__13), 
             .S0 (nx24713)) ;
    mux21_ni ix57799 (.Y (nx57798), .A0 (inputs_202__13), .A1 (inputs_203__13), 
             .S0 (nx24713)) ;
    mux21_ni ix57831 (.Y (nx57830), .A0 (nx57814), .A1 (nx57826), .S0 (nx23813)
             ) ;
    mux21_ni ix57815 (.Y (nx57814), .A0 (inputs_204__13), .A1 (inputs_205__13), 
             .S0 (nx24713)) ;
    mux21_ni ix57827 (.Y (nx57826), .A0 (inputs_206__13), .A1 (inputs_207__13), 
             .S0 (nx24713)) ;
    mux21_ni ix57895 (.Y (nx57894), .A0 (nx57862), .A1 (nx57890), .S0 (nx23317)
             ) ;
    mux21_ni ix57863 (.Y (nx57862), .A0 (nx57846), .A1 (nx57858), .S0 (nx23813)
             ) ;
    mux21_ni ix57847 (.Y (nx57846), .A0 (inputs_216__13), .A1 (inputs_217__13), 
             .S0 (nx24713)) ;
    mux21_ni ix57859 (.Y (nx57858), .A0 (inputs_218__13), .A1 (inputs_219__13), 
             .S0 (nx24713)) ;
    mux21_ni ix57891 (.Y (nx57890), .A0 (nx57874), .A1 (nx57886), .S0 (nx23813)
             ) ;
    mux21_ni ix57875 (.Y (nx57874), .A0 (inputs_220__13), .A1 (inputs_221__13), 
             .S0 (nx24713)) ;
    mux21_ni ix57887 (.Y (nx57886), .A0 (inputs_222__13), .A1 (inputs_223__13), 
             .S0 (nx24715)) ;
    mux21_ni ix58191 (.Y (nx58190), .A0 (nx58184), .A1 (nx58106), .S0 (nx23179)
             ) ;
    oai21 ix58185 (.Y (nx58184), .A0 (nx22357), .A1 (nx20421), .B0 (nx20433)) ;
    mux21 ix20422 (.Y (nx20421), .A0 (nx58148), .A1 (nx58176), .S0 (nx23059)) ;
    mux21_ni ix58149 (.Y (nx58148), .A0 (nx58132), .A1 (nx58144), .S0 (nx23815)
             ) ;
    mux21_ni ix58133 (.Y (nx58132), .A0 (inputs_228__13), .A1 (inputs_229__13), 
             .S0 (nx24715)) ;
    mux21_ni ix58145 (.Y (nx58144), .A0 (inputs_230__13), .A1 (inputs_231__13), 
             .S0 (nx24715)) ;
    mux21_ni ix58177 (.Y (nx58176), .A0 (nx58160), .A1 (nx58172), .S0 (nx23815)
             ) ;
    mux21_ni ix58161 (.Y (nx58160), .A0 (inputs_244__13), .A1 (inputs_245__13), 
             .S0 (nx24715)) ;
    mux21_ni ix58173 (.Y (nx58172), .A0 (inputs_246__13), .A1 (inputs_247__13), 
             .S0 (nx24715)) ;
    nand04 ix20434 (.Y (nx20433), .A0 (nx22357), .A1 (nx23815), .A2 (nx24715), .A3 (
           nx58120)) ;
    mux21_ni ix58121 (.Y (nx58120), .A0 (inputs_227__13), .A1 (inputs_243__13), 
             .S0 (nx23059)) ;
    mux21_ni ix58107 (.Y (nx58106), .A0 (nx58042), .A1 (nx58102), .S0 (nx23059)
             ) ;
    mux21_ni ix58043 (.Y (nx58042), .A0 (nx58010), .A1 (nx58038), .S0 (nx23317)
             ) ;
    mux21_ni ix58011 (.Y (nx58010), .A0 (nx57994), .A1 (nx58006), .S0 (nx23815)
             ) ;
    mux21_ni ix57995 (.Y (nx57994), .A0 (inputs_232__13), .A1 (inputs_233__13), 
             .S0 (nx24715)) ;
    mux21_ni ix58007 (.Y (nx58006), .A0 (inputs_234__13), .A1 (inputs_235__13), 
             .S0 (nx24717)) ;
    mux21_ni ix58039 (.Y (nx58038), .A0 (nx58022), .A1 (nx58034), .S0 (nx23815)
             ) ;
    mux21_ni ix58023 (.Y (nx58022), .A0 (inputs_236__13), .A1 (inputs_237__13), 
             .S0 (nx24717)) ;
    mux21_ni ix58035 (.Y (nx58034), .A0 (inputs_238__13), .A1 (inputs_239__13), 
             .S0 (nx24717)) ;
    mux21_ni ix58103 (.Y (nx58102), .A0 (nx58070), .A1 (nx58098), .S0 (nx23317)
             ) ;
    mux21_ni ix58071 (.Y (nx58070), .A0 (nx58054), .A1 (nx58066), .S0 (nx23815)
             ) ;
    mux21_ni ix58055 (.Y (nx58054), .A0 (inputs_248__13), .A1 (inputs_249__13), 
             .S0 (nx24717)) ;
    mux21_ni ix58067 (.Y (nx58066), .A0 (inputs_250__13), .A1 (inputs_251__13), 
             .S0 (nx24717)) ;
    mux21_ni ix58099 (.Y (nx58098), .A0 (nx58082), .A1 (nx58094), .S0 (nx23815)
             ) ;
    mux21_ni ix58083 (.Y (nx58082), .A0 (inputs_252__13), .A1 (inputs_253__13), 
             .S0 (nx24717)) ;
    mux21_ni ix58095 (.Y (nx58094), .A0 (inputs_254__13), .A1 (inputs_255__13), 
             .S0 (nx24717)) ;
    oai21 ix62369 (.Y (\output [14]), .A0 (nx22225), .A1 (nx20461), .B0 (nx20821
          )) ;
    mux21 ix20462 (.Y (nx20461), .A0 (nx59050), .A1 (nx59894), .S0 (nx22443)) ;
    mux21_ni ix59051 (.Y (nx59050), .A0 (nx58626), .A1 (nx59046), .S0 (nx22515)
             ) ;
    mux21_ni ix58627 (.Y (nx58626), .A0 (nx58414), .A1 (nx58622), .S0 (nx22655)
             ) ;
    mux21_ni ix58415 (.Y (nx58414), .A0 (nx58408), .A1 (nx58330), .S0 (nx23181)
             ) ;
    oai21 ix58409 (.Y (nx58408), .A0 (nx22359), .A1 (nx20471), .B0 (nx20483)) ;
    mux21 ix20472 (.Y (nx20471), .A0 (nx58372), .A1 (nx58400), .S0 (nx23061)) ;
    mux21_ni ix58373 (.Y (nx58372), .A0 (nx58356), .A1 (nx58368), .S0 (nx23817)
             ) ;
    mux21_ni ix58357 (.Y (nx58356), .A0 (inputs_260__14), .A1 (inputs_261__14), 
             .S0 (nx24719)) ;
    mux21_ni ix58369 (.Y (nx58368), .A0 (inputs_262__14), .A1 (inputs_263__14), 
             .S0 (nx24719)) ;
    mux21_ni ix58401 (.Y (nx58400), .A0 (nx58384), .A1 (nx58396), .S0 (nx23817)
             ) ;
    mux21_ni ix58385 (.Y (nx58384), .A0 (inputs_276__14), .A1 (inputs_277__14), 
             .S0 (nx24719)) ;
    mux21_ni ix58397 (.Y (nx58396), .A0 (inputs_278__14), .A1 (inputs_279__14), 
             .S0 (nx24719)) ;
    nand04 ix20484 (.Y (nx20483), .A0 (nx22359), .A1 (nx23817), .A2 (nx24719), .A3 (
           nx58344)) ;
    mux21_ni ix58345 (.Y (nx58344), .A0 (inputs_259__14), .A1 (inputs_275__14), 
             .S0 (nx23061)) ;
    mux21_ni ix58331 (.Y (nx58330), .A0 (nx58266), .A1 (nx58326), .S0 (nx23061)
             ) ;
    mux21_ni ix58267 (.Y (nx58266), .A0 (nx58234), .A1 (nx58262), .S0 (nx23319)
             ) ;
    mux21_ni ix58235 (.Y (nx58234), .A0 (nx58218), .A1 (nx58230), .S0 (nx23817)
             ) ;
    mux21_ni ix58219 (.Y (nx58218), .A0 (inputs_264__14), .A1 (inputs_265__14), 
             .S0 (nx24719)) ;
    mux21_ni ix58231 (.Y (nx58230), .A0 (inputs_266__14), .A1 (inputs_267__14), 
             .S0 (nx24719)) ;
    mux21_ni ix58263 (.Y (nx58262), .A0 (nx58246), .A1 (nx58258), .S0 (nx23817)
             ) ;
    mux21_ni ix58247 (.Y (nx58246), .A0 (inputs_268__14), .A1 (inputs_269__14), 
             .S0 (nx24721)) ;
    mux21_ni ix58259 (.Y (nx58258), .A0 (inputs_270__14), .A1 (inputs_271__14), 
             .S0 (nx24721)) ;
    mux21_ni ix58327 (.Y (nx58326), .A0 (nx58294), .A1 (nx58322), .S0 (nx23319)
             ) ;
    mux21_ni ix58295 (.Y (nx58294), .A0 (nx58278), .A1 (nx58290), .S0 (nx23817)
             ) ;
    mux21_ni ix58279 (.Y (nx58278), .A0 (inputs_280__14), .A1 (inputs_281__14), 
             .S0 (nx24721)) ;
    mux21_ni ix58291 (.Y (nx58290), .A0 (inputs_282__14), .A1 (inputs_283__14), 
             .S0 (nx24721)) ;
    mux21_ni ix58323 (.Y (nx58322), .A0 (nx58306), .A1 (nx58318), .S0 (nx23817)
             ) ;
    mux21_ni ix58307 (.Y (nx58306), .A0 (inputs_284__14), .A1 (inputs_285__14), 
             .S0 (nx24721)) ;
    mux21_ni ix58319 (.Y (nx58318), .A0 (inputs_286__14), .A1 (inputs_287__14), 
             .S0 (nx24721)) ;
    mux21_ni ix58623 (.Y (nx58622), .A0 (nx58616), .A1 (nx58538), .S0 (nx23181)
             ) ;
    oai21 ix58617 (.Y (nx58616), .A0 (nx22359), .A1 (nx20513), .B0 (nx20525)) ;
    mux21 ix20514 (.Y (nx20513), .A0 (nx58580), .A1 (nx58608), .S0 (nx23061)) ;
    mux21_ni ix58581 (.Y (nx58580), .A0 (nx58564), .A1 (nx58576), .S0 (nx23819)
             ) ;
    mux21_ni ix58565 (.Y (nx58564), .A0 (inputs_292__14), .A1 (inputs_293__14), 
             .S0 (nx24721)) ;
    mux21_ni ix58577 (.Y (nx58576), .A0 (inputs_294__14), .A1 (inputs_295__14), 
             .S0 (nx24723)) ;
    mux21_ni ix58609 (.Y (nx58608), .A0 (nx58592), .A1 (nx58604), .S0 (nx23819)
             ) ;
    mux21_ni ix58593 (.Y (nx58592), .A0 (inputs_308__14), .A1 (inputs_309__14), 
             .S0 (nx24723)) ;
    mux21_ni ix58605 (.Y (nx58604), .A0 (inputs_310__14), .A1 (inputs_311__14), 
             .S0 (nx24723)) ;
    nand04 ix20526 (.Y (nx20525), .A0 (nx22359), .A1 (nx23819), .A2 (nx24723), .A3 (
           nx58552)) ;
    mux21_ni ix58553 (.Y (nx58552), .A0 (inputs_291__14), .A1 (inputs_307__14), 
             .S0 (nx23061)) ;
    mux21_ni ix58539 (.Y (nx58538), .A0 (nx58474), .A1 (nx58534), .S0 (nx23061)
             ) ;
    mux21_ni ix58475 (.Y (nx58474), .A0 (nx58442), .A1 (nx58470), .S0 (nx23319)
             ) ;
    mux21_ni ix58443 (.Y (nx58442), .A0 (nx58426), .A1 (nx58438), .S0 (nx23819)
             ) ;
    mux21_ni ix58427 (.Y (nx58426), .A0 (inputs_296__14), .A1 (inputs_297__14), 
             .S0 (nx24723)) ;
    mux21_ni ix58439 (.Y (nx58438), .A0 (inputs_298__14), .A1 (inputs_299__14), 
             .S0 (nx24723)) ;
    mux21_ni ix58471 (.Y (nx58470), .A0 (nx58454), .A1 (nx58466), .S0 (nx23819)
             ) ;
    mux21_ni ix58455 (.Y (nx58454), .A0 (inputs_300__14), .A1 (inputs_301__14), 
             .S0 (nx24723)) ;
    mux21_ni ix58467 (.Y (nx58466), .A0 (inputs_302__14), .A1 (inputs_303__14), 
             .S0 (nx24725)) ;
    mux21_ni ix58535 (.Y (nx58534), .A0 (nx58502), .A1 (nx58530), .S0 (nx23319)
             ) ;
    mux21_ni ix58503 (.Y (nx58502), .A0 (nx58486), .A1 (nx58498), .S0 (nx23819)
             ) ;
    mux21_ni ix58487 (.Y (nx58486), .A0 (inputs_312__14), .A1 (inputs_313__14), 
             .S0 (nx24725)) ;
    mux21_ni ix58499 (.Y (nx58498), .A0 (inputs_314__14), .A1 (inputs_315__14), 
             .S0 (nx24725)) ;
    mux21_ni ix58531 (.Y (nx58530), .A0 (nx58514), .A1 (nx58526), .S0 (nx23819)
             ) ;
    mux21_ni ix58515 (.Y (nx58514), .A0 (inputs_316__14), .A1 (inputs_317__14), 
             .S0 (nx24725)) ;
    mux21_ni ix58527 (.Y (nx58526), .A0 (inputs_318__14), .A1 (inputs_319__14), 
             .S0 (nx24725)) ;
    mux21_ni ix59047 (.Y (nx59046), .A0 (nx58834), .A1 (nx59042), .S0 (nx22655)
             ) ;
    mux21_ni ix58835 (.Y (nx58834), .A0 (nx58828), .A1 (nx58750), .S0 (nx23181)
             ) ;
    oai21 ix58829 (.Y (nx58828), .A0 (nx22359), .A1 (nx20559), .B0 (nx20569)) ;
    mux21 ix20560 (.Y (nx20559), .A0 (nx58792), .A1 (nx58820), .S0 (nx23061)) ;
    mux21_ni ix58793 (.Y (nx58792), .A0 (nx58776), .A1 (nx58788), .S0 (nx23821)
             ) ;
    mux21_ni ix58777 (.Y (nx58776), .A0 (inputs_324__14), .A1 (inputs_325__14), 
             .S0 (nx24725)) ;
    mux21_ni ix58789 (.Y (nx58788), .A0 (inputs_326__14), .A1 (inputs_327__14), 
             .S0 (nx24725)) ;
    mux21_ni ix58821 (.Y (nx58820), .A0 (nx58804), .A1 (nx58816), .S0 (nx23821)
             ) ;
    mux21_ni ix58805 (.Y (nx58804), .A0 (inputs_340__14), .A1 (inputs_341__14), 
             .S0 (nx24727)) ;
    mux21_ni ix58817 (.Y (nx58816), .A0 (inputs_342__14), .A1 (inputs_343__14), 
             .S0 (nx24727)) ;
    nand04 ix20570 (.Y (nx20569), .A0 (nx22359), .A1 (nx23821), .A2 (nx24727), .A3 (
           nx58764)) ;
    mux21_ni ix58765 (.Y (nx58764), .A0 (inputs_323__14), .A1 (inputs_339__14), 
             .S0 (nx23063)) ;
    mux21_ni ix58751 (.Y (nx58750), .A0 (nx58686), .A1 (nx58746), .S0 (nx23063)
             ) ;
    mux21_ni ix58687 (.Y (nx58686), .A0 (nx58654), .A1 (nx58682), .S0 (nx23319)
             ) ;
    mux21_ni ix58655 (.Y (nx58654), .A0 (nx58638), .A1 (nx58650), .S0 (nx23821)
             ) ;
    mux21_ni ix58639 (.Y (nx58638), .A0 (inputs_328__14), .A1 (inputs_329__14), 
             .S0 (nx24727)) ;
    mux21_ni ix58651 (.Y (nx58650), .A0 (inputs_330__14), .A1 (inputs_331__14), 
             .S0 (nx24727)) ;
    mux21_ni ix58683 (.Y (nx58682), .A0 (nx58666), .A1 (nx58678), .S0 (nx23821)
             ) ;
    mux21_ni ix58667 (.Y (nx58666), .A0 (inputs_332__14), .A1 (inputs_333__14), 
             .S0 (nx24727)) ;
    mux21_ni ix58679 (.Y (nx58678), .A0 (inputs_334__14), .A1 (inputs_335__14), 
             .S0 (nx24727)) ;
    mux21_ni ix58747 (.Y (nx58746), .A0 (nx58714), .A1 (nx58742), .S0 (nx23319)
             ) ;
    mux21_ni ix58715 (.Y (nx58714), .A0 (nx58698), .A1 (nx58710), .S0 (nx23821)
             ) ;
    mux21_ni ix58699 (.Y (nx58698), .A0 (inputs_344__14), .A1 (inputs_345__14), 
             .S0 (nx24729)) ;
    mux21_ni ix58711 (.Y (nx58710), .A0 (inputs_346__14), .A1 (inputs_347__14), 
             .S0 (nx24729)) ;
    mux21_ni ix58743 (.Y (nx58742), .A0 (nx58726), .A1 (nx58738), .S0 (nx23821)
             ) ;
    mux21_ni ix58727 (.Y (nx58726), .A0 (inputs_348__14), .A1 (inputs_349__14), 
             .S0 (nx24729)) ;
    mux21_ni ix58739 (.Y (nx58738), .A0 (inputs_350__14), .A1 (inputs_351__14), 
             .S0 (nx24729)) ;
    mux21_ni ix59043 (.Y (nx59042), .A0 (nx59036), .A1 (nx58958), .S0 (nx23181)
             ) ;
    oai21 ix59037 (.Y (nx59036), .A0 (nx22359), .A1 (nx20599), .B0 (nx20609)) ;
    mux21 ix20600 (.Y (nx20599), .A0 (nx59000), .A1 (nx59028), .S0 (nx23063)) ;
    mux21_ni ix59001 (.Y (nx59000), .A0 (nx58984), .A1 (nx58996), .S0 (nx23823)
             ) ;
    mux21_ni ix58985 (.Y (nx58984), .A0 (inputs_356__14), .A1 (inputs_357__14), 
             .S0 (nx24729)) ;
    mux21_ni ix58997 (.Y (nx58996), .A0 (inputs_358__14), .A1 (inputs_359__14), 
             .S0 (nx24729)) ;
    mux21_ni ix59029 (.Y (nx59028), .A0 (nx59012), .A1 (nx59024), .S0 (nx23823)
             ) ;
    mux21_ni ix59013 (.Y (nx59012), .A0 (inputs_372__14), .A1 (inputs_373__14), 
             .S0 (nx24729)) ;
    mux21_ni ix59025 (.Y (nx59024), .A0 (inputs_374__14), .A1 (inputs_375__14), 
             .S0 (nx24731)) ;
    nand04 ix20610 (.Y (nx20609), .A0 (nx22361), .A1 (nx23823), .A2 (nx24731), .A3 (
           nx58972)) ;
    mux21_ni ix58973 (.Y (nx58972), .A0 (inputs_355__14), .A1 (inputs_371__14), 
             .S0 (nx23063)) ;
    mux21_ni ix58959 (.Y (nx58958), .A0 (nx58894), .A1 (nx58954), .S0 (nx23063)
             ) ;
    mux21_ni ix58895 (.Y (nx58894), .A0 (nx58862), .A1 (nx58890), .S0 (nx23319)
             ) ;
    mux21_ni ix58863 (.Y (nx58862), .A0 (nx58846), .A1 (nx58858), .S0 (nx23823)
             ) ;
    mux21_ni ix58847 (.Y (nx58846), .A0 (inputs_360__14), .A1 (inputs_361__14), 
             .S0 (nx24731)) ;
    mux21_ni ix58859 (.Y (nx58858), .A0 (inputs_362__14), .A1 (inputs_363__14), 
             .S0 (nx24731)) ;
    mux21_ni ix58891 (.Y (nx58890), .A0 (nx58874), .A1 (nx58886), .S0 (nx23823)
             ) ;
    mux21_ni ix58875 (.Y (nx58874), .A0 (inputs_364__14), .A1 (inputs_365__14), 
             .S0 (nx24731)) ;
    mux21_ni ix58887 (.Y (nx58886), .A0 (inputs_366__14), .A1 (inputs_367__14), 
             .S0 (nx24731)) ;
    mux21_ni ix58955 (.Y (nx58954), .A0 (nx58922), .A1 (nx58950), .S0 (nx23321)
             ) ;
    mux21_ni ix58923 (.Y (nx58922), .A0 (nx58906), .A1 (nx58918), .S0 (nx23823)
             ) ;
    mux21_ni ix58907 (.Y (nx58906), .A0 (inputs_376__14), .A1 (inputs_377__14), 
             .S0 (nx24731)) ;
    mux21_ni ix58919 (.Y (nx58918), .A0 (inputs_378__14), .A1 (inputs_379__14), 
             .S0 (nx24733)) ;
    mux21_ni ix58951 (.Y (nx58950), .A0 (nx58934), .A1 (nx58946), .S0 (nx23823)
             ) ;
    mux21_ni ix58935 (.Y (nx58934), .A0 (inputs_380__14), .A1 (inputs_381__14), 
             .S0 (nx24733)) ;
    mux21_ni ix58947 (.Y (nx58946), .A0 (inputs_382__14), .A1 (inputs_383__14), 
             .S0 (nx24733)) ;
    mux21_ni ix59895 (.Y (nx59894), .A0 (nx59470), .A1 (nx59890), .S0 (nx22515)
             ) ;
    mux21_ni ix59471 (.Y (nx59470), .A0 (nx59258), .A1 (nx59466), .S0 (nx22655)
             ) ;
    mux21_ni ix59259 (.Y (nx59258), .A0 (nx59252), .A1 (nx59174), .S0 (nx23181)
             ) ;
    oai21 ix59253 (.Y (nx59252), .A0 (nx22361), .A1 (nx20643), .B0 (nx20655)) ;
    mux21 ix20644 (.Y (nx20643), .A0 (nx59216), .A1 (nx59244), .S0 (nx23063)) ;
    mux21_ni ix59217 (.Y (nx59216), .A0 (nx59200), .A1 (nx59212), .S0 (nx23825)
             ) ;
    mux21_ni ix59201 (.Y (nx59200), .A0 (inputs_388__14), .A1 (inputs_389__14), 
             .S0 (nx24733)) ;
    mux21_ni ix59213 (.Y (nx59212), .A0 (inputs_390__14), .A1 (inputs_391__14), 
             .S0 (nx24733)) ;
    mux21_ni ix59245 (.Y (nx59244), .A0 (nx59228), .A1 (nx59240), .S0 (nx23825)
             ) ;
    mux21_ni ix59229 (.Y (nx59228), .A0 (inputs_404__14), .A1 (inputs_405__14), 
             .S0 (nx24733)) ;
    mux21_ni ix59241 (.Y (nx59240), .A0 (inputs_406__14), .A1 (inputs_407__14), 
             .S0 (nx24733)) ;
    nand04 ix20656 (.Y (nx20655), .A0 (nx22361), .A1 (nx23825), .A2 (nx24735), .A3 (
           nx59188)) ;
    mux21_ni ix59189 (.Y (nx59188), .A0 (inputs_387__14), .A1 (inputs_403__14), 
             .S0 (nx23063)) ;
    mux21_ni ix59175 (.Y (nx59174), .A0 (nx59110), .A1 (nx59170), .S0 (nx23065)
             ) ;
    mux21_ni ix59111 (.Y (nx59110), .A0 (nx59078), .A1 (nx59106), .S0 (nx23321)
             ) ;
    mux21_ni ix59079 (.Y (nx59078), .A0 (nx59062), .A1 (nx59074), .S0 (nx23825)
             ) ;
    mux21_ni ix59063 (.Y (nx59062), .A0 (inputs_392__14), .A1 (inputs_393__14), 
             .S0 (nx24735)) ;
    mux21_ni ix59075 (.Y (nx59074), .A0 (inputs_394__14), .A1 (inputs_395__14), 
             .S0 (nx24735)) ;
    mux21_ni ix59107 (.Y (nx59106), .A0 (nx59090), .A1 (nx59102), .S0 (nx23825)
             ) ;
    mux21_ni ix59091 (.Y (nx59090), .A0 (inputs_396__14), .A1 (inputs_397__14), 
             .S0 (nx24735)) ;
    mux21_ni ix59103 (.Y (nx59102), .A0 (inputs_398__14), .A1 (inputs_399__14), 
             .S0 (nx24735)) ;
    mux21_ni ix59171 (.Y (nx59170), .A0 (nx59138), .A1 (nx59166), .S0 (nx23321)
             ) ;
    mux21_ni ix59139 (.Y (nx59138), .A0 (nx59122), .A1 (nx59134), .S0 (nx23825)
             ) ;
    mux21_ni ix59123 (.Y (nx59122), .A0 (inputs_408__14), .A1 (inputs_409__14), 
             .S0 (nx24735)) ;
    mux21_ni ix59135 (.Y (nx59134), .A0 (inputs_410__14), .A1 (inputs_411__14), 
             .S0 (nx24735)) ;
    mux21_ni ix59167 (.Y (nx59166), .A0 (nx59150), .A1 (nx59162), .S0 (nx23825)
             ) ;
    mux21_ni ix59151 (.Y (nx59150), .A0 (inputs_412__14), .A1 (inputs_413__14), 
             .S0 (nx24737)) ;
    mux21_ni ix59163 (.Y (nx59162), .A0 (inputs_414__14), .A1 (inputs_415__14), 
             .S0 (nx24737)) ;
    mux21_ni ix59467 (.Y (nx59466), .A0 (nx59460), .A1 (nx59382), .S0 (nx23181)
             ) ;
    oai21 ix59461 (.Y (nx59460), .A0 (nx22361), .A1 (nx20689), .B0 (nx20701)) ;
    mux21 ix20690 (.Y (nx20689), .A0 (nx59424), .A1 (nx59452), .S0 (nx23065)) ;
    mux21_ni ix59425 (.Y (nx59424), .A0 (nx59408), .A1 (nx59420), .S0 (nx23827)
             ) ;
    mux21_ni ix59409 (.Y (nx59408), .A0 (inputs_420__14), .A1 (inputs_421__14), 
             .S0 (nx24737)) ;
    mux21_ni ix59421 (.Y (nx59420), .A0 (inputs_422__14), .A1 (inputs_423__14), 
             .S0 (nx24737)) ;
    mux21_ni ix59453 (.Y (nx59452), .A0 (nx59436), .A1 (nx59448), .S0 (nx23827)
             ) ;
    mux21_ni ix59437 (.Y (nx59436), .A0 (inputs_436__14), .A1 (inputs_437__14), 
             .S0 (nx24737)) ;
    mux21_ni ix59449 (.Y (nx59448), .A0 (inputs_438__14), .A1 (inputs_439__14), 
             .S0 (nx24737)) ;
    nand04 ix20702 (.Y (nx20701), .A0 (nx22361), .A1 (nx23827), .A2 (nx24737), .A3 (
           nx59396)) ;
    mux21_ni ix59397 (.Y (nx59396), .A0 (inputs_419__14), .A1 (inputs_435__14), 
             .S0 (nx23065)) ;
    mux21_ni ix59383 (.Y (nx59382), .A0 (nx59318), .A1 (nx59378), .S0 (nx23065)
             ) ;
    mux21_ni ix59319 (.Y (nx59318), .A0 (nx59286), .A1 (nx59314), .S0 (nx23321)
             ) ;
    mux21_ni ix59287 (.Y (nx59286), .A0 (nx59270), .A1 (nx59282), .S0 (nx23827)
             ) ;
    mux21_ni ix59271 (.Y (nx59270), .A0 (inputs_424__14), .A1 (inputs_425__14), 
             .S0 (nx24739)) ;
    mux21_ni ix59283 (.Y (nx59282), .A0 (inputs_426__14), .A1 (inputs_427__14), 
             .S0 (nx24739)) ;
    mux21_ni ix59315 (.Y (nx59314), .A0 (nx59298), .A1 (nx59310), .S0 (nx23827)
             ) ;
    mux21_ni ix59299 (.Y (nx59298), .A0 (inputs_428__14), .A1 (inputs_429__14), 
             .S0 (nx24739)) ;
    mux21_ni ix59311 (.Y (nx59310), .A0 (inputs_430__14), .A1 (inputs_431__14), 
             .S0 (nx24739)) ;
    mux21_ni ix59379 (.Y (nx59378), .A0 (nx59346), .A1 (nx59374), .S0 (nx23321)
             ) ;
    mux21_ni ix59347 (.Y (nx59346), .A0 (nx59330), .A1 (nx59342), .S0 (nx23827)
             ) ;
    mux21_ni ix59331 (.Y (nx59330), .A0 (inputs_440__14), .A1 (inputs_441__14), 
             .S0 (nx24739)) ;
    mux21_ni ix59343 (.Y (nx59342), .A0 (inputs_442__14), .A1 (inputs_443__14), 
             .S0 (nx24739)) ;
    mux21_ni ix59375 (.Y (nx59374), .A0 (nx59358), .A1 (nx59370), .S0 (nx23827)
             ) ;
    mux21_ni ix59359 (.Y (nx59358), .A0 (inputs_444__14), .A1 (inputs_445__14), 
             .S0 (nx24739)) ;
    mux21_ni ix59371 (.Y (nx59370), .A0 (inputs_446__14), .A1 (inputs_447__14), 
             .S0 (nx24741)) ;
    mux21_ni ix59891 (.Y (nx59890), .A0 (nx59678), .A1 (nx59886), .S0 (nx22655)
             ) ;
    mux21_ni ix59679 (.Y (nx59678), .A0 (nx59672), .A1 (nx59594), .S0 (nx23181)
             ) ;
    oai21 ix59673 (.Y (nx59672), .A0 (nx22361), .A1 (nx20733), .B0 (nx20745)) ;
    mux21 ix20734 (.Y (nx20733), .A0 (nx59636), .A1 (nx59664), .S0 (nx23065)) ;
    mux21_ni ix59637 (.Y (nx59636), .A0 (nx59620), .A1 (nx59632), .S0 (nx23829)
             ) ;
    mux21_ni ix59621 (.Y (nx59620), .A0 (inputs_452__14), .A1 (inputs_453__14), 
             .S0 (nx24741)) ;
    mux21_ni ix59633 (.Y (nx59632), .A0 (inputs_454__14), .A1 (inputs_455__14), 
             .S0 (nx24741)) ;
    mux21_ni ix59665 (.Y (nx59664), .A0 (nx59648), .A1 (nx59660), .S0 (nx23829)
             ) ;
    mux21_ni ix59649 (.Y (nx59648), .A0 (inputs_468__14), .A1 (inputs_469__14), 
             .S0 (nx24741)) ;
    mux21_ni ix59661 (.Y (nx59660), .A0 (inputs_470__14), .A1 (inputs_471__14), 
             .S0 (nx24741)) ;
    nand04 ix20746 (.Y (nx20745), .A0 (nx22361), .A1 (nx23829), .A2 (nx24741), .A3 (
           nx59608)) ;
    mux21_ni ix59609 (.Y (nx59608), .A0 (inputs_451__14), .A1 (inputs_467__14), 
             .S0 (nx23065)) ;
    mux21_ni ix59595 (.Y (nx59594), .A0 (nx59530), .A1 (nx59590), .S0 (nx23065)
             ) ;
    mux21_ni ix59531 (.Y (nx59530), .A0 (nx59498), .A1 (nx59526), .S0 (nx23321)
             ) ;
    mux21_ni ix59499 (.Y (nx59498), .A0 (nx59482), .A1 (nx59494), .S0 (nx23829)
             ) ;
    mux21_ni ix59483 (.Y (nx59482), .A0 (inputs_456__14), .A1 (inputs_457__14), 
             .S0 (nx24741)) ;
    mux21_ni ix59495 (.Y (nx59494), .A0 (inputs_458__14), .A1 (inputs_459__14), 
             .S0 (nx24743)) ;
    mux21_ni ix59527 (.Y (nx59526), .A0 (nx59510), .A1 (nx59522), .S0 (nx23829)
             ) ;
    mux21_ni ix59511 (.Y (nx59510), .A0 (inputs_460__14), .A1 (inputs_461__14), 
             .S0 (nx24743)) ;
    mux21_ni ix59523 (.Y (nx59522), .A0 (inputs_462__14), .A1 (inputs_463__14), 
             .S0 (nx24743)) ;
    mux21_ni ix59591 (.Y (nx59590), .A0 (nx59558), .A1 (nx59586), .S0 (nx23321)
             ) ;
    mux21_ni ix59559 (.Y (nx59558), .A0 (nx59542), .A1 (nx59554), .S0 (nx23829)
             ) ;
    mux21_ni ix59543 (.Y (nx59542), .A0 (inputs_472__14), .A1 (inputs_473__14), 
             .S0 (nx24743)) ;
    mux21_ni ix59555 (.Y (nx59554), .A0 (inputs_474__14), .A1 (inputs_475__14), 
             .S0 (nx24743)) ;
    mux21_ni ix59587 (.Y (nx59586), .A0 (nx59570), .A1 (nx59582), .S0 (nx23829)
             ) ;
    mux21_ni ix59571 (.Y (nx59570), .A0 (inputs_476__14), .A1 (inputs_477__14), 
             .S0 (nx24743)) ;
    mux21_ni ix59583 (.Y (nx59582), .A0 (inputs_478__14), .A1 (inputs_479__14), 
             .S0 (nx24743)) ;
    mux21_ni ix59887 (.Y (nx59886), .A0 (nx59880), .A1 (nx59802), .S0 (nx23183)
             ) ;
    oai21 ix59881 (.Y (nx59880), .A0 (nx22363), .A1 (nx20781), .B0 (nx20793)) ;
    mux21 ix20782 (.Y (nx20781), .A0 (nx59844), .A1 (nx59872), .S0 (nx23067)) ;
    mux21_ni ix59845 (.Y (nx59844), .A0 (nx59828), .A1 (nx59840), .S0 (nx23831)
             ) ;
    mux21_ni ix59829 (.Y (nx59828), .A0 (inputs_484__14), .A1 (inputs_485__14), 
             .S0 (nx24745)) ;
    mux21_ni ix59841 (.Y (nx59840), .A0 (inputs_486__14), .A1 (inputs_487__14), 
             .S0 (nx24745)) ;
    mux21_ni ix59873 (.Y (nx59872), .A0 (nx59856), .A1 (nx59868), .S0 (nx23831)
             ) ;
    mux21_ni ix59857 (.Y (nx59856), .A0 (inputs_500__14), .A1 (inputs_501__14), 
             .S0 (nx24745)) ;
    mux21_ni ix59869 (.Y (nx59868), .A0 (inputs_502__14), .A1 (inputs_503__14), 
             .S0 (nx24745)) ;
    nand04 ix20794 (.Y (nx20793), .A0 (nx22363), .A1 (nx23831), .A2 (nx24745), .A3 (
           nx59816)) ;
    mux21_ni ix59817 (.Y (nx59816), .A0 (inputs_483__14), .A1 (inputs_499__14), 
             .S0 (nx23067)) ;
    mux21_ni ix59803 (.Y (nx59802), .A0 (nx59738), .A1 (nx59798), .S0 (nx23067)
             ) ;
    mux21_ni ix59739 (.Y (nx59738), .A0 (nx59706), .A1 (nx59734), .S0 (nx23323)
             ) ;
    mux21_ni ix59707 (.Y (nx59706), .A0 (nx59690), .A1 (nx59702), .S0 (nx23831)
             ) ;
    mux21_ni ix59691 (.Y (nx59690), .A0 (inputs_488__14), .A1 (inputs_489__14), 
             .S0 (nx24745)) ;
    mux21_ni ix59703 (.Y (nx59702), .A0 (inputs_490__14), .A1 (inputs_491__14), 
             .S0 (nx24745)) ;
    mux21_ni ix59735 (.Y (nx59734), .A0 (nx59718), .A1 (nx59730), .S0 (nx23831)
             ) ;
    mux21_ni ix59719 (.Y (nx59718), .A0 (inputs_492__14), .A1 (inputs_493__14), 
             .S0 (nx24747)) ;
    mux21_ni ix59731 (.Y (nx59730), .A0 (inputs_494__14), .A1 (inputs_495__14), 
             .S0 (nx24747)) ;
    mux21_ni ix59799 (.Y (nx59798), .A0 (nx59766), .A1 (nx59794), .S0 (nx23323)
             ) ;
    mux21_ni ix59767 (.Y (nx59766), .A0 (nx59750), .A1 (nx59762), .S0 (nx23831)
             ) ;
    mux21_ni ix59751 (.Y (nx59750), .A0 (inputs_504__14), .A1 (inputs_505__14), 
             .S0 (nx24747)) ;
    mux21_ni ix59763 (.Y (nx59762), .A0 (inputs_506__14), .A1 (inputs_507__14), 
             .S0 (nx24747)) ;
    mux21_ni ix59795 (.Y (nx59794), .A0 (nx59778), .A1 (nx59790), .S0 (nx23831)
             ) ;
    mux21_ni ix59779 (.Y (nx59778), .A0 (inputs_508__14), .A1 (inputs_509__14), 
             .S0 (nx24747)) ;
    mux21_ni ix59791 (.Y (nx59790), .A0 (inputs_510__14), .A1 (inputs_511__14), 
             .S0 (nx24747)) ;
    aoi32 ix20822 (.Y (nx20821), .A0 (nx60664), .A1 (nx24839), .A2 (nx22363), .B0 (
          nx22225), .B1 (nx62360)) ;
    oai21 ix60665 (.Y (nx60664), .A0 (nx23833), .A1 (nx20825), .B0 (nx20927)) ;
    mux21 ix20826 (.Y (nx20825), .A0 (nx60402), .A1 (nx60654), .S0 (nx24747)) ;
    mux21_ni ix60403 (.Y (nx60402), .A0 (nx60274), .A1 (nx60398), .S0 (nx22405)
             ) ;
    mux21_ni ix60275 (.Y (nx60274), .A0 (nx60210), .A1 (nx60270), .S0 (nx22443)
             ) ;
    mux21_ni ix60211 (.Y (nx60210), .A0 (nx60178), .A1 (nx60206), .S0 (nx22515)
             ) ;
    mux21_ni ix60179 (.Y (nx60178), .A0 (nx60162), .A1 (nx60174), .S0 (nx22655)
             ) ;
    mux21_ni ix60163 (.Y (nx60162), .A0 (inputs_0__14), .A1 (inputs_16__14), .S0 (
             nx23067)) ;
    mux21_ni ix60175 (.Y (nx60174), .A0 (inputs_32__14), .A1 (inputs_48__14), .S0 (
             nx23067)) ;
    mux21_ni ix60207 (.Y (nx60206), .A0 (nx60190), .A1 (nx60202), .S0 (nx22655)
             ) ;
    mux21_ni ix60191 (.Y (nx60190), .A0 (inputs_64__14), .A1 (inputs_80__14), .S0 (
             nx23067)) ;
    mux21_ni ix60203 (.Y (nx60202), .A0 (inputs_96__14), .A1 (inputs_112__14), .S0 (
             nx23067)) ;
    mux21_ni ix60271 (.Y (nx60270), .A0 (nx60238), .A1 (nx60266), .S0 (nx22515)
             ) ;
    mux21_ni ix60239 (.Y (nx60238), .A0 (nx60222), .A1 (nx60234), .S0 (nx22655)
             ) ;
    mux21_ni ix60223 (.Y (nx60222), .A0 (inputs_128__14), .A1 (inputs_144__14), 
             .S0 (nx23069)) ;
    mux21_ni ix60235 (.Y (nx60234), .A0 (inputs_160__14), .A1 (inputs_176__14), 
             .S0 (nx23069)) ;
    mux21_ni ix60267 (.Y (nx60266), .A0 (nx60250), .A1 (nx60262), .S0 (nx22657)
             ) ;
    mux21_ni ix60251 (.Y (nx60250), .A0 (inputs_192__14), .A1 (inputs_208__14), 
             .S0 (nx23069)) ;
    mux21_ni ix60263 (.Y (nx60262), .A0 (inputs_224__14), .A1 (inputs_240__14), 
             .S0 (nx23069)) ;
    mux21_ni ix60399 (.Y (nx60398), .A0 (nx60334), .A1 (nx60394), .S0 (nx22443)
             ) ;
    mux21_ni ix60335 (.Y (nx60334), .A0 (nx60302), .A1 (nx60330), .S0 (nx22515)
             ) ;
    mux21_ni ix60303 (.Y (nx60302), .A0 (nx60286), .A1 (nx60298), .S0 (nx22657)
             ) ;
    mux21_ni ix60287 (.Y (nx60286), .A0 (inputs_256__14), .A1 (inputs_272__14), 
             .S0 (nx23069)) ;
    mux21_ni ix60299 (.Y (nx60298), .A0 (inputs_288__14), .A1 (inputs_304__14), 
             .S0 (nx23069)) ;
    mux21_ni ix60331 (.Y (nx60330), .A0 (nx60314), .A1 (nx60326), .S0 (nx22657)
             ) ;
    mux21_ni ix60315 (.Y (nx60314), .A0 (inputs_320__14), .A1 (inputs_336__14), 
             .S0 (nx23069)) ;
    mux21_ni ix60327 (.Y (nx60326), .A0 (inputs_352__14), .A1 (inputs_368__14), 
             .S0 (nx23071)) ;
    mux21_ni ix60395 (.Y (nx60394), .A0 (nx60362), .A1 (nx60390), .S0 (nx22515)
             ) ;
    mux21_ni ix60363 (.Y (nx60362), .A0 (nx60346), .A1 (nx60358), .S0 (nx22657)
             ) ;
    mux21_ni ix60347 (.Y (nx60346), .A0 (inputs_384__14), .A1 (inputs_400__14), 
             .S0 (nx23071)) ;
    mux21_ni ix60359 (.Y (nx60358), .A0 (inputs_416__14), .A1 (inputs_432__14), 
             .S0 (nx23071)) ;
    mux21_ni ix60391 (.Y (nx60390), .A0 (nx60374), .A1 (nx60386), .S0 (nx22657)
             ) ;
    mux21_ni ix60375 (.Y (nx60374), .A0 (inputs_448__14), .A1 (inputs_464__14), 
             .S0 (nx23071)) ;
    mux21_ni ix60387 (.Y (nx60386), .A0 (inputs_480__14), .A1 (inputs_496__14), 
             .S0 (nx23071)) ;
    mux21_ni ix60655 (.Y (nx60654), .A0 (nx60526), .A1 (nx60650), .S0 (nx22405)
             ) ;
    mux21_ni ix60527 (.Y (nx60526), .A0 (nx60462), .A1 (nx60522), .S0 (nx22443)
             ) ;
    mux21_ni ix60463 (.Y (nx60462), .A0 (nx60430), .A1 (nx60458), .S0 (nx22515)
             ) ;
    mux21_ni ix60431 (.Y (nx60430), .A0 (nx60414), .A1 (nx60426), .S0 (nx22657)
             ) ;
    mux21_ni ix60415 (.Y (nx60414), .A0 (inputs_1__14), .A1 (inputs_17__14), .S0 (
             nx23071)) ;
    mux21_ni ix60427 (.Y (nx60426), .A0 (inputs_33__14), .A1 (inputs_49__14), .S0 (
             nx23071)) ;
    mux21_ni ix60459 (.Y (nx60458), .A0 (nx60442), .A1 (nx60454), .S0 (nx22657)
             ) ;
    mux21_ni ix60443 (.Y (nx60442), .A0 (inputs_65__14), .A1 (inputs_81__14), .S0 (
             nx23073)) ;
    mux21_ni ix60455 (.Y (nx60454), .A0 (inputs_97__14), .A1 (inputs_113__14), .S0 (
             nx23073)) ;
    mux21_ni ix60523 (.Y (nx60522), .A0 (nx60490), .A1 (nx60518), .S0 (nx22517)
             ) ;
    mux21_ni ix60491 (.Y (nx60490), .A0 (nx60474), .A1 (nx60486), .S0 (nx22659)
             ) ;
    mux21_ni ix60475 (.Y (nx60474), .A0 (inputs_129__14), .A1 (inputs_145__14), 
             .S0 (nx23073)) ;
    mux21_ni ix60487 (.Y (nx60486), .A0 (inputs_161__14), .A1 (inputs_177__14), 
             .S0 (nx23073)) ;
    mux21_ni ix60519 (.Y (nx60518), .A0 (nx60502), .A1 (nx60514), .S0 (nx22659)
             ) ;
    mux21_ni ix60503 (.Y (nx60502), .A0 (inputs_193__14), .A1 (inputs_209__14), 
             .S0 (nx23073)) ;
    mux21_ni ix60515 (.Y (nx60514), .A0 (inputs_225__14), .A1 (inputs_241__14), 
             .S0 (nx23073)) ;
    mux21_ni ix60651 (.Y (nx60650), .A0 (nx60586), .A1 (nx60646), .S0 (nx22443)
             ) ;
    mux21_ni ix60587 (.Y (nx60586), .A0 (nx60554), .A1 (nx60582), .S0 (nx22517)
             ) ;
    mux21_ni ix60555 (.Y (nx60554), .A0 (nx60538), .A1 (nx60550), .S0 (nx22659)
             ) ;
    mux21_ni ix60539 (.Y (nx60538), .A0 (inputs_257__14), .A1 (inputs_273__14), 
             .S0 (nx23073)) ;
    mux21_ni ix60551 (.Y (nx60550), .A0 (inputs_289__14), .A1 (inputs_305__14), 
             .S0 (nx23075)) ;
    mux21_ni ix60583 (.Y (nx60582), .A0 (nx60566), .A1 (nx60578), .S0 (nx22659)
             ) ;
    mux21_ni ix60567 (.Y (nx60566), .A0 (inputs_321__14), .A1 (inputs_337__14), 
             .S0 (nx23075)) ;
    mux21_ni ix60579 (.Y (nx60578), .A0 (inputs_353__14), .A1 (inputs_369__14), 
             .S0 (nx23075)) ;
    mux21_ni ix60647 (.Y (nx60646), .A0 (nx60614), .A1 (nx60642), .S0 (nx22517)
             ) ;
    mux21_ni ix60615 (.Y (nx60614), .A0 (nx60598), .A1 (nx60610), .S0 (nx22659)
             ) ;
    mux21_ni ix60599 (.Y (nx60598), .A0 (inputs_385__14), .A1 (inputs_401__14), 
             .S0 (nx23075)) ;
    mux21_ni ix60611 (.Y (nx60610), .A0 (inputs_417__14), .A1 (inputs_433__14), 
             .S0 (nx23075)) ;
    mux21_ni ix60643 (.Y (nx60642), .A0 (nx60626), .A1 (nx60638), .S0 (nx22659)
             ) ;
    mux21_ni ix60627 (.Y (nx60626), .A0 (inputs_449__14), .A1 (inputs_465__14), 
             .S0 (nx23075)) ;
    mux21_ni ix60639 (.Y (nx60638), .A0 (inputs_481__14), .A1 (inputs_497__14), 
             .S0 (nx23075)) ;
    nand03 ix20928 (.Y (nx20927), .A0 (nx60148), .A1 (nx23833), .A2 (nx22383)) ;
    mux21_ni ix60149 (.Y (nx60148), .A0 (nx60020), .A1 (nx60144), .S0 (nx22405)
             ) ;
    mux21_ni ix60021 (.Y (nx60020), .A0 (nx59956), .A1 (nx60016), .S0 (nx22443)
             ) ;
    mux21_ni ix59957 (.Y (nx59956), .A0 (nx59924), .A1 (nx59952), .S0 (nx22517)
             ) ;
    mux21_ni ix59925 (.Y (nx59924), .A0 (nx59908), .A1 (nx59920), .S0 (nx22659)
             ) ;
    mux21_ni ix59909 (.Y (nx59908), .A0 (inputs_2__14), .A1 (inputs_18__14), .S0 (
             nx23077)) ;
    mux21_ni ix59921 (.Y (nx59920), .A0 (inputs_34__14), .A1 (inputs_50__14), .S0 (
             nx23077)) ;
    mux21_ni ix59953 (.Y (nx59952), .A0 (nx59936), .A1 (nx59948), .S0 (nx22661)
             ) ;
    mux21_ni ix59937 (.Y (nx59936), .A0 (inputs_66__14), .A1 (inputs_82__14), .S0 (
             nx23077)) ;
    mux21_ni ix59949 (.Y (nx59948), .A0 (inputs_98__14), .A1 (inputs_114__14), .S0 (
             nx23077)) ;
    mux21_ni ix60017 (.Y (nx60016), .A0 (nx59984), .A1 (nx60012), .S0 (nx22517)
             ) ;
    mux21_ni ix59985 (.Y (nx59984), .A0 (nx59968), .A1 (nx59980), .S0 (nx22661)
             ) ;
    mux21_ni ix59969 (.Y (nx59968), .A0 (inputs_130__14), .A1 (inputs_146__14), 
             .S0 (nx23077)) ;
    mux21_ni ix59981 (.Y (nx59980), .A0 (inputs_162__14), .A1 (inputs_178__14), 
             .S0 (nx23077)) ;
    mux21_ni ix60013 (.Y (nx60012), .A0 (nx59996), .A1 (nx60008), .S0 (nx22661)
             ) ;
    mux21_ni ix59997 (.Y (nx59996), .A0 (inputs_194__14), .A1 (inputs_210__14), 
             .S0 (nx23077)) ;
    mux21_ni ix60009 (.Y (nx60008), .A0 (inputs_226__14), .A1 (inputs_242__14), 
             .S0 (nx23079)) ;
    mux21_ni ix60145 (.Y (nx60144), .A0 (nx60080), .A1 (nx60140), .S0 (nx22443)
             ) ;
    mux21_ni ix60081 (.Y (nx60080), .A0 (nx60048), .A1 (nx60076), .S0 (nx22517)
             ) ;
    mux21_ni ix60049 (.Y (nx60048), .A0 (nx60032), .A1 (nx60044), .S0 (nx22661)
             ) ;
    mux21_ni ix60033 (.Y (nx60032), .A0 (inputs_258__14), .A1 (inputs_274__14), 
             .S0 (nx23079)) ;
    mux21_ni ix60045 (.Y (nx60044), .A0 (inputs_290__14), .A1 (inputs_306__14), 
             .S0 (nx23079)) ;
    mux21_ni ix60077 (.Y (nx60076), .A0 (nx60060), .A1 (nx60072), .S0 (nx22661)
             ) ;
    mux21_ni ix60061 (.Y (nx60060), .A0 (inputs_322__14), .A1 (inputs_338__14), 
             .S0 (nx23079)) ;
    mux21_ni ix60073 (.Y (nx60072), .A0 (inputs_354__14), .A1 (inputs_370__14), 
             .S0 (nx23079)) ;
    mux21_ni ix60141 (.Y (nx60140), .A0 (nx60108), .A1 (nx60136), .S0 (nx22517)
             ) ;
    mux21_ni ix60109 (.Y (nx60108), .A0 (nx60092), .A1 (nx60104), .S0 (nx22661)
             ) ;
    mux21_ni ix60093 (.Y (nx60092), .A0 (inputs_386__14), .A1 (inputs_402__14), 
             .S0 (nx23079)) ;
    mux21_ni ix60105 (.Y (nx60104), .A0 (inputs_418__14), .A1 (inputs_434__14), 
             .S0 (nx23079)) ;
    mux21_ni ix60137 (.Y (nx60136), .A0 (nx60120), .A1 (nx60132), .S0 (nx22661)
             ) ;
    mux21_ni ix60121 (.Y (nx60120), .A0 (inputs_450__14), .A1 (inputs_466__14), 
             .S0 (nx23081)) ;
    mux21_ni ix60133 (.Y (nx60132), .A0 (inputs_482__14), .A1 (inputs_498__14), 
             .S0 (nx23081)) ;
    mux21_ni ix62361 (.Y (nx62360), .A0 (nx61512), .A1 (nx62356), .S0 (nx22445)
             ) ;
    mux21_ni ix61513 (.Y (nx61512), .A0 (nx61088), .A1 (nx61508), .S0 (nx22519)
             ) ;
    mux21_ni ix61089 (.Y (nx61088), .A0 (nx60876), .A1 (nx61084), .S0 (nx22663)
             ) ;
    mux21_ni ix60877 (.Y (nx60876), .A0 (nx60870), .A1 (nx60792), .S0 (nx23183)
             ) ;
    oai21 ix60871 (.Y (nx60870), .A0 (nx22363), .A1 (nx20987), .B0 (nx20997)) ;
    mux21 ix20988 (.Y (nx20987), .A0 (nx60834), .A1 (nx60862), .S0 (nx23081)) ;
    mux21_ni ix60835 (.Y (nx60834), .A0 (nx60818), .A1 (nx60830), .S0 (nx23833)
             ) ;
    mux21_ni ix60819 (.Y (nx60818), .A0 (inputs_4__14), .A1 (inputs_5__14), .S0 (
             nx24749)) ;
    mux21_ni ix60831 (.Y (nx60830), .A0 (inputs_6__14), .A1 (inputs_7__14), .S0 (
             nx24749)) ;
    mux21_ni ix60863 (.Y (nx60862), .A0 (nx60846), .A1 (nx60858), .S0 (nx23833)
             ) ;
    mux21_ni ix60847 (.Y (nx60846), .A0 (inputs_20__14), .A1 (inputs_21__14), .S0 (
             nx24749)) ;
    mux21_ni ix60859 (.Y (nx60858), .A0 (inputs_22__14), .A1 (inputs_23__14), .S0 (
             nx24749)) ;
    nand04 ix20998 (.Y (nx20997), .A0 (nx22363), .A1 (nx23833), .A2 (nx24749), .A3 (
           nx60806)) ;
    mux21_ni ix60807 (.Y (nx60806), .A0 (inputs_3__14), .A1 (inputs_19__14), .S0 (
             nx23081)) ;
    mux21_ni ix60793 (.Y (nx60792), .A0 (nx60728), .A1 (nx60788), .S0 (nx23081)
             ) ;
    mux21_ni ix60729 (.Y (nx60728), .A0 (nx60696), .A1 (nx60724), .S0 (nx23323)
             ) ;
    mux21_ni ix60697 (.Y (nx60696), .A0 (nx60680), .A1 (nx60692), .S0 (nx23833)
             ) ;
    mux21_ni ix60681 (.Y (nx60680), .A0 (inputs_8__14), .A1 (inputs_9__14), .S0 (
             nx24749)) ;
    mux21_ni ix60693 (.Y (nx60692), .A0 (inputs_10__14), .A1 (inputs_11__14), .S0 (
             nx24749)) ;
    mux21_ni ix60725 (.Y (nx60724), .A0 (nx60708), .A1 (nx60720), .S0 (nx23833)
             ) ;
    mux21_ni ix60709 (.Y (nx60708), .A0 (inputs_12__14), .A1 (inputs_13__14), .S0 (
             nx24751)) ;
    mux21_ni ix60721 (.Y (nx60720), .A0 (inputs_14__14), .A1 (inputs_15__14), .S0 (
             nx24751)) ;
    mux21_ni ix60789 (.Y (nx60788), .A0 (nx60756), .A1 (nx60784), .S0 (nx23323)
             ) ;
    mux21_ni ix60757 (.Y (nx60756), .A0 (nx60740), .A1 (nx60752), .S0 (nx23835)
             ) ;
    mux21_ni ix60741 (.Y (nx60740), .A0 (inputs_24__14), .A1 (inputs_25__14), .S0 (
             nx24751)) ;
    mux21_ni ix60753 (.Y (nx60752), .A0 (inputs_26__14), .A1 (inputs_27__14), .S0 (
             nx24751)) ;
    mux21_ni ix60785 (.Y (nx60784), .A0 (nx60768), .A1 (nx60780), .S0 (nx23835)
             ) ;
    mux21_ni ix60769 (.Y (nx60768), .A0 (inputs_28__14), .A1 (inputs_29__14), .S0 (
             nx24751)) ;
    mux21_ni ix60781 (.Y (nx60780), .A0 (inputs_30__14), .A1 (inputs_31__14), .S0 (
             nx24751)) ;
    mux21_ni ix61085 (.Y (nx61084), .A0 (nx61078), .A1 (nx61000), .S0 (nx23183)
             ) ;
    oai21 ix61079 (.Y (nx61078), .A0 (nx22363), .A1 (nx21027), .B0 (nx21039)) ;
    mux21 ix21028 (.Y (nx21027), .A0 (nx61042), .A1 (nx61070), .S0 (nx23081)) ;
    mux21_ni ix61043 (.Y (nx61042), .A0 (nx61026), .A1 (nx61038), .S0 (nx23835)
             ) ;
    mux21_ni ix61027 (.Y (nx61026), .A0 (inputs_36__14), .A1 (inputs_37__14), .S0 (
             nx24751)) ;
    mux21_ni ix61039 (.Y (nx61038), .A0 (inputs_38__14), .A1 (inputs_39__14), .S0 (
             nx24753)) ;
    mux21_ni ix61071 (.Y (nx61070), .A0 (nx61054), .A1 (nx61066), .S0 (nx23835)
             ) ;
    mux21_ni ix61055 (.Y (nx61054), .A0 (inputs_52__14), .A1 (inputs_53__14), .S0 (
             nx24753)) ;
    mux21_ni ix61067 (.Y (nx61066), .A0 (inputs_54__14), .A1 (inputs_55__14), .S0 (
             nx24753)) ;
    nand04 ix21040 (.Y (nx21039), .A0 (nx22363), .A1 (nx23835), .A2 (nx24753), .A3 (
           nx61014)) ;
    mux21_ni ix61015 (.Y (nx61014), .A0 (inputs_35__14), .A1 (inputs_51__14), .S0 (
             nx23081)) ;
    mux21_ni ix61001 (.Y (nx61000), .A0 (nx60936), .A1 (nx60996), .S0 (nx23083)
             ) ;
    mux21_ni ix60937 (.Y (nx60936), .A0 (nx60904), .A1 (nx60932), .S0 (nx23323)
             ) ;
    mux21_ni ix60905 (.Y (nx60904), .A0 (nx60888), .A1 (nx60900), .S0 (nx23835)
             ) ;
    mux21_ni ix60889 (.Y (nx60888), .A0 (inputs_40__14), .A1 (inputs_41__14), .S0 (
             nx24753)) ;
    mux21_ni ix60901 (.Y (nx60900), .A0 (inputs_42__14), .A1 (inputs_43__14), .S0 (
             nx24753)) ;
    mux21_ni ix60933 (.Y (nx60932), .A0 (nx60916), .A1 (nx60928), .S0 (nx23835)
             ) ;
    mux21_ni ix60917 (.Y (nx60916), .A0 (inputs_44__14), .A1 (inputs_45__14), .S0 (
             nx24753)) ;
    mux21_ni ix60929 (.Y (nx60928), .A0 (inputs_46__14), .A1 (inputs_47__14), .S0 (
             nx24755)) ;
    mux21_ni ix60997 (.Y (nx60996), .A0 (nx60964), .A1 (nx60992), .S0 (nx23323)
             ) ;
    mux21_ni ix60965 (.Y (nx60964), .A0 (nx60948), .A1 (nx60960), .S0 (nx23837)
             ) ;
    mux21_ni ix60949 (.Y (nx60948), .A0 (inputs_56__14), .A1 (inputs_57__14), .S0 (
             nx24755)) ;
    mux21_ni ix60961 (.Y (nx60960), .A0 (inputs_58__14), .A1 (inputs_59__14), .S0 (
             nx24755)) ;
    mux21_ni ix60993 (.Y (nx60992), .A0 (nx60976), .A1 (nx60988), .S0 (nx23837)
             ) ;
    mux21_ni ix60977 (.Y (nx60976), .A0 (inputs_60__14), .A1 (inputs_61__14), .S0 (
             nx24755)) ;
    mux21_ni ix60989 (.Y (nx60988), .A0 (inputs_62__14), .A1 (inputs_63__14), .S0 (
             nx24755)) ;
    mux21_ni ix61509 (.Y (nx61508), .A0 (nx61296), .A1 (nx61504), .S0 (nx22663)
             ) ;
    mux21_ni ix61297 (.Y (nx61296), .A0 (nx61290), .A1 (nx61212), .S0 (nx23183)
             ) ;
    oai21 ix61291 (.Y (nx61290), .A0 (nx22365), .A1 (nx21073), .B0 (nx21085)) ;
    mux21 ix21074 (.Y (nx21073), .A0 (nx61254), .A1 (nx61282), .S0 (nx23083)) ;
    mux21_ni ix61255 (.Y (nx61254), .A0 (nx61238), .A1 (nx61250), .S0 (nx23837)
             ) ;
    mux21_ni ix61239 (.Y (nx61238), .A0 (inputs_68__14), .A1 (inputs_69__14), .S0 (
             nx24755)) ;
    mux21_ni ix61251 (.Y (nx61250), .A0 (inputs_70__14), .A1 (inputs_71__14), .S0 (
             nx24755)) ;
    mux21_ni ix61283 (.Y (nx61282), .A0 (nx61266), .A1 (nx61278), .S0 (nx23837)
             ) ;
    mux21_ni ix61267 (.Y (nx61266), .A0 (inputs_84__14), .A1 (inputs_85__14), .S0 (
             nx24757)) ;
    mux21_ni ix61279 (.Y (nx61278), .A0 (inputs_86__14), .A1 (inputs_87__14), .S0 (
             nx24757)) ;
    nand04 ix21086 (.Y (nx21085), .A0 (nx22365), .A1 (nx23837), .A2 (nx24757), .A3 (
           nx61226)) ;
    mux21_ni ix61227 (.Y (nx61226), .A0 (inputs_67__14), .A1 (inputs_83__14), .S0 (
             nx23083)) ;
    mux21_ni ix61213 (.Y (nx61212), .A0 (nx61148), .A1 (nx61208), .S0 (nx23083)
             ) ;
    mux21_ni ix61149 (.Y (nx61148), .A0 (nx61116), .A1 (nx61144), .S0 (nx23323)
             ) ;
    mux21_ni ix61117 (.Y (nx61116), .A0 (nx61100), .A1 (nx61112), .S0 (nx23837)
             ) ;
    mux21_ni ix61101 (.Y (nx61100), .A0 (inputs_72__14), .A1 (inputs_73__14), .S0 (
             nx24757)) ;
    mux21_ni ix61113 (.Y (nx61112), .A0 (inputs_74__14), .A1 (inputs_75__14), .S0 (
             nx24757)) ;
    mux21_ni ix61145 (.Y (nx61144), .A0 (nx61128), .A1 (nx61140), .S0 (nx23837)
             ) ;
    mux21_ni ix61129 (.Y (nx61128), .A0 (inputs_76__14), .A1 (inputs_77__14), .S0 (
             nx24757)) ;
    mux21_ni ix61141 (.Y (nx61140), .A0 (inputs_78__14), .A1 (inputs_79__14), .S0 (
             nx24757)) ;
    mux21_ni ix61209 (.Y (nx61208), .A0 (nx61176), .A1 (nx61204), .S0 (nx23325)
             ) ;
    mux21_ni ix61177 (.Y (nx61176), .A0 (nx61160), .A1 (nx61172), .S0 (nx23839)
             ) ;
    mux21_ni ix61161 (.Y (nx61160), .A0 (inputs_88__14), .A1 (inputs_89__14), .S0 (
             nx24759)) ;
    mux21_ni ix61173 (.Y (nx61172), .A0 (inputs_90__14), .A1 (inputs_91__14), .S0 (
             nx24759)) ;
    mux21_ni ix61205 (.Y (nx61204), .A0 (nx61188), .A1 (nx61200), .S0 (nx23839)
             ) ;
    mux21_ni ix61189 (.Y (nx61188), .A0 (inputs_92__14), .A1 (inputs_93__14), .S0 (
             nx24759)) ;
    mux21_ni ix61201 (.Y (nx61200), .A0 (inputs_94__14), .A1 (inputs_95__14), .S0 (
             nx24759)) ;
    mux21_ni ix61505 (.Y (nx61504), .A0 (nx61498), .A1 (nx61420), .S0 (nx23183)
             ) ;
    oai21 ix61499 (.Y (nx61498), .A0 (nx22365), .A1 (nx21117), .B0 (nx21127)) ;
    mux21 ix21118 (.Y (nx21117), .A0 (nx61462), .A1 (nx61490), .S0 (nx23083)) ;
    mux21_ni ix61463 (.Y (nx61462), .A0 (nx61446), .A1 (nx61458), .S0 (nx23839)
             ) ;
    mux21_ni ix61447 (.Y (nx61446), .A0 (inputs_100__14), .A1 (inputs_101__14), 
             .S0 (nx24759)) ;
    mux21_ni ix61459 (.Y (nx61458), .A0 (inputs_102__14), .A1 (inputs_103__14), 
             .S0 (nx24759)) ;
    mux21_ni ix61491 (.Y (nx61490), .A0 (nx61474), .A1 (nx61486), .S0 (nx23839)
             ) ;
    mux21_ni ix61475 (.Y (nx61474), .A0 (inputs_116__14), .A1 (inputs_117__14), 
             .S0 (nx24759)) ;
    mux21_ni ix61487 (.Y (nx61486), .A0 (inputs_118__14), .A1 (inputs_119__14), 
             .S0 (nx24761)) ;
    nand04 ix21128 (.Y (nx21127), .A0 (nx22365), .A1 (nx23839), .A2 (nx24761), .A3 (
           nx61434)) ;
    mux21_ni ix61435 (.Y (nx61434), .A0 (inputs_99__14), .A1 (inputs_115__14), .S0 (
             nx23083)) ;
    mux21_ni ix61421 (.Y (nx61420), .A0 (nx61356), .A1 (nx61416), .S0 (nx23083)
             ) ;
    mux21_ni ix61357 (.Y (nx61356), .A0 (nx61324), .A1 (nx61352), .S0 (nx23325)
             ) ;
    mux21_ni ix61325 (.Y (nx61324), .A0 (nx61308), .A1 (nx61320), .S0 (nx23839)
             ) ;
    mux21_ni ix61309 (.Y (nx61308), .A0 (inputs_104__14), .A1 (inputs_105__14), 
             .S0 (nx24761)) ;
    mux21_ni ix61321 (.Y (nx61320), .A0 (inputs_106__14), .A1 (inputs_107__14), 
             .S0 (nx24761)) ;
    mux21_ni ix61353 (.Y (nx61352), .A0 (nx61336), .A1 (nx61348), .S0 (nx23839)
             ) ;
    mux21_ni ix61337 (.Y (nx61336), .A0 (inputs_108__14), .A1 (inputs_109__14), 
             .S0 (nx24761)) ;
    mux21_ni ix61349 (.Y (nx61348), .A0 (inputs_110__14), .A1 (inputs_111__14), 
             .S0 (nx24761)) ;
    mux21_ni ix61417 (.Y (nx61416), .A0 (nx61384), .A1 (nx61412), .S0 (nx23325)
             ) ;
    mux21_ni ix61385 (.Y (nx61384), .A0 (nx61368), .A1 (nx61380), .S0 (nx23841)
             ) ;
    mux21_ni ix61369 (.Y (nx61368), .A0 (inputs_120__14), .A1 (inputs_121__14), 
             .S0 (nx24761)) ;
    mux21_ni ix61381 (.Y (nx61380), .A0 (inputs_122__14), .A1 (inputs_123__14), 
             .S0 (nx24763)) ;
    mux21_ni ix61413 (.Y (nx61412), .A0 (nx61396), .A1 (nx61408), .S0 (nx23841)
             ) ;
    mux21_ni ix61397 (.Y (nx61396), .A0 (inputs_124__14), .A1 (inputs_125__14), 
             .S0 (nx24763)) ;
    mux21_ni ix61409 (.Y (nx61408), .A0 (inputs_126__14), .A1 (inputs_127__14), 
             .S0 (nx24763)) ;
    mux21_ni ix62357 (.Y (nx62356), .A0 (nx61932), .A1 (nx62352), .S0 (nx22519)
             ) ;
    mux21_ni ix61933 (.Y (nx61932), .A0 (nx61720), .A1 (nx61928), .S0 (nx22663)
             ) ;
    mux21_ni ix61721 (.Y (nx61720), .A0 (nx61714), .A1 (nx61636), .S0 (nx23183)
             ) ;
    oai21 ix61715 (.Y (nx61714), .A0 (nx22365), .A1 (nx21163), .B0 (nx21175)) ;
    mux21 ix21164 (.Y (nx21163), .A0 (nx61678), .A1 (nx61706), .S0 (nx23085)) ;
    mux21_ni ix61679 (.Y (nx61678), .A0 (nx61662), .A1 (nx61674), .S0 (nx23841)
             ) ;
    mux21_ni ix61663 (.Y (nx61662), .A0 (inputs_132__14), .A1 (inputs_133__14), 
             .S0 (nx24763)) ;
    mux21_ni ix61675 (.Y (nx61674), .A0 (inputs_134__14), .A1 (inputs_135__14), 
             .S0 (nx24763)) ;
    mux21_ni ix61707 (.Y (nx61706), .A0 (nx61690), .A1 (nx61702), .S0 (nx23841)
             ) ;
    mux21_ni ix61691 (.Y (nx61690), .A0 (inputs_148__14), .A1 (inputs_149__14), 
             .S0 (nx24763)) ;
    mux21_ni ix61703 (.Y (nx61702), .A0 (inputs_150__14), .A1 (inputs_151__14), 
             .S0 (nx24763)) ;
    nand04 ix21176 (.Y (nx21175), .A0 (nx22365), .A1 (nx23841), .A2 (nx24765), .A3 (
           nx61650)) ;
    mux21_ni ix61651 (.Y (nx61650), .A0 (inputs_131__14), .A1 (inputs_147__14), 
             .S0 (nx23085)) ;
    mux21_ni ix61637 (.Y (nx61636), .A0 (nx61572), .A1 (nx61632), .S0 (nx23085)
             ) ;
    mux21_ni ix61573 (.Y (nx61572), .A0 (nx61540), .A1 (nx61568), .S0 (nx23325)
             ) ;
    mux21_ni ix61541 (.Y (nx61540), .A0 (nx61524), .A1 (nx61536), .S0 (nx23841)
             ) ;
    mux21_ni ix61525 (.Y (nx61524), .A0 (inputs_136__14), .A1 (inputs_137__14), 
             .S0 (nx24765)) ;
    mux21_ni ix61537 (.Y (nx61536), .A0 (inputs_138__14), .A1 (inputs_139__14), 
             .S0 (nx24765)) ;
    mux21_ni ix61569 (.Y (nx61568), .A0 (nx61552), .A1 (nx61564), .S0 (nx23841)
             ) ;
    mux21_ni ix61553 (.Y (nx61552), .A0 (inputs_140__14), .A1 (inputs_141__14), 
             .S0 (nx24765)) ;
    mux21_ni ix61565 (.Y (nx61564), .A0 (inputs_142__14), .A1 (inputs_143__14), 
             .S0 (nx24765)) ;
    mux21_ni ix61633 (.Y (nx61632), .A0 (nx61600), .A1 (nx61628), .S0 (nx23325)
             ) ;
    mux21_ni ix61601 (.Y (nx61600), .A0 (nx61584), .A1 (nx61596), .S0 (nx23843)
             ) ;
    mux21_ni ix61585 (.Y (nx61584), .A0 (inputs_152__14), .A1 (inputs_153__14), 
             .S0 (nx24765)) ;
    mux21_ni ix61597 (.Y (nx61596), .A0 (inputs_154__14), .A1 (inputs_155__14), 
             .S0 (nx24765)) ;
    mux21_ni ix61629 (.Y (nx61628), .A0 (nx61612), .A1 (nx61624), .S0 (nx23843)
             ) ;
    mux21_ni ix61613 (.Y (nx61612), .A0 (inputs_156__14), .A1 (inputs_157__14), 
             .S0 (nx24767)) ;
    mux21_ni ix61625 (.Y (nx61624), .A0 (inputs_158__14), .A1 (inputs_159__14), 
             .S0 (nx24767)) ;
    mux21_ni ix61929 (.Y (nx61928), .A0 (nx61922), .A1 (nx61844), .S0 (nx23183)
             ) ;
    oai21 ix61923 (.Y (nx61922), .A0 (nx22365), .A1 (nx21209), .B0 (nx21221)) ;
    mux21 ix21210 (.Y (nx21209), .A0 (nx61886), .A1 (nx61914), .S0 (nx23085)) ;
    mux21_ni ix61887 (.Y (nx61886), .A0 (nx61870), .A1 (nx61882), .S0 (nx23843)
             ) ;
    mux21_ni ix61871 (.Y (nx61870), .A0 (inputs_164__14), .A1 (inputs_165__14), 
             .S0 (nx24767)) ;
    mux21_ni ix61883 (.Y (nx61882), .A0 (inputs_166__14), .A1 (inputs_167__14), 
             .S0 (nx24767)) ;
    mux21_ni ix61915 (.Y (nx61914), .A0 (nx61898), .A1 (nx61910), .S0 (nx23843)
             ) ;
    mux21_ni ix61899 (.Y (nx61898), .A0 (inputs_180__14), .A1 (inputs_181__14), 
             .S0 (nx24767)) ;
    mux21_ni ix61911 (.Y (nx61910), .A0 (inputs_182__14), .A1 (inputs_183__14), 
             .S0 (nx24767)) ;
    nand04 ix21222 (.Y (nx21221), .A0 (nx22367), .A1 (nx23843), .A2 (nx24767), .A3 (
           nx61858)) ;
    mux21_ni ix61859 (.Y (nx61858), .A0 (inputs_163__14), .A1 (inputs_179__14), 
             .S0 (nx23085)) ;
    mux21_ni ix61845 (.Y (nx61844), .A0 (nx61780), .A1 (nx61840), .S0 (nx23085)
             ) ;
    mux21_ni ix61781 (.Y (nx61780), .A0 (nx61748), .A1 (nx61776), .S0 (nx23325)
             ) ;
    mux21_ni ix61749 (.Y (nx61748), .A0 (nx61732), .A1 (nx61744), .S0 (nx23843)
             ) ;
    mux21_ni ix61733 (.Y (nx61732), .A0 (inputs_168__14), .A1 (inputs_169__14), 
             .S0 (nx24769)) ;
    mux21_ni ix61745 (.Y (nx61744), .A0 (inputs_170__14), .A1 (inputs_171__14), 
             .S0 (nx24769)) ;
    mux21_ni ix61777 (.Y (nx61776), .A0 (nx61760), .A1 (nx61772), .S0 (nx23843)
             ) ;
    mux21_ni ix61761 (.Y (nx61760), .A0 (inputs_172__14), .A1 (inputs_173__14), 
             .S0 (nx24769)) ;
    mux21_ni ix61773 (.Y (nx61772), .A0 (inputs_174__14), .A1 (inputs_175__14), 
             .S0 (nx24769)) ;
    mux21_ni ix61841 (.Y (nx61840), .A0 (nx61808), .A1 (nx61836), .S0 (nx23325)
             ) ;
    mux21_ni ix61809 (.Y (nx61808), .A0 (nx61792), .A1 (nx61804), .S0 (nx23845)
             ) ;
    mux21_ni ix61793 (.Y (nx61792), .A0 (inputs_184__14), .A1 (inputs_185__14), 
             .S0 (nx24769)) ;
    mux21_ni ix61805 (.Y (nx61804), .A0 (inputs_186__14), .A1 (inputs_187__14), 
             .S0 (nx24769)) ;
    mux21_ni ix61837 (.Y (nx61836), .A0 (nx61820), .A1 (nx61832), .S0 (nx23845)
             ) ;
    mux21_ni ix61821 (.Y (nx61820), .A0 (inputs_188__14), .A1 (inputs_189__14), 
             .S0 (nx24769)) ;
    mux21_ni ix61833 (.Y (nx61832), .A0 (inputs_190__14), .A1 (inputs_191__14), 
             .S0 (nx24771)) ;
    mux21_ni ix62353 (.Y (nx62352), .A0 (nx62140), .A1 (nx62348), .S0 (nx22663)
             ) ;
    mux21_ni ix62141 (.Y (nx62140), .A0 (nx62134), .A1 (nx62056), .S0 (nx23185)
             ) ;
    oai21 ix62135 (.Y (nx62134), .A0 (nx22367), .A1 (nx21253), .B0 (nx21267)) ;
    mux21 ix21254 (.Y (nx21253), .A0 (nx62098), .A1 (nx62126), .S0 (nx23085)) ;
    mux21_ni ix62099 (.Y (nx62098), .A0 (nx62082), .A1 (nx62094), .S0 (nx23845)
             ) ;
    mux21_ni ix62083 (.Y (nx62082), .A0 (inputs_196__14), .A1 (inputs_197__14), 
             .S0 (nx24771)) ;
    mux21_ni ix62095 (.Y (nx62094), .A0 (inputs_198__14), .A1 (inputs_199__14), 
             .S0 (nx24771)) ;
    mux21_ni ix62127 (.Y (nx62126), .A0 (nx62110), .A1 (nx62122), .S0 (nx23845)
             ) ;
    mux21_ni ix62111 (.Y (nx62110), .A0 (inputs_212__14), .A1 (inputs_213__14), 
             .S0 (nx24771)) ;
    mux21_ni ix62123 (.Y (nx62122), .A0 (inputs_214__14), .A1 (inputs_215__14), 
             .S0 (nx24771)) ;
    nand04 ix21268 (.Y (nx21267), .A0 (nx22367), .A1 (nx23845), .A2 (nx24771), .A3 (
           nx62070)) ;
    mux21_ni ix62071 (.Y (nx62070), .A0 (inputs_195__14), .A1 (inputs_211__14), 
             .S0 (nx23087)) ;
    mux21_ni ix62057 (.Y (nx62056), .A0 (nx61992), .A1 (nx62052), .S0 (nx23087)
             ) ;
    mux21_ni ix61993 (.Y (nx61992), .A0 (nx61960), .A1 (nx61988), .S0 (nx23327)
             ) ;
    mux21_ni ix61961 (.Y (nx61960), .A0 (nx61944), .A1 (nx61956), .S0 (nx23845)
             ) ;
    mux21_ni ix61945 (.Y (nx61944), .A0 (inputs_200__14), .A1 (inputs_201__14), 
             .S0 (nx24771)) ;
    mux21_ni ix61957 (.Y (nx61956), .A0 (inputs_202__14), .A1 (inputs_203__14), 
             .S0 (nx24773)) ;
    mux21_ni ix61989 (.Y (nx61988), .A0 (nx61972), .A1 (nx61984), .S0 (nx23845)
             ) ;
    mux21_ni ix61973 (.Y (nx61972), .A0 (inputs_204__14), .A1 (inputs_205__14), 
             .S0 (nx24773)) ;
    mux21_ni ix61985 (.Y (nx61984), .A0 (inputs_206__14), .A1 (inputs_207__14), 
             .S0 (nx24773)) ;
    mux21_ni ix62053 (.Y (nx62052), .A0 (nx62020), .A1 (nx62048), .S0 (nx23327)
             ) ;
    mux21_ni ix62021 (.Y (nx62020), .A0 (nx62004), .A1 (nx62016), .S0 (nx23847)
             ) ;
    mux21_ni ix62005 (.Y (nx62004), .A0 (inputs_216__14), .A1 (inputs_217__14), 
             .S0 (nx24773)) ;
    mux21_ni ix62017 (.Y (nx62016), .A0 (inputs_218__14), .A1 (inputs_219__14), 
             .S0 (nx24773)) ;
    mux21_ni ix62049 (.Y (nx62048), .A0 (nx62032), .A1 (nx62044), .S0 (nx23847)
             ) ;
    mux21_ni ix62033 (.Y (nx62032), .A0 (inputs_220__14), .A1 (inputs_221__14), 
             .S0 (nx24773)) ;
    mux21_ni ix62045 (.Y (nx62044), .A0 (inputs_222__14), .A1 (inputs_223__14), 
             .S0 (nx24773)) ;
    mux21_ni ix62349 (.Y (nx62348), .A0 (nx62342), .A1 (nx62264), .S0 (nx23185)
             ) ;
    oai21 ix62343 (.Y (nx62342), .A0 (nx22367), .A1 (nx21297), .B0 (nx21309)) ;
    mux21 ix21298 (.Y (nx21297), .A0 (nx62306), .A1 (nx62334), .S0 (nx23087)) ;
    mux21_ni ix62307 (.Y (nx62306), .A0 (nx62290), .A1 (nx62302), .S0 (nx23847)
             ) ;
    mux21_ni ix62291 (.Y (nx62290), .A0 (inputs_228__14), .A1 (inputs_229__14), 
             .S0 (nx24775)) ;
    mux21_ni ix62303 (.Y (nx62302), .A0 (inputs_230__14), .A1 (inputs_231__14), 
             .S0 (nx24775)) ;
    mux21_ni ix62335 (.Y (nx62334), .A0 (nx62318), .A1 (nx62330), .S0 (nx23847)
             ) ;
    mux21_ni ix62319 (.Y (nx62318), .A0 (inputs_244__14), .A1 (inputs_245__14), 
             .S0 (nx24775)) ;
    mux21_ni ix62331 (.Y (nx62330), .A0 (inputs_246__14), .A1 (inputs_247__14), 
             .S0 (nx24775)) ;
    nand04 ix21310 (.Y (nx21309), .A0 (nx22367), .A1 (nx23847), .A2 (nx24775), .A3 (
           nx62278)) ;
    mux21_ni ix62279 (.Y (nx62278), .A0 (inputs_227__14), .A1 (inputs_243__14), 
             .S0 (nx23087)) ;
    mux21_ni ix62265 (.Y (nx62264), .A0 (nx62200), .A1 (nx62260), .S0 (nx23087)
             ) ;
    mux21_ni ix62201 (.Y (nx62200), .A0 (nx62168), .A1 (nx62196), .S0 (nx23327)
             ) ;
    mux21_ni ix62169 (.Y (nx62168), .A0 (nx62152), .A1 (nx62164), .S0 (nx23847)
             ) ;
    mux21_ni ix62153 (.Y (nx62152), .A0 (inputs_232__14), .A1 (inputs_233__14), 
             .S0 (nx24775)) ;
    mux21_ni ix62165 (.Y (nx62164), .A0 (inputs_234__14), .A1 (inputs_235__14), 
             .S0 (nx24775)) ;
    mux21_ni ix62197 (.Y (nx62196), .A0 (nx62180), .A1 (nx62192), .S0 (nx23847)
             ) ;
    mux21_ni ix62181 (.Y (nx62180), .A0 (inputs_236__14), .A1 (inputs_237__14), 
             .S0 (nx24777)) ;
    mux21_ni ix62193 (.Y (nx62192), .A0 (inputs_238__14), .A1 (inputs_239__14), 
             .S0 (nx24777)) ;
    mux21_ni ix62261 (.Y (nx62260), .A0 (nx62228), .A1 (nx62256), .S0 (nx23327)
             ) ;
    mux21_ni ix62229 (.Y (nx62228), .A0 (nx62212), .A1 (nx62224), .S0 (nx23849)
             ) ;
    mux21_ni ix62213 (.Y (nx62212), .A0 (inputs_248__14), .A1 (inputs_249__14), 
             .S0 (nx24777)) ;
    mux21_ni ix62225 (.Y (nx62224), .A0 (inputs_250__14), .A1 (inputs_251__14), 
             .S0 (nx24777)) ;
    mux21_ni ix62257 (.Y (nx62256), .A0 (nx62240), .A1 (nx62252), .S0 (nx23849)
             ) ;
    mux21_ni ix62241 (.Y (nx62240), .A0 (inputs_252__14), .A1 (inputs_253__14), 
             .S0 (nx24777)) ;
    mux21_ni ix62253 (.Y (nx62252), .A0 (inputs_254__14), .A1 (inputs_255__14), 
             .S0 (nx24777)) ;
    oai21 ix66527 (.Y (\output [15]), .A0 (nx22225), .A1 (nx21339), .B0 (nx21701
          )) ;
    mux21 ix21340 (.Y (nx21339), .A0 (nx63208), .A1 (nx64052), .S0 (nx22445)) ;
    mux21_ni ix63209 (.Y (nx63208), .A0 (nx62784), .A1 (nx63204), .S0 (nx22519)
             ) ;
    mux21_ni ix62785 (.Y (nx62784), .A0 (nx62572), .A1 (nx62780), .S0 (nx22663)
             ) ;
    mux21_ni ix62573 (.Y (nx62572), .A0 (nx62566), .A1 (nx62488), .S0 (nx23185)
             ) ;
    oai21 ix62567 (.Y (nx62566), .A0 (nx22367), .A1 (nx21349), .B0 (nx21361)) ;
    mux21 ix21350 (.Y (nx21349), .A0 (nx62530), .A1 (nx62558), .S0 (nx23087)) ;
    mux21_ni ix62531 (.Y (nx62530), .A0 (nx62514), .A1 (nx62526), .S0 (nx23849)
             ) ;
    mux21_ni ix62515 (.Y (nx62514), .A0 (inputs_260__15), .A1 (inputs_261__15), 
             .S0 (nx24777)) ;
    mux21_ni ix62527 (.Y (nx62526), .A0 (inputs_262__15), .A1 (inputs_263__15), 
             .S0 (nx24779)) ;
    mux21_ni ix62559 (.Y (nx62558), .A0 (nx62542), .A1 (nx62554), .S0 (nx23849)
             ) ;
    mux21_ni ix62543 (.Y (nx62542), .A0 (inputs_276__15), .A1 (inputs_277__15), 
             .S0 (nx24779)) ;
    mux21_ni ix62555 (.Y (nx62554), .A0 (inputs_278__15), .A1 (inputs_279__15), 
             .S0 (nx24779)) ;
    nand04 ix21362 (.Y (nx21361), .A0 (nx22367), .A1 (nx23849), .A2 (nx24779), .A3 (
           nx62502)) ;
    mux21_ni ix62503 (.Y (nx62502), .A0 (inputs_259__15), .A1 (inputs_275__15), 
             .S0 (nx23087)) ;
    mux21_ni ix62489 (.Y (nx62488), .A0 (nx62424), .A1 (nx62484), .S0 (nx23089)
             ) ;
    mux21_ni ix62425 (.Y (nx62424), .A0 (nx62392), .A1 (nx62420), .S0 (nx23327)
             ) ;
    mux21_ni ix62393 (.Y (nx62392), .A0 (nx62376), .A1 (nx62388), .S0 (nx23849)
             ) ;
    mux21_ni ix62377 (.Y (nx62376), .A0 (inputs_264__15), .A1 (inputs_265__15), 
             .S0 (nx24779)) ;
    mux21_ni ix62389 (.Y (nx62388), .A0 (inputs_266__15), .A1 (inputs_267__15), 
             .S0 (nx24779)) ;
    mux21_ni ix62421 (.Y (nx62420), .A0 (nx62404), .A1 (nx62416), .S0 (nx23849)
             ) ;
    mux21_ni ix62405 (.Y (nx62404), .A0 (inputs_268__15), .A1 (inputs_269__15), 
             .S0 (nx24779)) ;
    mux21_ni ix62417 (.Y (nx62416), .A0 (inputs_270__15), .A1 (inputs_271__15), 
             .S0 (nx24781)) ;
    mux21_ni ix62485 (.Y (nx62484), .A0 (nx62452), .A1 (nx62480), .S0 (nx23327)
             ) ;
    mux21_ni ix62453 (.Y (nx62452), .A0 (nx62436), .A1 (nx62448), .S0 (nx23851)
             ) ;
    mux21_ni ix62437 (.Y (nx62436), .A0 (inputs_280__15), .A1 (inputs_281__15), 
             .S0 (nx24781)) ;
    mux21_ni ix62449 (.Y (nx62448), .A0 (inputs_282__15), .A1 (inputs_283__15), 
             .S0 (nx24781)) ;
    mux21_ni ix62481 (.Y (nx62480), .A0 (nx62464), .A1 (nx62476), .S0 (nx23851)
             ) ;
    mux21_ni ix62465 (.Y (nx62464), .A0 (inputs_284__15), .A1 (inputs_285__15), 
             .S0 (nx24781)) ;
    mux21_ni ix62477 (.Y (nx62476), .A0 (inputs_286__15), .A1 (inputs_287__15), 
             .S0 (nx24781)) ;
    mux21_ni ix62781 (.Y (nx62780), .A0 (nx62774), .A1 (nx62696), .S0 (nx23185)
             ) ;
    oai21 ix62775 (.Y (nx62774), .A0 (nx22369), .A1 (nx21391), .B0 (nx21405)) ;
    mux21 ix21392 (.Y (nx21391), .A0 (nx62738), .A1 (nx62766), .S0 (nx23089)) ;
    mux21_ni ix62739 (.Y (nx62738), .A0 (nx62722), .A1 (nx62734), .S0 (nx23851)
             ) ;
    mux21_ni ix62723 (.Y (nx62722), .A0 (inputs_292__15), .A1 (inputs_293__15), 
             .S0 (nx24781)) ;
    mux21_ni ix62735 (.Y (nx62734), .A0 (inputs_294__15), .A1 (inputs_295__15), 
             .S0 (nx24781)) ;
    mux21_ni ix62767 (.Y (nx62766), .A0 (nx62750), .A1 (nx62762), .S0 (nx23851)
             ) ;
    mux21_ni ix62751 (.Y (nx62750), .A0 (inputs_308__15), .A1 (inputs_309__15), 
             .S0 (nx24783)) ;
    mux21_ni ix62763 (.Y (nx62762), .A0 (inputs_310__15), .A1 (inputs_311__15), 
             .S0 (nx24783)) ;
    nand04 ix21406 (.Y (nx21405), .A0 (nx22369), .A1 (nx23851), .A2 (nx24783), .A3 (
           nx62710)) ;
    mux21_ni ix62711 (.Y (nx62710), .A0 (inputs_291__15), .A1 (inputs_307__15), 
             .S0 (nx23089)) ;
    mux21_ni ix62697 (.Y (nx62696), .A0 (nx62632), .A1 (nx62692), .S0 (nx23089)
             ) ;
    mux21_ni ix62633 (.Y (nx62632), .A0 (nx62600), .A1 (nx62628), .S0 (nx23327)
             ) ;
    mux21_ni ix62601 (.Y (nx62600), .A0 (nx62584), .A1 (nx62596), .S0 (nx23851)
             ) ;
    mux21_ni ix62585 (.Y (nx62584), .A0 (inputs_296__15), .A1 (inputs_297__15), 
             .S0 (nx24783)) ;
    mux21_ni ix62597 (.Y (nx62596), .A0 (inputs_298__15), .A1 (inputs_299__15), 
             .S0 (nx24783)) ;
    mux21_ni ix62629 (.Y (nx62628), .A0 (nx62612), .A1 (nx62624), .S0 (nx23851)
             ) ;
    mux21_ni ix62613 (.Y (nx62612), .A0 (inputs_300__15), .A1 (inputs_301__15), 
             .S0 (nx24783)) ;
    mux21_ni ix62625 (.Y (nx62624), .A0 (inputs_302__15), .A1 (inputs_303__15), 
             .S0 (nx24783)) ;
    mux21_ni ix62693 (.Y (nx62692), .A0 (nx62660), .A1 (nx62688), .S0 (nx23329)
             ) ;
    mux21_ni ix62661 (.Y (nx62660), .A0 (nx62644), .A1 (nx62656), .S0 (nx23853)
             ) ;
    mux21_ni ix62645 (.Y (nx62644), .A0 (inputs_312__15), .A1 (inputs_313__15), 
             .S0 (nx24785)) ;
    mux21_ni ix62657 (.Y (nx62656), .A0 (inputs_314__15), .A1 (inputs_315__15), 
             .S0 (nx24785)) ;
    mux21_ni ix62689 (.Y (nx62688), .A0 (nx62672), .A1 (nx62684), .S0 (nx23853)
             ) ;
    mux21_ni ix62673 (.Y (nx62672), .A0 (inputs_316__15), .A1 (inputs_317__15), 
             .S0 (nx24785)) ;
    mux21_ni ix62685 (.Y (nx62684), .A0 (inputs_318__15), .A1 (inputs_319__15), 
             .S0 (nx24785)) ;
    mux21_ni ix63205 (.Y (nx63204), .A0 (nx62992), .A1 (nx63200), .S0 (nx22663)
             ) ;
    mux21_ni ix62993 (.Y (nx62992), .A0 (nx62986), .A1 (nx62908), .S0 (nx23185)
             ) ;
    oai21 ix62987 (.Y (nx62986), .A0 (nx22369), .A1 (nx21435), .B0 (nx21447)) ;
    mux21 ix21436 (.Y (nx21435), .A0 (nx62950), .A1 (nx62978), .S0 (nx23089)) ;
    mux21_ni ix62951 (.Y (nx62950), .A0 (nx62934), .A1 (nx62946), .S0 (nx23853)
             ) ;
    mux21_ni ix62935 (.Y (nx62934), .A0 (inputs_324__15), .A1 (inputs_325__15), 
             .S0 (nx24785)) ;
    mux21_ni ix62947 (.Y (nx62946), .A0 (inputs_326__15), .A1 (inputs_327__15), 
             .S0 (nx24785)) ;
    mux21_ni ix62979 (.Y (nx62978), .A0 (nx62962), .A1 (nx62974), .S0 (nx23853)
             ) ;
    mux21_ni ix62963 (.Y (nx62962), .A0 (inputs_340__15), .A1 (inputs_341__15), 
             .S0 (nx24785)) ;
    mux21_ni ix62975 (.Y (nx62974), .A0 (inputs_342__15), .A1 (inputs_343__15), 
             .S0 (nx24787)) ;
    nand04 ix21448 (.Y (nx21447), .A0 (nx22369), .A1 (nx23853), .A2 (nx24787), .A3 (
           nx62922)) ;
    mux21_ni ix62923 (.Y (nx62922), .A0 (inputs_323__15), .A1 (inputs_339__15), 
             .S0 (nx23089)) ;
    mux21_ni ix62909 (.Y (nx62908), .A0 (nx62844), .A1 (nx62904), .S0 (nx23089)
             ) ;
    mux21_ni ix62845 (.Y (nx62844), .A0 (nx62812), .A1 (nx62840), .S0 (nx23329)
             ) ;
    mux21_ni ix62813 (.Y (nx62812), .A0 (nx62796), .A1 (nx62808), .S0 (nx23853)
             ) ;
    mux21_ni ix62797 (.Y (nx62796), .A0 (inputs_328__15), .A1 (inputs_329__15), 
             .S0 (nx24787)) ;
    mux21_ni ix62809 (.Y (nx62808), .A0 (inputs_330__15), .A1 (inputs_331__15), 
             .S0 (nx24787)) ;
    mux21_ni ix62841 (.Y (nx62840), .A0 (nx62824), .A1 (nx62836), .S0 (nx23853)
             ) ;
    mux21_ni ix62825 (.Y (nx62824), .A0 (inputs_332__15), .A1 (inputs_333__15), 
             .S0 (nx24787)) ;
    mux21_ni ix62837 (.Y (nx62836), .A0 (inputs_334__15), .A1 (inputs_335__15), 
             .S0 (nx24787)) ;
    mux21_ni ix62905 (.Y (nx62904), .A0 (nx62872), .A1 (nx62900), .S0 (nx23329)
             ) ;
    mux21_ni ix62873 (.Y (nx62872), .A0 (nx62856), .A1 (nx62868), .S0 (nx23855)
             ) ;
    mux21_ni ix62857 (.Y (nx62856), .A0 (inputs_344__15), .A1 (inputs_345__15), 
             .S0 (nx24787)) ;
    mux21_ni ix62869 (.Y (nx62868), .A0 (inputs_346__15), .A1 (inputs_347__15), 
             .S0 (nx24789)) ;
    mux21_ni ix62901 (.Y (nx62900), .A0 (nx62884), .A1 (nx62896), .S0 (nx23855)
             ) ;
    mux21_ni ix62885 (.Y (nx62884), .A0 (inputs_348__15), .A1 (inputs_349__15), 
             .S0 (nx24789)) ;
    mux21_ni ix62897 (.Y (nx62896), .A0 (inputs_350__15), .A1 (inputs_351__15), 
             .S0 (nx24789)) ;
    mux21_ni ix63201 (.Y (nx63200), .A0 (nx63194), .A1 (nx63116), .S0 (nx23185)
             ) ;
    oai21 ix63195 (.Y (nx63194), .A0 (nx22369), .A1 (nx21479), .B0 (nx21491)) ;
    mux21 ix21480 (.Y (nx21479), .A0 (nx63158), .A1 (nx63186), .S0 (nx23091)) ;
    mux21_ni ix63159 (.Y (nx63158), .A0 (nx63142), .A1 (nx63154), .S0 (nx23855)
             ) ;
    mux21_ni ix63143 (.Y (nx63142), .A0 (inputs_356__15), .A1 (inputs_357__15), 
             .S0 (nx24789)) ;
    mux21_ni ix63155 (.Y (nx63154), .A0 (inputs_358__15), .A1 (inputs_359__15), 
             .S0 (nx24789)) ;
    mux21_ni ix63187 (.Y (nx63186), .A0 (nx63170), .A1 (nx63182), .S0 (nx23855)
             ) ;
    mux21_ni ix63171 (.Y (nx63170), .A0 (inputs_372__15), .A1 (inputs_373__15), 
             .S0 (nx24789)) ;
    mux21_ni ix63183 (.Y (nx63182), .A0 (inputs_374__15), .A1 (inputs_375__15), 
             .S0 (nx24789)) ;
    nand04 ix21492 (.Y (nx21491), .A0 (nx22369), .A1 (nx23855), .A2 (nx24791), .A3 (
           nx63130)) ;
    mux21_ni ix63131 (.Y (nx63130), .A0 (inputs_355__15), .A1 (inputs_371__15), 
             .S0 (nx23091)) ;
    mux21_ni ix63117 (.Y (nx63116), .A0 (nx63052), .A1 (nx63112), .S0 (nx23091)
             ) ;
    mux21_ni ix63053 (.Y (nx63052), .A0 (nx63020), .A1 (nx63048), .S0 (nx23329)
             ) ;
    mux21_ni ix63021 (.Y (nx63020), .A0 (nx63004), .A1 (nx63016), .S0 (nx23855)
             ) ;
    mux21_ni ix63005 (.Y (nx63004), .A0 (inputs_360__15), .A1 (inputs_361__15), 
             .S0 (nx24791)) ;
    mux21_ni ix63017 (.Y (nx63016), .A0 (inputs_362__15), .A1 (inputs_363__15), 
             .S0 (nx24791)) ;
    mux21_ni ix63049 (.Y (nx63048), .A0 (nx63032), .A1 (nx63044), .S0 (nx23855)
             ) ;
    mux21_ni ix63033 (.Y (nx63032), .A0 (inputs_364__15), .A1 (inputs_365__15), 
             .S0 (nx24791)) ;
    mux21_ni ix63045 (.Y (nx63044), .A0 (inputs_366__15), .A1 (inputs_367__15), 
             .S0 (nx24791)) ;
    mux21_ni ix63113 (.Y (nx63112), .A0 (nx63080), .A1 (nx63108), .S0 (nx23329)
             ) ;
    mux21_ni ix63081 (.Y (nx63080), .A0 (nx63064), .A1 (nx63076), .S0 (nx23857)
             ) ;
    mux21_ni ix63065 (.Y (nx63064), .A0 (inputs_376__15), .A1 (inputs_377__15), 
             .S0 (nx24791)) ;
    mux21_ni ix63077 (.Y (nx63076), .A0 (inputs_378__15), .A1 (inputs_379__15), 
             .S0 (nx24791)) ;
    mux21_ni ix63109 (.Y (nx63108), .A0 (nx63092), .A1 (nx63104), .S0 (nx23857)
             ) ;
    mux21_ni ix63093 (.Y (nx63092), .A0 (inputs_380__15), .A1 (inputs_381__15), 
             .S0 (nx24793)) ;
    mux21_ni ix63105 (.Y (nx63104), .A0 (inputs_382__15), .A1 (inputs_383__15), 
             .S0 (nx24793)) ;
    mux21_ni ix64053 (.Y (nx64052), .A0 (nx63628), .A1 (nx64048), .S0 (nx22519)
             ) ;
    mux21_ni ix63629 (.Y (nx63628), .A0 (nx63416), .A1 (nx63624), .S0 (nx22663)
             ) ;
    mux21_ni ix63417 (.Y (nx63416), .A0 (nx63410), .A1 (nx63332), .S0 (nx23185)
             ) ;
    oai21 ix63411 (.Y (nx63410), .A0 (nx22369), .A1 (nx21525), .B0 (nx21539)) ;
    mux21 ix21526 (.Y (nx21525), .A0 (nx63374), .A1 (nx63402), .S0 (nx23091)) ;
    mux21_ni ix63375 (.Y (nx63374), .A0 (nx63358), .A1 (nx63370), .S0 (nx23857)
             ) ;
    mux21_ni ix63359 (.Y (nx63358), .A0 (inputs_388__15), .A1 (inputs_389__15), 
             .S0 (nx24793)) ;
    mux21_ni ix63371 (.Y (nx63370), .A0 (inputs_390__15), .A1 (inputs_391__15), 
             .S0 (nx24793)) ;
    mux21_ni ix63403 (.Y (nx63402), .A0 (nx63386), .A1 (nx63398), .S0 (nx23857)
             ) ;
    mux21_ni ix63387 (.Y (nx63386), .A0 (inputs_404__15), .A1 (inputs_405__15), 
             .S0 (nx24793)) ;
    mux21_ni ix63399 (.Y (nx63398), .A0 (inputs_406__15), .A1 (inputs_407__15), 
             .S0 (nx24793)) ;
    nand04 ix21540 (.Y (nx21539), .A0 (nx22371), .A1 (nx23857), .A2 (nx24793), .A3 (
           nx63346)) ;
    mux21_ni ix63347 (.Y (nx63346), .A0 (inputs_387__15), .A1 (inputs_403__15), 
             .S0 (nx23091)) ;
    mux21_ni ix63333 (.Y (nx63332), .A0 (nx63268), .A1 (nx63328), .S0 (nx23091)
             ) ;
    mux21_ni ix63269 (.Y (nx63268), .A0 (nx63236), .A1 (nx63264), .S0 (nx23329)
             ) ;
    mux21_ni ix63237 (.Y (nx63236), .A0 (nx63220), .A1 (nx63232), .S0 (nx23857)
             ) ;
    mux21_ni ix63221 (.Y (nx63220), .A0 (inputs_392__15), .A1 (inputs_393__15), 
             .S0 (nx24795)) ;
    mux21_ni ix63233 (.Y (nx63232), .A0 (inputs_394__15), .A1 (inputs_395__15), 
             .S0 (nx24795)) ;
    mux21_ni ix63265 (.Y (nx63264), .A0 (nx63248), .A1 (nx63260), .S0 (nx23857)
             ) ;
    mux21_ni ix63249 (.Y (nx63248), .A0 (inputs_396__15), .A1 (inputs_397__15), 
             .S0 (nx24795)) ;
    mux21_ni ix63261 (.Y (nx63260), .A0 (inputs_398__15), .A1 (inputs_399__15), 
             .S0 (nx24795)) ;
    mux21_ni ix63329 (.Y (nx63328), .A0 (nx63296), .A1 (nx63324), .S0 (nx23329)
             ) ;
    mux21_ni ix63297 (.Y (nx63296), .A0 (nx63280), .A1 (nx63292), .S0 (nx23859)
             ) ;
    mux21_ni ix63281 (.Y (nx63280), .A0 (inputs_408__15), .A1 (inputs_409__15), 
             .S0 (nx24795)) ;
    mux21_ni ix63293 (.Y (nx63292), .A0 (inputs_410__15), .A1 (inputs_411__15), 
             .S0 (nx24795)) ;
    mux21_ni ix63325 (.Y (nx63324), .A0 (nx63308), .A1 (nx63320), .S0 (nx23859)
             ) ;
    mux21_ni ix63309 (.Y (nx63308), .A0 (inputs_412__15), .A1 (inputs_413__15), 
             .S0 (nx24795)) ;
    mux21_ni ix63321 (.Y (nx63320), .A0 (inputs_414__15), .A1 (inputs_415__15), 
             .S0 (nx24797)) ;
    mux21_ni ix63625 (.Y (nx63624), .A0 (nx63618), .A1 (nx63540), .S0 (nx23187)
             ) ;
    oai21 ix63619 (.Y (nx63618), .A0 (nx22371), .A1 (nx21569), .B0 (nx21583)) ;
    mux21 ix21570 (.Y (nx21569), .A0 (nx63582), .A1 (nx63610), .S0 (nx23091)) ;
    mux21_ni ix63583 (.Y (nx63582), .A0 (nx63566), .A1 (nx63578), .S0 (nx23859)
             ) ;
    mux21_ni ix63567 (.Y (nx63566), .A0 (inputs_420__15), .A1 (inputs_421__15), 
             .S0 (nx24797)) ;
    mux21_ni ix63579 (.Y (nx63578), .A0 (inputs_422__15), .A1 (inputs_423__15), 
             .S0 (nx24797)) ;
    mux21_ni ix63611 (.Y (nx63610), .A0 (nx63594), .A1 (nx63606), .S0 (nx23859)
             ) ;
    mux21_ni ix63595 (.Y (nx63594), .A0 (inputs_436__15), .A1 (inputs_437__15), 
             .S0 (nx24797)) ;
    mux21_ni ix63607 (.Y (nx63606), .A0 (inputs_438__15), .A1 (inputs_439__15), 
             .S0 (nx24797)) ;
    nand04 ix21584 (.Y (nx21583), .A0 (nx22371), .A1 (nx23859), .A2 (nx24797), .A3 (
           nx63554)) ;
    mux21_ni ix63555 (.Y (nx63554), .A0 (inputs_419__15), .A1 (inputs_435__15), 
             .S0 (nx23093)) ;
    mux21_ni ix63541 (.Y (nx63540), .A0 (nx63476), .A1 (nx63536), .S0 (nx23093)
             ) ;
    mux21_ni ix63477 (.Y (nx63476), .A0 (nx63444), .A1 (nx63472), .S0 (nx23331)
             ) ;
    mux21_ni ix63445 (.Y (nx63444), .A0 (nx63428), .A1 (nx63440), .S0 (nx23859)
             ) ;
    mux21_ni ix63429 (.Y (nx63428), .A0 (inputs_424__15), .A1 (inputs_425__15), 
             .S0 (nx24797)) ;
    mux21_ni ix63441 (.Y (nx63440), .A0 (inputs_426__15), .A1 (inputs_427__15), 
             .S0 (nx24799)) ;
    mux21_ni ix63473 (.Y (nx63472), .A0 (nx63456), .A1 (nx63468), .S0 (nx23859)
             ) ;
    mux21_ni ix63457 (.Y (nx63456), .A0 (inputs_428__15), .A1 (inputs_429__15), 
             .S0 (nx24799)) ;
    mux21_ni ix63469 (.Y (nx63468), .A0 (inputs_430__15), .A1 (inputs_431__15), 
             .S0 (nx24799)) ;
    mux21_ni ix63537 (.Y (nx63536), .A0 (nx63504), .A1 (nx63532), .S0 (nx23331)
             ) ;
    mux21_ni ix63505 (.Y (nx63504), .A0 (nx63488), .A1 (nx63500), .S0 (nx23861)
             ) ;
    mux21_ni ix63489 (.Y (nx63488), .A0 (inputs_440__15), .A1 (inputs_441__15), 
             .S0 (nx24799)) ;
    mux21_ni ix63501 (.Y (nx63500), .A0 (inputs_442__15), .A1 (inputs_443__15), 
             .S0 (nx24799)) ;
    mux21_ni ix63533 (.Y (nx63532), .A0 (nx63516), .A1 (nx63528), .S0 (nx23861)
             ) ;
    mux21_ni ix63517 (.Y (nx63516), .A0 (inputs_444__15), .A1 (inputs_445__15), 
             .S0 (nx24799)) ;
    mux21_ni ix63529 (.Y (nx63528), .A0 (inputs_446__15), .A1 (inputs_447__15), 
             .S0 (nx24799)) ;
    mux21_ni ix64049 (.Y (nx64048), .A0 (nx63836), .A1 (nx64044), .S0 (nx22665)
             ) ;
    mux21_ni ix63837 (.Y (nx63836), .A0 (nx63830), .A1 (nx63752), .S0 (nx23187)
             ) ;
    oai21 ix63831 (.Y (nx63830), .A0 (nx22371), .A1 (nx21617), .B0 (nx21631)) ;
    mux21 ix21618 (.Y (nx21617), .A0 (nx63794), .A1 (nx63822), .S0 (nx23093)) ;
    mux21_ni ix63795 (.Y (nx63794), .A0 (nx63778), .A1 (nx63790), .S0 (nx23861)
             ) ;
    mux21_ni ix63779 (.Y (nx63778), .A0 (inputs_452__15), .A1 (inputs_453__15), 
             .S0 (nx24801)) ;
    mux21_ni ix63791 (.Y (nx63790), .A0 (inputs_454__15), .A1 (inputs_455__15), 
             .S0 (nx24801)) ;
    mux21_ni ix63823 (.Y (nx63822), .A0 (nx63806), .A1 (nx63818), .S0 (nx23861)
             ) ;
    mux21_ni ix63807 (.Y (nx63806), .A0 (inputs_468__15), .A1 (inputs_469__15), 
             .S0 (nx24801)) ;
    mux21_ni ix63819 (.Y (nx63818), .A0 (inputs_470__15), .A1 (inputs_471__15), 
             .S0 (nx24801)) ;
    nand04 ix21632 (.Y (nx21631), .A0 (nx22371), .A1 (nx23861), .A2 (nx24801), .A3 (
           nx63766)) ;
    mux21_ni ix63767 (.Y (nx63766), .A0 (inputs_451__15), .A1 (inputs_467__15), 
             .S0 (nx23093)) ;
    mux21_ni ix63753 (.Y (nx63752), .A0 (nx63688), .A1 (nx63748), .S0 (nx23093)
             ) ;
    mux21_ni ix63689 (.Y (nx63688), .A0 (nx63656), .A1 (nx63684), .S0 (nx23331)
             ) ;
    mux21_ni ix63657 (.Y (nx63656), .A0 (nx63640), .A1 (nx63652), .S0 (nx23861)
             ) ;
    mux21_ni ix63641 (.Y (nx63640), .A0 (inputs_456__15), .A1 (inputs_457__15), 
             .S0 (nx24801)) ;
    mux21_ni ix63653 (.Y (nx63652), .A0 (inputs_458__15), .A1 (inputs_459__15), 
             .S0 (nx24801)) ;
    mux21_ni ix63685 (.Y (nx63684), .A0 (nx63668), .A1 (nx63680), .S0 (nx23861)
             ) ;
    mux21_ni ix63669 (.Y (nx63668), .A0 (inputs_460__15), .A1 (inputs_461__15), 
             .S0 (nx24803)) ;
    mux21_ni ix63681 (.Y (nx63680), .A0 (inputs_462__15), .A1 (inputs_463__15), 
             .S0 (nx24803)) ;
    mux21_ni ix63749 (.Y (nx63748), .A0 (nx63716), .A1 (nx63744), .S0 (nx23331)
             ) ;
    mux21_ni ix63717 (.Y (nx63716), .A0 (nx63700), .A1 (nx63712), .S0 (nx23863)
             ) ;
    mux21_ni ix63701 (.Y (nx63700), .A0 (inputs_472__15), .A1 (inputs_473__15), 
             .S0 (nx24803)) ;
    mux21_ni ix63713 (.Y (nx63712), .A0 (inputs_474__15), .A1 (inputs_475__15), 
             .S0 (nx24803)) ;
    mux21_ni ix63745 (.Y (nx63744), .A0 (nx63728), .A1 (nx63740), .S0 (nx23863)
             ) ;
    mux21_ni ix63729 (.Y (nx63728), .A0 (inputs_476__15), .A1 (inputs_477__15), 
             .S0 (nx24803)) ;
    mux21_ni ix63741 (.Y (nx63740), .A0 (inputs_478__15), .A1 (inputs_479__15), 
             .S0 (nx24803)) ;
    mux21_ni ix64045 (.Y (nx64044), .A0 (nx64038), .A1 (nx63960), .S0 (nx23187)
             ) ;
    oai21 ix64039 (.Y (nx64038), .A0 (nx22371), .A1 (nx21661), .B0 (nx21673)) ;
    mux21 ix21662 (.Y (nx21661), .A0 (nx64002), .A1 (nx64030), .S0 (nx23093)) ;
    mux21_ni ix64003 (.Y (nx64002), .A0 (nx63986), .A1 (nx63998), .S0 (nx23863)
             ) ;
    mux21_ni ix63987 (.Y (nx63986), .A0 (inputs_484__15), .A1 (inputs_485__15), 
             .S0 (nx24803)) ;
    mux21_ni ix63999 (.Y (nx63998), .A0 (inputs_486__15), .A1 (inputs_487__15), 
             .S0 (nx24805)) ;
    mux21_ni ix64031 (.Y (nx64030), .A0 (nx64014), .A1 (nx64026), .S0 (nx23863)
             ) ;
    mux21_ni ix64015 (.Y (nx64014), .A0 (inputs_500__15), .A1 (inputs_501__15), 
             .S0 (nx24805)) ;
    mux21_ni ix64027 (.Y (nx64026), .A0 (inputs_502__15), .A1 (inputs_503__15), 
             .S0 (nx24805)) ;
    nand04 ix21674 (.Y (nx21673), .A0 (nx22371), .A1 (nx23863), .A2 (nx24805), .A3 (
           nx63974)) ;
    mux21_ni ix63975 (.Y (nx63974), .A0 (inputs_483__15), .A1 (inputs_499__15), 
             .S0 (nx23093)) ;
    mux21_ni ix63961 (.Y (nx63960), .A0 (nx63896), .A1 (nx63956), .S0 (nx23095)
             ) ;
    mux21_ni ix63897 (.Y (nx63896), .A0 (nx63864), .A1 (nx63892), .S0 (nx23331)
             ) ;
    mux21_ni ix63865 (.Y (nx63864), .A0 (nx63848), .A1 (nx63860), .S0 (nx23863)
             ) ;
    mux21_ni ix63849 (.Y (nx63848), .A0 (inputs_488__15), .A1 (inputs_489__15), 
             .S0 (nx24805)) ;
    mux21_ni ix63861 (.Y (nx63860), .A0 (inputs_490__15), .A1 (inputs_491__15), 
             .S0 (nx24805)) ;
    mux21_ni ix63893 (.Y (nx63892), .A0 (nx63876), .A1 (nx63888), .S0 (nx23863)
             ) ;
    mux21_ni ix63877 (.Y (nx63876), .A0 (inputs_492__15), .A1 (inputs_493__15), 
             .S0 (nx24805)) ;
    mux21_ni ix63889 (.Y (nx63888), .A0 (inputs_494__15), .A1 (inputs_495__15), 
             .S0 (nx24807)) ;
    mux21_ni ix63957 (.Y (nx63956), .A0 (nx63924), .A1 (nx63952), .S0 (nx23331)
             ) ;
    mux21_ni ix63925 (.Y (nx63924), .A0 (nx63908), .A1 (nx63920), .S0 (nx23865)
             ) ;
    mux21_ni ix63909 (.Y (nx63908), .A0 (inputs_504__15), .A1 (inputs_505__15), 
             .S0 (nx24807)) ;
    mux21_ni ix63921 (.Y (nx63920), .A0 (inputs_506__15), .A1 (inputs_507__15), 
             .S0 (nx24807)) ;
    mux21_ni ix63953 (.Y (nx63952), .A0 (nx63936), .A1 (nx63948), .S0 (nx23865)
             ) ;
    mux21_ni ix63937 (.Y (nx63936), .A0 (inputs_508__15), .A1 (inputs_509__15), 
             .S0 (nx24807)) ;
    mux21_ni ix63949 (.Y (nx63948), .A0 (inputs_510__15), .A1 (inputs_511__15), 
             .S0 (nx24807)) ;
    aoi32 ix21702 (.Y (nx21701), .A0 (nx64822), .A1 (nx24839), .A2 (nx22373), .B0 (
          nx22225), .B1 (nx66518)) ;
    oai21 ix64823 (.Y (nx64822), .A0 (nx23865), .A1 (nx21705), .B0 (nx21807)) ;
    mux21 ix21706 (.Y (nx21705), .A0 (nx64810), .A1 (nx64560), .S0 (nx24807)) ;
    mux21_ni ix64811 (.Y (nx64810), .A0 (nx64682), .A1 (nx64806), .S0 (nx22405)
             ) ;
    mux21_ni ix64683 (.Y (nx64682), .A0 (nx64618), .A1 (nx64678), .S0 (nx22445)
             ) ;
    mux21_ni ix64619 (.Y (nx64618), .A0 (nx64586), .A1 (nx64614), .S0 (nx22519)
             ) ;
    mux21_ni ix64587 (.Y (nx64586), .A0 (nx64570), .A1 (nx64582), .S0 (nx22665)
             ) ;
    mux21_ni ix64571 (.Y (nx64570), .A0 (inputs_0__15), .A1 (inputs_16__15), .S0 (
             nx23095)) ;
    mux21_ni ix64583 (.Y (nx64582), .A0 (inputs_32__15), .A1 (inputs_48__15), .S0 (
             nx23095)) ;
    mux21_ni ix64615 (.Y (nx64614), .A0 (nx64598), .A1 (nx64610), .S0 (nx22665)
             ) ;
    mux21_ni ix64599 (.Y (nx64598), .A0 (inputs_64__15), .A1 (inputs_80__15), .S0 (
             nx23095)) ;
    mux21_ni ix64611 (.Y (nx64610), .A0 (inputs_96__15), .A1 (inputs_112__15), .S0 (
             nx23095)) ;
    mux21_ni ix64679 (.Y (nx64678), .A0 (nx64646), .A1 (nx64674), .S0 (nx22519)
             ) ;
    mux21_ni ix64647 (.Y (nx64646), .A0 (nx64630), .A1 (nx64642), .S0 (nx22665)
             ) ;
    mux21_ni ix64631 (.Y (nx64630), .A0 (inputs_128__15), .A1 (inputs_144__15), 
             .S0 (nx23095)) ;
    mux21_ni ix64643 (.Y (nx64642), .A0 (inputs_160__15), .A1 (inputs_176__15), 
             .S0 (nx23095)) ;
    mux21_ni ix64675 (.Y (nx64674), .A0 (nx64658), .A1 (nx64670), .S0 (nx22665)
             ) ;
    mux21_ni ix64659 (.Y (nx64658), .A0 (inputs_192__15), .A1 (inputs_208__15), 
             .S0 (nx23097)) ;
    mux21_ni ix64671 (.Y (nx64670), .A0 (inputs_224__15), .A1 (inputs_240__15), 
             .S0 (nx23097)) ;
    mux21_ni ix64807 (.Y (nx64806), .A0 (nx64742), .A1 (nx64802), .S0 (nx22445)
             ) ;
    mux21_ni ix64743 (.Y (nx64742), .A0 (nx64710), .A1 (nx64738), .S0 (nx22519)
             ) ;
    mux21_ni ix64711 (.Y (nx64710), .A0 (nx64694), .A1 (nx64706), .S0 (nx22665)
             ) ;
    mux21_ni ix64695 (.Y (nx64694), .A0 (inputs_256__15), .A1 (inputs_272__15), 
             .S0 (nx23097)) ;
    mux21_ni ix64707 (.Y (nx64706), .A0 (inputs_288__15), .A1 (inputs_304__15), 
             .S0 (nx23097)) ;
    mux21_ni ix64739 (.Y (nx64738), .A0 (nx64722), .A1 (nx64734), .S0 (nx22665)
             ) ;
    mux21_ni ix64723 (.Y (nx64722), .A0 (inputs_320__15), .A1 (inputs_336__15), 
             .S0 (nx23097)) ;
    mux21_ni ix64735 (.Y (nx64734), .A0 (inputs_352__15), .A1 (inputs_368__15), 
             .S0 (nx23097)) ;
    mux21_ni ix64803 (.Y (nx64802), .A0 (nx64770), .A1 (nx64798), .S0 (nx22521)
             ) ;
    mux21_ni ix64771 (.Y (nx64770), .A0 (nx64754), .A1 (nx64766), .S0 (nx22667)
             ) ;
    mux21_ni ix64755 (.Y (nx64754), .A0 (inputs_384__15), .A1 (inputs_400__15), 
             .S0 (nx23097)) ;
    mux21_ni ix64767 (.Y (nx64766), .A0 (inputs_416__15), .A1 (inputs_432__15), 
             .S0 (nx23099)) ;
    mux21_ni ix64799 (.Y (nx64798), .A0 (nx64782), .A1 (nx64794), .S0 (nx22667)
             ) ;
    mux21_ni ix64783 (.Y (nx64782), .A0 (inputs_448__15), .A1 (inputs_464__15), 
             .S0 (nx23099)) ;
    mux21_ni ix64795 (.Y (nx64794), .A0 (inputs_480__15), .A1 (inputs_496__15), 
             .S0 (nx23099)) ;
    mux21_ni ix64561 (.Y (nx64560), .A0 (nx64432), .A1 (nx64556), .S0 (nx22405)
             ) ;
    mux21_ni ix64433 (.Y (nx64432), .A0 (nx64368), .A1 (nx64428), .S0 (nx22445)
             ) ;
    mux21_ni ix64369 (.Y (nx64368), .A0 (nx64336), .A1 (nx64364), .S0 (nx22521)
             ) ;
    mux21_ni ix64337 (.Y (nx64336), .A0 (nx64320), .A1 (nx64332), .S0 (nx22667)
             ) ;
    mux21_ni ix64321 (.Y (nx64320), .A0 (inputs_1__15), .A1 (inputs_17__15), .S0 (
             nx23099)) ;
    mux21_ni ix64333 (.Y (nx64332), .A0 (inputs_33__15), .A1 (inputs_49__15), .S0 (
             nx23099)) ;
    mux21_ni ix64365 (.Y (nx64364), .A0 (nx64348), .A1 (nx64360), .S0 (nx22667)
             ) ;
    mux21_ni ix64349 (.Y (nx64348), .A0 (inputs_65__15), .A1 (inputs_81__15), .S0 (
             nx23099)) ;
    mux21_ni ix64361 (.Y (nx64360), .A0 (inputs_97__15), .A1 (inputs_113__15), .S0 (
             nx23099)) ;
    mux21_ni ix64429 (.Y (nx64428), .A0 (nx64396), .A1 (nx64424), .S0 (nx22521)
             ) ;
    mux21_ni ix64397 (.Y (nx64396), .A0 (nx64380), .A1 (nx64392), .S0 (nx22667)
             ) ;
    mux21_ni ix64381 (.Y (nx64380), .A0 (inputs_129__15), .A1 (inputs_145__15), 
             .S0 (nx23101)) ;
    mux21_ni ix64393 (.Y (nx64392), .A0 (inputs_161__15), .A1 (inputs_177__15), 
             .S0 (nx23101)) ;
    mux21_ni ix64425 (.Y (nx64424), .A0 (nx64408), .A1 (nx64420), .S0 (nx22667)
             ) ;
    mux21_ni ix64409 (.Y (nx64408), .A0 (inputs_193__15), .A1 (inputs_209__15), 
             .S0 (nx23101)) ;
    mux21_ni ix64421 (.Y (nx64420), .A0 (inputs_225__15), .A1 (inputs_241__15), 
             .S0 (nx23101)) ;
    mux21_ni ix64557 (.Y (nx64556), .A0 (nx64492), .A1 (nx64552), .S0 (nx22445)
             ) ;
    mux21_ni ix64493 (.Y (nx64492), .A0 (nx64460), .A1 (nx64488), .S0 (nx22521)
             ) ;
    mux21_ni ix64461 (.Y (nx64460), .A0 (nx64444), .A1 (nx64456), .S0 (nx22667)
             ) ;
    mux21_ni ix64445 (.Y (nx64444), .A0 (inputs_257__15), .A1 (inputs_273__15), 
             .S0 (nx23101)) ;
    mux21_ni ix64457 (.Y (nx64456), .A0 (inputs_289__15), .A1 (inputs_305__15), 
             .S0 (nx23101)) ;
    mux21_ni ix64489 (.Y (nx64488), .A0 (nx64472), .A1 (nx64484), .S0 (nx22669)
             ) ;
    mux21_ni ix64473 (.Y (nx64472), .A0 (inputs_321__15), .A1 (inputs_337__15), 
             .S0 (nx23101)) ;
    mux21_ni ix64485 (.Y (nx64484), .A0 (inputs_353__15), .A1 (inputs_369__15), 
             .S0 (nx23103)) ;
    mux21_ni ix64553 (.Y (nx64552), .A0 (nx64520), .A1 (nx64548), .S0 (nx22521)
             ) ;
    mux21_ni ix64521 (.Y (nx64520), .A0 (nx64504), .A1 (nx64516), .S0 (nx22669)
             ) ;
    mux21_ni ix64505 (.Y (nx64504), .A0 (inputs_385__15), .A1 (inputs_401__15), 
             .S0 (nx23103)) ;
    mux21_ni ix64517 (.Y (nx64516), .A0 (inputs_417__15), .A1 (inputs_433__15), 
             .S0 (nx23103)) ;
    mux21_ni ix64549 (.Y (nx64548), .A0 (nx64532), .A1 (nx64544), .S0 (nx22669)
             ) ;
    mux21_ni ix64533 (.Y (nx64532), .A0 (inputs_449__15), .A1 (inputs_465__15), 
             .S0 (nx23103)) ;
    mux21_ni ix64545 (.Y (nx64544), .A0 (inputs_481__15), .A1 (inputs_497__15), 
             .S0 (nx23103)) ;
    nand03 ix21808 (.Y (nx21807), .A0 (nx64306), .A1 (nx23865), .A2 (nx22383)) ;
    mux21_ni ix64307 (.Y (nx64306), .A0 (nx64178), .A1 (nx64302), .S0 (nx22405)
             ) ;
    mux21_ni ix64179 (.Y (nx64178), .A0 (nx64114), .A1 (nx64174), .S0 (nx22445)
             ) ;
    mux21_ni ix64115 (.Y (nx64114), .A0 (nx64082), .A1 (nx64110), .S0 (nx22521)
             ) ;
    mux21_ni ix64083 (.Y (nx64082), .A0 (nx64066), .A1 (nx64078), .S0 (nx22669)
             ) ;
    mux21_ni ix64067 (.Y (nx64066), .A0 (inputs_2__15), .A1 (inputs_18__15), .S0 (
             nx23103)) ;
    mux21_ni ix64079 (.Y (nx64078), .A0 (inputs_34__15), .A1 (inputs_50__15), .S0 (
             nx23103)) ;
    mux21_ni ix64111 (.Y (nx64110), .A0 (nx64094), .A1 (nx64106), .S0 (nx22669)
             ) ;
    mux21_ni ix64095 (.Y (nx64094), .A0 (inputs_66__15), .A1 (inputs_82__15), .S0 (
             nx23105)) ;
    mux21_ni ix64107 (.Y (nx64106), .A0 (inputs_98__15), .A1 (inputs_114__15), .S0 (
             nx23105)) ;
    mux21_ni ix64175 (.Y (nx64174), .A0 (nx64142), .A1 (nx64170), .S0 (nx22521)
             ) ;
    mux21_ni ix64143 (.Y (nx64142), .A0 (nx64126), .A1 (nx64138), .S0 (nx22669)
             ) ;
    mux21_ni ix64127 (.Y (nx64126), .A0 (inputs_130__15), .A1 (inputs_146__15), 
             .S0 (nx23105)) ;
    mux21_ni ix64139 (.Y (nx64138), .A0 (inputs_162__15), .A1 (inputs_178__15), 
             .S0 (nx23105)) ;
    mux21_ni ix64171 (.Y (nx64170), .A0 (nx64154), .A1 (nx64166), .S0 (nx22669)
             ) ;
    mux21_ni ix64155 (.Y (nx64154), .A0 (inputs_194__15), .A1 (inputs_210__15), 
             .S0 (nx23105)) ;
    mux21_ni ix64167 (.Y (nx64166), .A0 (inputs_226__15), .A1 (inputs_242__15), 
             .S0 (nx23105)) ;
    mux21_ni ix64303 (.Y (nx64302), .A0 (nx64238), .A1 (nx64298), .S0 (nx22447)
             ) ;
    mux21_ni ix64239 (.Y (nx64238), .A0 (nx64206), .A1 (nx64234), .S0 (nx22523)
             ) ;
    mux21_ni ix64207 (.Y (nx64206), .A0 (nx64190), .A1 (nx64202), .S0 (nx22671)
             ) ;
    mux21_ni ix64191 (.Y (nx64190), .A0 (inputs_258__15), .A1 (inputs_274__15), 
             .S0 (nx23105)) ;
    mux21_ni ix64203 (.Y (nx64202), .A0 (inputs_290__15), .A1 (inputs_306__15), 
             .S0 (nx23107)) ;
    mux21_ni ix64235 (.Y (nx64234), .A0 (nx64218), .A1 (nx64230), .S0 (nx22671)
             ) ;
    mux21_ni ix64219 (.Y (nx64218), .A0 (inputs_322__15), .A1 (inputs_338__15), 
             .S0 (nx23107)) ;
    mux21_ni ix64231 (.Y (nx64230), .A0 (inputs_354__15), .A1 (inputs_370__15), 
             .S0 (nx23107)) ;
    mux21_ni ix64299 (.Y (nx64298), .A0 (nx64266), .A1 (nx64294), .S0 (nx22523)
             ) ;
    mux21_ni ix64267 (.Y (nx64266), .A0 (nx64250), .A1 (nx64262), .S0 (nx22671)
             ) ;
    mux21_ni ix64251 (.Y (nx64250), .A0 (inputs_386__15), .A1 (inputs_402__15), 
             .S0 (nx23107)) ;
    mux21_ni ix64263 (.Y (nx64262), .A0 (inputs_418__15), .A1 (inputs_434__15), 
             .S0 (nx23107)) ;
    mux21_ni ix64295 (.Y (nx64294), .A0 (nx64278), .A1 (nx64290), .S0 (nx22671)
             ) ;
    mux21_ni ix64279 (.Y (nx64278), .A0 (inputs_450__15), .A1 (inputs_466__15), 
             .S0 (nx23107)) ;
    mux21_ni ix64291 (.Y (nx64290), .A0 (inputs_482__15), .A1 (inputs_498__15), 
             .S0 (nx23107)) ;
    mux21_ni ix66519 (.Y (nx66518), .A0 (nx65670), .A1 (nx66514), .S0 (nx22447)
             ) ;
    mux21_ni ix65671 (.Y (nx65670), .A0 (nx65246), .A1 (nx65666), .S0 (nx22523)
             ) ;
    mux21_ni ix65247 (.Y (nx65246), .A0 (nx65034), .A1 (nx65242), .S0 (nx22671)
             ) ;
    mux21_ni ix65035 (.Y (nx65034), .A0 (nx65028), .A1 (nx64950), .S0 (nx23187)
             ) ;
    oai21 ix65029 (.Y (nx65028), .A0 (nx22373), .A1 (nx21867), .B0 (nx21879)) ;
    mux21 ix21868 (.Y (nx21867), .A0 (nx64992), .A1 (nx65020), .S0 (nx23109)) ;
    mux21_ni ix64993 (.Y (nx64992), .A0 (nx64976), .A1 (nx64988), .S0 (nx23865)
             ) ;
    mux21_ni ix64977 (.Y (nx64976), .A0 (inputs_4__15), .A1 (inputs_5__15), .S0 (
             nx24807)) ;
    mux21_ni ix64989 (.Y (nx64988), .A0 (inputs_6__15), .A1 (inputs_7__15), .S0 (
             nx24809)) ;
    mux21_ni ix65021 (.Y (nx65020), .A0 (nx65004), .A1 (nx65016), .S0 (nx23865)
             ) ;
    mux21_ni ix65005 (.Y (nx65004), .A0 (inputs_20__15), .A1 (inputs_21__15), .S0 (
             nx24809)) ;
    mux21_ni ix65017 (.Y (nx65016), .A0 (inputs_22__15), .A1 (inputs_23__15), .S0 (
             nx24809)) ;
    nand04 ix21880 (.Y (nx21879), .A0 (nx22373), .A1 (nx23865), .A2 (nx24809), .A3 (
           nx64964)) ;
    mux21_ni ix64965 (.Y (nx64964), .A0 (inputs_3__15), .A1 (inputs_19__15), .S0 (
             nx23109)) ;
    mux21_ni ix64951 (.Y (nx64950), .A0 (nx64886), .A1 (nx64946), .S0 (nx23109)
             ) ;
    mux21_ni ix64887 (.Y (nx64886), .A0 (nx64854), .A1 (nx64882), .S0 (nx23331)
             ) ;
    mux21_ni ix64855 (.Y (nx64854), .A0 (nx64838), .A1 (nx64850), .S0 (nx23867)
             ) ;
    mux21_ni ix64839 (.Y (nx64838), .A0 (inputs_8__15), .A1 (inputs_9__15), .S0 (
             nx24809)) ;
    mux21_ni ix64851 (.Y (nx64850), .A0 (inputs_10__15), .A1 (inputs_11__15), .S0 (
             nx24809)) ;
    mux21_ni ix64883 (.Y (nx64882), .A0 (nx64866), .A1 (nx64878), .S0 (nx23867)
             ) ;
    mux21_ni ix64867 (.Y (nx64866), .A0 (inputs_12__15), .A1 (inputs_13__15), .S0 (
             nx24809)) ;
    mux21_ni ix64879 (.Y (nx64878), .A0 (inputs_14__15), .A1 (inputs_15__15), .S0 (
             nx24811)) ;
    mux21_ni ix64947 (.Y (nx64946), .A0 (nx64914), .A1 (nx64942), .S0 (nx23333)
             ) ;
    mux21_ni ix64915 (.Y (nx64914), .A0 (nx64898), .A1 (nx64910), .S0 (nx23867)
             ) ;
    mux21_ni ix64899 (.Y (nx64898), .A0 (inputs_24__15), .A1 (inputs_25__15), .S0 (
             nx24811)) ;
    mux21_ni ix64911 (.Y (nx64910), .A0 (inputs_26__15), .A1 (inputs_27__15), .S0 (
             nx24811)) ;
    mux21_ni ix64943 (.Y (nx64942), .A0 (nx64926), .A1 (nx64938), .S0 (nx23867)
             ) ;
    mux21_ni ix64927 (.Y (nx64926), .A0 (inputs_28__15), .A1 (inputs_29__15), .S0 (
             nx24811)) ;
    mux21_ni ix64939 (.Y (nx64938), .A0 (inputs_30__15), .A1 (inputs_31__15), .S0 (
             nx24811)) ;
    mux21_ni ix65243 (.Y (nx65242), .A0 (nx65236), .A1 (nx65158), .S0 (nx23187)
             ) ;
    oai21 ix65237 (.Y (nx65236), .A0 (nx22373), .A1 (nx21911), .B0 (nx21923)) ;
    mux21 ix21912 (.Y (nx21911), .A0 (nx65200), .A1 (nx65228), .S0 (nx23109)) ;
    mux21_ni ix65201 (.Y (nx65200), .A0 (nx65184), .A1 (nx65196), .S0 (nx23867)
             ) ;
    mux21_ni ix65185 (.Y (nx65184), .A0 (inputs_36__15), .A1 (inputs_37__15), .S0 (
             nx24811)) ;
    mux21_ni ix65197 (.Y (nx65196), .A0 (inputs_38__15), .A1 (inputs_39__15), .S0 (
             nx24811)) ;
    mux21_ni ix65229 (.Y (nx65228), .A0 (nx65212), .A1 (nx65224), .S0 (nx23867)
             ) ;
    mux21_ni ix65213 (.Y (nx65212), .A0 (inputs_52__15), .A1 (inputs_53__15), .S0 (
             nx24813)) ;
    mux21_ni ix65225 (.Y (nx65224), .A0 (inputs_54__15), .A1 (inputs_55__15), .S0 (
             nx24813)) ;
    nand04 ix21924 (.Y (nx21923), .A0 (nx22373), .A1 (nx23867), .A2 (nx24813), .A3 (
           nx65172)) ;
    mux21_ni ix65173 (.Y (nx65172), .A0 (inputs_35__15), .A1 (inputs_51__15), .S0 (
             nx23109)) ;
    mux21_ni ix65159 (.Y (nx65158), .A0 (nx65094), .A1 (nx65154), .S0 (nx23109)
             ) ;
    mux21_ni ix65095 (.Y (nx65094), .A0 (nx65062), .A1 (nx65090), .S0 (nx23333)
             ) ;
    mux21_ni ix65063 (.Y (nx65062), .A0 (nx65046), .A1 (nx65058), .S0 (nx23869)
             ) ;
    mux21_ni ix65047 (.Y (nx65046), .A0 (inputs_40__15), .A1 (inputs_41__15), .S0 (
             nx24813)) ;
    mux21_ni ix65059 (.Y (nx65058), .A0 (inputs_42__15), .A1 (inputs_43__15), .S0 (
             nx24813)) ;
    mux21_ni ix65091 (.Y (nx65090), .A0 (nx65074), .A1 (nx65086), .S0 (nx23869)
             ) ;
    mux21_ni ix65075 (.Y (nx65074), .A0 (inputs_44__15), .A1 (inputs_45__15), .S0 (
             nx24813)) ;
    mux21_ni ix65087 (.Y (nx65086), .A0 (inputs_46__15), .A1 (inputs_47__15), .S0 (
             nx24813)) ;
    mux21_ni ix65155 (.Y (nx65154), .A0 (nx65122), .A1 (nx65150), .S0 (nx23333)
             ) ;
    mux21_ni ix65123 (.Y (nx65122), .A0 (nx65106), .A1 (nx65118), .S0 (nx23869)
             ) ;
    mux21_ni ix65107 (.Y (nx65106), .A0 (inputs_56__15), .A1 (inputs_57__15), .S0 (
             nx24815)) ;
    mux21_ni ix65119 (.Y (nx65118), .A0 (inputs_58__15), .A1 (inputs_59__15), .S0 (
             nx24815)) ;
    mux21_ni ix65151 (.Y (nx65150), .A0 (nx65134), .A1 (nx65146), .S0 (nx23869)
             ) ;
    mux21_ni ix65135 (.Y (nx65134), .A0 (inputs_60__15), .A1 (inputs_61__15), .S0 (
             nx24815)) ;
    mux21_ni ix65147 (.Y (nx65146), .A0 (inputs_62__15), .A1 (inputs_63__15), .S0 (
             nx24815)) ;
    mux21_ni ix65667 (.Y (nx65666), .A0 (nx65454), .A1 (nx65662), .S0 (nx22671)
             ) ;
    mux21_ni ix65455 (.Y (nx65454), .A0 (nx65448), .A1 (nx65370), .S0 (nx23187)
             ) ;
    oai21 ix65449 (.Y (nx65448), .A0 (nx22373), .A1 (nx21955), .B0 (nx21967)) ;
    mux21 ix21956 (.Y (nx21955), .A0 (nx65412), .A1 (nx65440), .S0 (nx23109)) ;
    mux21_ni ix65413 (.Y (nx65412), .A0 (nx65396), .A1 (nx65408), .S0 (nx23869)
             ) ;
    mux21_ni ix65397 (.Y (nx65396), .A0 (inputs_68__15), .A1 (inputs_69__15), .S0 (
             nx24815)) ;
    mux21_ni ix65409 (.Y (nx65408), .A0 (inputs_70__15), .A1 (inputs_71__15), .S0 (
             nx24815)) ;
    mux21_ni ix65441 (.Y (nx65440), .A0 (nx65424), .A1 (nx65436), .S0 (nx23869)
             ) ;
    mux21_ni ix65425 (.Y (nx65424), .A0 (inputs_84__15), .A1 (inputs_85__15), .S0 (
             nx24815)) ;
    mux21_ni ix65437 (.Y (nx65436), .A0 (inputs_86__15), .A1 (inputs_87__15), .S0 (
             nx24817)) ;
    nand04 ix21968 (.Y (nx21967), .A0 (nx22373), .A1 (nx23869), .A2 (nx24817), .A3 (
           nx65384)) ;
    mux21_ni ix65385 (.Y (nx65384), .A0 (inputs_67__15), .A1 (inputs_83__15), .S0 (
             nx23111)) ;
    mux21_ni ix65371 (.Y (nx65370), .A0 (nx65306), .A1 (nx65366), .S0 (nx23111)
             ) ;
    mux21_ni ix65307 (.Y (nx65306), .A0 (nx65274), .A1 (nx65302), .S0 (nx23333)
             ) ;
    mux21_ni ix65275 (.Y (nx65274), .A0 (nx65258), .A1 (nx65270), .S0 (nx23871)
             ) ;
    mux21_ni ix65259 (.Y (nx65258), .A0 (inputs_72__15), .A1 (inputs_73__15), .S0 (
             nx24817)) ;
    mux21_ni ix65271 (.Y (nx65270), .A0 (inputs_74__15), .A1 (inputs_75__15), .S0 (
             nx24817)) ;
    mux21_ni ix65303 (.Y (nx65302), .A0 (nx65286), .A1 (nx65298), .S0 (nx23871)
             ) ;
    mux21_ni ix65287 (.Y (nx65286), .A0 (inputs_76__15), .A1 (inputs_77__15), .S0 (
             nx24817)) ;
    mux21_ni ix65299 (.Y (nx65298), .A0 (inputs_78__15), .A1 (inputs_79__15), .S0 (
             nx24817)) ;
    mux21_ni ix65367 (.Y (nx65366), .A0 (nx65334), .A1 (nx65362), .S0 (nx23333)
             ) ;
    mux21_ni ix65335 (.Y (nx65334), .A0 (nx65318), .A1 (nx65330), .S0 (nx23871)
             ) ;
    mux21_ni ix65319 (.Y (nx65318), .A0 (inputs_88__15), .A1 (inputs_89__15), .S0 (
             nx24817)) ;
    mux21_ni ix65331 (.Y (nx65330), .A0 (inputs_90__15), .A1 (inputs_91__15), .S0 (
             nx24819)) ;
    mux21_ni ix65363 (.Y (nx65362), .A0 (nx65346), .A1 (nx65358), .S0 (nx23871)
             ) ;
    mux21_ni ix65347 (.Y (nx65346), .A0 (inputs_92__15), .A1 (inputs_93__15), .S0 (
             nx24819)) ;
    mux21_ni ix65359 (.Y (nx65358), .A0 (inputs_94__15), .A1 (inputs_95__15), .S0 (
             nx24819)) ;
    mux21_ni ix65663 (.Y (nx65662), .A0 (nx65656), .A1 (nx65578), .S0 (nx23187)
             ) ;
    oai21 ix65657 (.Y (nx65656), .A0 (nx22375), .A1 (nx21997), .B0 (nx22009)) ;
    mux21 ix21998 (.Y (nx21997), .A0 (nx65620), .A1 (nx65648), .S0 (nx23111)) ;
    mux21_ni ix65621 (.Y (nx65620), .A0 (nx65604), .A1 (nx65616), .S0 (nx23871)
             ) ;
    mux21_ni ix65605 (.Y (nx65604), .A0 (inputs_100__15), .A1 (inputs_101__15), 
             .S0 (nx24819)) ;
    mux21_ni ix65617 (.Y (nx65616), .A0 (inputs_102__15), .A1 (inputs_103__15), 
             .S0 (nx24819)) ;
    mux21_ni ix65649 (.Y (nx65648), .A0 (nx65632), .A1 (nx65644), .S0 (nx23871)
             ) ;
    mux21_ni ix65633 (.Y (nx65632), .A0 (inputs_116__15), .A1 (inputs_117__15), 
             .S0 (nx24819)) ;
    mux21_ni ix65645 (.Y (nx65644), .A0 (inputs_118__15), .A1 (inputs_119__15), 
             .S0 (nx24819)) ;
    nand04 ix22010 (.Y (nx22009), .A0 (nx22375), .A1 (nx23871), .A2 (nx24821), .A3 (
           nx65592)) ;
    mux21_ni ix65593 (.Y (nx65592), .A0 (inputs_99__15), .A1 (inputs_115__15), .S0 (
             nx23111)) ;
    mux21_ni ix65579 (.Y (nx65578), .A0 (nx65514), .A1 (nx65574), .S0 (nx23111)
             ) ;
    mux21_ni ix65515 (.Y (nx65514), .A0 (nx65482), .A1 (nx65510), .S0 (nx23333)
             ) ;
    mux21_ni ix65483 (.Y (nx65482), .A0 (nx65466), .A1 (nx65478), .S0 (nx23873)
             ) ;
    mux21_ni ix65467 (.Y (nx65466), .A0 (inputs_104__15), .A1 (inputs_105__15), 
             .S0 (nx24821)) ;
    mux21_ni ix65479 (.Y (nx65478), .A0 (inputs_106__15), .A1 (inputs_107__15), 
             .S0 (nx24821)) ;
    mux21_ni ix65511 (.Y (nx65510), .A0 (nx65494), .A1 (nx65506), .S0 (nx23873)
             ) ;
    mux21_ni ix65495 (.Y (nx65494), .A0 (inputs_108__15), .A1 (inputs_109__15), 
             .S0 (nx24821)) ;
    mux21_ni ix65507 (.Y (nx65506), .A0 (inputs_110__15), .A1 (inputs_111__15), 
             .S0 (nx24821)) ;
    mux21_ni ix65575 (.Y (nx65574), .A0 (nx65542), .A1 (nx65570), .S0 (nx23333)
             ) ;
    mux21_ni ix65543 (.Y (nx65542), .A0 (nx65526), .A1 (nx65538), .S0 (nx23873)
             ) ;
    mux21_ni ix65527 (.Y (nx65526), .A0 (inputs_120__15), .A1 (inputs_121__15), 
             .S0 (nx24821)) ;
    mux21_ni ix65539 (.Y (nx65538), .A0 (inputs_122__15), .A1 (inputs_123__15), 
             .S0 (nx24821)) ;
    mux21_ni ix65571 (.Y (nx65570), .A0 (nx65554), .A1 (nx65566), .S0 (nx23873)
             ) ;
    mux21_ni ix65555 (.Y (nx65554), .A0 (inputs_124__15), .A1 (inputs_125__15), 
             .S0 (nx24823)) ;
    mux21_ni ix65567 (.Y (nx65566), .A0 (inputs_126__15), .A1 (inputs_127__15), 
             .S0 (nx24823)) ;
    mux21_ni ix66515 (.Y (nx66514), .A0 (nx66090), .A1 (nx66510), .S0 (nx22523)
             ) ;
    mux21_ni ix66091 (.Y (nx66090), .A0 (nx65878), .A1 (nx66086), .S0 (nx22671)
             ) ;
    mux21_ni ix65879 (.Y (nx65878), .A0 (nx65872), .A1 (nx65794), .S0 (nx23189)
             ) ;
    oai21 ix65873 (.Y (nx65872), .A0 (nx22375), .A1 (nx22045), .B0 (nx22057)) ;
    mux21 ix22046 (.Y (nx22045), .A0 (nx65836), .A1 (nx65864), .S0 (nx23111)) ;
    mux21_ni ix65837 (.Y (nx65836), .A0 (nx65820), .A1 (nx65832), .S0 (nx23873)
             ) ;
    mux21_ni ix65821 (.Y (nx65820), .A0 (inputs_132__15), .A1 (inputs_133__15), 
             .S0 (nx24823)) ;
    mux21_ni ix65833 (.Y (nx65832), .A0 (inputs_134__15), .A1 (inputs_135__15), 
             .S0 (nx24823)) ;
    mux21_ni ix65865 (.Y (nx65864), .A0 (nx65848), .A1 (nx65860), .S0 (nx23873)
             ) ;
    mux21_ni ix65849 (.Y (nx65848), .A0 (inputs_148__15), .A1 (inputs_149__15), 
             .S0 (nx24823)) ;
    mux21_ni ix65861 (.Y (nx65860), .A0 (inputs_150__15), .A1 (inputs_151__15), 
             .S0 (nx24823)) ;
    nand04 ix22058 (.Y (nx22057), .A0 (nx22375), .A1 (nx23873), .A2 (nx24823), .A3 (
           nx65808)) ;
    mux21_ni ix65809 (.Y (nx65808), .A0 (inputs_131__15), .A1 (inputs_147__15), 
             .S0 (nx23111)) ;
    mux21_ni ix65795 (.Y (nx65794), .A0 (nx65730), .A1 (nx65790), .S0 (nx23113)
             ) ;
    mux21_ni ix65731 (.Y (nx65730), .A0 (nx65698), .A1 (nx65726), .S0 (nx23335)
             ) ;
    mux21_ni ix65699 (.Y (nx65698), .A0 (nx65682), .A1 (nx65694), .S0 (nx23875)
             ) ;
    mux21_ni ix65683 (.Y (nx65682), .A0 (inputs_136__15), .A1 (inputs_137__15), 
             .S0 (nx24825)) ;
    mux21_ni ix65695 (.Y (nx65694), .A0 (inputs_138__15), .A1 (inputs_139__15), 
             .S0 (nx24825)) ;
    mux21_ni ix65727 (.Y (nx65726), .A0 (nx65710), .A1 (nx65722), .S0 (nx23875)
             ) ;
    mux21_ni ix65711 (.Y (nx65710), .A0 (inputs_140__15), .A1 (inputs_141__15), 
             .S0 (nx24825)) ;
    mux21_ni ix65723 (.Y (nx65722), .A0 (inputs_142__15), .A1 (inputs_143__15), 
             .S0 (nx24825)) ;
    mux21_ni ix65791 (.Y (nx65790), .A0 (nx65758), .A1 (nx65786), .S0 (nx23335)
             ) ;
    mux21_ni ix65759 (.Y (nx65758), .A0 (nx65742), .A1 (nx65754), .S0 (nx23875)
             ) ;
    mux21_ni ix65743 (.Y (nx65742), .A0 (inputs_152__15), .A1 (inputs_153__15), 
             .S0 (nx24825)) ;
    mux21_ni ix65755 (.Y (nx65754), .A0 (inputs_154__15), .A1 (inputs_155__15), 
             .S0 (nx24825)) ;
    mux21_ni ix65787 (.Y (nx65786), .A0 (nx65770), .A1 (nx65782), .S0 (nx23875)
             ) ;
    mux21_ni ix65771 (.Y (nx65770), .A0 (inputs_156__15), .A1 (inputs_157__15), 
             .S0 (nx24825)) ;
    mux21_ni ix65783 (.Y (nx65782), .A0 (inputs_158__15), .A1 (inputs_159__15), 
             .S0 (nx24827)) ;
    mux21_ni ix66087 (.Y (nx66086), .A0 (nx66080), .A1 (nx66002), .S0 (nx23189)
             ) ;
    oai21 ix66081 (.Y (nx66080), .A0 (nx22375), .A1 (nx22087), .B0 (nx22097)) ;
    mux21 ix22088 (.Y (nx22087), .A0 (nx66044), .A1 (nx66072), .S0 (nx23113)) ;
    mux21_ni ix66045 (.Y (nx66044), .A0 (nx66028), .A1 (nx66040), .S0 (nx23875)
             ) ;
    mux21_ni ix66029 (.Y (nx66028), .A0 (inputs_164__15), .A1 (inputs_165__15), 
             .S0 (nx24827)) ;
    mux21_ni ix66041 (.Y (nx66040), .A0 (inputs_166__15), .A1 (inputs_167__15), 
             .S0 (nx24827)) ;
    mux21_ni ix66073 (.Y (nx66072), .A0 (nx66056), .A1 (nx66068), .S0 (nx23875)
             ) ;
    mux21_ni ix66057 (.Y (nx66056), .A0 (inputs_180__15), .A1 (inputs_181__15), 
             .S0 (nx24827)) ;
    mux21_ni ix66069 (.Y (nx66068), .A0 (inputs_182__15), .A1 (inputs_183__15), 
             .S0 (nx24827)) ;
    nand04 ix22098 (.Y (nx22097), .A0 (nx22375), .A1 (nx23875), .A2 (nx24827), .A3 (
           nx66016)) ;
    mux21_ni ix66017 (.Y (nx66016), .A0 (inputs_163__15), .A1 (inputs_179__15), 
             .S0 (nx23113)) ;
    mux21_ni ix66003 (.Y (nx66002), .A0 (nx65938), .A1 (nx65998), .S0 (nx23113)
             ) ;
    mux21_ni ix65939 (.Y (nx65938), .A0 (nx65906), .A1 (nx65934), .S0 (nx23335)
             ) ;
    mux21_ni ix65907 (.Y (nx65906), .A0 (nx65890), .A1 (nx65902), .S0 (nx23877)
             ) ;
    mux21_ni ix65891 (.Y (nx65890), .A0 (inputs_168__15), .A1 (inputs_169__15), 
             .S0 (nx24827)) ;
    mux21_ni ix65903 (.Y (nx65902), .A0 (inputs_170__15), .A1 (inputs_171__15), 
             .S0 (nx24829)) ;
    mux21_ni ix65935 (.Y (nx65934), .A0 (nx65918), .A1 (nx65930), .S0 (nx23877)
             ) ;
    mux21_ni ix65919 (.Y (nx65918), .A0 (inputs_172__15), .A1 (inputs_173__15), 
             .S0 (nx24829)) ;
    mux21_ni ix65931 (.Y (nx65930), .A0 (inputs_174__15), .A1 (inputs_175__15), 
             .S0 (nx24829)) ;
    mux21_ni ix65999 (.Y (nx65998), .A0 (nx65966), .A1 (nx65994), .S0 (nx23335)
             ) ;
    mux21_ni ix65967 (.Y (nx65966), .A0 (nx65950), .A1 (nx65962), .S0 (nx23877)
             ) ;
    mux21_ni ix65951 (.Y (nx65950), .A0 (inputs_184__15), .A1 (inputs_185__15), 
             .S0 (nx24829)) ;
    mux21_ni ix65963 (.Y (nx65962), .A0 (inputs_186__15), .A1 (inputs_187__15), 
             .S0 (nx24829)) ;
    mux21_ni ix65995 (.Y (nx65994), .A0 (nx65978), .A1 (nx65990), .S0 (nx23877)
             ) ;
    mux21_ni ix65979 (.Y (nx65978), .A0 (inputs_188__15), .A1 (inputs_189__15), 
             .S0 (nx24829)) ;
    mux21_ni ix65991 (.Y (nx65990), .A0 (inputs_190__15), .A1 (inputs_191__15), 
             .S0 (nx24829)) ;
    mux21_ni ix66511 (.Y (nx66510), .A0 (nx66298), .A1 (nx66506), .S0 (nx22673)
             ) ;
    mux21_ni ix66299 (.Y (nx66298), .A0 (nx66292), .A1 (nx66214), .S0 (nx23189)
             ) ;
    oai21 ix66293 (.Y (nx66292), .A0 (nx22375), .A1 (nx22129), .B0 (nx22141)) ;
    mux21 ix22130 (.Y (nx22129), .A0 (nx66256), .A1 (nx66284), .S0 (nx23113)) ;
    mux21_ni ix66257 (.Y (nx66256), .A0 (nx66240), .A1 (nx66252), .S0 (nx23877)
             ) ;
    mux21_ni ix66241 (.Y (nx66240), .A0 (inputs_196__15), .A1 (inputs_197__15), 
             .S0 (nx24831)) ;
    mux21_ni ix66253 (.Y (nx66252), .A0 (inputs_198__15), .A1 (inputs_199__15), 
             .S0 (nx24831)) ;
    mux21_ni ix66285 (.Y (nx66284), .A0 (nx66268), .A1 (nx66280), .S0 (nx23877)
             ) ;
    mux21_ni ix66269 (.Y (nx66268), .A0 (inputs_212__15), .A1 (inputs_213__15), 
             .S0 (nx24831)) ;
    mux21_ni ix66281 (.Y (nx66280), .A0 (inputs_214__15), .A1 (inputs_215__15), 
             .S0 (nx24831)) ;
    nand04 ix22142 (.Y (nx22141), .A0 (nx22377), .A1 (nx23877), .A2 (nx24831), .A3 (
           nx66228)) ;
    mux21_ni ix66229 (.Y (nx66228), .A0 (inputs_195__15), .A1 (inputs_211__15), 
             .S0 (nx23113)) ;
    mux21_ni ix66215 (.Y (nx66214), .A0 (nx66150), .A1 (nx66210), .S0 (nx23113)
             ) ;
    mux21_ni ix66151 (.Y (nx66150), .A0 (nx66118), .A1 (nx66146), .S0 (nx23335)
             ) ;
    mux21_ni ix66119 (.Y (nx66118), .A0 (nx66102), .A1 (nx66114), .S0 (nx23879)
             ) ;
    mux21_ni ix66103 (.Y (nx66102), .A0 (inputs_200__15), .A1 (inputs_201__15), 
             .S0 (nx24831)) ;
    mux21_ni ix66115 (.Y (nx66114), .A0 (inputs_202__15), .A1 (inputs_203__15), 
             .S0 (nx24831)) ;
    mux21_ni ix66147 (.Y (nx66146), .A0 (nx66130), .A1 (nx66142), .S0 (nx23879)
             ) ;
    mux21_ni ix66131 (.Y (nx66130), .A0 (inputs_204__15), .A1 (inputs_205__15), 
             .S0 (nx24833)) ;
    mux21_ni ix66143 (.Y (nx66142), .A0 (inputs_206__15), .A1 (inputs_207__15), 
             .S0 (nx24833)) ;
    mux21_ni ix66211 (.Y (nx66210), .A0 (nx66178), .A1 (nx66206), .S0 (nx23335)
             ) ;
    mux21_ni ix66179 (.Y (nx66178), .A0 (nx66162), .A1 (nx66174), .S0 (nx23879)
             ) ;
    mux21_ni ix66163 (.Y (nx66162), .A0 (inputs_216__15), .A1 (inputs_217__15), 
             .S0 (nx24833)) ;
    mux21_ni ix66175 (.Y (nx66174), .A0 (inputs_218__15), .A1 (inputs_219__15), 
             .S0 (nx24833)) ;
    mux21_ni ix66207 (.Y (nx66206), .A0 (nx66190), .A1 (nx66202), .S0 (nx23879)
             ) ;
    mux21_ni ix66191 (.Y (nx66190), .A0 (inputs_220__15), .A1 (inputs_221__15), 
             .S0 (nx24833)) ;
    mux21_ni ix66203 (.Y (nx66202), .A0 (inputs_222__15), .A1 (inputs_223__15), 
             .S0 (nx24833)) ;
    mux21_ni ix66507 (.Y (nx66506), .A0 (nx66500), .A1 (nx66422), .S0 (nx23189)
             ) ;
    oai21 ix66501 (.Y (nx66500), .A0 (nx22377), .A1 (nx22173), .B0 (nx22183)) ;
    mux21 ix22174 (.Y (nx22173), .A0 (nx66464), .A1 (nx66492), .S0 (nx23115)) ;
    mux21_ni ix66465 (.Y (nx66464), .A0 (nx66448), .A1 (nx66460), .S0 (nx23879)
             ) ;
    mux21_ni ix66449 (.Y (nx66448), .A0 (inputs_228__15), .A1 (inputs_229__15), 
             .S0 (nx24833)) ;
    mux21_ni ix66461 (.Y (nx66460), .A0 (inputs_230__15), .A1 (inputs_231__15), 
             .S0 (nx24835)) ;
    mux21_ni ix66493 (.Y (nx66492), .A0 (nx66476), .A1 (nx66488), .S0 (nx23879)
             ) ;
    mux21_ni ix66477 (.Y (nx66476), .A0 (inputs_244__15), .A1 (inputs_245__15), 
             .S0 (nx24835)) ;
    mux21_ni ix66489 (.Y (nx66488), .A0 (inputs_246__15), .A1 (inputs_247__15), 
             .S0 (nx24835)) ;
    nand04 ix22184 (.Y (nx22183), .A0 (nx22377), .A1 (nx23879), .A2 (nx24835), .A3 (
           nx66436)) ;
    mux21_ni ix66437 (.Y (nx66436), .A0 (inputs_227__15), .A1 (inputs_243__15), 
             .S0 (nx23115)) ;
    mux21_ni ix66423 (.Y (nx66422), .A0 (nx66358), .A1 (nx66418), .S0 (nx23115)
             ) ;
    mux21_ni ix66359 (.Y (nx66358), .A0 (nx66326), .A1 (nx66354), .S0 (nx23335)
             ) ;
    mux21_ni ix66327 (.Y (nx66326), .A0 (nx66310), .A1 (nx66322), .S0 (nx23881)
             ) ;
    mux21_ni ix66311 (.Y (nx66310), .A0 (inputs_232__15), .A1 (inputs_233__15), 
             .S0 (nx24835)) ;
    mux21_ni ix66323 (.Y (nx66322), .A0 (inputs_234__15), .A1 (inputs_235__15), 
             .S0 (nx24835)) ;
    mux21_ni ix66355 (.Y (nx66354), .A0 (nx66338), .A1 (nx66350), .S0 (nx23881)
             ) ;
    mux21_ni ix66339 (.Y (nx66338), .A0 (inputs_236__15), .A1 (inputs_237__15), 
             .S0 (nx24835)) ;
    mux21_ni ix66351 (.Y (nx66350), .A0 (inputs_238__15), .A1 (inputs_239__15), 
             .S0 (nx24837)) ;
    mux21_ni ix66419 (.Y (nx66418), .A0 (nx66386), .A1 (nx66414), .S0 (nx23337)
             ) ;
    mux21_ni ix66387 (.Y (nx66386), .A0 (nx66370), .A1 (nx66382), .S0 (nx23881)
             ) ;
    mux21_ni ix66371 (.Y (nx66370), .A0 (inputs_248__15), .A1 (inputs_249__15), 
             .S0 (nx24837)) ;
    mux21_ni ix66383 (.Y (nx66382), .A0 (inputs_250__15), .A1 (inputs_251__15), 
             .S0 (nx24837)) ;
    mux21_ni ix66415 (.Y (nx66414), .A0 (nx66398), .A1 (nx66410), .S0 (nx23881)
             ) ;
    mux21_ni ix66399 (.Y (nx66398), .A0 (inputs_252__15), .A1 (inputs_253__15), 
             .S0 (nx24837)) ;
    mux21_ni ix66411 (.Y (nx66410), .A0 (inputs_254__15), .A1 (inputs_255__15), 
             .S0 (nx24837)) ;
    inv02 ix22216 (.Y (nx22217), .A (selectionLines[8])) ;
    inv02 ix22218 (.Y (nx22219), .A (nx22405)) ;
    inv02 ix22220 (.Y (nx22221), .A (nx22407)) ;
    inv02 ix22222 (.Y (nx22223), .A (nx22407)) ;
    inv02 ix22224 (.Y (nx22225), .A (nx22407)) ;
    inv02 ix22226 (.Y (nx22227), .A (selectionLines[2])) ;
    inv02 ix22228 (.Y (nx22229), .A (nx23337)) ;
    inv02 ix22230 (.Y (nx22231), .A (nx23337)) ;
    inv02 ix22232 (.Y (nx22233), .A (nx23337)) ;
    inv02 ix22234 (.Y (nx22235), .A (nx23337)) ;
    inv02 ix22236 (.Y (nx22237), .A (nx23337)) ;
    inv02 ix22238 (.Y (nx22239), .A (nx23337)) ;
    inv02 ix22240 (.Y (nx22241), .A (nx23339)) ;
    inv02 ix22242 (.Y (nx22243), .A (nx23339)) ;
    inv02 ix22244 (.Y (nx22245), .A (nx23339)) ;
    inv02 ix22246 (.Y (nx22247), .A (nx23339)) ;
    inv02 ix22248 (.Y (nx22249), .A (nx23339)) ;
    inv02 ix22250 (.Y (nx22251), .A (nx23339)) ;
    inv02 ix22252 (.Y (nx22253), .A (nx23339)) ;
    inv02 ix22254 (.Y (nx22255), .A (nx23341)) ;
    inv02 ix22256 (.Y (nx22257), .A (nx23341)) ;
    inv02 ix22258 (.Y (nx22259), .A (nx23341)) ;
    inv02 ix22260 (.Y (nx22261), .A (nx23341)) ;
    inv02 ix22262 (.Y (nx22263), .A (nx23341)) ;
    inv02 ix22264 (.Y (nx22265), .A (nx23341)) ;
    inv02 ix22266 (.Y (nx22267), .A (nx23341)) ;
    inv02 ix22268 (.Y (nx22269), .A (nx23343)) ;
    inv02 ix22270 (.Y (nx22271), .A (nx23343)) ;
    inv02 ix22272 (.Y (nx22273), .A (nx23343)) ;
    inv02 ix22274 (.Y (nx22275), .A (nx23343)) ;
    inv02 ix22276 (.Y (nx22277), .A (nx23343)) ;
    inv02 ix22278 (.Y (nx22279), .A (nx23343)) ;
    inv02 ix22280 (.Y (nx22281), .A (nx23343)) ;
    inv02 ix22282 (.Y (nx22283), .A (nx23345)) ;
    inv02 ix22284 (.Y (nx22285), .A (nx23345)) ;
    inv02 ix22286 (.Y (nx22287), .A (nx23345)) ;
    inv02 ix22288 (.Y (nx22289), .A (nx23345)) ;
    inv02 ix22290 (.Y (nx22291), .A (nx23345)) ;
    inv02 ix22292 (.Y (nx22293), .A (nx23345)) ;
    inv02 ix22294 (.Y (nx22295), .A (nx23345)) ;
    inv02 ix22296 (.Y (nx22297), .A (nx23347)) ;
    inv02 ix22298 (.Y (nx22299), .A (nx23347)) ;
    inv02 ix22300 (.Y (nx22301), .A (nx23347)) ;
    inv02 ix22302 (.Y (nx22303), .A (nx23347)) ;
    inv02 ix22304 (.Y (nx22305), .A (nx23347)) ;
    inv02 ix22306 (.Y (nx22307), .A (nx23347)) ;
    inv02 ix22308 (.Y (nx22309), .A (nx23347)) ;
    inv02 ix22310 (.Y (nx22311), .A (nx23349)) ;
    inv02 ix22312 (.Y (nx22313), .A (nx23349)) ;
    inv02 ix22314 (.Y (nx22315), .A (nx23349)) ;
    inv02 ix22316 (.Y (nx22317), .A (nx23349)) ;
    inv02 ix22318 (.Y (nx22319), .A (nx23349)) ;
    inv02 ix22320 (.Y (nx22321), .A (nx23349)) ;
    inv02 ix22322 (.Y (nx22323), .A (nx23349)) ;
    inv02 ix22324 (.Y (nx22325), .A (nx23351)) ;
    inv02 ix22326 (.Y (nx22327), .A (nx23351)) ;
    inv02 ix22328 (.Y (nx22329), .A (nx23351)) ;
    inv02 ix22330 (.Y (nx22331), .A (nx23351)) ;
    inv02 ix22332 (.Y (nx22333), .A (nx23351)) ;
    inv02 ix22334 (.Y (nx22335), .A (nx23351)) ;
    inv02 ix22336 (.Y (nx22337), .A (nx23351)) ;
    inv02 ix22338 (.Y (nx22339), .A (nx23353)) ;
    inv02 ix22340 (.Y (nx22341), .A (nx23353)) ;
    inv02 ix22342 (.Y (nx22343), .A (nx23353)) ;
    inv02 ix22344 (.Y (nx22345), .A (nx23353)) ;
    inv02 ix22346 (.Y (nx22347), .A (nx23353)) ;
    inv02 ix22348 (.Y (nx22349), .A (nx23353)) ;
    inv02 ix22350 (.Y (nx22351), .A (nx23353)) ;
    inv02 ix22352 (.Y (nx22353), .A (nx23355)) ;
    inv02 ix22354 (.Y (nx22355), .A (nx23355)) ;
    inv02 ix22356 (.Y (nx22357), .A (nx23355)) ;
    inv02 ix22358 (.Y (nx22359), .A (nx23355)) ;
    inv02 ix22360 (.Y (nx22361), .A (nx23355)) ;
    inv02 ix22362 (.Y (nx22363), .A (nx23355)) ;
    inv02 ix22364 (.Y (nx22365), .A (nx23355)) ;
    inv02 ix22366 (.Y (nx22367), .A (nx23357)) ;
    inv02 ix22368 (.Y (nx22369), .A (nx23357)) ;
    inv02 ix22370 (.Y (nx22371), .A (nx23357)) ;
    inv02 ix22372 (.Y (nx22373), .A (nx23357)) ;
    inv02 ix22374 (.Y (nx22375), .A (nx23357)) ;
    inv02 ix22376 (.Y (nx22377), .A (nx23357)) ;
    inv02 ix22378 (.Y (nx22379), .A (selectionLines[0])) ;
    inv02 ix22380 (.Y (nx22381), .A (nx24837)) ;
    inv02 ix22382 (.Y (nx22383), .A (nx24837)) ;
    inv01 ix22384 (.Y (nx22385), .A (nx23189)) ;
    inv01 ix22386 (.Y (nx22387), .A (nx23189)) ;
    inv02 ix22392 (.Y (nx22393), .A (nx24853)) ;
    inv02 ix22394 (.Y (nx22395), .A (nx24853)) ;
    inv02 ix22396 (.Y (nx22397), .A (nx24853)) ;
    inv02 ix22398 (.Y (nx22399), .A (nx24853)) ;
    inv02 ix22400 (.Y (nx22401), .A (nx24853)) ;
    inv02 ix22402 (.Y (nx22403), .A (nx24853)) ;
    inv02 ix22404 (.Y (nx22405), .A (nx24853)) ;
    inv02 ix22406 (.Y (nx22407), .A (nx22217)) ;
    inv02 ix22410 (.Y (nx22411), .A (nx25017)) ;
    inv02 ix22412 (.Y (nx22413), .A (nx25017)) ;
    inv02 ix22414 (.Y (nx22415), .A (nx25017)) ;
    inv02 ix22416 (.Y (nx22417), .A (nx25017)) ;
    inv02 ix22418 (.Y (nx22419), .A (nx25017)) ;
    inv02 ix22420 (.Y (nx22421), .A (nx25017)) ;
    inv02 ix22422 (.Y (nx22423), .A (nx25017)) ;
    inv02 ix22424 (.Y (nx22425), .A (nx25019)) ;
    inv02 ix22426 (.Y (nx22427), .A (nx25019)) ;
    inv02 ix22428 (.Y (nx22429), .A (nx25019)) ;
    inv02 ix22430 (.Y (nx22431), .A (nx25019)) ;
    inv02 ix22432 (.Y (nx22433), .A (nx25019)) ;
    inv02 ix22434 (.Y (nx22435), .A (nx25019)) ;
    inv02 ix22436 (.Y (nx22437), .A (nx25019)) ;
    inv02 ix22438 (.Y (nx22439), .A (nx25021)) ;
    inv02 ix22440 (.Y (nx22441), .A (nx25021)) ;
    inv02 ix22442 (.Y (nx22443), .A (nx25021)) ;
    inv02 ix22444 (.Y (nx22445), .A (nx25021)) ;
    inv02 ix22446 (.Y (nx22447), .A (nx25021)) ;
    inv02 ix22450 (.Y (nx22451), .A (nx25023)) ;
    inv02 ix22452 (.Y (nx22453), .A (nx25023)) ;
    inv02 ix22454 (.Y (nx22455), .A (nx25023)) ;
    inv02 ix22456 (.Y (nx22457), .A (nx25023)) ;
    inv02 ix22458 (.Y (nx22459), .A (nx25023)) ;
    inv02 ix22460 (.Y (nx22461), .A (nx25023)) ;
    inv02 ix22462 (.Y (nx22463), .A (nx25023)) ;
    inv02 ix22464 (.Y (nx22465), .A (nx25025)) ;
    inv02 ix22466 (.Y (nx22467), .A (nx25025)) ;
    inv02 ix22468 (.Y (nx22469), .A (nx25025)) ;
    inv02 ix22470 (.Y (nx22471), .A (nx25025)) ;
    inv02 ix22472 (.Y (nx22473), .A (nx25025)) ;
    inv02 ix22474 (.Y (nx22475), .A (nx25025)) ;
    inv02 ix22476 (.Y (nx22477), .A (nx25025)) ;
    inv02 ix22478 (.Y (nx22479), .A (nx25027)) ;
    inv02 ix22480 (.Y (nx22481), .A (nx25027)) ;
    inv02 ix22482 (.Y (nx22483), .A (nx25027)) ;
    inv02 ix22484 (.Y (nx22485), .A (nx25027)) ;
    inv02 ix22486 (.Y (nx22487), .A (nx25027)) ;
    inv02 ix22488 (.Y (nx22489), .A (nx25027)) ;
    inv02 ix22490 (.Y (nx22491), .A (nx25027)) ;
    inv02 ix22492 (.Y (nx22493), .A (nx25029)) ;
    inv02 ix22494 (.Y (nx22495), .A (nx25029)) ;
    inv02 ix22496 (.Y (nx22497), .A (nx25029)) ;
    inv02 ix22498 (.Y (nx22499), .A (nx25029)) ;
    inv02 ix22500 (.Y (nx22501), .A (nx25029)) ;
    inv02 ix22502 (.Y (nx22503), .A (nx25029)) ;
    inv02 ix22504 (.Y (nx22505), .A (nx25029)) ;
    inv02 ix22506 (.Y (nx22507), .A (nx25031)) ;
    inv02 ix22508 (.Y (nx22509), .A (nx25031)) ;
    inv02 ix22510 (.Y (nx22511), .A (nx25031)) ;
    inv02 ix22512 (.Y (nx22513), .A (nx25031)) ;
    inv02 ix22514 (.Y (nx22515), .A (nx25031)) ;
    inv02 ix22516 (.Y (nx22517), .A (nx25031)) ;
    inv02 ix22518 (.Y (nx22519), .A (nx25031)) ;
    inv02 ix22520 (.Y (nx22521), .A (nx25033)) ;
    inv02 ix22522 (.Y (nx22523), .A (nx25033)) ;
    inv02 ix22526 (.Y (nx22527), .A (nx25035)) ;
    inv02 ix22528 (.Y (nx22529), .A (nx25035)) ;
    inv02 ix22530 (.Y (nx22531), .A (nx25035)) ;
    inv02 ix22532 (.Y (nx22533), .A (nx25035)) ;
    inv02 ix22534 (.Y (nx22535), .A (nx25035)) ;
    inv02 ix22536 (.Y (nx22537), .A (nx25035)) ;
    inv02 ix22538 (.Y (nx22539), .A (nx25035)) ;
    inv02 ix22540 (.Y (nx22541), .A (nx25037)) ;
    inv02 ix22542 (.Y (nx22543), .A (nx25037)) ;
    inv02 ix22544 (.Y (nx22545), .A (nx25037)) ;
    inv02 ix22546 (.Y (nx22547), .A (nx25037)) ;
    inv02 ix22548 (.Y (nx22549), .A (nx25037)) ;
    inv02 ix22550 (.Y (nx22551), .A (nx25037)) ;
    inv02 ix22552 (.Y (nx22553), .A (nx25037)) ;
    inv02 ix22554 (.Y (nx22555), .A (nx25039)) ;
    inv02 ix22556 (.Y (nx22557), .A (nx25039)) ;
    inv02 ix22558 (.Y (nx22559), .A (nx25039)) ;
    inv02 ix22560 (.Y (nx22561), .A (nx25039)) ;
    inv02 ix22562 (.Y (nx22563), .A (nx25039)) ;
    inv02 ix22564 (.Y (nx22565), .A (nx25039)) ;
    inv02 ix22566 (.Y (nx22567), .A (nx25039)) ;
    inv02 ix22568 (.Y (nx22569), .A (nx25041)) ;
    inv02 ix22570 (.Y (nx22571), .A (nx25041)) ;
    inv02 ix22572 (.Y (nx22573), .A (nx25041)) ;
    inv02 ix22574 (.Y (nx22575), .A (nx25041)) ;
    inv02 ix22576 (.Y (nx22577), .A (nx25041)) ;
    inv02 ix22578 (.Y (nx22579), .A (nx25041)) ;
    inv02 ix22580 (.Y (nx22581), .A (nx25041)) ;
    inv02 ix22582 (.Y (nx22583), .A (nx25043)) ;
    inv02 ix22584 (.Y (nx22585), .A (nx25043)) ;
    inv02 ix22586 (.Y (nx22587), .A (nx25043)) ;
    inv02 ix22588 (.Y (nx22589), .A (nx25043)) ;
    inv02 ix22590 (.Y (nx22591), .A (nx25043)) ;
    inv02 ix22592 (.Y (nx22593), .A (nx25043)) ;
    inv02 ix22594 (.Y (nx22595), .A (nx25043)) ;
    inv02 ix22596 (.Y (nx22597), .A (nx25045)) ;
    inv02 ix22598 (.Y (nx22599), .A (nx25045)) ;
    inv02 ix22600 (.Y (nx22601), .A (nx25045)) ;
    inv02 ix22602 (.Y (nx22603), .A (nx25045)) ;
    inv02 ix22604 (.Y (nx22605), .A (nx25045)) ;
    inv02 ix22606 (.Y (nx22607), .A (nx25045)) ;
    inv02 ix22608 (.Y (nx22609), .A (nx25045)) ;
    inv02 ix22610 (.Y (nx22611), .A (nx25047)) ;
    inv02 ix22612 (.Y (nx22613), .A (nx25047)) ;
    inv02 ix22614 (.Y (nx22615), .A (nx25047)) ;
    inv02 ix22616 (.Y (nx22617), .A (nx25047)) ;
    inv02 ix22618 (.Y (nx22619), .A (nx25047)) ;
    inv02 ix22620 (.Y (nx22621), .A (nx25047)) ;
    inv02 ix22622 (.Y (nx22623), .A (nx25047)) ;
    inv02 ix22624 (.Y (nx22625), .A (nx25049)) ;
    inv02 ix22626 (.Y (nx22627), .A (nx25049)) ;
    inv02 ix22628 (.Y (nx22629), .A (nx25049)) ;
    inv02 ix22630 (.Y (nx22631), .A (nx25049)) ;
    inv02 ix22632 (.Y (nx22633), .A (nx25049)) ;
    inv02 ix22634 (.Y (nx22635), .A (nx25049)) ;
    inv02 ix22636 (.Y (nx22637), .A (nx25049)) ;
    inv02 ix22638 (.Y (nx22639), .A (nx25051)) ;
    inv02 ix22640 (.Y (nx22641), .A (nx25051)) ;
    inv02 ix22642 (.Y (nx22643), .A (nx25051)) ;
    inv02 ix22644 (.Y (nx22645), .A (nx25051)) ;
    inv02 ix22646 (.Y (nx22647), .A (nx25051)) ;
    inv02 ix22648 (.Y (nx22649), .A (nx25051)) ;
    inv02 ix22650 (.Y (nx22651), .A (nx25051)) ;
    inv02 ix22652 (.Y (nx22653), .A (nx25053)) ;
    inv02 ix22654 (.Y (nx22655), .A (nx25053)) ;
    inv02 ix22656 (.Y (nx22657), .A (nx25053)) ;
    inv02 ix22658 (.Y (nx22659), .A (nx25053)) ;
    inv02 ix22660 (.Y (nx22661), .A (nx25053)) ;
    inv02 ix22662 (.Y (nx22663), .A (nx25053)) ;
    inv02 ix22664 (.Y (nx22665), .A (nx25053)) ;
    inv02 ix22666 (.Y (nx22667), .A (nx25055)) ;
    inv02 ix22668 (.Y (nx22669), .A (nx25055)) ;
    inv02 ix22670 (.Y (nx22671), .A (nx25055)) ;
    inv02 ix22672 (.Y (nx22673), .A (nx25055)) ;
    inv02 ix22676 (.Y (nx22677), .A (nx25057)) ;
    inv02 ix22678 (.Y (nx22679), .A (nx25057)) ;
    inv02 ix22680 (.Y (nx22681), .A (nx25057)) ;
    inv02 ix22682 (.Y (nx22683), .A (nx25057)) ;
    inv02 ix22684 (.Y (nx22685), .A (nx25057)) ;
    inv02 ix22686 (.Y (nx22687), .A (nx25057)) ;
    inv02 ix22688 (.Y (nx22689), .A (nx25057)) ;
    inv02 ix22690 (.Y (nx22691), .A (nx25059)) ;
    inv02 ix22692 (.Y (nx22693), .A (nx25059)) ;
    inv02 ix22694 (.Y (nx22695), .A (nx25059)) ;
    inv02 ix22696 (.Y (nx22697), .A (nx25059)) ;
    inv02 ix22698 (.Y (nx22699), .A (nx25059)) ;
    inv02 ix22700 (.Y (nx22701), .A (nx25059)) ;
    inv02 ix22702 (.Y (nx22703), .A (nx25059)) ;
    inv02 ix22704 (.Y (nx22705), .A (nx25061)) ;
    inv02 ix22706 (.Y (nx22707), .A (nx25061)) ;
    inv02 ix22708 (.Y (nx22709), .A (nx25061)) ;
    inv02 ix22710 (.Y (nx22711), .A (nx25061)) ;
    inv02 ix22712 (.Y (nx22713), .A (nx25061)) ;
    inv02 ix22714 (.Y (nx22715), .A (nx25061)) ;
    inv02 ix22716 (.Y (nx22717), .A (nx25061)) ;
    inv02 ix22718 (.Y (nx22719), .A (nx25063)) ;
    inv02 ix22720 (.Y (nx22721), .A (nx25063)) ;
    inv02 ix22722 (.Y (nx22723), .A (nx25063)) ;
    inv02 ix22724 (.Y (nx22725), .A (nx25063)) ;
    inv02 ix22726 (.Y (nx22727), .A (nx25063)) ;
    inv02 ix22728 (.Y (nx22729), .A (nx25063)) ;
    inv02 ix22730 (.Y (nx22731), .A (nx25063)) ;
    inv02 ix22732 (.Y (nx22733), .A (nx25065)) ;
    inv02 ix22734 (.Y (nx22735), .A (nx25065)) ;
    inv02 ix22736 (.Y (nx22737), .A (nx25065)) ;
    inv02 ix22738 (.Y (nx22739), .A (nx25065)) ;
    inv02 ix22740 (.Y (nx22741), .A (nx25065)) ;
    inv02 ix22742 (.Y (nx22743), .A (nx25065)) ;
    inv02 ix22744 (.Y (nx22745), .A (nx25065)) ;
    inv02 ix22746 (.Y (nx22747), .A (nx25067)) ;
    inv02 ix22748 (.Y (nx22749), .A (nx25067)) ;
    inv02 ix22750 (.Y (nx22751), .A (nx25067)) ;
    inv02 ix22752 (.Y (nx22753), .A (nx25067)) ;
    inv02 ix22754 (.Y (nx22755), .A (nx25067)) ;
    inv02 ix22756 (.Y (nx22757), .A (nx25067)) ;
    inv02 ix22758 (.Y (nx22759), .A (nx25067)) ;
    inv02 ix22760 (.Y (nx22761), .A (nx25069)) ;
    inv02 ix22762 (.Y (nx22763), .A (nx25069)) ;
    inv02 ix22764 (.Y (nx22765), .A (nx25069)) ;
    inv02 ix22766 (.Y (nx22767), .A (nx25069)) ;
    inv02 ix22768 (.Y (nx22769), .A (nx25069)) ;
    inv02 ix22770 (.Y (nx22771), .A (nx25069)) ;
    inv02 ix22772 (.Y (nx22773), .A (nx25069)) ;
    inv02 ix22774 (.Y (nx22775), .A (nx25071)) ;
    inv02 ix22776 (.Y (nx22777), .A (nx25071)) ;
    inv02 ix22778 (.Y (nx22779), .A (nx25071)) ;
    inv02 ix22780 (.Y (nx22781), .A (nx25071)) ;
    inv02 ix22782 (.Y (nx22783), .A (nx25071)) ;
    inv02 ix22784 (.Y (nx22785), .A (nx25071)) ;
    inv02 ix22786 (.Y (nx22787), .A (nx25071)) ;
    inv02 ix22788 (.Y (nx22789), .A (nx25073)) ;
    inv02 ix22790 (.Y (nx22791), .A (nx25073)) ;
    inv02 ix22792 (.Y (nx22793), .A (nx25073)) ;
    inv02 ix22794 (.Y (nx22795), .A (nx25073)) ;
    inv02 ix22796 (.Y (nx22797), .A (nx25073)) ;
    inv02 ix22798 (.Y (nx22799), .A (nx25073)) ;
    inv02 ix22800 (.Y (nx22801), .A (nx25073)) ;
    inv02 ix22802 (.Y (nx22803), .A (nx25075)) ;
    inv02 ix22804 (.Y (nx22805), .A (nx25075)) ;
    inv02 ix22806 (.Y (nx22807), .A (nx25075)) ;
    inv02 ix22808 (.Y (nx22809), .A (nx25075)) ;
    inv02 ix22810 (.Y (nx22811), .A (nx25075)) ;
    inv02 ix22812 (.Y (nx22813), .A (nx25075)) ;
    inv02 ix22814 (.Y (nx22815), .A (nx25075)) ;
    inv02 ix22816 (.Y (nx22817), .A (nx25077)) ;
    inv02 ix22818 (.Y (nx22819), .A (nx25077)) ;
    inv02 ix22820 (.Y (nx22821), .A (nx25077)) ;
    inv02 ix22822 (.Y (nx22823), .A (nx25077)) ;
    inv02 ix22824 (.Y (nx22825), .A (nx25077)) ;
    inv02 ix22826 (.Y (nx22827), .A (nx25077)) ;
    inv02 ix22828 (.Y (nx22829), .A (nx25077)) ;
    inv02 ix22830 (.Y (nx22831), .A (nx25079)) ;
    inv02 ix22832 (.Y (nx22833), .A (nx25079)) ;
    inv02 ix22834 (.Y (nx22835), .A (nx25079)) ;
    inv02 ix22836 (.Y (nx22837), .A (nx25079)) ;
    inv02 ix22838 (.Y (nx22839), .A (nx25079)) ;
    inv02 ix22840 (.Y (nx22841), .A (nx25079)) ;
    inv02 ix22842 (.Y (nx22843), .A (nx25079)) ;
    inv02 ix22844 (.Y (nx22845), .A (nx25081)) ;
    inv02 ix22846 (.Y (nx22847), .A (nx25081)) ;
    inv02 ix22848 (.Y (nx22849), .A (nx25081)) ;
    inv02 ix22850 (.Y (nx22851), .A (nx25081)) ;
    inv02 ix22852 (.Y (nx22853), .A (nx25081)) ;
    inv02 ix22854 (.Y (nx22855), .A (nx25081)) ;
    inv02 ix22856 (.Y (nx22857), .A (nx25081)) ;
    inv02 ix22858 (.Y (nx22859), .A (nx25083)) ;
    inv02 ix22860 (.Y (nx22861), .A (nx25083)) ;
    inv02 ix22862 (.Y (nx22863), .A (nx25083)) ;
    inv02 ix22864 (.Y (nx22865), .A (nx25083)) ;
    inv02 ix22866 (.Y (nx22867), .A (nx25083)) ;
    inv02 ix22868 (.Y (nx22869), .A (nx25083)) ;
    inv02 ix22870 (.Y (nx22871), .A (nx25083)) ;
    inv02 ix22872 (.Y (nx22873), .A (nx25085)) ;
    inv02 ix22874 (.Y (nx22875), .A (nx25085)) ;
    inv02 ix22876 (.Y (nx22877), .A (nx25085)) ;
    inv02 ix22878 (.Y (nx22879), .A (nx25085)) ;
    inv02 ix22880 (.Y (nx22881), .A (nx25085)) ;
    inv02 ix22882 (.Y (nx22883), .A (nx25085)) ;
    inv02 ix22884 (.Y (nx22885), .A (nx25085)) ;
    inv02 ix22886 (.Y (nx22887), .A (nx25087)) ;
    inv02 ix22888 (.Y (nx22889), .A (nx25087)) ;
    inv02 ix22890 (.Y (nx22891), .A (nx25087)) ;
    inv02 ix22892 (.Y (nx22893), .A (nx25087)) ;
    inv02 ix22894 (.Y (nx22895), .A (nx25087)) ;
    inv02 ix22896 (.Y (nx22897), .A (nx25087)) ;
    inv02 ix22898 (.Y (nx22899), .A (nx25087)) ;
    inv02 ix22900 (.Y (nx22901), .A (nx25089)) ;
    inv02 ix22902 (.Y (nx22903), .A (nx25089)) ;
    inv02 ix22904 (.Y (nx22905), .A (nx25089)) ;
    inv02 ix22906 (.Y (nx22907), .A (nx25089)) ;
    inv02 ix22908 (.Y (nx22909), .A (nx25089)) ;
    inv02 ix22910 (.Y (nx22911), .A (nx25089)) ;
    inv02 ix22912 (.Y (nx22913), .A (nx25089)) ;
    inv02 ix22914 (.Y (nx22915), .A (nx25091)) ;
    inv02 ix22916 (.Y (nx22917), .A (nx25091)) ;
    inv02 ix22918 (.Y (nx22919), .A (nx25091)) ;
    inv02 ix22920 (.Y (nx22921), .A (nx25091)) ;
    inv02 ix22922 (.Y (nx22923), .A (nx25091)) ;
    inv02 ix22924 (.Y (nx22925), .A (nx25091)) ;
    inv02 ix22926 (.Y (nx22927), .A (nx25091)) ;
    inv02 ix22928 (.Y (nx22929), .A (nx25093)) ;
    inv02 ix22930 (.Y (nx22931), .A (nx25093)) ;
    inv02 ix22932 (.Y (nx22933), .A (nx25093)) ;
    inv02 ix22934 (.Y (nx22935), .A (nx25093)) ;
    inv02 ix22936 (.Y (nx22937), .A (nx25093)) ;
    inv02 ix22938 (.Y (nx22939), .A (nx25093)) ;
    inv02 ix22940 (.Y (nx22941), .A (nx25093)) ;
    inv02 ix22942 (.Y (nx22943), .A (nx25095)) ;
    inv02 ix22944 (.Y (nx22945), .A (nx25095)) ;
    inv02 ix22946 (.Y (nx22947), .A (nx25095)) ;
    inv02 ix22948 (.Y (nx22949), .A (nx25095)) ;
    inv02 ix22950 (.Y (nx22951), .A (nx25095)) ;
    inv02 ix22952 (.Y (nx22953), .A (nx25095)) ;
    inv02 ix22954 (.Y (nx22955), .A (nx25095)) ;
    inv02 ix22956 (.Y (nx22957), .A (nx25097)) ;
    inv02 ix22958 (.Y (nx22959), .A (nx25097)) ;
    inv02 ix22960 (.Y (nx22961), .A (nx25097)) ;
    inv02 ix22962 (.Y (nx22963), .A (nx25097)) ;
    inv02 ix22964 (.Y (nx22965), .A (nx25097)) ;
    inv02 ix22966 (.Y (nx22967), .A (nx25097)) ;
    inv02 ix22968 (.Y (nx22969), .A (nx25097)) ;
    inv02 ix22970 (.Y (nx22971), .A (nx25099)) ;
    inv02 ix22972 (.Y (nx22973), .A (nx25099)) ;
    inv02 ix22974 (.Y (nx22975), .A (nx25099)) ;
    inv02 ix22976 (.Y (nx22977), .A (nx25099)) ;
    inv02 ix22978 (.Y (nx22979), .A (nx25099)) ;
    inv02 ix22980 (.Y (nx22981), .A (nx25099)) ;
    inv02 ix22982 (.Y (nx22983), .A (nx25099)) ;
    inv02 ix22984 (.Y (nx22985), .A (nx25101)) ;
    inv02 ix22986 (.Y (nx22987), .A (nx25101)) ;
    inv02 ix22988 (.Y (nx22989), .A (nx25101)) ;
    inv02 ix22990 (.Y (nx22991), .A (nx25101)) ;
    inv02 ix22992 (.Y (nx22993), .A (nx25101)) ;
    inv02 ix22994 (.Y (nx22995), .A (nx25101)) ;
    inv02 ix22996 (.Y (nx22997), .A (nx25101)) ;
    inv02 ix22998 (.Y (nx22999), .A (nx25103)) ;
    inv02 ix23000 (.Y (nx23001), .A (nx25103)) ;
    inv02 ix23002 (.Y (nx23003), .A (nx25103)) ;
    inv02 ix23004 (.Y (nx23005), .A (nx25103)) ;
    inv02 ix23006 (.Y (nx23007), .A (nx25103)) ;
    inv02 ix23008 (.Y (nx23009), .A (nx25103)) ;
    inv02 ix23010 (.Y (nx23011), .A (nx25103)) ;
    inv02 ix23012 (.Y (nx23013), .A (nx25105)) ;
    inv02 ix23014 (.Y (nx23015), .A (nx25105)) ;
    inv02 ix23016 (.Y (nx23017), .A (nx25105)) ;
    inv02 ix23018 (.Y (nx23019), .A (nx25105)) ;
    inv02 ix23020 (.Y (nx23021), .A (nx25105)) ;
    inv02 ix23022 (.Y (nx23023), .A (nx25105)) ;
    inv02 ix23024 (.Y (nx23025), .A (nx25105)) ;
    inv02 ix23026 (.Y (nx23027), .A (nx25107)) ;
    inv02 ix23028 (.Y (nx23029), .A (nx25107)) ;
    inv02 ix23030 (.Y (nx23031), .A (nx25107)) ;
    inv02 ix23032 (.Y (nx23033), .A (nx25107)) ;
    inv02 ix23034 (.Y (nx23035), .A (nx25107)) ;
    inv02 ix23036 (.Y (nx23037), .A (nx25107)) ;
    inv02 ix23038 (.Y (nx23039), .A (nx25107)) ;
    inv02 ix23040 (.Y (nx23041), .A (nx25109)) ;
    inv02 ix23042 (.Y (nx23043), .A (nx25109)) ;
    inv02 ix23044 (.Y (nx23045), .A (nx25109)) ;
    inv02 ix23046 (.Y (nx23047), .A (nx25109)) ;
    inv02 ix23048 (.Y (nx23049), .A (nx25109)) ;
    inv02 ix23050 (.Y (nx23051), .A (nx25109)) ;
    inv02 ix23052 (.Y (nx23053), .A (nx25109)) ;
    inv02 ix23054 (.Y (nx23055), .A (nx25111)) ;
    inv02 ix23056 (.Y (nx23057), .A (nx25111)) ;
    inv02 ix23058 (.Y (nx23059), .A (nx25111)) ;
    inv02 ix23060 (.Y (nx23061), .A (nx25111)) ;
    inv02 ix23062 (.Y (nx23063), .A (nx25111)) ;
    inv02 ix23064 (.Y (nx23065), .A (nx25111)) ;
    inv02 ix23066 (.Y (nx23067), .A (nx25111)) ;
    inv02 ix23068 (.Y (nx23069), .A (nx25113)) ;
    inv02 ix23070 (.Y (nx23071), .A (nx25113)) ;
    inv02 ix23072 (.Y (nx23073), .A (nx25113)) ;
    inv02 ix23074 (.Y (nx23075), .A (nx25113)) ;
    inv02 ix23076 (.Y (nx23077), .A (nx25113)) ;
    inv02 ix23078 (.Y (nx23079), .A (nx25113)) ;
    inv02 ix23080 (.Y (nx23081), .A (nx25113)) ;
    inv02 ix23082 (.Y (nx23083), .A (nx25115)) ;
    inv02 ix23084 (.Y (nx23085), .A (nx25115)) ;
    inv02 ix23086 (.Y (nx23087), .A (nx25115)) ;
    inv02 ix23088 (.Y (nx23089), .A (nx25115)) ;
    inv02 ix23090 (.Y (nx23091), .A (nx25115)) ;
    inv02 ix23092 (.Y (nx23093), .A (nx25115)) ;
    inv02 ix23094 (.Y (nx23095), .A (nx25115)) ;
    inv02 ix23096 (.Y (nx23097), .A (nx25117)) ;
    inv02 ix23098 (.Y (nx23099), .A (nx25117)) ;
    inv02 ix23100 (.Y (nx23101), .A (nx25117)) ;
    inv02 ix23102 (.Y (nx23103), .A (nx25117)) ;
    inv02 ix23104 (.Y (nx23105), .A (nx25117)) ;
    inv02 ix23106 (.Y (nx23107), .A (nx25117)) ;
    inv02 ix23108 (.Y (nx23109), .A (nx25117)) ;
    inv02 ix23110 (.Y (nx23111), .A (nx25119)) ;
    inv02 ix23112 (.Y (nx23113), .A (nx25119)) ;
    inv02 ix23114 (.Y (nx23115), .A (nx25119)) ;
    inv02 ix23116 (.Y (nx23117), .A (nx24839)) ;
    inv02 ix23118 (.Y (nx23119), .A (nx24839)) ;
    inv02 ix23120 (.Y (nx23121), .A (nx24839)) ;
    inv02 ix23122 (.Y (nx23123), .A (nx24841)) ;
    inv02 ix23124 (.Y (nx23125), .A (nx24841)) ;
    inv02 ix23126 (.Y (nx23127), .A (nx24841)) ;
    inv02 ix23128 (.Y (nx23129), .A (nx24841)) ;
    inv02 ix23130 (.Y (nx23131), .A (nx24841)) ;
    inv02 ix23132 (.Y (nx23133), .A (nx24841)) ;
    inv02 ix23134 (.Y (nx23135), .A (nx24841)) ;
    inv02 ix23136 (.Y (nx23137), .A (nx24843)) ;
    inv02 ix23138 (.Y (nx23139), .A (nx24843)) ;
    inv02 ix23140 (.Y (nx23141), .A (nx24843)) ;
    inv02 ix23142 (.Y (nx23143), .A (nx24843)) ;
    inv02 ix23144 (.Y (nx23145), .A (nx24843)) ;
    inv02 ix23146 (.Y (nx23147), .A (nx24843)) ;
    inv02 ix23148 (.Y (nx23149), .A (nx24843)) ;
    inv02 ix23150 (.Y (nx23151), .A (nx24845)) ;
    inv02 ix23152 (.Y (nx23153), .A (nx24845)) ;
    inv02 ix23154 (.Y (nx23155), .A (nx24845)) ;
    inv02 ix23156 (.Y (nx23157), .A (nx24845)) ;
    inv02 ix23158 (.Y (nx23159), .A (nx24845)) ;
    inv02 ix23160 (.Y (nx23161), .A (nx24845)) ;
    inv02 ix23162 (.Y (nx23163), .A (nx24845)) ;
    inv02 ix23164 (.Y (nx23165), .A (nx24847)) ;
    inv02 ix23166 (.Y (nx23167), .A (nx24847)) ;
    inv02 ix23168 (.Y (nx23169), .A (nx24847)) ;
    inv02 ix23170 (.Y (nx23171), .A (nx24847)) ;
    inv02 ix23172 (.Y (nx23173), .A (nx24847)) ;
    inv02 ix23174 (.Y (nx23175), .A (nx24847)) ;
    inv02 ix23176 (.Y (nx23177), .A (nx24847)) ;
    inv02 ix23178 (.Y (nx23179), .A (nx24849)) ;
    inv02 ix23180 (.Y (nx23181), .A (nx24849)) ;
    inv02 ix23182 (.Y (nx23183), .A (nx24849)) ;
    inv02 ix23184 (.Y (nx23185), .A (nx24849)) ;
    inv02 ix23186 (.Y (nx23187), .A (nx24849)) ;
    inv02 ix23188 (.Y (nx23189), .A (nx24849)) ;
    inv02 ix23190 (.Y (nx23191), .A (nx24857)) ;
    inv02 ix23192 (.Y (nx23193), .A (nx24857)) ;
    inv02 ix23194 (.Y (nx23195), .A (nx24857)) ;
    inv02 ix23196 (.Y (nx23197), .A (nx24857)) ;
    inv02 ix23198 (.Y (nx23199), .A (nx24857)) ;
    inv02 ix23200 (.Y (nx23201), .A (nx24857)) ;
    inv02 ix23202 (.Y (nx23203), .A (nx24857)) ;
    inv02 ix23204 (.Y (nx23205), .A (nx24859)) ;
    inv02 ix23206 (.Y (nx23207), .A (nx24859)) ;
    inv02 ix23208 (.Y (nx23209), .A (nx24859)) ;
    inv02 ix23210 (.Y (nx23211), .A (nx24859)) ;
    inv02 ix23212 (.Y (nx23213), .A (nx24859)) ;
    inv02 ix23214 (.Y (nx23215), .A (nx24859)) ;
    inv02 ix23216 (.Y (nx23217), .A (nx24859)) ;
    inv02 ix23218 (.Y (nx23219), .A (nx24861)) ;
    inv02 ix23220 (.Y (nx23221), .A (nx24861)) ;
    inv02 ix23222 (.Y (nx23223), .A (nx24861)) ;
    inv02 ix23224 (.Y (nx23225), .A (nx24861)) ;
    inv02 ix23226 (.Y (nx23227), .A (nx24861)) ;
    inv02 ix23228 (.Y (nx23229), .A (nx24861)) ;
    inv02 ix23230 (.Y (nx23231), .A (nx24861)) ;
    inv02 ix23232 (.Y (nx23233), .A (nx24863)) ;
    inv02 ix23234 (.Y (nx23235), .A (nx24863)) ;
    inv02 ix23236 (.Y (nx23237), .A (nx24863)) ;
    inv02 ix23238 (.Y (nx23239), .A (nx24863)) ;
    inv02 ix23240 (.Y (nx23241), .A (nx24863)) ;
    inv02 ix23242 (.Y (nx23243), .A (nx24863)) ;
    inv02 ix23244 (.Y (nx23245), .A (nx24863)) ;
    inv02 ix23246 (.Y (nx23247), .A (nx24865)) ;
    inv02 ix23248 (.Y (nx23249), .A (nx24865)) ;
    inv02 ix23250 (.Y (nx23251), .A (nx24865)) ;
    inv02 ix23252 (.Y (nx23253), .A (nx24865)) ;
    inv02 ix23254 (.Y (nx23255), .A (nx24865)) ;
    inv02 ix23256 (.Y (nx23257), .A (nx24865)) ;
    inv02 ix23258 (.Y (nx23259), .A (nx24865)) ;
    inv02 ix23260 (.Y (nx23261), .A (nx24867)) ;
    inv02 ix23262 (.Y (nx23263), .A (nx24867)) ;
    inv02 ix23264 (.Y (nx23265), .A (nx24867)) ;
    inv02 ix23266 (.Y (nx23267), .A (nx24867)) ;
    inv02 ix23268 (.Y (nx23269), .A (nx24867)) ;
    inv02 ix23270 (.Y (nx23271), .A (nx24867)) ;
    inv02 ix23272 (.Y (nx23273), .A (nx24867)) ;
    inv02 ix23274 (.Y (nx23275), .A (nx24869)) ;
    inv02 ix23276 (.Y (nx23277), .A (nx24869)) ;
    inv02 ix23278 (.Y (nx23279), .A (nx24869)) ;
    inv02 ix23280 (.Y (nx23281), .A (nx24869)) ;
    inv02 ix23282 (.Y (nx23283), .A (nx24869)) ;
    inv02 ix23284 (.Y (nx23285), .A (nx24869)) ;
    inv02 ix23286 (.Y (nx23287), .A (nx24869)) ;
    inv02 ix23288 (.Y (nx23289), .A (nx24871)) ;
    inv02 ix23290 (.Y (nx23291), .A (nx24871)) ;
    inv02 ix23292 (.Y (nx23293), .A (nx24871)) ;
    inv02 ix23294 (.Y (nx23295), .A (nx24871)) ;
    inv02 ix23296 (.Y (nx23297), .A (nx24871)) ;
    inv02 ix23298 (.Y (nx23299), .A (nx24871)) ;
    inv02 ix23300 (.Y (nx23301), .A (nx24871)) ;
    inv02 ix23302 (.Y (nx23303), .A (nx24873)) ;
    inv02 ix23304 (.Y (nx23305), .A (nx24873)) ;
    inv02 ix23306 (.Y (nx23307), .A (nx24873)) ;
    inv02 ix23308 (.Y (nx23309), .A (nx24873)) ;
    inv02 ix23310 (.Y (nx23311), .A (nx24873)) ;
    inv02 ix23312 (.Y (nx23313), .A (nx24873)) ;
    inv02 ix23314 (.Y (nx23315), .A (nx24873)) ;
    inv02 ix23316 (.Y (nx23317), .A (nx24875)) ;
    inv02 ix23318 (.Y (nx23319), .A (nx24875)) ;
    inv02 ix23320 (.Y (nx23321), .A (nx24875)) ;
    inv02 ix23322 (.Y (nx23323), .A (nx24875)) ;
    inv02 ix23324 (.Y (nx23325), .A (nx24875)) ;
    inv02 ix23326 (.Y (nx23327), .A (nx24875)) ;
    inv02 ix23328 (.Y (nx23329), .A (nx24875)) ;
    inv02 ix23330 (.Y (nx23331), .A (nx24877)) ;
    inv02 ix23332 (.Y (nx23333), .A (nx24877)) ;
    inv02 ix23334 (.Y (nx23335), .A (nx24877)) ;
    inv02 ix23336 (.Y (nx23337), .A (nx24877)) ;
    inv02 ix23338 (.Y (nx23339), .A (nx24877)) ;
    inv02 ix23340 (.Y (nx23341), .A (nx24877)) ;
    inv02 ix23342 (.Y (nx23343), .A (nx24877)) ;
    inv02 ix23344 (.Y (nx23345), .A (nx22227)) ;
    inv02 ix23346 (.Y (nx23347), .A (nx22227)) ;
    inv02 ix23348 (.Y (nx23349), .A (nx22227)) ;
    inv02 ix23350 (.Y (nx23351), .A (nx22227)) ;
    inv02 ix23352 (.Y (nx23353), .A (nx22227)) ;
    inv02 ix23354 (.Y (nx23355), .A (nx22227)) ;
    inv02 ix23356 (.Y (nx23357), .A (nx22227)) ;
    inv02 ix23360 (.Y (nx23361), .A (nx25121)) ;
    inv02 ix23362 (.Y (nx23363), .A (nx25121)) ;
    inv02 ix23364 (.Y (nx23365), .A (nx25121)) ;
    inv02 ix23366 (.Y (nx23367), .A (nx25121)) ;
    inv02 ix23368 (.Y (nx23369), .A (nx25121)) ;
    inv02 ix23370 (.Y (nx23371), .A (nx25121)) ;
    inv02 ix23372 (.Y (nx23373), .A (nx25121)) ;
    inv02 ix23374 (.Y (nx23375), .A (nx25123)) ;
    inv02 ix23376 (.Y (nx23377), .A (nx25123)) ;
    inv02 ix23378 (.Y (nx23379), .A (nx25123)) ;
    inv02 ix23380 (.Y (nx23381), .A (nx25123)) ;
    inv02 ix23382 (.Y (nx23383), .A (nx25123)) ;
    inv02 ix23384 (.Y (nx23385), .A (nx25123)) ;
    inv02 ix23386 (.Y (nx23387), .A (nx25123)) ;
    inv02 ix23388 (.Y (nx23389), .A (nx25125)) ;
    inv02 ix23390 (.Y (nx23391), .A (nx25125)) ;
    inv02 ix23392 (.Y (nx23393), .A (nx25125)) ;
    inv02 ix23394 (.Y (nx23395), .A (nx25125)) ;
    inv02 ix23396 (.Y (nx23397), .A (nx25125)) ;
    inv02 ix23398 (.Y (nx23399), .A (nx25125)) ;
    inv02 ix23400 (.Y (nx23401), .A (nx25125)) ;
    inv02 ix23402 (.Y (nx23403), .A (nx25127)) ;
    inv02 ix23404 (.Y (nx23405), .A (nx25127)) ;
    inv02 ix23406 (.Y (nx23407), .A (nx25127)) ;
    inv02 ix23408 (.Y (nx23409), .A (nx25127)) ;
    inv02 ix23410 (.Y (nx23411), .A (nx25127)) ;
    inv02 ix23412 (.Y (nx23413), .A (nx25127)) ;
    inv02 ix23414 (.Y (nx23415), .A (nx25127)) ;
    inv02 ix23416 (.Y (nx23417), .A (nx25129)) ;
    inv02 ix23418 (.Y (nx23419), .A (nx25129)) ;
    inv02 ix23420 (.Y (nx23421), .A (nx25129)) ;
    inv02 ix23422 (.Y (nx23423), .A (nx25129)) ;
    inv02 ix23424 (.Y (nx23425), .A (nx25129)) ;
    inv02 ix23426 (.Y (nx23427), .A (nx25129)) ;
    inv02 ix23428 (.Y (nx23429), .A (nx25129)) ;
    inv02 ix23430 (.Y (nx23431), .A (nx25131)) ;
    inv02 ix23432 (.Y (nx23433), .A (nx25131)) ;
    inv02 ix23434 (.Y (nx23435), .A (nx25131)) ;
    inv02 ix23436 (.Y (nx23437), .A (nx25131)) ;
    inv02 ix23438 (.Y (nx23439), .A (nx25131)) ;
    inv02 ix23440 (.Y (nx23441), .A (nx25131)) ;
    inv02 ix23442 (.Y (nx23443), .A (nx25131)) ;
    inv02 ix23444 (.Y (nx23445), .A (nx25133)) ;
    inv02 ix23446 (.Y (nx23447), .A (nx25133)) ;
    inv02 ix23448 (.Y (nx23449), .A (nx25133)) ;
    inv02 ix23450 (.Y (nx23451), .A (nx25133)) ;
    inv02 ix23452 (.Y (nx23453), .A (nx25133)) ;
    inv02 ix23454 (.Y (nx23455), .A (nx25133)) ;
    inv02 ix23456 (.Y (nx23457), .A (nx25133)) ;
    inv02 ix23458 (.Y (nx23459), .A (nx25135)) ;
    inv02 ix23460 (.Y (nx23461), .A (nx25135)) ;
    inv02 ix23462 (.Y (nx23463), .A (nx25135)) ;
    inv02 ix23464 (.Y (nx23465), .A (nx25135)) ;
    inv02 ix23466 (.Y (nx23467), .A (nx25135)) ;
    inv02 ix23468 (.Y (nx23469), .A (nx25135)) ;
    inv02 ix23470 (.Y (nx23471), .A (nx25135)) ;
    inv02 ix23472 (.Y (nx23473), .A (nx25137)) ;
    inv02 ix23474 (.Y (nx23475), .A (nx25137)) ;
    inv02 ix23476 (.Y (nx23477), .A (nx25137)) ;
    inv02 ix23478 (.Y (nx23479), .A (nx25137)) ;
    inv02 ix23480 (.Y (nx23481), .A (nx25137)) ;
    inv02 ix23482 (.Y (nx23483), .A (nx25137)) ;
    inv02 ix23484 (.Y (nx23485), .A (nx25137)) ;
    inv02 ix23486 (.Y (nx23487), .A (nx25139)) ;
    inv02 ix23488 (.Y (nx23489), .A (nx25139)) ;
    inv02 ix23490 (.Y (nx23491), .A (nx25139)) ;
    inv02 ix23492 (.Y (nx23493), .A (nx25139)) ;
    inv02 ix23494 (.Y (nx23495), .A (nx25139)) ;
    inv02 ix23496 (.Y (nx23497), .A (nx25139)) ;
    inv02 ix23498 (.Y (nx23499), .A (nx25139)) ;
    inv02 ix23500 (.Y (nx23501), .A (nx25141)) ;
    inv02 ix23502 (.Y (nx23503), .A (nx25141)) ;
    inv02 ix23504 (.Y (nx23505), .A (nx25141)) ;
    inv02 ix23506 (.Y (nx23507), .A (nx25141)) ;
    inv02 ix23508 (.Y (nx23509), .A (nx25141)) ;
    inv02 ix23510 (.Y (nx23511), .A (nx25141)) ;
    inv02 ix23512 (.Y (nx23513), .A (nx25141)) ;
    inv02 ix23514 (.Y (nx23515), .A (nx25143)) ;
    inv02 ix23516 (.Y (nx23517), .A (nx25143)) ;
    inv02 ix23518 (.Y (nx23519), .A (nx25143)) ;
    inv02 ix23520 (.Y (nx23521), .A (nx25143)) ;
    inv02 ix23522 (.Y (nx23523), .A (nx25143)) ;
    inv02 ix23524 (.Y (nx23525), .A (nx25143)) ;
    inv02 ix23526 (.Y (nx23527), .A (nx25143)) ;
    inv02 ix23528 (.Y (nx23529), .A (nx25145)) ;
    inv02 ix23530 (.Y (nx23531), .A (nx25145)) ;
    inv02 ix23532 (.Y (nx23533), .A (nx25145)) ;
    inv02 ix23534 (.Y (nx23535), .A (nx25145)) ;
    inv02 ix23536 (.Y (nx23537), .A (nx25145)) ;
    inv02 ix23538 (.Y (nx23539), .A (nx25145)) ;
    inv02 ix23540 (.Y (nx23541), .A (nx25145)) ;
    inv02 ix23542 (.Y (nx23543), .A (nx25147)) ;
    inv02 ix23544 (.Y (nx23545), .A (nx25147)) ;
    inv02 ix23546 (.Y (nx23547), .A (nx25147)) ;
    inv02 ix23548 (.Y (nx23549), .A (nx25147)) ;
    inv02 ix23550 (.Y (nx23551), .A (nx25147)) ;
    inv02 ix23552 (.Y (nx23553), .A (nx25147)) ;
    inv02 ix23554 (.Y (nx23555), .A (nx25147)) ;
    inv02 ix23556 (.Y (nx23557), .A (nx25149)) ;
    inv02 ix23558 (.Y (nx23559), .A (nx25149)) ;
    inv02 ix23560 (.Y (nx23561), .A (nx25149)) ;
    inv02 ix23562 (.Y (nx23563), .A (nx25149)) ;
    inv02 ix23564 (.Y (nx23565), .A (nx25149)) ;
    inv02 ix23566 (.Y (nx23567), .A (nx25149)) ;
    inv02 ix23568 (.Y (nx23569), .A (nx25149)) ;
    inv02 ix23570 (.Y (nx23571), .A (nx25151)) ;
    inv02 ix23572 (.Y (nx23573), .A (nx25151)) ;
    inv02 ix23574 (.Y (nx23575), .A (nx25151)) ;
    inv02 ix23576 (.Y (nx23577), .A (nx25151)) ;
    inv02 ix23578 (.Y (nx23579), .A (nx25151)) ;
    inv02 ix23580 (.Y (nx23581), .A (nx25151)) ;
    inv02 ix23582 (.Y (nx23583), .A (nx25151)) ;
    inv02 ix23584 (.Y (nx23585), .A (nx25153)) ;
    inv02 ix23586 (.Y (nx23587), .A (nx25153)) ;
    inv02 ix23588 (.Y (nx23589), .A (nx25153)) ;
    inv02 ix23590 (.Y (nx23591), .A (nx25153)) ;
    inv02 ix23592 (.Y (nx23593), .A (nx25153)) ;
    inv02 ix23594 (.Y (nx23595), .A (nx25153)) ;
    inv02 ix23596 (.Y (nx23597), .A (nx25153)) ;
    inv02 ix23598 (.Y (nx23599), .A (nx25155)) ;
    inv02 ix23600 (.Y (nx23601), .A (nx25155)) ;
    inv02 ix23602 (.Y (nx23603), .A (nx25155)) ;
    inv02 ix23604 (.Y (nx23605), .A (nx25155)) ;
    inv02 ix23606 (.Y (nx23607), .A (nx25155)) ;
    inv02 ix23608 (.Y (nx23609), .A (nx25155)) ;
    inv02 ix23610 (.Y (nx23611), .A (nx25155)) ;
    inv02 ix23612 (.Y (nx23613), .A (nx25157)) ;
    inv02 ix23614 (.Y (nx23615), .A (nx25157)) ;
    inv02 ix23616 (.Y (nx23617), .A (nx25157)) ;
    inv02 ix23618 (.Y (nx23619), .A (nx25157)) ;
    inv02 ix23620 (.Y (nx23621), .A (nx25157)) ;
    inv02 ix23622 (.Y (nx23623), .A (nx25157)) ;
    inv02 ix23624 (.Y (nx23625), .A (nx25157)) ;
    inv02 ix23626 (.Y (nx23627), .A (nx25159)) ;
    inv02 ix23628 (.Y (nx23629), .A (nx25159)) ;
    inv02 ix23630 (.Y (nx23631), .A (nx25159)) ;
    inv02 ix23632 (.Y (nx23633), .A (nx25159)) ;
    inv02 ix23634 (.Y (nx23635), .A (nx25159)) ;
    inv02 ix23636 (.Y (nx23637), .A (nx25159)) ;
    inv02 ix23638 (.Y (nx23639), .A (nx25159)) ;
    inv02 ix23640 (.Y (nx23641), .A (nx25161)) ;
    inv02 ix23642 (.Y (nx23643), .A (nx25161)) ;
    inv02 ix23644 (.Y (nx23645), .A (nx25161)) ;
    inv02 ix23646 (.Y (nx23647), .A (nx25161)) ;
    inv02 ix23648 (.Y (nx23649), .A (nx25161)) ;
    inv02 ix23650 (.Y (nx23651), .A (nx25161)) ;
    inv02 ix23652 (.Y (nx23653), .A (nx25161)) ;
    inv02 ix23654 (.Y (nx23655), .A (nx25163)) ;
    inv02 ix23656 (.Y (nx23657), .A (nx25163)) ;
    inv02 ix23658 (.Y (nx23659), .A (nx25163)) ;
    inv02 ix23660 (.Y (nx23661), .A (nx25163)) ;
    inv02 ix23662 (.Y (nx23663), .A (nx25163)) ;
    inv02 ix23664 (.Y (nx23665), .A (nx25163)) ;
    inv02 ix23666 (.Y (nx23667), .A (nx25163)) ;
    inv02 ix23668 (.Y (nx23669), .A (nx25165)) ;
    inv02 ix23670 (.Y (nx23671), .A (nx25165)) ;
    inv02 ix23672 (.Y (nx23673), .A (nx25165)) ;
    inv02 ix23674 (.Y (nx23675), .A (nx25165)) ;
    inv02 ix23676 (.Y (nx23677), .A (nx25165)) ;
    inv02 ix23678 (.Y (nx23679), .A (nx25165)) ;
    inv02 ix23680 (.Y (nx23681), .A (nx25165)) ;
    inv02 ix23682 (.Y (nx23683), .A (nx25167)) ;
    inv02 ix23684 (.Y (nx23685), .A (nx25167)) ;
    inv02 ix23686 (.Y (nx23687), .A (nx25167)) ;
    inv02 ix23688 (.Y (nx23689), .A (nx25167)) ;
    inv02 ix23690 (.Y (nx23691), .A (nx25167)) ;
    inv02 ix23692 (.Y (nx23693), .A (nx25167)) ;
    inv02 ix23694 (.Y (nx23695), .A (nx25167)) ;
    inv02 ix23696 (.Y (nx23697), .A (nx25169)) ;
    inv02 ix23698 (.Y (nx23699), .A (nx25169)) ;
    inv02 ix23700 (.Y (nx23701), .A (nx25169)) ;
    inv02 ix23702 (.Y (nx23703), .A (nx25169)) ;
    inv02 ix23704 (.Y (nx23705), .A (nx25169)) ;
    inv02 ix23706 (.Y (nx23707), .A (nx25169)) ;
    inv02 ix23708 (.Y (nx23709), .A (nx25169)) ;
    inv02 ix23710 (.Y (nx23711), .A (nx25171)) ;
    inv02 ix23712 (.Y (nx23713), .A (nx25171)) ;
    inv02 ix23714 (.Y (nx23715), .A (nx25171)) ;
    inv02 ix23716 (.Y (nx23717), .A (nx25171)) ;
    inv02 ix23718 (.Y (nx23719), .A (nx25171)) ;
    inv02 ix23720 (.Y (nx23721), .A (nx25171)) ;
    inv02 ix23722 (.Y (nx23723), .A (nx25171)) ;
    inv02 ix23724 (.Y (nx23725), .A (nx25173)) ;
    inv02 ix23726 (.Y (nx23727), .A (nx25173)) ;
    inv02 ix23728 (.Y (nx23729), .A (nx25173)) ;
    inv02 ix23730 (.Y (nx23731), .A (nx25173)) ;
    inv02 ix23732 (.Y (nx23733), .A (nx25173)) ;
    inv02 ix23734 (.Y (nx23735), .A (nx25173)) ;
    inv02 ix23736 (.Y (nx23737), .A (nx25173)) ;
    inv02 ix23738 (.Y (nx23739), .A (nx25175)) ;
    inv02 ix23740 (.Y (nx23741), .A (nx25175)) ;
    inv02 ix23742 (.Y (nx23743), .A (nx25175)) ;
    inv02 ix23744 (.Y (nx23745), .A (nx25175)) ;
    inv02 ix23746 (.Y (nx23747), .A (nx25175)) ;
    inv02 ix23748 (.Y (nx23749), .A (nx25175)) ;
    inv02 ix23750 (.Y (nx23751), .A (nx25175)) ;
    inv02 ix23752 (.Y (nx23753), .A (nx25177)) ;
    inv02 ix23754 (.Y (nx23755), .A (nx25177)) ;
    inv02 ix23756 (.Y (nx23757), .A (nx25177)) ;
    inv02 ix23758 (.Y (nx23759), .A (nx25177)) ;
    inv02 ix23760 (.Y (nx23761), .A (nx25177)) ;
    inv02 ix23762 (.Y (nx23763), .A (nx25177)) ;
    inv02 ix23764 (.Y (nx23765), .A (nx25177)) ;
    inv02 ix23766 (.Y (nx23767), .A (nx25179)) ;
    inv02 ix23768 (.Y (nx23769), .A (nx25179)) ;
    inv02 ix23770 (.Y (nx23771), .A (nx25179)) ;
    inv02 ix23772 (.Y (nx23773), .A (nx25179)) ;
    inv02 ix23774 (.Y (nx23775), .A (nx25179)) ;
    inv02 ix23776 (.Y (nx23777), .A (nx25179)) ;
    inv02 ix23778 (.Y (nx23779), .A (nx25179)) ;
    inv02 ix23780 (.Y (nx23781), .A (nx25181)) ;
    inv02 ix23782 (.Y (nx23783), .A (nx25181)) ;
    inv02 ix23784 (.Y (nx23785), .A (nx25181)) ;
    inv02 ix23786 (.Y (nx23787), .A (nx25181)) ;
    inv02 ix23788 (.Y (nx23789), .A (nx25181)) ;
    inv02 ix23790 (.Y (nx23791), .A (nx25181)) ;
    inv02 ix23792 (.Y (nx23793), .A (nx25181)) ;
    inv02 ix23794 (.Y (nx23795), .A (nx25183)) ;
    inv02 ix23796 (.Y (nx23797), .A (nx25183)) ;
    inv02 ix23798 (.Y (nx23799), .A (nx25183)) ;
    inv02 ix23800 (.Y (nx23801), .A (nx25183)) ;
    inv02 ix23802 (.Y (nx23803), .A (nx25183)) ;
    inv02 ix23804 (.Y (nx23805), .A (nx25183)) ;
    inv02 ix23806 (.Y (nx23807), .A (nx25183)) ;
    inv02 ix23808 (.Y (nx23809), .A (nx25185)) ;
    inv02 ix23810 (.Y (nx23811), .A (nx25185)) ;
    inv02 ix23812 (.Y (nx23813), .A (nx25185)) ;
    inv02 ix23814 (.Y (nx23815), .A (nx25185)) ;
    inv02 ix23816 (.Y (nx23817), .A (nx25185)) ;
    inv02 ix23818 (.Y (nx23819), .A (nx25185)) ;
    inv02 ix23820 (.Y (nx23821), .A (nx25185)) ;
    inv02 ix23822 (.Y (nx23823), .A (nx25187)) ;
    inv02 ix23824 (.Y (nx23825), .A (nx25187)) ;
    inv02 ix23826 (.Y (nx23827), .A (nx25187)) ;
    inv02 ix23828 (.Y (nx23829), .A (nx25187)) ;
    inv02 ix23830 (.Y (nx23831), .A (nx25187)) ;
    inv02 ix23832 (.Y (nx23833), .A (nx25187)) ;
    inv02 ix23834 (.Y (nx23835), .A (nx25187)) ;
    inv02 ix23836 (.Y (nx23837), .A (nx25189)) ;
    inv02 ix23838 (.Y (nx23839), .A (nx25189)) ;
    inv02 ix23840 (.Y (nx23841), .A (nx25189)) ;
    inv02 ix23842 (.Y (nx23843), .A (nx25189)) ;
    inv02 ix23844 (.Y (nx23845), .A (nx25189)) ;
    inv02 ix23846 (.Y (nx23847), .A (nx25189)) ;
    inv02 ix23848 (.Y (nx23849), .A (nx25189)) ;
    inv02 ix23850 (.Y (nx23851), .A (nx25191)) ;
    inv02 ix23852 (.Y (nx23853), .A (nx25191)) ;
    inv02 ix23854 (.Y (nx23855), .A (nx25191)) ;
    inv02 ix23856 (.Y (nx23857), .A (nx25191)) ;
    inv02 ix23858 (.Y (nx23859), .A (nx25191)) ;
    inv02 ix23860 (.Y (nx23861), .A (nx25191)) ;
    inv02 ix23862 (.Y (nx23863), .A (nx25191)) ;
    inv02 ix23864 (.Y (nx23865), .A (nx25193)) ;
    inv02 ix23866 (.Y (nx23867), .A (nx25193)) ;
    inv02 ix23868 (.Y (nx23869), .A (nx25193)) ;
    inv02 ix23870 (.Y (nx23871), .A (nx25193)) ;
    inv02 ix23872 (.Y (nx23873), .A (nx25193)) ;
    inv02 ix23874 (.Y (nx23875), .A (nx25193)) ;
    inv02 ix23876 (.Y (nx23877), .A (nx25193)) ;
    inv02 ix23878 (.Y (nx23879), .A (nx25195)) ;
    inv02 ix23880 (.Y (nx23881), .A (nx25195)) ;
    inv02 ix23882 (.Y (nx23883), .A (nx24881)) ;
    inv02 ix23884 (.Y (nx23885), .A (nx24881)) ;
    inv02 ix23886 (.Y (nx23887), .A (nx24881)) ;
    inv02 ix23888 (.Y (nx23889), .A (nx24881)) ;
    inv02 ix23890 (.Y (nx23891), .A (nx24881)) ;
    inv02 ix23892 (.Y (nx23893), .A (nx24881)) ;
    inv02 ix23894 (.Y (nx23895), .A (nx24881)) ;
    inv02 ix23896 (.Y (nx23897), .A (nx24883)) ;
    inv02 ix23898 (.Y (nx23899), .A (nx24883)) ;
    inv02 ix23900 (.Y (nx23901), .A (nx24883)) ;
    inv02 ix23902 (.Y (nx23903), .A (nx24883)) ;
    inv02 ix23904 (.Y (nx23905), .A (nx24883)) ;
    inv02 ix23906 (.Y (nx23907), .A (nx24883)) ;
    inv02 ix23908 (.Y (nx23909), .A (nx24883)) ;
    inv02 ix23910 (.Y (nx23911), .A (nx24885)) ;
    inv02 ix23912 (.Y (nx23913), .A (nx24885)) ;
    inv02 ix23914 (.Y (nx23915), .A (nx24885)) ;
    inv02 ix23916 (.Y (nx23917), .A (nx24885)) ;
    inv02 ix23918 (.Y (nx23919), .A (nx24885)) ;
    inv02 ix23920 (.Y (nx23921), .A (nx24885)) ;
    inv02 ix23922 (.Y (nx23923), .A (nx24885)) ;
    inv02 ix23924 (.Y (nx23925), .A (nx24887)) ;
    inv02 ix23926 (.Y (nx23927), .A (nx24887)) ;
    inv02 ix23928 (.Y (nx23929), .A (nx24887)) ;
    inv02 ix23930 (.Y (nx23931), .A (nx24887)) ;
    inv02 ix23932 (.Y (nx23933), .A (nx24887)) ;
    inv02 ix23934 (.Y (nx23935), .A (nx24887)) ;
    inv02 ix23936 (.Y (nx23937), .A (nx24887)) ;
    inv02 ix23938 (.Y (nx23939), .A (nx24889)) ;
    inv02 ix23940 (.Y (nx23941), .A (nx24889)) ;
    inv02 ix23942 (.Y (nx23943), .A (nx24889)) ;
    inv02 ix23944 (.Y (nx23945), .A (nx24889)) ;
    inv02 ix23946 (.Y (nx23947), .A (nx24889)) ;
    inv02 ix23948 (.Y (nx23949), .A (nx24889)) ;
    inv02 ix23950 (.Y (nx23951), .A (nx24889)) ;
    inv02 ix23952 (.Y (nx23953), .A (nx24891)) ;
    inv02 ix23954 (.Y (nx23955), .A (nx24891)) ;
    inv02 ix23956 (.Y (nx23957), .A (nx24891)) ;
    inv02 ix23958 (.Y (nx23959), .A (nx24891)) ;
    inv02 ix23960 (.Y (nx23961), .A (nx24891)) ;
    inv02 ix23962 (.Y (nx23963), .A (nx24891)) ;
    inv02 ix23964 (.Y (nx23965), .A (nx24891)) ;
    inv02 ix23966 (.Y (nx23967), .A (nx24893)) ;
    inv02 ix23968 (.Y (nx23969), .A (nx24893)) ;
    inv02 ix23970 (.Y (nx23971), .A (nx24893)) ;
    inv02 ix23972 (.Y (nx23973), .A (nx24893)) ;
    inv02 ix23974 (.Y (nx23975), .A (nx24893)) ;
    inv02 ix23976 (.Y (nx23977), .A (nx24893)) ;
    inv02 ix23978 (.Y (nx23979), .A (nx24893)) ;
    inv02 ix23980 (.Y (nx23981), .A (nx24895)) ;
    inv02 ix23982 (.Y (nx23983), .A (nx24895)) ;
    inv02 ix23984 (.Y (nx23985), .A (nx24895)) ;
    inv02 ix23986 (.Y (nx23987), .A (nx24895)) ;
    inv02 ix23988 (.Y (nx23989), .A (nx24895)) ;
    inv02 ix23990 (.Y (nx23991), .A (nx24895)) ;
    inv02 ix23992 (.Y (nx23993), .A (nx24895)) ;
    inv02 ix23994 (.Y (nx23995), .A (nx24897)) ;
    inv02 ix23996 (.Y (nx23997), .A (nx24897)) ;
    inv02 ix23998 (.Y (nx23999), .A (nx24897)) ;
    inv02 ix24000 (.Y (nx24001), .A (nx24897)) ;
    inv02 ix24002 (.Y (nx24003), .A (nx24897)) ;
    inv02 ix24004 (.Y (nx24005), .A (nx24897)) ;
    inv02 ix24006 (.Y (nx24007), .A (nx24897)) ;
    inv02 ix24008 (.Y (nx24009), .A (nx24899)) ;
    inv02 ix24010 (.Y (nx24011), .A (nx24899)) ;
    inv02 ix24012 (.Y (nx24013), .A (nx24899)) ;
    inv02 ix24014 (.Y (nx24015), .A (nx24899)) ;
    inv02 ix24016 (.Y (nx24017), .A (nx24899)) ;
    inv02 ix24018 (.Y (nx24019), .A (nx24899)) ;
    inv02 ix24020 (.Y (nx24021), .A (nx24899)) ;
    inv02 ix24022 (.Y (nx24023), .A (nx24901)) ;
    inv02 ix24024 (.Y (nx24025), .A (nx24901)) ;
    inv02 ix24026 (.Y (nx24027), .A (nx24901)) ;
    inv02 ix24028 (.Y (nx24029), .A (nx24901)) ;
    inv02 ix24030 (.Y (nx24031), .A (nx24901)) ;
    inv02 ix24032 (.Y (nx24033), .A (nx24901)) ;
    inv02 ix24034 (.Y (nx24035), .A (nx24901)) ;
    inv02 ix24036 (.Y (nx24037), .A (nx24903)) ;
    inv02 ix24038 (.Y (nx24039), .A (nx24903)) ;
    inv02 ix24040 (.Y (nx24041), .A (nx24903)) ;
    inv02 ix24042 (.Y (nx24043), .A (nx24903)) ;
    inv02 ix24044 (.Y (nx24045), .A (nx24903)) ;
    inv02 ix24046 (.Y (nx24047), .A (nx24903)) ;
    inv02 ix24048 (.Y (nx24049), .A (nx24903)) ;
    inv02 ix24050 (.Y (nx24051), .A (nx24905)) ;
    inv02 ix24052 (.Y (nx24053), .A (nx24905)) ;
    inv02 ix24054 (.Y (nx24055), .A (nx24905)) ;
    inv02 ix24056 (.Y (nx24057), .A (nx24905)) ;
    inv02 ix24058 (.Y (nx24059), .A (nx24905)) ;
    inv02 ix24060 (.Y (nx24061), .A (nx24905)) ;
    inv02 ix24062 (.Y (nx24063), .A (nx24905)) ;
    inv02 ix24064 (.Y (nx24065), .A (nx24907)) ;
    inv02 ix24066 (.Y (nx24067), .A (nx24907)) ;
    inv02 ix24068 (.Y (nx24069), .A (nx24907)) ;
    inv02 ix24070 (.Y (nx24071), .A (nx24907)) ;
    inv02 ix24072 (.Y (nx24073), .A (nx24907)) ;
    inv02 ix24074 (.Y (nx24075), .A (nx24907)) ;
    inv02 ix24076 (.Y (nx24077), .A (nx24907)) ;
    inv02 ix24078 (.Y (nx24079), .A (nx24909)) ;
    inv02 ix24080 (.Y (nx24081), .A (nx24909)) ;
    inv02 ix24082 (.Y (nx24083), .A (nx24909)) ;
    inv02 ix24084 (.Y (nx24085), .A (nx24909)) ;
    inv02 ix24086 (.Y (nx24087), .A (nx24909)) ;
    inv02 ix24088 (.Y (nx24089), .A (nx24909)) ;
    inv02 ix24090 (.Y (nx24091), .A (nx24909)) ;
    inv02 ix24092 (.Y (nx24093), .A (nx24911)) ;
    inv02 ix24094 (.Y (nx24095), .A (nx24911)) ;
    inv02 ix24096 (.Y (nx24097), .A (nx24911)) ;
    inv02 ix24098 (.Y (nx24099), .A (nx24911)) ;
    inv02 ix24100 (.Y (nx24101), .A (nx24911)) ;
    inv02 ix24102 (.Y (nx24103), .A (nx24911)) ;
    inv02 ix24104 (.Y (nx24105), .A (nx24911)) ;
    inv02 ix24106 (.Y (nx24107), .A (nx24913)) ;
    inv02 ix24108 (.Y (nx24109), .A (nx24913)) ;
    inv02 ix24110 (.Y (nx24111), .A (nx24913)) ;
    inv02 ix24112 (.Y (nx24113), .A (nx24913)) ;
    inv02 ix24114 (.Y (nx24115), .A (nx24913)) ;
    inv02 ix24116 (.Y (nx24117), .A (nx24913)) ;
    inv02 ix24118 (.Y (nx24119), .A (nx24913)) ;
    inv02 ix24120 (.Y (nx24121), .A (nx24915)) ;
    inv02 ix24122 (.Y (nx24123), .A (nx24915)) ;
    inv02 ix24124 (.Y (nx24125), .A (nx24915)) ;
    inv02 ix24126 (.Y (nx24127), .A (nx24915)) ;
    inv02 ix24128 (.Y (nx24129), .A (nx24915)) ;
    inv02 ix24130 (.Y (nx24131), .A (nx24915)) ;
    inv02 ix24132 (.Y (nx24133), .A (nx24915)) ;
    inv02 ix24134 (.Y (nx24135), .A (nx24917)) ;
    inv02 ix24136 (.Y (nx24137), .A (nx24917)) ;
    inv02 ix24138 (.Y (nx24139), .A (nx24917)) ;
    inv02 ix24140 (.Y (nx24141), .A (nx24917)) ;
    inv02 ix24142 (.Y (nx24143), .A (nx24917)) ;
    inv02 ix24144 (.Y (nx24145), .A (nx24917)) ;
    inv02 ix24146 (.Y (nx24147), .A (nx24917)) ;
    inv02 ix24148 (.Y (nx24149), .A (nx24919)) ;
    inv02 ix24150 (.Y (nx24151), .A (nx24919)) ;
    inv02 ix24152 (.Y (nx24153), .A (nx24919)) ;
    inv02 ix24154 (.Y (nx24155), .A (nx24919)) ;
    inv02 ix24156 (.Y (nx24157), .A (nx24919)) ;
    inv02 ix24158 (.Y (nx24159), .A (nx24919)) ;
    inv02 ix24160 (.Y (nx24161), .A (nx24919)) ;
    inv02 ix24162 (.Y (nx24163), .A (nx24921)) ;
    inv02 ix24164 (.Y (nx24165), .A (nx24921)) ;
    inv02 ix24166 (.Y (nx24167), .A (nx24921)) ;
    inv02 ix24168 (.Y (nx24169), .A (nx24921)) ;
    inv02 ix24170 (.Y (nx24171), .A (nx24921)) ;
    inv02 ix24172 (.Y (nx24173), .A (nx24921)) ;
    inv02 ix24174 (.Y (nx24175), .A (nx24921)) ;
    inv02 ix24176 (.Y (nx24177), .A (nx24923)) ;
    inv02 ix24178 (.Y (nx24179), .A (nx24923)) ;
    inv02 ix24180 (.Y (nx24181), .A (nx24923)) ;
    inv02 ix24182 (.Y (nx24183), .A (nx24923)) ;
    inv02 ix24184 (.Y (nx24185), .A (nx24923)) ;
    inv02 ix24186 (.Y (nx24187), .A (nx24923)) ;
    inv02 ix24188 (.Y (nx24189), .A (nx24923)) ;
    inv02 ix24190 (.Y (nx24191), .A (nx24925)) ;
    inv02 ix24192 (.Y (nx24193), .A (nx24925)) ;
    inv02 ix24194 (.Y (nx24195), .A (nx24925)) ;
    inv02 ix24196 (.Y (nx24197), .A (nx24925)) ;
    inv02 ix24198 (.Y (nx24199), .A (nx24925)) ;
    inv02 ix24200 (.Y (nx24201), .A (nx24925)) ;
    inv02 ix24202 (.Y (nx24203), .A (nx24925)) ;
    inv02 ix24204 (.Y (nx24205), .A (nx24927)) ;
    inv02 ix24206 (.Y (nx24207), .A (nx24927)) ;
    inv02 ix24208 (.Y (nx24209), .A (nx24927)) ;
    inv02 ix24210 (.Y (nx24211), .A (nx24927)) ;
    inv02 ix24212 (.Y (nx24213), .A (nx24927)) ;
    inv02 ix24214 (.Y (nx24215), .A (nx24927)) ;
    inv02 ix24216 (.Y (nx24217), .A (nx24927)) ;
    inv02 ix24218 (.Y (nx24219), .A (nx24929)) ;
    inv02 ix24220 (.Y (nx24221), .A (nx24929)) ;
    inv02 ix24222 (.Y (nx24223), .A (nx24929)) ;
    inv02 ix24224 (.Y (nx24225), .A (nx24929)) ;
    inv02 ix24226 (.Y (nx24227), .A (nx24929)) ;
    inv02 ix24228 (.Y (nx24229), .A (nx24929)) ;
    inv02 ix24230 (.Y (nx24231), .A (nx24929)) ;
    inv02 ix24232 (.Y (nx24233), .A (nx24931)) ;
    inv02 ix24234 (.Y (nx24235), .A (nx24931)) ;
    inv02 ix24236 (.Y (nx24237), .A (nx24931)) ;
    inv02 ix24238 (.Y (nx24239), .A (nx24931)) ;
    inv02 ix24240 (.Y (nx24241), .A (nx24931)) ;
    inv02 ix24242 (.Y (nx24243), .A (nx24931)) ;
    inv02 ix24244 (.Y (nx24245), .A (nx24931)) ;
    inv02 ix24246 (.Y (nx24247), .A (nx24933)) ;
    inv02 ix24248 (.Y (nx24249), .A (nx24933)) ;
    inv02 ix24250 (.Y (nx24251), .A (nx24933)) ;
    inv02 ix24252 (.Y (nx24253), .A (nx24933)) ;
    inv02 ix24254 (.Y (nx24255), .A (nx24933)) ;
    inv02 ix24256 (.Y (nx24257), .A (nx24933)) ;
    inv02 ix24258 (.Y (nx24259), .A (nx24933)) ;
    inv02 ix24260 (.Y (nx24261), .A (nx24935)) ;
    inv02 ix24262 (.Y (nx24263), .A (nx24935)) ;
    inv02 ix24264 (.Y (nx24265), .A (nx24935)) ;
    inv02 ix24266 (.Y (nx24267), .A (nx24935)) ;
    inv02 ix24268 (.Y (nx24269), .A (nx24935)) ;
    inv02 ix24270 (.Y (nx24271), .A (nx24935)) ;
    inv02 ix24272 (.Y (nx24273), .A (nx24935)) ;
    inv02 ix24274 (.Y (nx24275), .A (nx24937)) ;
    inv02 ix24276 (.Y (nx24277), .A (nx24937)) ;
    inv02 ix24278 (.Y (nx24279), .A (nx24937)) ;
    inv02 ix24280 (.Y (nx24281), .A (nx24937)) ;
    inv02 ix24282 (.Y (nx24283), .A (nx24937)) ;
    inv02 ix24284 (.Y (nx24285), .A (nx24937)) ;
    inv02 ix24286 (.Y (nx24287), .A (nx24937)) ;
    inv02 ix24288 (.Y (nx24289), .A (nx24939)) ;
    inv02 ix24290 (.Y (nx24291), .A (nx24939)) ;
    inv02 ix24292 (.Y (nx24293), .A (nx24939)) ;
    inv02 ix24294 (.Y (nx24295), .A (nx24939)) ;
    inv02 ix24296 (.Y (nx24297), .A (nx24939)) ;
    inv02 ix24298 (.Y (nx24299), .A (nx24939)) ;
    inv02 ix24300 (.Y (nx24301), .A (nx24939)) ;
    inv02 ix24302 (.Y (nx24303), .A (nx24941)) ;
    inv02 ix24304 (.Y (nx24305), .A (nx24941)) ;
    inv02 ix24306 (.Y (nx24307), .A (nx24941)) ;
    inv02 ix24308 (.Y (nx24309), .A (nx24941)) ;
    inv02 ix24310 (.Y (nx24311), .A (nx24941)) ;
    inv02 ix24312 (.Y (nx24313), .A (nx24941)) ;
    inv02 ix24314 (.Y (nx24315), .A (nx24941)) ;
    inv02 ix24316 (.Y (nx24317), .A (nx24943)) ;
    inv02 ix24318 (.Y (nx24319), .A (nx24943)) ;
    inv02 ix24320 (.Y (nx24321), .A (nx24943)) ;
    inv02 ix24322 (.Y (nx24323), .A (nx24943)) ;
    inv02 ix24324 (.Y (nx24325), .A (nx24943)) ;
    inv02 ix24326 (.Y (nx24327), .A (nx24943)) ;
    inv02 ix24328 (.Y (nx24329), .A (nx24943)) ;
    inv02 ix24330 (.Y (nx24331), .A (nx24945)) ;
    inv02 ix24332 (.Y (nx24333), .A (nx24945)) ;
    inv02 ix24334 (.Y (nx24335), .A (nx24945)) ;
    inv02 ix24336 (.Y (nx24337), .A (nx24945)) ;
    inv02 ix24338 (.Y (nx24339), .A (nx24945)) ;
    inv02 ix24340 (.Y (nx24341), .A (nx24945)) ;
    inv02 ix24342 (.Y (nx24343), .A (nx24945)) ;
    inv02 ix24344 (.Y (nx24345), .A (nx24947)) ;
    inv02 ix24346 (.Y (nx24347), .A (nx24947)) ;
    inv02 ix24348 (.Y (nx24349), .A (nx24947)) ;
    inv02 ix24350 (.Y (nx24351), .A (nx24947)) ;
    inv02 ix24352 (.Y (nx24353), .A (nx24947)) ;
    inv02 ix24354 (.Y (nx24355), .A (nx24947)) ;
    inv02 ix24356 (.Y (nx24357), .A (nx24947)) ;
    inv02 ix24358 (.Y (nx24359), .A (nx24949)) ;
    inv02 ix24360 (.Y (nx24361), .A (nx24949)) ;
    inv02 ix24362 (.Y (nx24363), .A (nx24949)) ;
    inv02 ix24364 (.Y (nx24365), .A (nx24949)) ;
    inv02 ix24366 (.Y (nx24367), .A (nx24949)) ;
    inv02 ix24368 (.Y (nx24369), .A (nx24949)) ;
    inv02 ix24370 (.Y (nx24371), .A (nx24949)) ;
    inv02 ix24372 (.Y (nx24373), .A (nx24951)) ;
    inv02 ix24374 (.Y (nx24375), .A (nx24951)) ;
    inv02 ix24376 (.Y (nx24377), .A (nx24951)) ;
    inv02 ix24378 (.Y (nx24379), .A (nx24951)) ;
    inv02 ix24380 (.Y (nx24381), .A (nx24951)) ;
    inv02 ix24382 (.Y (nx24383), .A (nx24951)) ;
    inv02 ix24384 (.Y (nx24385), .A (nx24951)) ;
    inv02 ix24386 (.Y (nx24387), .A (nx24953)) ;
    inv02 ix24388 (.Y (nx24389), .A (nx24953)) ;
    inv02 ix24390 (.Y (nx24391), .A (nx24953)) ;
    inv02 ix24392 (.Y (nx24393), .A (nx24953)) ;
    inv02 ix24394 (.Y (nx24395), .A (nx24953)) ;
    inv02 ix24396 (.Y (nx24397), .A (nx24953)) ;
    inv02 ix24398 (.Y (nx24399), .A (nx24953)) ;
    inv02 ix24400 (.Y (nx24401), .A (nx24955)) ;
    inv02 ix24402 (.Y (nx24403), .A (nx24955)) ;
    inv02 ix24404 (.Y (nx24405), .A (nx24955)) ;
    inv02 ix24406 (.Y (nx24407), .A (nx24955)) ;
    inv02 ix24408 (.Y (nx24409), .A (nx24955)) ;
    inv02 ix24410 (.Y (nx24411), .A (nx24955)) ;
    inv02 ix24412 (.Y (nx24413), .A (nx24955)) ;
    inv02 ix24414 (.Y (nx24415), .A (nx24957)) ;
    inv02 ix24416 (.Y (nx24417), .A (nx24957)) ;
    inv02 ix24418 (.Y (nx24419), .A (nx24957)) ;
    inv02 ix24420 (.Y (nx24421), .A (nx24957)) ;
    inv02 ix24422 (.Y (nx24423), .A (nx24957)) ;
    inv02 ix24424 (.Y (nx24425), .A (nx24957)) ;
    inv02 ix24426 (.Y (nx24427), .A (nx24957)) ;
    inv02 ix24428 (.Y (nx24429), .A (nx24959)) ;
    inv02 ix24430 (.Y (nx24431), .A (nx24959)) ;
    inv02 ix24432 (.Y (nx24433), .A (nx24959)) ;
    inv02 ix24434 (.Y (nx24435), .A (nx24959)) ;
    inv02 ix24436 (.Y (nx24437), .A (nx24959)) ;
    inv02 ix24438 (.Y (nx24439), .A (nx24959)) ;
    inv02 ix24440 (.Y (nx24441), .A (nx24959)) ;
    inv02 ix24442 (.Y (nx24443), .A (nx24961)) ;
    inv02 ix24444 (.Y (nx24445), .A (nx24961)) ;
    inv02 ix24446 (.Y (nx24447), .A (nx24961)) ;
    inv02 ix24448 (.Y (nx24449), .A (nx24961)) ;
    inv02 ix24450 (.Y (nx24451), .A (nx24961)) ;
    inv02 ix24452 (.Y (nx24453), .A (nx24961)) ;
    inv02 ix24454 (.Y (nx24455), .A (nx24961)) ;
    inv02 ix24456 (.Y (nx24457), .A (nx24963)) ;
    inv02 ix24458 (.Y (nx24459), .A (nx24963)) ;
    inv02 ix24460 (.Y (nx24461), .A (nx24963)) ;
    inv02 ix24462 (.Y (nx24463), .A (nx24963)) ;
    inv02 ix24464 (.Y (nx24465), .A (nx24963)) ;
    inv02 ix24466 (.Y (nx24467), .A (nx24963)) ;
    inv02 ix24468 (.Y (nx24469), .A (nx24963)) ;
    inv02 ix24470 (.Y (nx24471), .A (nx24965)) ;
    inv02 ix24472 (.Y (nx24473), .A (nx24965)) ;
    inv02 ix24474 (.Y (nx24475), .A (nx24965)) ;
    inv02 ix24476 (.Y (nx24477), .A (nx24965)) ;
    inv02 ix24478 (.Y (nx24479), .A (nx24965)) ;
    inv02 ix24480 (.Y (nx24481), .A (nx24965)) ;
    inv02 ix24482 (.Y (nx24483), .A (nx24965)) ;
    inv02 ix24484 (.Y (nx24485), .A (nx24967)) ;
    inv02 ix24486 (.Y (nx24487), .A (nx24967)) ;
    inv02 ix24488 (.Y (nx24489), .A (nx24967)) ;
    inv02 ix24490 (.Y (nx24491), .A (nx24967)) ;
    inv02 ix24492 (.Y (nx24493), .A (nx24967)) ;
    inv02 ix24494 (.Y (nx24495), .A (nx24967)) ;
    inv02 ix24496 (.Y (nx24497), .A (nx24967)) ;
    inv02 ix24498 (.Y (nx24499), .A (nx24969)) ;
    inv02 ix24500 (.Y (nx24501), .A (nx24969)) ;
    inv02 ix24502 (.Y (nx24503), .A (nx24969)) ;
    inv02 ix24504 (.Y (nx24505), .A (nx24969)) ;
    inv02 ix24506 (.Y (nx24507), .A (nx24969)) ;
    inv02 ix24508 (.Y (nx24509), .A (nx24969)) ;
    inv02 ix24510 (.Y (nx24511), .A (nx24969)) ;
    inv02 ix24512 (.Y (nx24513), .A (nx24971)) ;
    inv02 ix24514 (.Y (nx24515), .A (nx24971)) ;
    inv02 ix24516 (.Y (nx24517), .A (nx24971)) ;
    inv02 ix24518 (.Y (nx24519), .A (nx24971)) ;
    inv02 ix24520 (.Y (nx24521), .A (nx24971)) ;
    inv02 ix24522 (.Y (nx24523), .A (nx24971)) ;
    inv02 ix24524 (.Y (nx24525), .A (nx24971)) ;
    inv02 ix24526 (.Y (nx24527), .A (nx24973)) ;
    inv02 ix24528 (.Y (nx24529), .A (nx24973)) ;
    inv02 ix24530 (.Y (nx24531), .A (nx24973)) ;
    inv02 ix24532 (.Y (nx24533), .A (nx24973)) ;
    inv02 ix24534 (.Y (nx24535), .A (nx24973)) ;
    inv02 ix24536 (.Y (nx24537), .A (nx24973)) ;
    inv02 ix24538 (.Y (nx24539), .A (nx24973)) ;
    inv02 ix24540 (.Y (nx24541), .A (nx24975)) ;
    inv02 ix24542 (.Y (nx24543), .A (nx24975)) ;
    inv02 ix24544 (.Y (nx24545), .A (nx24975)) ;
    inv02 ix24546 (.Y (nx24547), .A (nx24975)) ;
    inv02 ix24548 (.Y (nx24549), .A (nx24975)) ;
    inv02 ix24550 (.Y (nx24551), .A (nx24975)) ;
    inv02 ix24552 (.Y (nx24553), .A (nx24975)) ;
    inv02 ix24554 (.Y (nx24555), .A (nx24977)) ;
    inv02 ix24556 (.Y (nx24557), .A (nx24977)) ;
    inv02 ix24558 (.Y (nx24559), .A (nx24977)) ;
    inv02 ix24560 (.Y (nx24561), .A (nx24977)) ;
    inv02 ix24562 (.Y (nx24563), .A (nx24977)) ;
    inv02 ix24564 (.Y (nx24565), .A (nx24977)) ;
    inv02 ix24566 (.Y (nx24567), .A (nx24977)) ;
    inv02 ix24568 (.Y (nx24569), .A (nx24979)) ;
    inv02 ix24570 (.Y (nx24571), .A (nx24979)) ;
    inv02 ix24572 (.Y (nx24573), .A (nx24979)) ;
    inv02 ix24574 (.Y (nx24575), .A (nx24979)) ;
    inv02 ix24576 (.Y (nx24577), .A (nx24979)) ;
    inv02 ix24578 (.Y (nx24579), .A (nx24979)) ;
    inv02 ix24580 (.Y (nx24581), .A (nx24979)) ;
    inv02 ix24582 (.Y (nx24583), .A (nx24981)) ;
    inv02 ix24584 (.Y (nx24585), .A (nx24981)) ;
    inv02 ix24586 (.Y (nx24587), .A (nx24981)) ;
    inv02 ix24588 (.Y (nx24589), .A (nx24981)) ;
    inv02 ix24590 (.Y (nx24591), .A (nx24981)) ;
    inv02 ix24592 (.Y (nx24593), .A (nx24981)) ;
    inv02 ix24594 (.Y (nx24595), .A (nx24981)) ;
    inv02 ix24596 (.Y (nx24597), .A (nx24983)) ;
    inv02 ix24598 (.Y (nx24599), .A (nx24983)) ;
    inv02 ix24600 (.Y (nx24601), .A (nx24983)) ;
    inv02 ix24602 (.Y (nx24603), .A (nx24983)) ;
    inv02 ix24604 (.Y (nx24605), .A (nx24983)) ;
    inv02 ix24606 (.Y (nx24607), .A (nx24983)) ;
    inv02 ix24608 (.Y (nx24609), .A (nx24983)) ;
    inv02 ix24610 (.Y (nx24611), .A (nx24985)) ;
    inv02 ix24612 (.Y (nx24613), .A (nx24985)) ;
    inv02 ix24614 (.Y (nx24615), .A (nx24985)) ;
    inv02 ix24616 (.Y (nx24617), .A (nx24985)) ;
    inv02 ix24618 (.Y (nx24619), .A (nx24985)) ;
    inv02 ix24620 (.Y (nx24621), .A (nx24985)) ;
    inv02 ix24622 (.Y (nx24623), .A (nx24985)) ;
    inv02 ix24624 (.Y (nx24625), .A (nx24987)) ;
    inv02 ix24626 (.Y (nx24627), .A (nx24987)) ;
    inv02 ix24628 (.Y (nx24629), .A (nx24987)) ;
    inv02 ix24630 (.Y (nx24631), .A (nx24987)) ;
    inv02 ix24632 (.Y (nx24633), .A (nx24987)) ;
    inv02 ix24634 (.Y (nx24635), .A (nx24987)) ;
    inv02 ix24636 (.Y (nx24637), .A (nx24987)) ;
    inv02 ix24638 (.Y (nx24639), .A (nx24989)) ;
    inv02 ix24640 (.Y (nx24641), .A (nx24989)) ;
    inv02 ix24642 (.Y (nx24643), .A (nx24989)) ;
    inv02 ix24644 (.Y (nx24645), .A (nx24989)) ;
    inv02 ix24646 (.Y (nx24647), .A (nx24989)) ;
    inv02 ix24648 (.Y (nx24649), .A (nx24989)) ;
    inv02 ix24650 (.Y (nx24651), .A (nx24989)) ;
    inv02 ix24652 (.Y (nx24653), .A (nx24991)) ;
    inv02 ix24654 (.Y (nx24655), .A (nx24991)) ;
    inv02 ix24656 (.Y (nx24657), .A (nx24991)) ;
    inv02 ix24658 (.Y (nx24659), .A (nx24991)) ;
    inv02 ix24660 (.Y (nx24661), .A (nx24991)) ;
    inv02 ix24662 (.Y (nx24663), .A (nx24991)) ;
    inv02 ix24664 (.Y (nx24665), .A (nx24991)) ;
    inv02 ix24666 (.Y (nx24667), .A (nx24993)) ;
    inv02 ix24668 (.Y (nx24669), .A (nx24993)) ;
    inv02 ix24670 (.Y (nx24671), .A (nx24993)) ;
    inv02 ix24672 (.Y (nx24673), .A (nx24993)) ;
    inv02 ix24674 (.Y (nx24675), .A (nx24993)) ;
    inv02 ix24676 (.Y (nx24677), .A (nx24993)) ;
    inv02 ix24678 (.Y (nx24679), .A (nx24993)) ;
    inv02 ix24680 (.Y (nx24681), .A (nx24995)) ;
    inv02 ix24682 (.Y (nx24683), .A (nx24995)) ;
    inv02 ix24684 (.Y (nx24685), .A (nx24995)) ;
    inv02 ix24686 (.Y (nx24687), .A (nx24995)) ;
    inv02 ix24688 (.Y (nx24689), .A (nx24995)) ;
    inv02 ix24690 (.Y (nx24691), .A (nx24995)) ;
    inv02 ix24692 (.Y (nx24693), .A (nx24995)) ;
    inv02 ix24694 (.Y (nx24695), .A (nx24997)) ;
    inv02 ix24696 (.Y (nx24697), .A (nx24997)) ;
    inv02 ix24698 (.Y (nx24699), .A (nx24997)) ;
    inv02 ix24700 (.Y (nx24701), .A (nx24997)) ;
    inv02 ix24702 (.Y (nx24703), .A (nx24997)) ;
    inv02 ix24704 (.Y (nx24705), .A (nx24997)) ;
    inv02 ix24706 (.Y (nx24707), .A (nx24997)) ;
    inv02 ix24708 (.Y (nx24709), .A (nx24999)) ;
    inv02 ix24710 (.Y (nx24711), .A (nx24999)) ;
    inv02 ix24712 (.Y (nx24713), .A (nx24999)) ;
    inv02 ix24714 (.Y (nx24715), .A (nx24999)) ;
    inv02 ix24716 (.Y (nx24717), .A (nx24999)) ;
    inv02 ix24718 (.Y (nx24719), .A (nx24999)) ;
    inv02 ix24720 (.Y (nx24721), .A (nx24999)) ;
    inv02 ix24722 (.Y (nx24723), .A (nx25001)) ;
    inv02 ix24724 (.Y (nx24725), .A (nx25001)) ;
    inv02 ix24726 (.Y (nx24727), .A (nx25001)) ;
    inv02 ix24728 (.Y (nx24729), .A (nx25001)) ;
    inv02 ix24730 (.Y (nx24731), .A (nx25001)) ;
    inv02 ix24732 (.Y (nx24733), .A (nx25001)) ;
    inv02 ix24734 (.Y (nx24735), .A (nx25001)) ;
    inv02 ix24736 (.Y (nx24737), .A (nx25003)) ;
    inv02 ix24738 (.Y (nx24739), .A (nx25003)) ;
    inv02 ix24740 (.Y (nx24741), .A (nx25003)) ;
    inv02 ix24742 (.Y (nx24743), .A (nx25003)) ;
    inv02 ix24744 (.Y (nx24745), .A (nx25003)) ;
    inv02 ix24746 (.Y (nx24747), .A (nx25003)) ;
    inv02 ix24748 (.Y (nx24749), .A (nx25003)) ;
    inv02 ix24750 (.Y (nx24751), .A (nx25005)) ;
    inv02 ix24752 (.Y (nx24753), .A (nx25005)) ;
    inv02 ix24754 (.Y (nx24755), .A (nx25005)) ;
    inv02 ix24756 (.Y (nx24757), .A (nx25005)) ;
    inv02 ix24758 (.Y (nx24759), .A (nx25005)) ;
    inv02 ix24760 (.Y (nx24761), .A (nx25005)) ;
    inv02 ix24762 (.Y (nx24763), .A (nx25005)) ;
    inv02 ix24764 (.Y (nx24765), .A (nx25007)) ;
    inv02 ix24766 (.Y (nx24767), .A (nx25007)) ;
    inv02 ix24768 (.Y (nx24769), .A (nx25007)) ;
    inv02 ix24770 (.Y (nx24771), .A (nx25007)) ;
    inv02 ix24772 (.Y (nx24773), .A (nx25007)) ;
    inv02 ix24774 (.Y (nx24775), .A (nx25007)) ;
    inv02 ix24776 (.Y (nx24777), .A (nx25007)) ;
    inv02 ix24778 (.Y (nx24779), .A (nx25009)) ;
    inv02 ix24780 (.Y (nx24781), .A (nx25009)) ;
    inv02 ix24782 (.Y (nx24783), .A (nx25009)) ;
    inv02 ix24784 (.Y (nx24785), .A (nx25009)) ;
    inv02 ix24786 (.Y (nx24787), .A (nx25009)) ;
    inv02 ix24788 (.Y (nx24789), .A (nx25009)) ;
    inv02 ix24790 (.Y (nx24791), .A (nx25009)) ;
    inv02 ix24792 (.Y (nx24793), .A (nx25011)) ;
    inv02 ix24794 (.Y (nx24795), .A (nx25011)) ;
    inv02 ix24796 (.Y (nx24797), .A (nx25011)) ;
    inv02 ix24798 (.Y (nx24799), .A (nx25011)) ;
    inv02 ix24800 (.Y (nx24801), .A (nx25011)) ;
    inv02 ix24802 (.Y (nx24803), .A (nx25011)) ;
    inv02 ix24804 (.Y (nx24805), .A (nx25011)) ;
    inv02 ix24806 (.Y (nx24807), .A (nx25013)) ;
    inv02 ix24808 (.Y (nx24809), .A (nx25013)) ;
    inv02 ix24810 (.Y (nx24811), .A (nx25013)) ;
    inv02 ix24812 (.Y (nx24813), .A (nx25013)) ;
    inv02 ix24814 (.Y (nx24815), .A (nx25013)) ;
    inv02 ix24816 (.Y (nx24817), .A (nx25013)) ;
    inv02 ix24818 (.Y (nx24819), .A (nx25013)) ;
    inv02 ix24820 (.Y (nx24821), .A (nx25015)) ;
    inv02 ix24822 (.Y (nx24823), .A (nx25015)) ;
    inv02 ix24824 (.Y (nx24825), .A (nx25015)) ;
    inv02 ix24826 (.Y (nx24827), .A (nx25015)) ;
    inv02 ix24828 (.Y (nx24829), .A (nx25015)) ;
    inv02 ix24830 (.Y (nx24831), .A (nx25015)) ;
    inv02 ix24832 (.Y (nx24833), .A (nx25015)) ;
    inv02 ix24834 (.Y (nx24835), .A (nx22379)) ;
    inv02 ix24836 (.Y (nx24837), .A (nx22379)) ;
    inv02 ix24838 (.Y (nx24839), .A (selectionLines[3])) ;
    inv02 ix24840 (.Y (nx24841), .A (selectionLines[3])) ;
    inv02 ix24842 (.Y (nx24843), .A (selectionLines[3])) ;
    inv02 ix24844 (.Y (nx24845), .A (selectionLines[3])) ;
    inv02 ix24846 (.Y (nx24847), .A (selectionLines[3])) ;
    inv02 ix24848 (.Y (nx24849), .A (selectionLines[3])) ;
    inv02 ix24850 (.Y (nx24851), .A (selectionLines[8])) ;
    inv02 ix24852 (.Y (nx24853), .A (selectionLines[8])) ;
    inv02 ix24854 (.Y (nx24855), .A (nx25227)) ;
    inv02 ix24856 (.Y (nx24857), .A (nx25227)) ;
    inv02 ix24858 (.Y (nx24859), .A (nx25227)) ;
    inv02 ix24860 (.Y (nx24861), .A (nx25227)) ;
    inv02 ix24862 (.Y (nx24863), .A (nx25227)) ;
    inv02 ix24864 (.Y (nx24865), .A (nx25227)) ;
    inv02 ix24866 (.Y (nx24867), .A (nx25227)) ;
    inv02 ix24868 (.Y (nx24869), .A (nx25229)) ;
    inv02 ix24870 (.Y (nx24871), .A (nx25229)) ;
    inv02 ix24872 (.Y (nx24873), .A (nx25229)) ;
    inv02 ix24874 (.Y (nx24875), .A (nx25229)) ;
    inv02 ix24876 (.Y (nx24877), .A (nx25229)) ;
    inv02 ix24878 (.Y (nx24879), .A (nx25231)) ;
    inv02 ix24880 (.Y (nx24881), .A (nx25231)) ;
    inv02 ix24882 (.Y (nx24883), .A (nx25231)) ;
    inv02 ix24884 (.Y (nx24885), .A (nx25231)) ;
    inv02 ix24886 (.Y (nx24887), .A (nx25231)) ;
    inv02 ix24888 (.Y (nx24889), .A (nx25231)) ;
    inv02 ix24890 (.Y (nx24891), .A (nx25231)) ;
    inv02 ix24892 (.Y (nx24893), .A (nx25233)) ;
    inv02 ix24894 (.Y (nx24895), .A (nx25233)) ;
    inv02 ix24896 (.Y (nx24897), .A (nx25233)) ;
    inv02 ix24898 (.Y (nx24899), .A (nx25233)) ;
    inv02 ix24900 (.Y (nx24901), .A (nx25233)) ;
    inv02 ix24902 (.Y (nx24903), .A (nx25233)) ;
    inv02 ix24904 (.Y (nx24905), .A (nx25233)) ;
    inv02 ix24906 (.Y (nx24907), .A (nx25235)) ;
    inv02 ix24908 (.Y (nx24909), .A (nx25235)) ;
    inv02 ix24910 (.Y (nx24911), .A (nx25235)) ;
    inv02 ix24912 (.Y (nx24913), .A (nx25235)) ;
    inv02 ix24914 (.Y (nx24915), .A (nx25235)) ;
    inv02 ix24916 (.Y (nx24917), .A (nx25235)) ;
    inv02 ix24918 (.Y (nx24919), .A (nx25235)) ;
    inv02 ix24920 (.Y (nx24921), .A (nx25237)) ;
    inv02 ix24922 (.Y (nx24923), .A (nx25237)) ;
    inv02 ix24924 (.Y (nx24925), .A (nx25237)) ;
    inv02 ix24926 (.Y (nx24927), .A (nx25237)) ;
    inv02 ix24928 (.Y (nx24929), .A (nx25237)) ;
    inv02 ix24930 (.Y (nx24931), .A (nx25237)) ;
    inv02 ix24932 (.Y (nx24933), .A (nx25237)) ;
    inv02 ix24934 (.Y (nx24935), .A (nx25239)) ;
    inv02 ix24936 (.Y (nx24937), .A (nx25239)) ;
    inv02 ix24938 (.Y (nx24939), .A (nx25239)) ;
    inv02 ix24940 (.Y (nx24941), .A (nx25239)) ;
    inv02 ix24942 (.Y (nx24943), .A (nx25239)) ;
    inv02 ix24944 (.Y (nx24945), .A (nx25239)) ;
    inv02 ix24946 (.Y (nx24947), .A (nx25239)) ;
    inv02 ix24948 (.Y (nx24949), .A (nx25241)) ;
    inv02 ix24950 (.Y (nx24951), .A (nx25241)) ;
    inv02 ix24952 (.Y (nx24953), .A (nx25241)) ;
    inv02 ix24954 (.Y (nx24955), .A (nx25241)) ;
    inv02 ix24956 (.Y (nx24957), .A (nx25241)) ;
    inv02 ix24958 (.Y (nx24959), .A (nx25241)) ;
    inv02 ix24960 (.Y (nx24961), .A (nx25241)) ;
    inv02 ix24962 (.Y (nx24963), .A (nx25243)) ;
    inv02 ix24964 (.Y (nx24965), .A (nx25243)) ;
    inv02 ix24966 (.Y (nx24967), .A (nx25243)) ;
    inv02 ix24968 (.Y (nx24969), .A (nx25243)) ;
    inv02 ix24970 (.Y (nx24971), .A (nx25243)) ;
    inv02 ix24972 (.Y (nx24973), .A (nx25243)) ;
    inv02 ix24974 (.Y (nx24975), .A (nx25243)) ;
    inv02 ix24976 (.Y (nx24977), .A (nx25245)) ;
    inv02 ix24978 (.Y (nx24979), .A (nx25245)) ;
    inv02 ix24980 (.Y (nx24981), .A (nx25245)) ;
    inv02 ix24982 (.Y (nx24983), .A (nx25245)) ;
    inv02 ix24984 (.Y (nx24985), .A (nx25245)) ;
    inv02 ix24986 (.Y (nx24987), .A (nx25245)) ;
    inv02 ix24988 (.Y (nx24989), .A (nx25245)) ;
    inv02 ix24990 (.Y (nx24991), .A (nx25247)) ;
    inv02 ix24992 (.Y (nx24993), .A (nx25247)) ;
    inv02 ix24994 (.Y (nx24995), .A (nx25247)) ;
    inv02 ix24996 (.Y (nx24997), .A (nx25247)) ;
    inv02 ix24998 (.Y (nx24999), .A (nx25247)) ;
    inv02 ix25000 (.Y (nx25001), .A (nx25247)) ;
    inv02 ix25002 (.Y (nx25003), .A (nx25247)) ;
    inv02 ix25004 (.Y (nx25005), .A (nx25249)) ;
    inv02 ix25006 (.Y (nx25007), .A (nx25249)) ;
    inv02 ix25008 (.Y (nx25009), .A (nx25249)) ;
    inv02 ix25010 (.Y (nx25011), .A (nx25249)) ;
    inv02 ix25012 (.Y (nx25013), .A (nx25249)) ;
    inv02 ix25014 (.Y (nx25015), .A (nx25249)) ;
    inv02 ix25016 (.Y (nx25017), .A (selectionLines[7])) ;
    inv02 ix25018 (.Y (nx25019), .A (selectionLines[7])) ;
    inv02 ix25020 (.Y (nx25021), .A (selectionLines[7])) ;
    inv02 ix25022 (.Y (nx25023), .A (selectionLines[6])) ;
    inv02 ix25024 (.Y (nx25025), .A (selectionLines[6])) ;
    inv02 ix25026 (.Y (nx25027), .A (selectionLines[6])) ;
    inv02 ix25028 (.Y (nx25029), .A (selectionLines[6])) ;
    inv02 ix25030 (.Y (nx25031), .A (selectionLines[6])) ;
    inv02 ix25032 (.Y (nx25033), .A (selectionLines[6])) ;
    inv02 ix25034 (.Y (nx25035), .A (selectionLines[5])) ;
    inv02 ix25036 (.Y (nx25037), .A (nx25201)) ;
    inv02 ix25038 (.Y (nx25039), .A (nx25201)) ;
    inv02 ix25040 (.Y (nx25041), .A (nx25201)) ;
    inv02 ix25042 (.Y (nx25043), .A (nx25201)) ;
    inv02 ix25044 (.Y (nx25045), .A (nx25201)) ;
    inv02 ix25046 (.Y (nx25047), .A (nx25201)) ;
    inv02 ix25048 (.Y (nx25049), .A (nx25201)) ;
    inv02 ix25050 (.Y (nx25051), .A (nx25203)) ;
    inv02 ix25052 (.Y (nx25053), .A (nx25203)) ;
    inv02 ix25054 (.Y (nx25055), .A (nx25203)) ;
    inv02 ix25056 (.Y (nx25057), .A (selectionLines[4])) ;
    inv02 ix25058 (.Y (nx25059), .A (nx25205)) ;
    inv02 ix25060 (.Y (nx25061), .A (nx25205)) ;
    inv02 ix25062 (.Y (nx25063), .A (nx25205)) ;
    inv02 ix25064 (.Y (nx25065), .A (nx25205)) ;
    inv02 ix25066 (.Y (nx25067), .A (nx25205)) ;
    inv02 ix25068 (.Y (nx25069), .A (nx25205)) ;
    inv02 ix25070 (.Y (nx25071), .A (nx25205)) ;
    inv02 ix25072 (.Y (nx25073), .A (nx25207)) ;
    inv02 ix25074 (.Y (nx25075), .A (nx25207)) ;
    inv02 ix25076 (.Y (nx25077), .A (nx25207)) ;
    inv02 ix25078 (.Y (nx25079), .A (nx25207)) ;
    inv02 ix25080 (.Y (nx25081), .A (nx25207)) ;
    inv02 ix25082 (.Y (nx25083), .A (nx25207)) ;
    inv02 ix25084 (.Y (nx25085), .A (nx25207)) ;
    inv02 ix25086 (.Y (nx25087), .A (nx25209)) ;
    inv02 ix25088 (.Y (nx25089), .A (nx25209)) ;
    inv02 ix25090 (.Y (nx25091), .A (nx25209)) ;
    inv02 ix25092 (.Y (nx25093), .A (nx25209)) ;
    inv02 ix25094 (.Y (nx25095), .A (nx25209)) ;
    inv02 ix25096 (.Y (nx25097), .A (nx25209)) ;
    inv02 ix25098 (.Y (nx25099), .A (nx25209)) ;
    inv02 ix25100 (.Y (nx25101), .A (nx25211)) ;
    inv02 ix25102 (.Y (nx25103), .A (nx25211)) ;
    inv02 ix25104 (.Y (nx25105), .A (nx25211)) ;
    inv02 ix25106 (.Y (nx25107), .A (nx25211)) ;
    inv02 ix25108 (.Y (nx25109), .A (nx25211)) ;
    inv02 ix25110 (.Y (nx25111), .A (nx25211)) ;
    inv02 ix25112 (.Y (nx25113), .A (nx25211)) ;
    inv02 ix25114 (.Y (nx25115), .A (nx25213)) ;
    inv02 ix25116 (.Y (nx25117), .A (nx25213)) ;
    inv02 ix25118 (.Y (nx25119), .A (nx25213)) ;
    inv02 ix25120 (.Y (nx25121), .A (selectionLines[1])) ;
    inv02 ix25122 (.Y (nx25123), .A (nx25215)) ;
    inv02 ix25124 (.Y (nx25125), .A (nx25215)) ;
    inv02 ix25126 (.Y (nx25127), .A (nx25215)) ;
    inv02 ix25128 (.Y (nx25129), .A (nx25215)) ;
    inv02 ix25130 (.Y (nx25131), .A (nx25215)) ;
    inv02 ix25132 (.Y (nx25133), .A (nx25215)) ;
    inv02 ix25134 (.Y (nx25135), .A (nx25215)) ;
    inv02 ix25136 (.Y (nx25137), .A (nx25217)) ;
    inv02 ix25138 (.Y (nx25139), .A (nx25217)) ;
    inv02 ix25140 (.Y (nx25141), .A (nx25217)) ;
    inv02 ix25142 (.Y (nx25143), .A (nx25217)) ;
    inv02 ix25144 (.Y (nx25145), .A (nx25217)) ;
    inv02 ix25146 (.Y (nx25147), .A (nx25217)) ;
    inv02 ix25148 (.Y (nx25149), .A (nx25217)) ;
    inv02 ix25150 (.Y (nx25151), .A (nx25219)) ;
    inv02 ix25152 (.Y (nx25153), .A (nx25219)) ;
    inv02 ix25154 (.Y (nx25155), .A (nx25219)) ;
    inv02 ix25156 (.Y (nx25157), .A (nx25219)) ;
    inv02 ix25158 (.Y (nx25159), .A (nx25219)) ;
    inv02 ix25160 (.Y (nx25161), .A (nx25219)) ;
    inv02 ix25162 (.Y (nx25163), .A (nx25219)) ;
    inv02 ix25164 (.Y (nx25165), .A (nx25221)) ;
    inv02 ix25166 (.Y (nx25167), .A (nx25221)) ;
    inv02 ix25168 (.Y (nx25169), .A (nx25221)) ;
    inv02 ix25170 (.Y (nx25171), .A (nx25221)) ;
    inv02 ix25172 (.Y (nx25173), .A (nx25221)) ;
    inv02 ix25174 (.Y (nx25175), .A (nx25221)) ;
    inv02 ix25176 (.Y (nx25177), .A (nx25221)) ;
    inv02 ix25178 (.Y (nx25179), .A (nx25223)) ;
    inv02 ix25180 (.Y (nx25181), .A (nx25223)) ;
    inv02 ix25182 (.Y (nx25183), .A (nx25223)) ;
    inv02 ix25184 (.Y (nx25185), .A (nx25223)) ;
    inv02 ix25186 (.Y (nx25187), .A (nx25223)) ;
    inv02 ix25188 (.Y (nx25189), .A (nx25223)) ;
    inv02 ix25190 (.Y (nx25191), .A (nx25223)) ;
    inv02 ix25192 (.Y (nx25193), .A (nx25225)) ;
    inv02 ix25194 (.Y (nx25195), .A (nx25225)) ;
    inv02 ix25200 (.Y (nx25201), .A (nx25035)) ;
    inv02 ix25202 (.Y (nx25203), .A (nx25035)) ;
    inv02 ix25204 (.Y (nx25205), .A (nx25057)) ;
    inv02 ix25206 (.Y (nx25207), .A (nx25057)) ;
    inv02 ix25208 (.Y (nx25209), .A (nx25057)) ;
    inv02 ix25210 (.Y (nx25211), .A (nx25057)) ;
    inv02 ix25212 (.Y (nx25213), .A (nx25057)) ;
    inv02 ix25214 (.Y (nx25215), .A (nx25121)) ;
    inv02 ix25216 (.Y (nx25217), .A (nx25121)) ;
    inv02 ix25218 (.Y (nx25219), .A (nx25121)) ;
    inv02 ix25220 (.Y (nx25221), .A (nx25121)) ;
    inv02 ix25222 (.Y (nx25223), .A (nx25121)) ;
    inv02 ix25224 (.Y (nx25225), .A (nx25121)) ;
    inv02 ix25226 (.Y (nx25227), .A (nx22227)) ;
    inv02 ix25228 (.Y (nx25229), .A (nx22227)) ;
    inv02 ix25230 (.Y (nx25231), .A (nx22379)) ;
    inv02 ix25232 (.Y (nx25233), .A (nx22379)) ;
    inv02 ix25234 (.Y (nx25235), .A (nx22379)) ;
    inv02 ix25236 (.Y (nx25237), .A (nx22379)) ;
    inv02 ix25238 (.Y (nx25239), .A (nx22379)) ;
    inv02 ix25240 (.Y (nx25241), .A (nx22379)) ;
    inv02 ix25242 (.Y (nx25243), .A (nx22379)) ;
    inv02 ix25244 (.Y (nx25245), .A (nx22379)) ;
    inv02 ix25246 (.Y (nx25247), .A (nx22379)) ;
    inv02 ix25248 (.Y (nx25249), .A (nx22379)) ;
endmodule


module Decoder_9 ( T, en, decoded ) ;

    input [8:0]T ;
    input en ;
    output [511:0]decoded ;

    wire nx12, nx18, nx38, nx48, nx56, nx66, nx72, nx78, nx84, nx94, nx100, 
         nx106, nx112, nx120, nx126, nx132, nx138, nx920, nx1196, nx3745, nx3748, 
         nx3752, nx3758, nx3764, nx3768, nx3780, nx3792, nx3803, nx3808, nx3810, 
         nx3812, nx3832, nx3854, nx3872, nx3874, nx3947, nx3949, nx4043, nx4061, 
         nx4079, nx4097, nx4099, nx4173, nx4175, nx4252, nx4254, nx4327, nx4329, 
         nx4406, nx4418, nx4430, nx4442, nx4454, nx4466, nx4478, nx4490, nx4502, 
         nx4514, nx4526, nx4538, nx4550, nx4562, nx4574, nx4586, nx4606, nx4614, 
         nx4622, nx4638, nx4646, nx4654, nx4670, nx4678, nx4686, nx4694, nx4734, 
         nx4742, nx4750, nx4766, nx4774, nx4782, nx4798, nx4806, nx4814, nx4830, 
         nx4838, nx4846, nx4858, nx4860, nx4862, nx4864, nx4866, nx4868, nx4870, 
         nx4872, nx4874, nx4876, nx4878, nx4880, nx4882, nx4884, nx4886, nx4888, 
         nx4890, nx4892, nx4894, nx4896, nx4898, nx4900, nx4902, nx4904, nx4906, 
         nx4908, nx4910, nx4912, nx4914, nx4916, nx4918, nx4920, nx4922, nx4924, 
         nx4926, nx4928, nx4930, nx4932, nx4934, nx4936, nx4938, nx4940, nx4942, 
         nx4944, nx4946, nx4948, nx4950, nx4952, nx4954, nx4956, nx4958, nx4960, 
         nx4962, nx4964, nx4966, nx4968, nx4970, nx4972, nx4974, nx4976, nx4978, 
         nx4980, nx4982, nx4984, nx4986, nx4988, nx4990, nx4992, nx4994, nx4996, 
         nx4998, nx5000, nx5002, nx5004, nx5006, nx5008, nx5010, nx5012, nx5014, 
         nx5016, nx5018, nx5020, nx5022, nx5024, nx5026, nx5028, nx5030, nx5032, 
         nx5034, nx5036, nx5038, nx5040, nx5042, nx5044, nx5046, nx5048, nx5050, 
         nx5052, nx5054, nx5056, nx5058, nx5060, nx5062, nx5064, nx5066, nx5068, 
         nx5070, nx5072, nx5074, nx5076, nx5078, nx5080, nx5082, nx5084, nx5086, 
         nx5088, nx5090, nx5092, nx5094, nx5096, nx5098, nx5100, nx5102, nx5104, 
         nx5106, nx5108, nx5110, nx5112, nx5114, nx5116, nx5118, nx5120, nx5122, 
         nx5124, nx5126, nx5128, nx5130, nx5132, nx5134, nx5136, nx5138, nx5140, 
         nx5142, nx5144, nx5146, nx5148, nx5150, nx5152, nx5154, nx5156, nx5158, 
         nx5160, nx5162, nx5164, nx5166, nx5168, nx5170, nx5172, nx5174, nx5176, 
         nx5178, nx5180, nx5182, nx5184, nx5186, nx5188, nx5190, nx5192, nx5194, 
         nx5196, nx5198, nx5200, nx5202, nx5204, nx5206, nx5208, nx5210, nx5212, 
         nx5214, nx5216, nx5218, nx5220, nx5222, nx5224, nx5226, nx5228;



    nand04 ix13 (.Y (nx12), .A0 (T[0]), .A1 (nx4864), .A2 (T[2]), .A3 (nx4862)
           ) ;
    or02 ix3746 (.Y (nx3745), .A0 (nx18), .A1 (nx3748)) ;
    nand02 ix19 (.Y (nx18), .A0 (T[4]), .A1 (T[5])) ;
    nand04 ix3749 (.Y (nx3748), .A0 (T[8]), .A1 (en), .A2 (nx4858), .A3 (nx4860)
           ) ;
    nand03 ix39 (.Y (nx38), .A0 (nx3752), .A1 (T[2]), .A2 (nx4862)) ;
    nand03 ix49 (.Y (nx48), .A0 (nx3758), .A1 (T[2]), .A2 (nx4862)) ;
    nand03 ix57 (.Y (nx56), .A0 (nx3764), .A1 (T[2]), .A2 (nx4862)) ;
    nor02_2x ix3765 (.Y (nx3764), .A0 (T[0]), .A1 (nx4864)) ;
    nand03 ix67 (.Y (nx66), .A0 (nx3768), .A1 (T[0]), .A2 (nx4864)) ;
    nand02 ix73 (.Y (nx72), .A0 (nx3768), .A1 (nx3752)) ;
    nand02 ix79 (.Y (nx78), .A0 (nx3768), .A1 (nx3758)) ;
    nand02 ix85 (.Y (nx84), .A0 (nx3768), .A1 (nx3764)) ;
    nand03 ix95 (.Y (nx94), .A0 (nx3780), .A1 (T[0]), .A2 (nx4864)) ;
    nand02 ix101 (.Y (nx100), .A0 (nx3780), .A1 (nx3752)) ;
    nand02 ix107 (.Y (nx106), .A0 (nx3780), .A1 (nx3758)) ;
    nand02 ix113 (.Y (nx112), .A0 (nx3780), .A1 (nx3764)) ;
    nand03 ix121 (.Y (nx120), .A0 (nx3792), .A1 (T[0]), .A2 (nx4864)) ;
    nor02_2x ix3793 (.Y (nx3792), .A0 (T[2]), .A1 (nx4862)) ;
    nand02 ix127 (.Y (nx126), .A0 (nx3792), .A1 (nx3752)) ;
    nand02 ix133 (.Y (nx132), .A0 (nx3792), .A1 (nx3758)) ;
    nand02 ix139 (.Y (nx138), .A0 (nx3792), .A1 (nx3764)) ;
    nand02 ix3809 (.Y (nx3808), .A0 (T[8]), .A1 (en)) ;
    inv01 ix3811 (.Y (nx3810), .A (T[7])) ;
    inv01 ix3813 (.Y (nx3812), .A (T[6])) ;
    nor02_2x ix3855 (.Y (nx3854), .A0 (T[4]), .A1 (T[5])) ;
    or02 ix3873 (.Y (nx3872), .A0 (nx18), .A1 (nx3874)) ;
    nand04 ix3875 (.Y (nx3874), .A0 (T[8]), .A1 (en), .A2 (nx4858), .A3 (nx3812)
           ) ;
    or02 ix3948 (.Y (nx3947), .A0 (nx18), .A1 (nx3949)) ;
    nand04 ix3950 (.Y (nx3949), .A0 (T[8]), .A1 (en), .A2 (nx3810), .A3 (nx4860)
           ) ;
    nor03_2x ix921 (.Y (nx920), .A0 (nx3808), .A1 (nx4858), .A2 (nx4860)) ;
    nand02 ix4044 (.Y (nx4043), .A0 (nx3803), .A1 (nx920)) ;
    nand02 ix4062 (.Y (nx4061), .A0 (nx3832), .A1 (nx920)) ;
    nand02 ix4080 (.Y (nx4079), .A0 (nx3854), .A1 (nx920)) ;
    or02 ix4098 (.Y (nx4097), .A0 (nx18), .A1 (nx4099)) ;
    nand03 ix4100 (.Y (nx4099), .A0 (nx1196), .A1 (nx4858), .A2 (nx4860)) ;
    nor02ii ix1197 (.Y (nx1196), .A0 (T[8]), .A1 (en)) ;
    or02 ix4174 (.Y (nx4173), .A0 (nx18), .A1 (nx4175)) ;
    nand03 ix4176 (.Y (nx4175), .A0 (nx1196), .A1 (nx4858), .A2 (nx3812)) ;
    or02 ix4253 (.Y (nx4252), .A0 (nx18), .A1 (nx4254)) ;
    nand03 ix4255 (.Y (nx4254), .A0 (nx1196), .A1 (nx3810), .A2 (nx4860)) ;
    or02 ix4328 (.Y (nx4327), .A0 (nx18), .A1 (nx4329)) ;
    nand03 ix4330 (.Y (nx4329), .A0 (nx1196), .A1 (nx3810), .A2 (nx3812)) ;
    inv01 ix4405 (.Y (nx4406), .A (nx12)) ;
    inv01 ix4417 (.Y (nx4418), .A (nx38)) ;
    inv01 ix4429 (.Y (nx4430), .A (nx48)) ;
    inv01 ix4441 (.Y (nx4442), .A (nx56)) ;
    inv01 ix4453 (.Y (nx4454), .A (nx66)) ;
    inv01 ix4465 (.Y (nx4466), .A (nx72)) ;
    inv01 ix4477 (.Y (nx4478), .A (nx78)) ;
    inv01 ix4489 (.Y (nx4490), .A (nx84)) ;
    inv01 ix4501 (.Y (nx4502), .A (nx94)) ;
    inv01 ix4513 (.Y (nx4514), .A (nx100)) ;
    inv01 ix4525 (.Y (nx4526), .A (nx106)) ;
    inv01 ix4537 (.Y (nx4538), .A (nx112)) ;
    inv01 ix4549 (.Y (nx4550), .A (nx120)) ;
    inv01 ix4561 (.Y (nx4562), .A (nx126)) ;
    inv01 ix4573 (.Y (nx4574), .A (nx132)) ;
    inv01 ix4585 (.Y (nx4586), .A (nx138)) ;
    and02 ix33 (.Y (decoded[511]), .A0 (nx4866), .A1 (nx4994)) ;
    and02 ix43 (.Y (decoded[510]), .A0 (nx4874), .A1 (nx4994)) ;
    nor02ii ix3753 (.Y (nx3752), .A0 (T[0]), .A1 (nx4864)) ;
    and02 ix53 (.Y (decoded[509]), .A0 (nx4882), .A1 (nx4994)) ;
    nor02ii ix3759 (.Y (nx3758), .A0 (nx4864), .A1 (T[0])) ;
    and02 ix61 (.Y (decoded[508]), .A0 (nx4890), .A1 (nx4994)) ;
    and02 ix71 (.Y (decoded[507]), .A0 (nx4898), .A1 (nx4994)) ;
    nor02ii ix3769 (.Y (nx3768), .A0 (T[2]), .A1 (nx4862)) ;
    and02 ix77 (.Y (decoded[506]), .A0 (nx4906), .A1 (nx4994)) ;
    and02 ix83 (.Y (decoded[505]), .A0 (nx4914), .A1 (nx4994)) ;
    and02 ix89 (.Y (decoded[504]), .A0 (nx4922), .A1 (nx4996)) ;
    and02 ix99 (.Y (decoded[503]), .A0 (nx4930), .A1 (nx4996)) ;
    nor02ii ix3781 (.Y (nx3780), .A0 (nx4862), .A1 (T[2])) ;
    and02 ix105 (.Y (decoded[502]), .A0 (nx4938), .A1 (nx4996)) ;
    and02 ix111 (.Y (decoded[501]), .A0 (nx4946), .A1 (nx4996)) ;
    and02 ix117 (.Y (decoded[500]), .A0 (nx4954), .A1 (nx4996)) ;
    and02 ix125 (.Y (decoded[499]), .A0 (nx4962), .A1 (nx4996)) ;
    and02 ix131 (.Y (decoded[498]), .A0 (nx4970), .A1 (nx4996)) ;
    and02 ix137 (.Y (decoded[497]), .A0 (nx4978), .A1 (nx4998)) ;
    and02 ix143 (.Y (decoded[496]), .A0 (nx4986), .A1 (nx4998)) ;
    and02 ix155 (.Y (decoded[495]), .A0 (nx4866), .A1 (nx5002)) ;
    nor02ii ix3802 (.Y (nx4606), .A0 (nx3748), .A1 (nx3803)) ;
    nor02ii ix3804 (.Y (nx3803), .A0 (T[4]), .A1 (T[5])) ;
    and02 ix159 (.Y (decoded[494]), .A0 (nx4874), .A1 (nx5002)) ;
    and02 ix163 (.Y (decoded[493]), .A0 (nx4882), .A1 (nx5002)) ;
    and02 ix167 (.Y (decoded[492]), .A0 (nx4890), .A1 (nx5002)) ;
    and02 ix171 (.Y (decoded[491]), .A0 (nx4898), .A1 (nx5002)) ;
    and02 ix175 (.Y (decoded[490]), .A0 (nx4906), .A1 (nx5002)) ;
    and02 ix179 (.Y (decoded[489]), .A0 (nx4914), .A1 (nx5002)) ;
    and02 ix183 (.Y (decoded[488]), .A0 (nx4922), .A1 (nx5004)) ;
    and02 ix187 (.Y (decoded[487]), .A0 (nx4930), .A1 (nx5004)) ;
    and02 ix191 (.Y (decoded[486]), .A0 (nx4938), .A1 (nx5004)) ;
    and02 ix195 (.Y (decoded[485]), .A0 (nx4946), .A1 (nx5004)) ;
    and02 ix199 (.Y (decoded[484]), .A0 (nx4954), .A1 (nx5004)) ;
    and02 ix203 (.Y (decoded[483]), .A0 (nx4962), .A1 (nx5004)) ;
    and02 ix207 (.Y (decoded[482]), .A0 (nx4970), .A1 (nx5004)) ;
    and02 ix211 (.Y (decoded[481]), .A0 (nx4978), .A1 (nx5006)) ;
    and02 ix215 (.Y (decoded[480]), .A0 (nx4986), .A1 (nx5006)) ;
    and02 ix227 (.Y (decoded[479]), .A0 (nx4866), .A1 (nx5010)) ;
    nor02ii ix3831 (.Y (nx4614), .A0 (nx3748), .A1 (nx3832)) ;
    nor02ii ix3833 (.Y (nx3832), .A0 (T[5]), .A1 (T[4])) ;
    and02 ix231 (.Y (decoded[478]), .A0 (nx4874), .A1 (nx5010)) ;
    and02 ix235 (.Y (decoded[477]), .A0 (nx4882), .A1 (nx5010)) ;
    and02 ix239 (.Y (decoded[476]), .A0 (nx4890), .A1 (nx5010)) ;
    and02 ix243 (.Y (decoded[475]), .A0 (nx4898), .A1 (nx5010)) ;
    and02 ix247 (.Y (decoded[474]), .A0 (nx4906), .A1 (nx5010)) ;
    and02 ix251 (.Y (decoded[473]), .A0 (nx4914), .A1 (nx5010)) ;
    and02 ix255 (.Y (decoded[472]), .A0 (nx4922), .A1 (nx5012)) ;
    and02 ix259 (.Y (decoded[471]), .A0 (nx4930), .A1 (nx5012)) ;
    and02 ix263 (.Y (decoded[470]), .A0 (nx4938), .A1 (nx5012)) ;
    and02 ix267 (.Y (decoded[469]), .A0 (nx4946), .A1 (nx5012)) ;
    and02 ix271 (.Y (decoded[468]), .A0 (nx4954), .A1 (nx5012)) ;
    and02 ix275 (.Y (decoded[467]), .A0 (nx4962), .A1 (nx5012)) ;
    and02 ix279 (.Y (decoded[466]), .A0 (nx4970), .A1 (nx5012)) ;
    and02 ix283 (.Y (decoded[465]), .A0 (nx4978), .A1 (nx5014)) ;
    and02 ix287 (.Y (decoded[464]), .A0 (nx4986), .A1 (nx5014)) ;
    and02 ix297 (.Y (decoded[463]), .A0 (nx4866), .A1 (nx5018)) ;
    nor02ii ix3853 (.Y (nx4622), .A0 (nx3748), .A1 (nx3854)) ;
    and02 ix301 (.Y (decoded[462]), .A0 (nx4874), .A1 (nx5018)) ;
    and02 ix305 (.Y (decoded[461]), .A0 (nx4882), .A1 (nx5018)) ;
    and02 ix309 (.Y (decoded[460]), .A0 (nx4890), .A1 (nx5018)) ;
    and02 ix313 (.Y (decoded[459]), .A0 (nx4898), .A1 (nx5018)) ;
    and02 ix317 (.Y (decoded[458]), .A0 (nx4906), .A1 (nx5018)) ;
    and02 ix321 (.Y (decoded[457]), .A0 (nx4914), .A1 (nx5018)) ;
    and02 ix325 (.Y (decoded[456]), .A0 (nx4922), .A1 (nx5020)) ;
    and02 ix329 (.Y (decoded[455]), .A0 (nx4930), .A1 (nx5020)) ;
    and02 ix333 (.Y (decoded[454]), .A0 (nx4938), .A1 (nx5020)) ;
    and02 ix337 (.Y (decoded[453]), .A0 (nx4946), .A1 (nx5020)) ;
    and02 ix341 (.Y (decoded[452]), .A0 (nx4954), .A1 (nx5020)) ;
    and02 ix345 (.Y (decoded[451]), .A0 (nx4962), .A1 (nx5020)) ;
    and02 ix349 (.Y (decoded[450]), .A0 (nx4970), .A1 (nx5020)) ;
    and02 ix353 (.Y (decoded[449]), .A0 (nx4978), .A1 (nx5022)) ;
    and02 ix357 (.Y (decoded[448]), .A0 (nx4986), .A1 (nx5022)) ;
    and02 ix371 (.Y (decoded[447]), .A0 (nx4866), .A1 (nx5024)) ;
    and02 ix375 (.Y (decoded[446]), .A0 (nx4874), .A1 (nx5024)) ;
    and02 ix379 (.Y (decoded[445]), .A0 (nx4882), .A1 (nx5024)) ;
    and02 ix383 (.Y (decoded[444]), .A0 (nx4890), .A1 (nx5024)) ;
    and02 ix387 (.Y (decoded[443]), .A0 (nx4898), .A1 (nx5024)) ;
    and02 ix391 (.Y (decoded[442]), .A0 (nx4906), .A1 (nx5024)) ;
    and02 ix395 (.Y (decoded[441]), .A0 (nx4914), .A1 (nx5024)) ;
    and02 ix399 (.Y (decoded[440]), .A0 (nx4922), .A1 (nx5026)) ;
    and02 ix403 (.Y (decoded[439]), .A0 (nx4930), .A1 (nx5026)) ;
    and02 ix407 (.Y (decoded[438]), .A0 (nx4938), .A1 (nx5026)) ;
    and02 ix411 (.Y (decoded[437]), .A0 (nx4946), .A1 (nx5026)) ;
    and02 ix415 (.Y (decoded[436]), .A0 (nx4954), .A1 (nx5026)) ;
    and02 ix419 (.Y (decoded[435]), .A0 (nx4962), .A1 (nx5026)) ;
    and02 ix423 (.Y (decoded[434]), .A0 (nx4970), .A1 (nx5026)) ;
    and02 ix427 (.Y (decoded[433]), .A0 (nx4978), .A1 (nx5028)) ;
    and02 ix431 (.Y (decoded[432]), .A0 (nx4986), .A1 (nx5028)) ;
    and02 ix439 (.Y (decoded[431]), .A0 (nx4866), .A1 (nx5032)) ;
    nor02ii ix3893 (.Y (nx4638), .A0 (nx3874), .A1 (nx3803)) ;
    and02 ix443 (.Y (decoded[430]), .A0 (nx4874), .A1 (nx5032)) ;
    and02 ix447 (.Y (decoded[429]), .A0 (nx4882), .A1 (nx5032)) ;
    and02 ix451 (.Y (decoded[428]), .A0 (nx4890), .A1 (nx5032)) ;
    and02 ix455 (.Y (decoded[427]), .A0 (nx4898), .A1 (nx5032)) ;
    and02 ix459 (.Y (decoded[426]), .A0 (nx4906), .A1 (nx5032)) ;
    and02 ix463 (.Y (decoded[425]), .A0 (nx4914), .A1 (nx5032)) ;
    and02 ix467 (.Y (decoded[424]), .A0 (nx4922), .A1 (nx5034)) ;
    and02 ix471 (.Y (decoded[423]), .A0 (nx4930), .A1 (nx5034)) ;
    and02 ix475 (.Y (decoded[422]), .A0 (nx4938), .A1 (nx5034)) ;
    and02 ix479 (.Y (decoded[421]), .A0 (nx4946), .A1 (nx5034)) ;
    and02 ix483 (.Y (decoded[420]), .A0 (nx4954), .A1 (nx5034)) ;
    and02 ix487 (.Y (decoded[419]), .A0 (nx4962), .A1 (nx5034)) ;
    and02 ix491 (.Y (decoded[418]), .A0 (nx4970), .A1 (nx5034)) ;
    and02 ix495 (.Y (decoded[417]), .A0 (nx4978), .A1 (nx5036)) ;
    and02 ix499 (.Y (decoded[416]), .A0 (nx4986), .A1 (nx5036)) ;
    and02 ix507 (.Y (decoded[415]), .A0 (nx4866), .A1 (nx5040)) ;
    nor02ii ix3912 (.Y (nx4646), .A0 (nx3874), .A1 (nx3832)) ;
    and02 ix511 (.Y (decoded[414]), .A0 (nx4874), .A1 (nx5040)) ;
    and02 ix515 (.Y (decoded[413]), .A0 (nx4882), .A1 (nx5040)) ;
    and02 ix519 (.Y (decoded[412]), .A0 (nx4890), .A1 (nx5040)) ;
    and02 ix523 (.Y (decoded[411]), .A0 (nx4898), .A1 (nx5040)) ;
    and02 ix527 (.Y (decoded[410]), .A0 (nx4906), .A1 (nx5040)) ;
    and02 ix531 (.Y (decoded[409]), .A0 (nx4914), .A1 (nx5040)) ;
    and02 ix535 (.Y (decoded[408]), .A0 (nx4922), .A1 (nx5042)) ;
    and02 ix539 (.Y (decoded[407]), .A0 (nx4930), .A1 (nx5042)) ;
    and02 ix543 (.Y (decoded[406]), .A0 (nx4938), .A1 (nx5042)) ;
    and02 ix547 (.Y (decoded[405]), .A0 (nx4946), .A1 (nx5042)) ;
    and02 ix551 (.Y (decoded[404]), .A0 (nx4954), .A1 (nx5042)) ;
    and02 ix555 (.Y (decoded[403]), .A0 (nx4962), .A1 (nx5042)) ;
    and02 ix559 (.Y (decoded[402]), .A0 (nx4970), .A1 (nx5042)) ;
    and02 ix563 (.Y (decoded[401]), .A0 (nx4978), .A1 (nx5044)) ;
    and02 ix567 (.Y (decoded[400]), .A0 (nx4986), .A1 (nx5044)) ;
    and02 ix575 (.Y (decoded[399]), .A0 (nx4868), .A1 (nx5048)) ;
    nor02ii ix3930 (.Y (nx4654), .A0 (nx3874), .A1 (nx3854)) ;
    and02 ix579 (.Y (decoded[398]), .A0 (nx4876), .A1 (nx5048)) ;
    and02 ix583 (.Y (decoded[397]), .A0 (nx4884), .A1 (nx5048)) ;
    and02 ix587 (.Y (decoded[396]), .A0 (nx4892), .A1 (nx5048)) ;
    and02 ix591 (.Y (decoded[395]), .A0 (nx4900), .A1 (nx5048)) ;
    and02 ix595 (.Y (decoded[394]), .A0 (nx4908), .A1 (nx5048)) ;
    and02 ix599 (.Y (decoded[393]), .A0 (nx4916), .A1 (nx5048)) ;
    and02 ix603 (.Y (decoded[392]), .A0 (nx4924), .A1 (nx5050)) ;
    and02 ix607 (.Y (decoded[391]), .A0 (nx4932), .A1 (nx5050)) ;
    and02 ix611 (.Y (decoded[390]), .A0 (nx4940), .A1 (nx5050)) ;
    and02 ix615 (.Y (decoded[389]), .A0 (nx4948), .A1 (nx5050)) ;
    and02 ix619 (.Y (decoded[388]), .A0 (nx4956), .A1 (nx5050)) ;
    and02 ix623 (.Y (decoded[387]), .A0 (nx4964), .A1 (nx5050)) ;
    and02 ix627 (.Y (decoded[386]), .A0 (nx4972), .A1 (nx5050)) ;
    and02 ix631 (.Y (decoded[385]), .A0 (nx4980), .A1 (nx5052)) ;
    and02 ix635 (.Y (decoded[384]), .A0 (nx4988), .A1 (nx5052)) ;
    and02 ix649 (.Y (decoded[383]), .A0 (nx4868), .A1 (nx5054)) ;
    and02 ix653 (.Y (decoded[382]), .A0 (nx4876), .A1 (nx5054)) ;
    and02 ix657 (.Y (decoded[381]), .A0 (nx4884), .A1 (nx5054)) ;
    and02 ix661 (.Y (decoded[380]), .A0 (nx4892), .A1 (nx5054)) ;
    and02 ix665 (.Y (decoded[379]), .A0 (nx4900), .A1 (nx5054)) ;
    and02 ix669 (.Y (decoded[378]), .A0 (nx4908), .A1 (nx5054)) ;
    and02 ix673 (.Y (decoded[377]), .A0 (nx4916), .A1 (nx5054)) ;
    and02 ix677 (.Y (decoded[376]), .A0 (nx4924), .A1 (nx5056)) ;
    and02 ix681 (.Y (decoded[375]), .A0 (nx4932), .A1 (nx5056)) ;
    and02 ix685 (.Y (decoded[374]), .A0 (nx4940), .A1 (nx5056)) ;
    and02 ix689 (.Y (decoded[373]), .A0 (nx4948), .A1 (nx5056)) ;
    and02 ix693 (.Y (decoded[372]), .A0 (nx4956), .A1 (nx5056)) ;
    and02 ix697 (.Y (decoded[371]), .A0 (nx4964), .A1 (nx5056)) ;
    and02 ix701 (.Y (decoded[370]), .A0 (nx4972), .A1 (nx5056)) ;
    and02 ix705 (.Y (decoded[369]), .A0 (nx4980), .A1 (nx5058)) ;
    and02 ix709 (.Y (decoded[368]), .A0 (nx4988), .A1 (nx5058)) ;
    and02 ix717 (.Y (decoded[367]), .A0 (nx4868), .A1 (nx5062)) ;
    nor02ii ix3968 (.Y (nx4670), .A0 (nx3949), .A1 (nx3803)) ;
    and02 ix721 (.Y (decoded[366]), .A0 (nx4876), .A1 (nx5062)) ;
    and02 ix725 (.Y (decoded[365]), .A0 (nx4884), .A1 (nx5062)) ;
    and02 ix729 (.Y (decoded[364]), .A0 (nx4892), .A1 (nx5062)) ;
    and02 ix733 (.Y (decoded[363]), .A0 (nx4900), .A1 (nx5062)) ;
    and02 ix737 (.Y (decoded[362]), .A0 (nx4908), .A1 (nx5062)) ;
    and02 ix741 (.Y (decoded[361]), .A0 (nx4916), .A1 (nx5062)) ;
    and02 ix745 (.Y (decoded[360]), .A0 (nx4924), .A1 (nx5064)) ;
    and02 ix749 (.Y (decoded[359]), .A0 (nx4932), .A1 (nx5064)) ;
    and02 ix753 (.Y (decoded[358]), .A0 (nx4940), .A1 (nx5064)) ;
    and02 ix757 (.Y (decoded[357]), .A0 (nx4948), .A1 (nx5064)) ;
    and02 ix761 (.Y (decoded[356]), .A0 (nx4956), .A1 (nx5064)) ;
    and02 ix765 (.Y (decoded[355]), .A0 (nx4964), .A1 (nx5064)) ;
    and02 ix769 (.Y (decoded[354]), .A0 (nx4972), .A1 (nx5064)) ;
    and02 ix773 (.Y (decoded[353]), .A0 (nx4980), .A1 (nx5066)) ;
    and02 ix777 (.Y (decoded[352]), .A0 (nx4988), .A1 (nx5066)) ;
    and02 ix785 (.Y (decoded[351]), .A0 (nx4868), .A1 (nx5070)) ;
    nor02ii ix3987 (.Y (nx4678), .A0 (nx3949), .A1 (nx3832)) ;
    and02 ix789 (.Y (decoded[350]), .A0 (nx4876), .A1 (nx5070)) ;
    and02 ix793 (.Y (decoded[349]), .A0 (nx4884), .A1 (nx5070)) ;
    and02 ix797 (.Y (decoded[348]), .A0 (nx4892), .A1 (nx5070)) ;
    and02 ix801 (.Y (decoded[347]), .A0 (nx4900), .A1 (nx5070)) ;
    and02 ix805 (.Y (decoded[346]), .A0 (nx4908), .A1 (nx5070)) ;
    and02 ix809 (.Y (decoded[345]), .A0 (nx4916), .A1 (nx5070)) ;
    and02 ix813 (.Y (decoded[344]), .A0 (nx4924), .A1 (nx5072)) ;
    and02 ix817 (.Y (decoded[343]), .A0 (nx4932), .A1 (nx5072)) ;
    and02 ix821 (.Y (decoded[342]), .A0 (nx4940), .A1 (nx5072)) ;
    and02 ix825 (.Y (decoded[341]), .A0 (nx4948), .A1 (nx5072)) ;
    and02 ix829 (.Y (decoded[340]), .A0 (nx4956), .A1 (nx5072)) ;
    and02 ix833 (.Y (decoded[339]), .A0 (nx4964), .A1 (nx5072)) ;
    and02 ix837 (.Y (decoded[338]), .A0 (nx4972), .A1 (nx5072)) ;
    and02 ix841 (.Y (decoded[337]), .A0 (nx4980), .A1 (nx5074)) ;
    and02 ix845 (.Y (decoded[336]), .A0 (nx4988), .A1 (nx5074)) ;
    and02 ix853 (.Y (decoded[335]), .A0 (nx4868), .A1 (nx5078)) ;
    nor02ii ix4005 (.Y (nx4686), .A0 (nx3949), .A1 (nx3854)) ;
    and02 ix857 (.Y (decoded[334]), .A0 (nx4876), .A1 (nx5078)) ;
    and02 ix861 (.Y (decoded[333]), .A0 (nx4884), .A1 (nx5078)) ;
    and02 ix865 (.Y (decoded[332]), .A0 (nx4892), .A1 (nx5078)) ;
    and02 ix869 (.Y (decoded[331]), .A0 (nx4900), .A1 (nx5078)) ;
    and02 ix873 (.Y (decoded[330]), .A0 (nx4908), .A1 (nx5078)) ;
    and02 ix877 (.Y (decoded[329]), .A0 (nx4916), .A1 (nx5078)) ;
    and02 ix881 (.Y (decoded[328]), .A0 (nx4924), .A1 (nx5080)) ;
    and02 ix885 (.Y (decoded[327]), .A0 (nx4932), .A1 (nx5080)) ;
    and02 ix889 (.Y (decoded[326]), .A0 (nx4940), .A1 (nx5080)) ;
    and02 ix893 (.Y (decoded[325]), .A0 (nx4948), .A1 (nx5080)) ;
    and02 ix897 (.Y (decoded[324]), .A0 (nx4956), .A1 (nx5080)) ;
    and02 ix901 (.Y (decoded[323]), .A0 (nx4964), .A1 (nx5080)) ;
    and02 ix905 (.Y (decoded[322]), .A0 (nx4972), .A1 (nx5080)) ;
    and02 ix909 (.Y (decoded[321]), .A0 (nx4980), .A1 (nx5082)) ;
    and02 ix913 (.Y (decoded[320]), .A0 (nx4988), .A1 (nx5082)) ;
    and02 ix929 (.Y (decoded[319]), .A0 (nx4868), .A1 (nx5086)) ;
    nor02ii ix4023 (.Y (nx4694), .A0 (nx18), .A1 (nx920)) ;
    and02 ix933 (.Y (decoded[318]), .A0 (nx4876), .A1 (nx5086)) ;
    and02 ix937 (.Y (decoded[317]), .A0 (nx4884), .A1 (nx5086)) ;
    and02 ix941 (.Y (decoded[316]), .A0 (nx4892), .A1 (nx5086)) ;
    and02 ix945 (.Y (decoded[315]), .A0 (nx4900), .A1 (nx5086)) ;
    and02 ix949 (.Y (decoded[314]), .A0 (nx4908), .A1 (nx5086)) ;
    and02 ix953 (.Y (decoded[313]), .A0 (nx4916), .A1 (nx5086)) ;
    and02 ix957 (.Y (decoded[312]), .A0 (nx4924), .A1 (nx5088)) ;
    and02 ix961 (.Y (decoded[311]), .A0 (nx4932), .A1 (nx5088)) ;
    and02 ix965 (.Y (decoded[310]), .A0 (nx4940), .A1 (nx5088)) ;
    and02 ix969 (.Y (decoded[309]), .A0 (nx4948), .A1 (nx5088)) ;
    and02 ix973 (.Y (decoded[308]), .A0 (nx4956), .A1 (nx5088)) ;
    and02 ix977 (.Y (decoded[307]), .A0 (nx4964), .A1 (nx5088)) ;
    and02 ix981 (.Y (decoded[306]), .A0 (nx4972), .A1 (nx5088)) ;
    and02 ix985 (.Y (decoded[305]), .A0 (nx4980), .A1 (nx5090)) ;
    and02 ix989 (.Y (decoded[304]), .A0 (nx4988), .A1 (nx5090)) ;
    and02 ix997 (.Y (decoded[303]), .A0 (nx4868), .A1 (nx5092)) ;
    and02 ix1001 (.Y (decoded[302]), .A0 (nx4876), .A1 (nx5092)) ;
    and02 ix1005 (.Y (decoded[301]), .A0 (nx4884), .A1 (nx5092)) ;
    and02 ix1009 (.Y (decoded[300]), .A0 (nx4892), .A1 (nx5092)) ;
    and02 ix1013 (.Y (decoded[299]), .A0 (nx4900), .A1 (nx5092)) ;
    and02 ix1017 (.Y (decoded[298]), .A0 (nx4908), .A1 (nx5092)) ;
    and02 ix1021 (.Y (decoded[297]), .A0 (nx4916), .A1 (nx5092)) ;
    and02 ix1025 (.Y (decoded[296]), .A0 (nx4924), .A1 (nx5094)) ;
    and02 ix1029 (.Y (decoded[295]), .A0 (nx4932), .A1 (nx5094)) ;
    and02 ix1033 (.Y (decoded[294]), .A0 (nx4940), .A1 (nx5094)) ;
    and02 ix1037 (.Y (decoded[293]), .A0 (nx4948), .A1 (nx5094)) ;
    and02 ix1041 (.Y (decoded[292]), .A0 (nx4956), .A1 (nx5094)) ;
    and02 ix1045 (.Y (decoded[291]), .A0 (nx4964), .A1 (nx5094)) ;
    and02 ix1049 (.Y (decoded[290]), .A0 (nx4972), .A1 (nx5094)) ;
    and02 ix1053 (.Y (decoded[289]), .A0 (nx4980), .A1 (nx5096)) ;
    and02 ix1057 (.Y (decoded[288]), .A0 (nx4988), .A1 (nx5096)) ;
    and02 ix1065 (.Y (decoded[287]), .A0 (nx4870), .A1 (nx5098)) ;
    and02 ix1069 (.Y (decoded[286]), .A0 (nx4878), .A1 (nx5098)) ;
    and02 ix1073 (.Y (decoded[285]), .A0 (nx4886), .A1 (nx5098)) ;
    and02 ix1077 (.Y (decoded[284]), .A0 (nx4894), .A1 (nx5098)) ;
    and02 ix1081 (.Y (decoded[283]), .A0 (nx4902), .A1 (nx5098)) ;
    and02 ix1085 (.Y (decoded[282]), .A0 (nx4910), .A1 (nx5098)) ;
    and02 ix1089 (.Y (decoded[281]), .A0 (nx4918), .A1 (nx5098)) ;
    and02 ix1093 (.Y (decoded[280]), .A0 (nx4926), .A1 (nx5100)) ;
    and02 ix1097 (.Y (decoded[279]), .A0 (nx4934), .A1 (nx5100)) ;
    and02 ix1101 (.Y (decoded[278]), .A0 (nx4942), .A1 (nx5100)) ;
    and02 ix1105 (.Y (decoded[277]), .A0 (nx4950), .A1 (nx5100)) ;
    and02 ix1109 (.Y (decoded[276]), .A0 (nx4958), .A1 (nx5100)) ;
    and02 ix1113 (.Y (decoded[275]), .A0 (nx4966), .A1 (nx5100)) ;
    and02 ix1117 (.Y (decoded[274]), .A0 (nx4974), .A1 (nx5100)) ;
    and02 ix1121 (.Y (decoded[273]), .A0 (nx4982), .A1 (nx5102)) ;
    and02 ix1125 (.Y (decoded[272]), .A0 (nx4990), .A1 (nx5102)) ;
    and02 ix1133 (.Y (decoded[271]), .A0 (nx4870), .A1 (nx5104)) ;
    and02 ix1137 (.Y (decoded[270]), .A0 (nx4878), .A1 (nx5104)) ;
    and02 ix1141 (.Y (decoded[269]), .A0 (nx4886), .A1 (nx5104)) ;
    and02 ix1145 (.Y (decoded[268]), .A0 (nx4894), .A1 (nx5104)) ;
    and02 ix1149 (.Y (decoded[267]), .A0 (nx4902), .A1 (nx5104)) ;
    and02 ix1153 (.Y (decoded[266]), .A0 (nx4910), .A1 (nx5104)) ;
    and02 ix1157 (.Y (decoded[265]), .A0 (nx4918), .A1 (nx5104)) ;
    and02 ix1161 (.Y (decoded[264]), .A0 (nx4926), .A1 (nx5106)) ;
    and02 ix1165 (.Y (decoded[263]), .A0 (nx4934), .A1 (nx5106)) ;
    and02 ix1169 (.Y (decoded[262]), .A0 (nx4942), .A1 (nx5106)) ;
    and02 ix1173 (.Y (decoded[261]), .A0 (nx4950), .A1 (nx5106)) ;
    and02 ix1177 (.Y (decoded[260]), .A0 (nx4958), .A1 (nx5106)) ;
    and02 ix1181 (.Y (decoded[259]), .A0 (nx4966), .A1 (nx5106)) ;
    and02 ix1185 (.Y (decoded[258]), .A0 (nx4974), .A1 (nx5106)) ;
    and02 ix1189 (.Y (decoded[257]), .A0 (nx4982), .A1 (nx5108)) ;
    and02 ix1193 (.Y (decoded[256]), .A0 (nx4990), .A1 (nx5108)) ;
    and02 ix1209 (.Y (decoded[255]), .A0 (nx4870), .A1 (nx5110)) ;
    and02 ix1213 (.Y (decoded[254]), .A0 (nx4878), .A1 (nx5110)) ;
    and02 ix1217 (.Y (decoded[253]), .A0 (nx4886), .A1 (nx5110)) ;
    and02 ix1221 (.Y (decoded[252]), .A0 (nx4894), .A1 (nx5110)) ;
    and02 ix1225 (.Y (decoded[251]), .A0 (nx4902), .A1 (nx5110)) ;
    and02 ix1229 (.Y (decoded[250]), .A0 (nx4910), .A1 (nx5110)) ;
    and02 ix1233 (.Y (decoded[249]), .A0 (nx4918), .A1 (nx5110)) ;
    and02 ix1237 (.Y (decoded[248]), .A0 (nx4926), .A1 (nx5112)) ;
    and02 ix1241 (.Y (decoded[247]), .A0 (nx4934), .A1 (nx5112)) ;
    and02 ix1245 (.Y (decoded[246]), .A0 (nx4942), .A1 (nx5112)) ;
    and02 ix1249 (.Y (decoded[245]), .A0 (nx4950), .A1 (nx5112)) ;
    and02 ix1253 (.Y (decoded[244]), .A0 (nx4958), .A1 (nx5112)) ;
    and02 ix1257 (.Y (decoded[243]), .A0 (nx4966), .A1 (nx5112)) ;
    and02 ix1261 (.Y (decoded[242]), .A0 (nx4974), .A1 (nx5112)) ;
    and02 ix1265 (.Y (decoded[241]), .A0 (nx4982), .A1 (nx5114)) ;
    and02 ix1269 (.Y (decoded[240]), .A0 (nx4990), .A1 (nx5114)) ;
    and02 ix1277 (.Y (decoded[239]), .A0 (nx4870), .A1 (nx5118)) ;
    nor02ii ix4119 (.Y (nx4734), .A0 (nx4099), .A1 (nx3803)) ;
    and02 ix1281 (.Y (decoded[238]), .A0 (nx4878), .A1 (nx5118)) ;
    and02 ix1285 (.Y (decoded[237]), .A0 (nx4886), .A1 (nx5118)) ;
    and02 ix1289 (.Y (decoded[236]), .A0 (nx4894), .A1 (nx5118)) ;
    and02 ix1293 (.Y (decoded[235]), .A0 (nx4902), .A1 (nx5118)) ;
    and02 ix1297 (.Y (decoded[234]), .A0 (nx4910), .A1 (nx5118)) ;
    and02 ix1301 (.Y (decoded[233]), .A0 (nx4918), .A1 (nx5118)) ;
    and02 ix1305 (.Y (decoded[232]), .A0 (nx4926), .A1 (nx5120)) ;
    and02 ix1309 (.Y (decoded[231]), .A0 (nx4934), .A1 (nx5120)) ;
    and02 ix1313 (.Y (decoded[230]), .A0 (nx4942), .A1 (nx5120)) ;
    and02 ix1317 (.Y (decoded[229]), .A0 (nx4950), .A1 (nx5120)) ;
    and02 ix1321 (.Y (decoded[228]), .A0 (nx4958), .A1 (nx5120)) ;
    and02 ix1325 (.Y (decoded[227]), .A0 (nx4966), .A1 (nx5120)) ;
    and02 ix1329 (.Y (decoded[226]), .A0 (nx4974), .A1 (nx5120)) ;
    and02 ix1333 (.Y (decoded[225]), .A0 (nx4982), .A1 (nx5122)) ;
    and02 ix1337 (.Y (decoded[224]), .A0 (nx4990), .A1 (nx5122)) ;
    and02 ix1345 (.Y (decoded[223]), .A0 (nx4870), .A1 (nx5126)) ;
    nor02ii ix4138 (.Y (nx4742), .A0 (nx4099), .A1 (nx3832)) ;
    and02 ix1349 (.Y (decoded[222]), .A0 (nx4878), .A1 (nx5126)) ;
    and02 ix1353 (.Y (decoded[221]), .A0 (nx4886), .A1 (nx5126)) ;
    and02 ix1357 (.Y (decoded[220]), .A0 (nx4894), .A1 (nx5126)) ;
    and02 ix1361 (.Y (decoded[219]), .A0 (nx4902), .A1 (nx5126)) ;
    and02 ix1365 (.Y (decoded[218]), .A0 (nx4910), .A1 (nx5126)) ;
    and02 ix1369 (.Y (decoded[217]), .A0 (nx4918), .A1 (nx5126)) ;
    and02 ix1373 (.Y (decoded[216]), .A0 (nx4926), .A1 (nx5128)) ;
    and02 ix1377 (.Y (decoded[215]), .A0 (nx4934), .A1 (nx5128)) ;
    and02 ix1381 (.Y (decoded[214]), .A0 (nx4942), .A1 (nx5128)) ;
    and02 ix1385 (.Y (decoded[213]), .A0 (nx4950), .A1 (nx5128)) ;
    and02 ix1389 (.Y (decoded[212]), .A0 (nx4958), .A1 (nx5128)) ;
    and02 ix1393 (.Y (decoded[211]), .A0 (nx4966), .A1 (nx5128)) ;
    and02 ix1397 (.Y (decoded[210]), .A0 (nx4974), .A1 (nx5128)) ;
    and02 ix1401 (.Y (decoded[209]), .A0 (nx4982), .A1 (nx5130)) ;
    and02 ix1405 (.Y (decoded[208]), .A0 (nx4990), .A1 (nx5130)) ;
    and02 ix1413 (.Y (decoded[207]), .A0 (nx4870), .A1 (nx5134)) ;
    nor02ii ix4156 (.Y (nx4750), .A0 (nx4099), .A1 (nx3854)) ;
    and02 ix1417 (.Y (decoded[206]), .A0 (nx4878), .A1 (nx5134)) ;
    and02 ix1421 (.Y (decoded[205]), .A0 (nx4886), .A1 (nx5134)) ;
    and02 ix1425 (.Y (decoded[204]), .A0 (nx4894), .A1 (nx5134)) ;
    and02 ix1429 (.Y (decoded[203]), .A0 (nx4902), .A1 (nx5134)) ;
    and02 ix1433 (.Y (decoded[202]), .A0 (nx4910), .A1 (nx5134)) ;
    and02 ix1437 (.Y (decoded[201]), .A0 (nx4918), .A1 (nx5134)) ;
    and02 ix1441 (.Y (decoded[200]), .A0 (nx4926), .A1 (nx5136)) ;
    and02 ix1445 (.Y (decoded[199]), .A0 (nx4934), .A1 (nx5136)) ;
    and02 ix1449 (.Y (decoded[198]), .A0 (nx4942), .A1 (nx5136)) ;
    and02 ix1453 (.Y (decoded[197]), .A0 (nx4950), .A1 (nx5136)) ;
    and02 ix1457 (.Y (decoded[196]), .A0 (nx4958), .A1 (nx5136)) ;
    and02 ix1461 (.Y (decoded[195]), .A0 (nx4966), .A1 (nx5136)) ;
    and02 ix1465 (.Y (decoded[194]), .A0 (nx4974), .A1 (nx5136)) ;
    and02 ix1469 (.Y (decoded[193]), .A0 (nx4982), .A1 (nx5138)) ;
    and02 ix1473 (.Y (decoded[192]), .A0 (nx4990), .A1 (nx5138)) ;
    and02 ix1487 (.Y (decoded[191]), .A0 (nx4870), .A1 (nx5140)) ;
    and02 ix1491 (.Y (decoded[190]), .A0 (nx4878), .A1 (nx5140)) ;
    and02 ix1495 (.Y (decoded[189]), .A0 (nx4886), .A1 (nx5140)) ;
    and02 ix1499 (.Y (decoded[188]), .A0 (nx4894), .A1 (nx5140)) ;
    and02 ix1503 (.Y (decoded[187]), .A0 (nx4902), .A1 (nx5140)) ;
    and02 ix1507 (.Y (decoded[186]), .A0 (nx4910), .A1 (nx5140)) ;
    and02 ix1511 (.Y (decoded[185]), .A0 (nx4918), .A1 (nx5140)) ;
    and02 ix1515 (.Y (decoded[184]), .A0 (nx4926), .A1 (nx5142)) ;
    and02 ix1519 (.Y (decoded[183]), .A0 (nx4934), .A1 (nx5142)) ;
    and02 ix1523 (.Y (decoded[182]), .A0 (nx4942), .A1 (nx5142)) ;
    and02 ix1527 (.Y (decoded[181]), .A0 (nx4950), .A1 (nx5142)) ;
    and02 ix1531 (.Y (decoded[180]), .A0 (nx4958), .A1 (nx5142)) ;
    and02 ix1535 (.Y (decoded[179]), .A0 (nx4966), .A1 (nx5142)) ;
    and02 ix1539 (.Y (decoded[178]), .A0 (nx4974), .A1 (nx5142)) ;
    and02 ix1543 (.Y (decoded[177]), .A0 (nx4982), .A1 (nx5144)) ;
    and02 ix1547 (.Y (decoded[176]), .A0 (nx4990), .A1 (nx5144)) ;
    and02 ix1555 (.Y (decoded[175]), .A0 (nx4872), .A1 (nx5148)) ;
    nor02ii ix4194 (.Y (nx4766), .A0 (nx4175), .A1 (nx3803)) ;
    and02 ix1559 (.Y (decoded[174]), .A0 (nx4880), .A1 (nx5148)) ;
    and02 ix1563 (.Y (decoded[173]), .A0 (nx4888), .A1 (nx5148)) ;
    and02 ix1567 (.Y (decoded[172]), .A0 (nx4896), .A1 (nx5148)) ;
    and02 ix1571 (.Y (decoded[171]), .A0 (nx4904), .A1 (nx5148)) ;
    and02 ix1575 (.Y (decoded[170]), .A0 (nx4912), .A1 (nx5148)) ;
    and02 ix1579 (.Y (decoded[169]), .A0 (nx4920), .A1 (nx5148)) ;
    and02 ix1583 (.Y (decoded[168]), .A0 (nx4928), .A1 (nx5150)) ;
    and02 ix1587 (.Y (decoded[167]), .A0 (nx4936), .A1 (nx5150)) ;
    and02 ix1591 (.Y (decoded[166]), .A0 (nx4944), .A1 (nx5150)) ;
    and02 ix1595 (.Y (decoded[165]), .A0 (nx4952), .A1 (nx5150)) ;
    and02 ix1599 (.Y (decoded[164]), .A0 (nx4960), .A1 (nx5150)) ;
    and02 ix1603 (.Y (decoded[163]), .A0 (nx4968), .A1 (nx5150)) ;
    and02 ix1607 (.Y (decoded[162]), .A0 (nx4976), .A1 (nx5150)) ;
    and02 ix1611 (.Y (decoded[161]), .A0 (nx4984), .A1 (nx5152)) ;
    and02 ix1615 (.Y (decoded[160]), .A0 (nx4992), .A1 (nx5152)) ;
    and02 ix1623 (.Y (decoded[159]), .A0 (nx4872), .A1 (nx5156)) ;
    nor02ii ix4217 (.Y (nx4774), .A0 (nx4175), .A1 (nx3832)) ;
    and02 ix1627 (.Y (decoded[158]), .A0 (nx4880), .A1 (nx5156)) ;
    and02 ix1631 (.Y (decoded[157]), .A0 (nx4888), .A1 (nx5156)) ;
    and02 ix1635 (.Y (decoded[156]), .A0 (nx4896), .A1 (nx5156)) ;
    and02 ix1639 (.Y (decoded[155]), .A0 (nx4904), .A1 (nx5156)) ;
    and02 ix1643 (.Y (decoded[154]), .A0 (nx4912), .A1 (nx5156)) ;
    and02 ix1647 (.Y (decoded[153]), .A0 (nx4920), .A1 (nx5156)) ;
    and02 ix1651 (.Y (decoded[152]), .A0 (nx4928), .A1 (nx5158)) ;
    and02 ix1655 (.Y (decoded[151]), .A0 (nx4936), .A1 (nx5158)) ;
    and02 ix1659 (.Y (decoded[150]), .A0 (nx4944), .A1 (nx5158)) ;
    and02 ix1663 (.Y (decoded[149]), .A0 (nx4952), .A1 (nx5158)) ;
    and02 ix1667 (.Y (decoded[148]), .A0 (nx4960), .A1 (nx5158)) ;
    and02 ix1671 (.Y (decoded[147]), .A0 (nx4968), .A1 (nx5158)) ;
    and02 ix1675 (.Y (decoded[146]), .A0 (nx4976), .A1 (nx5158)) ;
    and02 ix1679 (.Y (decoded[145]), .A0 (nx4984), .A1 (nx5160)) ;
    and02 ix1683 (.Y (decoded[144]), .A0 (nx4992), .A1 (nx5160)) ;
    and02 ix1691 (.Y (decoded[143]), .A0 (nx4872), .A1 (nx5164)) ;
    nor02ii ix4235 (.Y (nx4782), .A0 (nx4175), .A1 (nx3854)) ;
    and02 ix1695 (.Y (decoded[142]), .A0 (nx4880), .A1 (nx5164)) ;
    and02 ix1699 (.Y (decoded[141]), .A0 (nx4888), .A1 (nx5164)) ;
    and02 ix1703 (.Y (decoded[140]), .A0 (nx4896), .A1 (nx5164)) ;
    and02 ix1707 (.Y (decoded[139]), .A0 (nx4904), .A1 (nx5164)) ;
    and02 ix1711 (.Y (decoded[138]), .A0 (nx4912), .A1 (nx5164)) ;
    and02 ix1715 (.Y (decoded[137]), .A0 (nx4920), .A1 (nx5164)) ;
    and02 ix1719 (.Y (decoded[136]), .A0 (nx4928), .A1 (nx5166)) ;
    and02 ix1723 (.Y (decoded[135]), .A0 (nx4936), .A1 (nx5166)) ;
    and02 ix1727 (.Y (decoded[134]), .A0 (nx4944), .A1 (nx5166)) ;
    and02 ix1731 (.Y (decoded[133]), .A0 (nx4952), .A1 (nx5166)) ;
    and02 ix1735 (.Y (decoded[132]), .A0 (nx4960), .A1 (nx5166)) ;
    and02 ix1739 (.Y (decoded[131]), .A0 (nx4968), .A1 (nx5166)) ;
    and02 ix1743 (.Y (decoded[130]), .A0 (nx4976), .A1 (nx5166)) ;
    and02 ix1747 (.Y (decoded[129]), .A0 (nx4984), .A1 (nx5168)) ;
    and02 ix1751 (.Y (decoded[128]), .A0 (nx4992), .A1 (nx5168)) ;
    and02 ix1765 (.Y (decoded[127]), .A0 (nx4872), .A1 (nx5170)) ;
    and02 ix1769 (.Y (decoded[126]), .A0 (nx4880), .A1 (nx5170)) ;
    and02 ix1773 (.Y (decoded[125]), .A0 (nx4888), .A1 (nx5170)) ;
    and02 ix1777 (.Y (decoded[124]), .A0 (nx4896), .A1 (nx5170)) ;
    and02 ix1781 (.Y (decoded[123]), .A0 (nx4904), .A1 (nx5170)) ;
    and02 ix1785 (.Y (decoded[122]), .A0 (nx4912), .A1 (nx5170)) ;
    and02 ix1789 (.Y (decoded[121]), .A0 (nx4920), .A1 (nx5170)) ;
    and02 ix1793 (.Y (decoded[120]), .A0 (nx4928), .A1 (nx5172)) ;
    and02 ix1797 (.Y (decoded[119]), .A0 (nx4936), .A1 (nx5172)) ;
    and02 ix1801 (.Y (decoded[118]), .A0 (nx4944), .A1 (nx5172)) ;
    and02 ix1805 (.Y (decoded[117]), .A0 (nx4952), .A1 (nx5172)) ;
    and02 ix1809 (.Y (decoded[116]), .A0 (nx4960), .A1 (nx5172)) ;
    and02 ix1813 (.Y (decoded[115]), .A0 (nx4968), .A1 (nx5172)) ;
    and02 ix1817 (.Y (decoded[114]), .A0 (nx4976), .A1 (nx5172)) ;
    and02 ix1821 (.Y (decoded[113]), .A0 (nx4984), .A1 (nx5174)) ;
    and02 ix1825 (.Y (decoded[112]), .A0 (nx4992), .A1 (nx5174)) ;
    and02 ix1833 (.Y (decoded[111]), .A0 (nx4872), .A1 (nx5178)) ;
    nor02ii ix4273 (.Y (nx4798), .A0 (nx4254), .A1 (nx3803)) ;
    and02 ix1837 (.Y (decoded[110]), .A0 (nx4880), .A1 (nx5178)) ;
    and02 ix1841 (.Y (decoded[109]), .A0 (nx4888), .A1 (nx5178)) ;
    and02 ix1845 (.Y (decoded[108]), .A0 (nx4896), .A1 (nx5178)) ;
    and02 ix1849 (.Y (decoded[107]), .A0 (nx4904), .A1 (nx5178)) ;
    and02 ix1853 (.Y (decoded[106]), .A0 (nx4912), .A1 (nx5178)) ;
    and02 ix1857 (.Y (decoded[105]), .A0 (nx4920), .A1 (nx5178)) ;
    and02 ix1861 (.Y (decoded[104]), .A0 (nx4928), .A1 (nx5180)) ;
    and02 ix1865 (.Y (decoded[103]), .A0 (nx4936), .A1 (nx5180)) ;
    and02 ix1869 (.Y (decoded[102]), .A0 (nx4944), .A1 (nx5180)) ;
    and02 ix1873 (.Y (decoded[101]), .A0 (nx4952), .A1 (nx5180)) ;
    and02 ix1877 (.Y (decoded[100]), .A0 (nx4960), .A1 (nx5180)) ;
    and02 ix1881 (.Y (decoded[99]), .A0 (nx4968), .A1 (nx5180)) ;
    and02 ix1885 (.Y (decoded[98]), .A0 (nx4976), .A1 (nx5180)) ;
    and02 ix1889 (.Y (decoded[97]), .A0 (nx4984), .A1 (nx5182)) ;
    and02 ix1893 (.Y (decoded[96]), .A0 (nx4992), .A1 (nx5182)) ;
    and02 ix1901 (.Y (decoded[95]), .A0 (nx4872), .A1 (nx5186)) ;
    nor02ii ix4292 (.Y (nx4806), .A0 (nx4254), .A1 (nx3832)) ;
    and02 ix1905 (.Y (decoded[94]), .A0 (nx4880), .A1 (nx5186)) ;
    and02 ix1909 (.Y (decoded[93]), .A0 (nx4888), .A1 (nx5186)) ;
    and02 ix1913 (.Y (decoded[92]), .A0 (nx4896), .A1 (nx5186)) ;
    and02 ix1917 (.Y (decoded[91]), .A0 (nx4904), .A1 (nx5186)) ;
    and02 ix1921 (.Y (decoded[90]), .A0 (nx4912), .A1 (nx5186)) ;
    and02 ix1925 (.Y (decoded[89]), .A0 (nx4920), .A1 (nx5186)) ;
    and02 ix1929 (.Y (decoded[88]), .A0 (nx4928), .A1 (nx5188)) ;
    and02 ix1933 (.Y (decoded[87]), .A0 (nx4936), .A1 (nx5188)) ;
    and02 ix1937 (.Y (decoded[86]), .A0 (nx4944), .A1 (nx5188)) ;
    and02 ix1941 (.Y (decoded[85]), .A0 (nx4952), .A1 (nx5188)) ;
    and02 ix1945 (.Y (decoded[84]), .A0 (nx4960), .A1 (nx5188)) ;
    and02 ix1949 (.Y (decoded[83]), .A0 (nx4968), .A1 (nx5188)) ;
    and02 ix1953 (.Y (decoded[82]), .A0 (nx4976), .A1 (nx5188)) ;
    and02 ix1957 (.Y (decoded[81]), .A0 (nx4984), .A1 (nx5190)) ;
    and02 ix1961 (.Y (decoded[80]), .A0 (nx4992), .A1 (nx5190)) ;
    and02 ix1969 (.Y (decoded[79]), .A0 (nx4872), .A1 (nx5194)) ;
    nor02ii ix4310 (.Y (nx4814), .A0 (nx4254), .A1 (nx3854)) ;
    and02 ix1973 (.Y (decoded[78]), .A0 (nx4880), .A1 (nx5194)) ;
    and02 ix1977 (.Y (decoded[77]), .A0 (nx4888), .A1 (nx5194)) ;
    and02 ix1981 (.Y (decoded[76]), .A0 (nx4896), .A1 (nx5194)) ;
    and02 ix1985 (.Y (decoded[75]), .A0 (nx4904), .A1 (nx5194)) ;
    and02 ix1989 (.Y (decoded[74]), .A0 (nx4912), .A1 (nx5194)) ;
    and02 ix1993 (.Y (decoded[73]), .A0 (nx4920), .A1 (nx5194)) ;
    and02 ix1997 (.Y (decoded[72]), .A0 (nx4928), .A1 (nx5196)) ;
    and02 ix2001 (.Y (decoded[71]), .A0 (nx4936), .A1 (nx5196)) ;
    and02 ix2005 (.Y (decoded[70]), .A0 (nx4944), .A1 (nx5196)) ;
    and02 ix2009 (.Y (decoded[69]), .A0 (nx4952), .A1 (nx5196)) ;
    and02 ix2013 (.Y (decoded[68]), .A0 (nx4960), .A1 (nx5196)) ;
    and02 ix2017 (.Y (decoded[67]), .A0 (nx4968), .A1 (nx5196)) ;
    and02 ix2021 (.Y (decoded[66]), .A0 (nx4976), .A1 (nx5196)) ;
    and02 ix2025 (.Y (decoded[65]), .A0 (nx4984), .A1 (nx5198)) ;
    and02 ix2029 (.Y (decoded[64]), .A0 (nx4992), .A1 (nx5198)) ;
    and02 ix2045 (.Y (decoded[63]), .A0 (nx4406), .A1 (nx5200)) ;
    and02 ix2049 (.Y (decoded[62]), .A0 (nx4418), .A1 (nx5200)) ;
    and02 ix2053 (.Y (decoded[61]), .A0 (nx4430), .A1 (nx5200)) ;
    and02 ix2057 (.Y (decoded[60]), .A0 (nx4442), .A1 (nx5200)) ;
    and02 ix2061 (.Y (decoded[59]), .A0 (nx4454), .A1 (nx5200)) ;
    and02 ix2065 (.Y (decoded[58]), .A0 (nx4466), .A1 (nx5200)) ;
    and02 ix2069 (.Y (decoded[57]), .A0 (nx4478), .A1 (nx5200)) ;
    and02 ix2073 (.Y (decoded[56]), .A0 (nx4490), .A1 (nx5202)) ;
    and02 ix2077 (.Y (decoded[55]), .A0 (nx4502), .A1 (nx5202)) ;
    and02 ix2081 (.Y (decoded[54]), .A0 (nx4514), .A1 (nx5202)) ;
    and02 ix2085 (.Y (decoded[53]), .A0 (nx4526), .A1 (nx5202)) ;
    and02 ix2089 (.Y (decoded[52]), .A0 (nx4538), .A1 (nx5202)) ;
    and02 ix2093 (.Y (decoded[51]), .A0 (nx4550), .A1 (nx5202)) ;
    and02 ix2097 (.Y (decoded[50]), .A0 (nx4562), .A1 (nx5202)) ;
    and02 ix2101 (.Y (decoded[49]), .A0 (nx4574), .A1 (nx5204)) ;
    and02 ix2105 (.Y (decoded[48]), .A0 (nx4586), .A1 (nx5204)) ;
    and02 ix2113 (.Y (decoded[47]), .A0 (nx4406), .A1 (nx5208)) ;
    nor02ii ix4348 (.Y (nx4830), .A0 (nx4329), .A1 (nx3803)) ;
    and02 ix2117 (.Y (decoded[46]), .A0 (nx4418), .A1 (nx5208)) ;
    and02 ix2121 (.Y (decoded[45]), .A0 (nx4430), .A1 (nx5208)) ;
    and02 ix2125 (.Y (decoded[44]), .A0 (nx4442), .A1 (nx5208)) ;
    and02 ix2129 (.Y (decoded[43]), .A0 (nx4454), .A1 (nx5208)) ;
    and02 ix2133 (.Y (decoded[42]), .A0 (nx4466), .A1 (nx5208)) ;
    and02 ix2137 (.Y (decoded[41]), .A0 (nx4478), .A1 (nx5208)) ;
    and02 ix2141 (.Y (decoded[40]), .A0 (nx4490), .A1 (nx5210)) ;
    and02 ix2145 (.Y (decoded[39]), .A0 (nx4502), .A1 (nx5210)) ;
    and02 ix2149 (.Y (decoded[38]), .A0 (nx4514), .A1 (nx5210)) ;
    and02 ix2153 (.Y (decoded[37]), .A0 (nx4526), .A1 (nx5210)) ;
    and02 ix2157 (.Y (decoded[36]), .A0 (nx4538), .A1 (nx5210)) ;
    and02 ix2161 (.Y (decoded[35]), .A0 (nx4550), .A1 (nx5210)) ;
    and02 ix2165 (.Y (decoded[34]), .A0 (nx4562), .A1 (nx5210)) ;
    and02 ix2169 (.Y (decoded[33]), .A0 (nx4574), .A1 (nx5212)) ;
    and02 ix2173 (.Y (decoded[32]), .A0 (nx4586), .A1 (nx5212)) ;
    and02 ix2181 (.Y (decoded[31]), .A0 (nx4406), .A1 (nx5216)) ;
    nor02ii ix4367 (.Y (nx4838), .A0 (nx4329), .A1 (nx3832)) ;
    and02 ix2185 (.Y (decoded[30]), .A0 (nx4418), .A1 (nx5216)) ;
    and02 ix2189 (.Y (decoded[29]), .A0 (nx4430), .A1 (nx5216)) ;
    and02 ix2193 (.Y (decoded[28]), .A0 (nx4442), .A1 (nx5216)) ;
    and02 ix2197 (.Y (decoded[27]), .A0 (nx4454), .A1 (nx5216)) ;
    and02 ix2201 (.Y (decoded[26]), .A0 (nx4466), .A1 (nx5216)) ;
    and02 ix2205 (.Y (decoded[25]), .A0 (nx4478), .A1 (nx5216)) ;
    and02 ix2209 (.Y (decoded[24]), .A0 (nx4490), .A1 (nx5218)) ;
    and02 ix2213 (.Y (decoded[23]), .A0 (nx4502), .A1 (nx5218)) ;
    and02 ix2217 (.Y (decoded[22]), .A0 (nx4514), .A1 (nx5218)) ;
    and02 ix2221 (.Y (decoded[21]), .A0 (nx4526), .A1 (nx5218)) ;
    and02 ix2225 (.Y (decoded[20]), .A0 (nx4538), .A1 (nx5218)) ;
    and02 ix2229 (.Y (decoded[19]), .A0 (nx4550), .A1 (nx5218)) ;
    and02 ix2233 (.Y (decoded[18]), .A0 (nx4562), .A1 (nx5218)) ;
    and02 ix2237 (.Y (decoded[17]), .A0 (nx4574), .A1 (nx5220)) ;
    and02 ix2241 (.Y (decoded[16]), .A0 (nx4586), .A1 (nx5220)) ;
    and02 ix2249 (.Y (decoded[15]), .A0 (nx4406), .A1 (nx5224)) ;
    nor02ii ix4385 (.Y (nx4846), .A0 (nx4329), .A1 (nx3854)) ;
    and02 ix2253 (.Y (decoded[14]), .A0 (nx4418), .A1 (nx5224)) ;
    and02 ix2257 (.Y (decoded[13]), .A0 (nx4430), .A1 (nx5224)) ;
    and02 ix2261 (.Y (decoded[12]), .A0 (nx4442), .A1 (nx5224)) ;
    and02 ix2265 (.Y (decoded[11]), .A0 (nx4454), .A1 (nx5224)) ;
    and02 ix2269 (.Y (decoded[10]), .A0 (nx4466), .A1 (nx5224)) ;
    and02 ix2273 (.Y (decoded[9]), .A0 (nx4478), .A1 (nx5224)) ;
    and02 ix2277 (.Y (decoded[8]), .A0 (nx4490), .A1 (nx5226)) ;
    and02 ix2281 (.Y (decoded[7]), .A0 (nx4502), .A1 (nx5226)) ;
    and02 ix2285 (.Y (decoded[6]), .A0 (nx4514), .A1 (nx5226)) ;
    and02 ix2289 (.Y (decoded[5]), .A0 (nx4526), .A1 (nx5226)) ;
    and02 ix2293 (.Y (decoded[4]), .A0 (nx4538), .A1 (nx5226)) ;
    and02 ix2297 (.Y (decoded[3]), .A0 (nx4550), .A1 (nx5226)) ;
    and02 ix2301 (.Y (decoded[2]), .A0 (nx4562), .A1 (nx5226)) ;
    and02 ix2305 (.Y (decoded[1]), .A0 (nx4574), .A1 (nx5228)) ;
    and02 ix2309 (.Y (decoded[0]), .A0 (nx4586), .A1 (nx5228)) ;
    inv02 ix4857 (.Y (nx4858), .A (nx3810)) ;
    inv02 ix4859 (.Y (nx4860), .A (nx3812)) ;
    buf02 ix4861 (.Y (nx4862), .A (T[3])) ;
    buf02 ix4863 (.Y (nx4864), .A (T[1])) ;
    inv01 ix4865 (.Y (nx4866), .A (nx12)) ;
    inv01 ix4867 (.Y (nx4868), .A (nx12)) ;
    inv01 ix4869 (.Y (nx4870), .A (nx12)) ;
    inv01 ix4871 (.Y (nx4872), .A (nx12)) ;
    inv01 ix4873 (.Y (nx4874), .A (nx38)) ;
    inv01 ix4875 (.Y (nx4876), .A (nx38)) ;
    inv01 ix4877 (.Y (nx4878), .A (nx38)) ;
    inv01 ix4879 (.Y (nx4880), .A (nx38)) ;
    inv01 ix4881 (.Y (nx4882), .A (nx48)) ;
    inv01 ix4883 (.Y (nx4884), .A (nx48)) ;
    inv01 ix4885 (.Y (nx4886), .A (nx48)) ;
    inv01 ix4887 (.Y (nx4888), .A (nx48)) ;
    inv01 ix4889 (.Y (nx4890), .A (nx56)) ;
    inv01 ix4891 (.Y (nx4892), .A (nx56)) ;
    inv01 ix4893 (.Y (nx4894), .A (nx56)) ;
    inv01 ix4895 (.Y (nx4896), .A (nx56)) ;
    inv01 ix4897 (.Y (nx4898), .A (nx66)) ;
    inv01 ix4899 (.Y (nx4900), .A (nx66)) ;
    inv01 ix4901 (.Y (nx4902), .A (nx66)) ;
    inv01 ix4903 (.Y (nx4904), .A (nx66)) ;
    inv01 ix4905 (.Y (nx4906), .A (nx72)) ;
    inv01 ix4907 (.Y (nx4908), .A (nx72)) ;
    inv01 ix4909 (.Y (nx4910), .A (nx72)) ;
    inv01 ix4911 (.Y (nx4912), .A (nx72)) ;
    inv01 ix4913 (.Y (nx4914), .A (nx78)) ;
    inv01 ix4915 (.Y (nx4916), .A (nx78)) ;
    inv01 ix4917 (.Y (nx4918), .A (nx78)) ;
    inv01 ix4919 (.Y (nx4920), .A (nx78)) ;
    inv01 ix4921 (.Y (nx4922), .A (nx84)) ;
    inv01 ix4923 (.Y (nx4924), .A (nx84)) ;
    inv01 ix4925 (.Y (nx4926), .A (nx84)) ;
    inv01 ix4927 (.Y (nx4928), .A (nx84)) ;
    inv01 ix4929 (.Y (nx4930), .A (nx94)) ;
    inv01 ix4931 (.Y (nx4932), .A (nx94)) ;
    inv01 ix4933 (.Y (nx4934), .A (nx94)) ;
    inv01 ix4935 (.Y (nx4936), .A (nx94)) ;
    inv01 ix4937 (.Y (nx4938), .A (nx100)) ;
    inv01 ix4939 (.Y (nx4940), .A (nx100)) ;
    inv01 ix4941 (.Y (nx4942), .A (nx100)) ;
    inv01 ix4943 (.Y (nx4944), .A (nx100)) ;
    inv01 ix4945 (.Y (nx4946), .A (nx106)) ;
    inv01 ix4947 (.Y (nx4948), .A (nx106)) ;
    inv01 ix4949 (.Y (nx4950), .A (nx106)) ;
    inv01 ix4951 (.Y (nx4952), .A (nx106)) ;
    inv01 ix4953 (.Y (nx4954), .A (nx112)) ;
    inv01 ix4955 (.Y (nx4956), .A (nx112)) ;
    inv01 ix4957 (.Y (nx4958), .A (nx112)) ;
    inv01 ix4959 (.Y (nx4960), .A (nx112)) ;
    inv01 ix4961 (.Y (nx4962), .A (nx120)) ;
    inv01 ix4963 (.Y (nx4964), .A (nx120)) ;
    inv01 ix4965 (.Y (nx4966), .A (nx120)) ;
    inv01 ix4967 (.Y (nx4968), .A (nx120)) ;
    inv01 ix4969 (.Y (nx4970), .A (nx126)) ;
    inv01 ix4971 (.Y (nx4972), .A (nx126)) ;
    inv01 ix4973 (.Y (nx4974), .A (nx126)) ;
    inv01 ix4975 (.Y (nx4976), .A (nx126)) ;
    inv01 ix4977 (.Y (nx4978), .A (nx132)) ;
    inv01 ix4979 (.Y (nx4980), .A (nx132)) ;
    inv01 ix4981 (.Y (nx4982), .A (nx132)) ;
    inv01 ix4983 (.Y (nx4984), .A (nx132)) ;
    inv01 ix4985 (.Y (nx4986), .A (nx138)) ;
    inv01 ix4987 (.Y (nx4988), .A (nx138)) ;
    inv01 ix4989 (.Y (nx4990), .A (nx138)) ;
    inv01 ix4991 (.Y (nx4992), .A (nx138)) ;
    inv02 ix4993 (.Y (nx4994), .A (nx3745)) ;
    inv02 ix4995 (.Y (nx4996), .A (nx3745)) ;
    inv02 ix4997 (.Y (nx4998), .A (nx3745)) ;
    inv01 ix4999 (.Y (nx5000), .A (nx4606)) ;
    inv02 ix5001 (.Y (nx5002), .A (nx5000)) ;
    inv02 ix5003 (.Y (nx5004), .A (nx5000)) ;
    inv02 ix5005 (.Y (nx5006), .A (nx5000)) ;
    inv01 ix5007 (.Y (nx5008), .A (nx4614)) ;
    inv02 ix5009 (.Y (nx5010), .A (nx5008)) ;
    inv02 ix5011 (.Y (nx5012), .A (nx5008)) ;
    inv02 ix5013 (.Y (nx5014), .A (nx5008)) ;
    inv01 ix5015 (.Y (nx5016), .A (nx4622)) ;
    inv02 ix5017 (.Y (nx5018), .A (nx5016)) ;
    inv02 ix5019 (.Y (nx5020), .A (nx5016)) ;
    inv02 ix5021 (.Y (nx5022), .A (nx5016)) ;
    inv02 ix5023 (.Y (nx5024), .A (nx3872)) ;
    inv02 ix5025 (.Y (nx5026), .A (nx3872)) ;
    inv02 ix5027 (.Y (nx5028), .A (nx3872)) ;
    inv01 ix5029 (.Y (nx5030), .A (nx4638)) ;
    inv02 ix5031 (.Y (nx5032), .A (nx5030)) ;
    inv02 ix5033 (.Y (nx5034), .A (nx5030)) ;
    inv02 ix5035 (.Y (nx5036), .A (nx5030)) ;
    inv01 ix5037 (.Y (nx5038), .A (nx4646)) ;
    inv02 ix5039 (.Y (nx5040), .A (nx5038)) ;
    inv02 ix5041 (.Y (nx5042), .A (nx5038)) ;
    inv02 ix5043 (.Y (nx5044), .A (nx5038)) ;
    inv01 ix5045 (.Y (nx5046), .A (nx4654)) ;
    inv02 ix5047 (.Y (nx5048), .A (nx5046)) ;
    inv02 ix5049 (.Y (nx5050), .A (nx5046)) ;
    inv02 ix5051 (.Y (nx5052), .A (nx5046)) ;
    inv02 ix5053 (.Y (nx5054), .A (nx3947)) ;
    inv02 ix5055 (.Y (nx5056), .A (nx3947)) ;
    inv02 ix5057 (.Y (nx5058), .A (nx3947)) ;
    inv01 ix5059 (.Y (nx5060), .A (nx4670)) ;
    inv02 ix5061 (.Y (nx5062), .A (nx5060)) ;
    inv02 ix5063 (.Y (nx5064), .A (nx5060)) ;
    inv02 ix5065 (.Y (nx5066), .A (nx5060)) ;
    inv01 ix5067 (.Y (nx5068), .A (nx4678)) ;
    inv02 ix5069 (.Y (nx5070), .A (nx5068)) ;
    inv02 ix5071 (.Y (nx5072), .A (nx5068)) ;
    inv02 ix5073 (.Y (nx5074), .A (nx5068)) ;
    inv01 ix5075 (.Y (nx5076), .A (nx4686)) ;
    inv02 ix5077 (.Y (nx5078), .A (nx5076)) ;
    inv02 ix5079 (.Y (nx5080), .A (nx5076)) ;
    inv02 ix5081 (.Y (nx5082), .A (nx5076)) ;
    inv01 ix5083 (.Y (nx5084), .A (nx4694)) ;
    inv02 ix5085 (.Y (nx5086), .A (nx5084)) ;
    inv02 ix5087 (.Y (nx5088), .A (nx5084)) ;
    inv02 ix5089 (.Y (nx5090), .A (nx5084)) ;
    inv02 ix5091 (.Y (nx5092), .A (nx4043)) ;
    inv02 ix5093 (.Y (nx5094), .A (nx4043)) ;
    inv02 ix5095 (.Y (nx5096), .A (nx4043)) ;
    inv02 ix5097 (.Y (nx5098), .A (nx4061)) ;
    inv02 ix5099 (.Y (nx5100), .A (nx4061)) ;
    inv02 ix5101 (.Y (nx5102), .A (nx4061)) ;
    inv02 ix5103 (.Y (nx5104), .A (nx4079)) ;
    inv02 ix5105 (.Y (nx5106), .A (nx4079)) ;
    inv02 ix5107 (.Y (nx5108), .A (nx4079)) ;
    inv02 ix5109 (.Y (nx5110), .A (nx4097)) ;
    inv02 ix5111 (.Y (nx5112), .A (nx4097)) ;
    inv02 ix5113 (.Y (nx5114), .A (nx4097)) ;
    inv01 ix5115 (.Y (nx5116), .A (nx4734)) ;
    inv02 ix5117 (.Y (nx5118), .A (nx5116)) ;
    inv02 ix5119 (.Y (nx5120), .A (nx5116)) ;
    inv02 ix5121 (.Y (nx5122), .A (nx5116)) ;
    inv01 ix5123 (.Y (nx5124), .A (nx4742)) ;
    inv02 ix5125 (.Y (nx5126), .A (nx5124)) ;
    inv02 ix5127 (.Y (nx5128), .A (nx5124)) ;
    inv02 ix5129 (.Y (nx5130), .A (nx5124)) ;
    inv01 ix5131 (.Y (nx5132), .A (nx4750)) ;
    inv02 ix5133 (.Y (nx5134), .A (nx5132)) ;
    inv02 ix5135 (.Y (nx5136), .A (nx5132)) ;
    inv02 ix5137 (.Y (nx5138), .A (nx5132)) ;
    inv02 ix5139 (.Y (nx5140), .A (nx4173)) ;
    inv02 ix5141 (.Y (nx5142), .A (nx4173)) ;
    inv02 ix5143 (.Y (nx5144), .A (nx4173)) ;
    inv01 ix5145 (.Y (nx5146), .A (nx4766)) ;
    inv02 ix5147 (.Y (nx5148), .A (nx5146)) ;
    inv02 ix5149 (.Y (nx5150), .A (nx5146)) ;
    inv02 ix5151 (.Y (nx5152), .A (nx5146)) ;
    inv01 ix5153 (.Y (nx5154), .A (nx4774)) ;
    inv02 ix5155 (.Y (nx5156), .A (nx5154)) ;
    inv02 ix5157 (.Y (nx5158), .A (nx5154)) ;
    inv02 ix5159 (.Y (nx5160), .A (nx5154)) ;
    inv01 ix5161 (.Y (nx5162), .A (nx4782)) ;
    inv02 ix5163 (.Y (nx5164), .A (nx5162)) ;
    inv02 ix5165 (.Y (nx5166), .A (nx5162)) ;
    inv02 ix5167 (.Y (nx5168), .A (nx5162)) ;
    inv02 ix5169 (.Y (nx5170), .A (nx4252)) ;
    inv02 ix5171 (.Y (nx5172), .A (nx4252)) ;
    inv02 ix5173 (.Y (nx5174), .A (nx4252)) ;
    inv01 ix5175 (.Y (nx5176), .A (nx4798)) ;
    inv02 ix5177 (.Y (nx5178), .A (nx5176)) ;
    inv02 ix5179 (.Y (nx5180), .A (nx5176)) ;
    inv02 ix5181 (.Y (nx5182), .A (nx5176)) ;
    inv01 ix5183 (.Y (nx5184), .A (nx4806)) ;
    inv02 ix5185 (.Y (nx5186), .A (nx5184)) ;
    inv02 ix5187 (.Y (nx5188), .A (nx5184)) ;
    inv02 ix5189 (.Y (nx5190), .A (nx5184)) ;
    inv01 ix5191 (.Y (nx5192), .A (nx4814)) ;
    inv02 ix5193 (.Y (nx5194), .A (nx5192)) ;
    inv02 ix5195 (.Y (nx5196), .A (nx5192)) ;
    inv02 ix5197 (.Y (nx5198), .A (nx5192)) ;
    inv02 ix5199 (.Y (nx5200), .A (nx4327)) ;
    inv02 ix5201 (.Y (nx5202), .A (nx4327)) ;
    inv02 ix5203 (.Y (nx5204), .A (nx4327)) ;
    inv01 ix5205 (.Y (nx5206), .A (nx4830)) ;
    inv02 ix5207 (.Y (nx5208), .A (nx5206)) ;
    inv02 ix5209 (.Y (nx5210), .A (nx5206)) ;
    inv02 ix5211 (.Y (nx5212), .A (nx5206)) ;
    inv01 ix5213 (.Y (nx5214), .A (nx4838)) ;
    inv02 ix5215 (.Y (nx5216), .A (nx5214)) ;
    inv02 ix5217 (.Y (nx5218), .A (nx5214)) ;
    inv02 ix5219 (.Y (nx5220), .A (nx5214)) ;
    inv01 ix5221 (.Y (nx5222), .A (nx4846)) ;
    inv02 ix5223 (.Y (nx5224), .A (nx5222)) ;
    inv02 ix5225 (.Y (nx5226), .A (nx5222)) ;
    inv02 ix5227 (.Y (nx5228), .A (nx5222)) ;
endmodule


module DMAController_12_13_8_16_5 ( clk, reset, weightsInternalBus, 
                                    windowInternalBus, writeInternalBus, 
                                    weightsRamAddress, windowRamAddressRead, 
                                    windowRamAddressWrite, weightsRamDataInBus, 
                                    windowRamDataInBus, weightsRamRead, 
                                    windowRamRead, windowRamWrite, 
                                    windowRamDataOutBus, MFCWindowRam, 
                                    MFCWeightsRam, MFCWrite, loadNextFilter, 
                                    loadNextWindow, loadNextRow, loadOneWord, 
                                    loadThreeWord, filterFinished, sliceFinished, 
                                    layerFinished, layerType, write, 
                                    weightsSizeType, inputSize, outputSize, 
                                    windowRamBaseAddress1, windowRamBaseAddress2, 
                                    filterRamBaseAddress, windowReadOne, 
                                    windowReadFinal, weightsReadOne, 
                                    weightsReadFinal, writeDoneAll, writeDoneOne, 
                                    filterAluNumber, windowAluNumber ) ;

    input clk ;
    input reset ;
    output [39:0]weightsInternalBus ;
    output [79:0]windowInternalBus ;
    input [15:0]writeInternalBus ;
    output [11:0]weightsRamAddress ;
    output [12:0]windowRamAddressRead ;
    output [12:0]windowRamAddressWrite ;
    input [39:0]weightsRamDataInBus ;
    input [79:0]windowRamDataInBus ;
    output weightsRamRead ;
    output windowRamRead ;
    output windowRamWrite ;
    output [15:0]windowRamDataOutBus ;
    input MFCWindowRam ;
    input MFCWeightsRam ;
    input MFCWrite ;
    input loadNextFilter ;
    input loadNextWindow ;
    input loadNextRow ;
    input loadOneWord ;
    input loadThreeWord ;
    input filterFinished ;
    input sliceFinished ;
    input layerFinished ;
    input layerType ;
    input write ;
    input weightsSizeType ;
    input [12:0]inputSize ;
    input [12:0]outputSize ;
    input [12:0]windowRamBaseAddress1 ;
    input [12:0]windowRamBaseAddress2 ;
    input [11:0]filterRamBaseAddress ;
    output windowReadOne ;
    output windowReadFinal ;
    output weightsReadOne ;
    output weightsReadFinal ;
    output writeDoneAll ;
    output writeDoneOne ;
    output [2:0]filterAluNumber ;
    output [2:0]windowAluNumber ;

    wire currentReadRamBaseAddress_12, currentReadRamBaseAddress_11, 
         currentReadRamBaseAddress_10, currentReadRamBaseAddress_9, 
         currentReadRamBaseAddress_8, currentReadRamBaseAddress_7, 
         currentReadRamBaseAddress_6, currentReadRamBaseAddress_5, 
         currentReadRamBaseAddress_4, currentReadRamBaseAddress_3, 
         currentReadRamBaseAddress_2, currentReadRamBaseAddress_1, 
         currentReadRamBaseAddress_0, currentWriteRamBaseAddress_12, 
         currentWriteRamBaseAddress_11, currentWriteRamBaseAddress_10, 
         currentWriteRamBaseAddress_9, currentWriteRamBaseAddress_8, 
         currentWriteRamBaseAddress_7, currentWriteRamBaseAddress_6, 
         currentWriteRamBaseAddress_5, currentWriteRamBaseAddress_4, 
         currentWriteRamBaseAddress_3, currentWriteRamBaseAddress_2, 
         currentWriteRamBaseAddress_1, currentWriteRamBaseAddress_0, 
         ramBaseAddressSelector, windowInternalBusRLogic_79, 
         windowInternalBusRLogic_78, windowInternalBusRLogic_77, 
         windowInternalBusRLogic_76, windowInternalBusRLogic_75, 
         windowInternalBusRLogic_74, windowInternalBusRLogic_73, 
         windowInternalBusRLogic_72, windowInternalBusRLogic_71, 
         windowInternalBusRLogic_70, windowInternalBusRLogic_69, 
         windowInternalBusRLogic_68, windowInternalBusRLogic_67, 
         windowInternalBusRLogic_66, windowInternalBusRLogic_65, 
         windowInternalBusRLogic_64, windowInternalBusRLogic_63, 
         windowInternalBusRLogic_62, windowInternalBusRLogic_61, 
         windowInternalBusRLogic_60, windowInternalBusRLogic_59, 
         windowInternalBusRLogic_58, windowInternalBusRLogic_57, 
         windowInternalBusRLogic_56, windowInternalBusRLogic_55, 
         windowInternalBusRLogic_54, windowInternalBusRLogic_53, 
         windowInternalBusRLogic_52, windowInternalBusRLogic_51, 
         windowInternalBusRLogic_50, windowInternalBusRLogic_49, 
         windowInternalBusRLogic_48, windowInternalBusRLogic_47, 
         windowInternalBusRLogic_46, windowInternalBusRLogic_45, 
         windowInternalBusRLogic_44, windowInternalBusRLogic_43, 
         windowInternalBusRLogic_42, windowInternalBusRLogic_41, 
         windowInternalBusRLogic_40, windowInternalBusRLogic_39, 
         windowInternalBusRLogic_38, windowInternalBusRLogic_37, 
         windowInternalBusRLogic_36, windowInternalBusRLogic_35, 
         windowInternalBusRLogic_34, windowInternalBusRLogic_33, 
         windowInternalBusRLogic_32, windowInternalBusRLogic_31, 
         windowInternalBusRLogic_30, windowInternalBusRLogic_29, 
         windowInternalBusRLogic_28, windowInternalBusRLogic_27, 
         windowInternalBusRLogic_26, windowInternalBusRLogic_25, 
         windowInternalBusRLogic_24, windowInternalBusRLogic_23, 
         windowInternalBusRLogic_22, windowInternalBusRLogic_21, 
         windowInternalBusRLogic_20, windowInternalBusRLogic_19, 
         windowInternalBusRLogic_18, windowInternalBusRLogic_17, 
         windowInternalBusRLogic_16, windowInternalBusRLogic_15, 
         windowInternalBusRLogic_14, windowInternalBusRLogic_13, 
         windowInternalBusRLogic_12, windowInternalBusRLogic_11, 
         windowInternalBusRLogic_10, windowInternalBusRLogic_9, 
         windowInternalBusRLogic_8, windowInternalBusRLogic_7, 
         windowInternalBusRLogic_6, windowInternalBusRLogic_5, 
         windowInternalBusRLogic_4, windowInternalBusRLogic_3, 
         windowInternalBusRLogic_2, windowInternalBusRLogic_1, 
         windowInternalBusRLogic_0, switchRam, windowRLSwitchRam, filterStep_2, 
         filterStep_1, writeFinishFilter, loadWord, resetLogics, 
         weightsSizeForWindow_0, NOT_weightsSizeType_dup_606, NOT__4681, nx614;
    wire [15:0] \$dummy ;




    Mux2_13 readRamMux (.A ({windowRamBaseAddress1[12],windowRamBaseAddress1[11]
            ,windowRamBaseAddress1[10],windowRamBaseAddress1[9],
            windowRamBaseAddress1[8],windowRamBaseAddress1[7],
            windowRamBaseAddress1[6],windowRamBaseAddress1[5],
            windowRamBaseAddress1[4],windowRamBaseAddress1[3],
            windowRamBaseAddress1[2],windowRamBaseAddress1[1],
            windowRamBaseAddress1[0]}), .B ({windowRamBaseAddress2[12],
            windowRamBaseAddress2[11],windowRamBaseAddress2[10],
            windowRamBaseAddress2[9],windowRamBaseAddress2[8],
            windowRamBaseAddress2[7],windowRamBaseAddress2[6],
            windowRamBaseAddress2[5],windowRamBaseAddress2[4],
            windowRamBaseAddress2[3],windowRamBaseAddress2[2],
            windowRamBaseAddress2[1],windowRamBaseAddress2[0]}), .S (
            ramBaseAddressSelector), .C ({currentReadRamBaseAddress_12,
            currentReadRamBaseAddress_11,currentReadRamBaseAddress_10,
            currentReadRamBaseAddress_9,currentReadRamBaseAddress_8,
            currentReadRamBaseAddress_7,currentReadRamBaseAddress_6,
            currentReadRamBaseAddress_5,currentReadRamBaseAddress_4,
            currentReadRamBaseAddress_3,currentReadRamBaseAddress_2,
            currentReadRamBaseAddress_1,currentReadRamBaseAddress_0})) ;
    Mux2_13 writeRamMux (.A ({windowRamBaseAddress2[12],
            windowRamBaseAddress2[11],windowRamBaseAddress2[10],
            windowRamBaseAddress2[9],windowRamBaseAddress2[8],
            windowRamBaseAddress2[7],windowRamBaseAddress2[6],
            windowRamBaseAddress2[5],windowRamBaseAddress2[4],
            windowRamBaseAddress2[3],windowRamBaseAddress2[2],
            windowRamBaseAddress2[1],windowRamBaseAddress2[0]}), .B ({
            windowRamBaseAddress1[12],windowRamBaseAddress1[11],
            windowRamBaseAddress1[10],windowRamBaseAddress1[9],
            windowRamBaseAddress1[8],windowRamBaseAddress1[7],
            windowRamBaseAddress1[6],windowRamBaseAddress1[5],
            windowRamBaseAddress1[4],windowRamBaseAddress1[3],
            windowRamBaseAddress1[2],windowRamBaseAddress1[1],
            windowRamBaseAddress1[0]}), .S (ramBaseAddressSelector), .C ({
            currentWriteRamBaseAddress_12,currentWriteRamBaseAddress_11,
            currentWriteRamBaseAddress_10,currentWriteRamBaseAddress_9,
            currentWriteRamBaseAddress_8,currentWriteRamBaseAddress_7,
            currentWriteRamBaseAddress_6,currentWriteRamBaseAddress_5,
            currentWriteRamBaseAddress_4,currentWriteRamBaseAddress_3,
            currentWriteRamBaseAddress_2,currentWriteRamBaseAddress_1,
            currentWriteRamBaseAddress_0})) ;
    Tristate_80 readLogicTri (.\input  ({windowInternalBusRLogic_79,
                windowInternalBusRLogic_78,windowInternalBusRLogic_77,
                windowInternalBusRLogic_76,windowInternalBusRLogic_75,
                windowInternalBusRLogic_74,windowInternalBusRLogic_73,
                windowInternalBusRLogic_72,windowInternalBusRLogic_71,
                windowInternalBusRLogic_70,windowInternalBusRLogic_69,
                windowInternalBusRLogic_68,windowInternalBusRLogic_67,
                windowInternalBusRLogic_66,windowInternalBusRLogic_65,
                windowInternalBusRLogic_64,windowInternalBusRLogic_63,
                windowInternalBusRLogic_62,windowInternalBusRLogic_61,
                windowInternalBusRLogic_60,windowInternalBusRLogic_59,
                windowInternalBusRLogic_58,windowInternalBusRLogic_57,
                windowInternalBusRLogic_56,windowInternalBusRLogic_55,
                windowInternalBusRLogic_54,windowInternalBusRLogic_53,
                windowInternalBusRLogic_52,windowInternalBusRLogic_51,
                windowInternalBusRLogic_50,windowInternalBusRLogic_49,
                windowInternalBusRLogic_48,windowInternalBusRLogic_47,
                windowInternalBusRLogic_46,windowInternalBusRLogic_45,
                windowInternalBusRLogic_44,windowInternalBusRLogic_43,
                windowInternalBusRLogic_42,windowInternalBusRLogic_41,
                windowInternalBusRLogic_40,windowInternalBusRLogic_39,
                windowInternalBusRLogic_38,windowInternalBusRLogic_37,
                windowInternalBusRLogic_36,windowInternalBusRLogic_35,
                windowInternalBusRLogic_34,windowInternalBusRLogic_33,
                windowInternalBusRLogic_32,windowInternalBusRLogic_31,
                windowInternalBusRLogic_30,windowInternalBusRLogic_29,
                windowInternalBusRLogic_28,windowInternalBusRLogic_27,
                windowInternalBusRLogic_26,windowInternalBusRLogic_25,
                windowInternalBusRLogic_24,windowInternalBusRLogic_23,
                windowInternalBusRLogic_22,windowInternalBusRLogic_21,
                windowInternalBusRLogic_20,windowInternalBusRLogic_19,
                windowInternalBusRLogic_18,windowInternalBusRLogic_17,
                windowInternalBusRLogic_16,windowInternalBusRLogic_15,
                windowInternalBusRLogic_14,windowInternalBusRLogic_13,
                windowInternalBusRLogic_12,windowInternalBusRLogic_11,
                windowInternalBusRLogic_10,windowInternalBusRLogic_9,
                windowInternalBusRLogic_8,windowInternalBusRLogic_7,
                windowInternalBusRLogic_6,windowInternalBusRLogic_5,
                windowInternalBusRLogic_4,windowInternalBusRLogic_3,
                windowInternalBusRLogic_2,windowInternalBusRLogic_1,
                windowInternalBusRLogic_0}), .en (weightsSizeForWindow_0), .\output  (
                {windowInternalBus[79],windowInternalBus[78],
                windowInternalBus[77],windowInternalBus[76],
                windowInternalBus[75],windowInternalBus[74],
                windowInternalBus[73],windowInternalBus[72],
                windowInternalBus[71],windowInternalBus[70],
                windowInternalBus[69],windowInternalBus[68],
                windowInternalBus[67],windowInternalBus[66],
                windowInternalBus[65],windowInternalBus[64],
                windowInternalBus[63],windowInternalBus[62],
                windowInternalBus[61],windowInternalBus[60],
                windowInternalBus[59],windowInternalBus[58],
                windowInternalBus[57],windowInternalBus[56],
                windowInternalBus[55],windowInternalBus[54],
                windowInternalBus[53],windowInternalBus[52],
                windowInternalBus[51],windowInternalBus[50],
                windowInternalBus[49],windowInternalBus[48],
                windowInternalBus[47],windowInternalBus[46],
                windowInternalBus[45],windowInternalBus[44],
                windowInternalBus[43],windowInternalBus[42],
                windowInternalBus[41],windowInternalBus[40],
                windowInternalBus[39],windowInternalBus[38],
                windowInternalBus[37],windowInternalBus[36],
                windowInternalBus[35],windowInternalBus[34],
                windowInternalBus[33],windowInternalBus[32],
                windowInternalBus[31],windowInternalBus[30],
                windowInternalBus[29],windowInternalBus[28],
                windowInternalBus[27],windowInternalBus[26],
                windowInternalBus[25],windowInternalBus[24],
                windowInternalBus[23],windowInternalBus[22],
                windowInternalBus[21],windowInternalBus[20],
                windowInternalBus[19],windowInternalBus[18],
                windowInternalBus[17],windowInternalBus[16],
                windowInternalBus[15],windowInternalBus[14],
                windowInternalBus[13],windowInternalBus[12],
                windowInternalBus[11],windowInternalBus[10],windowInternalBus[9]
                ,windowInternalBus[8],windowInternalBus[7],windowInternalBus[6],
                windowInternalBus[5],windowInternalBus[4],windowInternalBus[3],
                windowInternalBus[2],windowInternalBus[1],windowInternalBus[0]})
                ) ;
    Tristate_16 writeLogicTri (.\input  ({writeInternalBus[15],
                writeInternalBus[14],writeInternalBus[13],writeInternalBus[12],
                writeInternalBus[11],writeInternalBus[10],writeInternalBus[9],
                writeInternalBus[8],writeInternalBus[7],writeInternalBus[6],
                writeInternalBus[5],writeInternalBus[4],writeInternalBus[3],
                writeInternalBus[2],writeInternalBus[1],writeInternalBus[0]}), .en (
                weightsSizeForWindow_0), .\output  ({windowRamDataOutBus[15],
                windowRamDataOutBus[14],windowRamDataOutBus[13],
                windowRamDataOutBus[12],windowRamDataOutBus[11],
                windowRamDataOutBus[10],windowRamDataOutBus[9],
                windowRamDataOutBus[8],windowRamDataOutBus[7],
                windowRamDataOutBus[6],windowRamDataOutBus[5],
                windowRamDataOutBus[4],windowRamDataOutBus[3],
                windowRamDataOutBus[2],windowRamDataOutBus[1],
                windowRamDataOutBus[0]})) ;
    ReadLogic_13_80_false windowReadLogicEnt (.clk (clk), .resetState (
                          resetLogics), .switchRam (windowRLSwitchRam), .ramBasedAddress (
                          {currentReadRamBaseAddress_12,
                          currentReadRamBaseAddress_11,
                          currentReadRamBaseAddress_10,
                          currentReadRamBaseAddress_9,
                          currentReadRamBaseAddress_8,
                          currentReadRamBaseAddress_7,
                          currentReadRamBaseAddress_6,
                          currentReadRamBaseAddress_5,
                          currentReadRamBaseAddress_4,
                          currentReadRamBaseAddress_3,
                          currentReadRamBaseAddress_2,
                          currentReadRamBaseAddress_1,
                          currentReadRamBaseAddress_0}), .internalBus ({
                          windowInternalBusRLogic_79,windowInternalBusRLogic_78,
                          windowInternalBusRLogic_77,windowInternalBusRLogic_76,
                          windowInternalBusRLogic_75,windowInternalBusRLogic_74,
                          windowInternalBusRLogic_73,windowInternalBusRLogic_72,
                          windowInternalBusRLogic_71,windowInternalBusRLogic_70,
                          windowInternalBusRLogic_69,windowInternalBusRLogic_68,
                          windowInternalBusRLogic_67,windowInternalBusRLogic_66,
                          windowInternalBusRLogic_65,windowInternalBusRLogic_64,
                          windowInternalBusRLogic_63,windowInternalBusRLogic_62,
                          windowInternalBusRLogic_61,windowInternalBusRLogic_60,
                          windowInternalBusRLogic_59,windowInternalBusRLogic_58,
                          windowInternalBusRLogic_57,windowInternalBusRLogic_56,
                          windowInternalBusRLogic_55,windowInternalBusRLogic_54,
                          windowInternalBusRLogic_53,windowInternalBusRLogic_52,
                          windowInternalBusRLogic_51,windowInternalBusRLogic_50,
                          windowInternalBusRLogic_49,windowInternalBusRLogic_48,
                          windowInternalBusRLogic_47,windowInternalBusRLogic_46,
                          windowInternalBusRLogic_45,windowInternalBusRLogic_44,
                          windowInternalBusRLogic_43,windowInternalBusRLogic_42,
                          windowInternalBusRLogic_41,windowInternalBusRLogic_40,
                          windowInternalBusRLogic_39,windowInternalBusRLogic_38,
                          windowInternalBusRLogic_37,windowInternalBusRLogic_36,
                          windowInternalBusRLogic_35,windowInternalBusRLogic_34,
                          windowInternalBusRLogic_33,windowInternalBusRLogic_32,
                          windowInternalBusRLogic_31,windowInternalBusRLogic_30,
                          windowInternalBusRLogic_29,windowInternalBusRLogic_28,
                          windowInternalBusRLogic_27,windowInternalBusRLogic_26,
                          windowInternalBusRLogic_25,windowInternalBusRLogic_24,
                          windowInternalBusRLogic_23,windowInternalBusRLogic_22,
                          windowInternalBusRLogic_21,windowInternalBusRLogic_20,
                          windowInternalBusRLogic_19,windowInternalBusRLogic_18,
                          windowInternalBusRLogic_17,windowInternalBusRLogic_16,
                          windowInternalBusRLogic_15,windowInternalBusRLogic_14,
                          windowInternalBusRLogic_13,windowInternalBusRLogic_12,
                          windowInternalBusRLogic_11,windowInternalBusRLogic_10,
                          windowInternalBusRLogic_9,windowInternalBusRLogic_8,
                          windowInternalBusRLogic_7,windowInternalBusRLogic_6,
                          windowInternalBusRLogic_5,windowInternalBusRLogic_4,
                          windowInternalBusRLogic_3,windowInternalBusRLogic_2,
                          windowInternalBusRLogic_1,windowInternalBusRLogic_0})
                          , .ramDataInBus ({windowRamDataInBus[79],
                          windowRamDataInBus[78],windowRamDataInBus[77],
                          windowRamDataInBus[76],windowRamDataInBus[75],
                          windowRamDataInBus[74],windowRamDataInBus[73],
                          windowRamDataInBus[72],windowRamDataInBus[71],
                          windowRamDataInBus[70],windowRamDataInBus[69],
                          windowRamDataInBus[68],windowRamDataInBus[67],
                          windowRamDataInBus[66],windowRamDataInBus[65],
                          windowRamDataInBus[64],windowRamDataInBus[63],
                          windowRamDataInBus[62],windowRamDataInBus[61],
                          windowRamDataInBus[60],windowRamDataInBus[59],
                          windowRamDataInBus[58],windowRamDataInBus[57],
                          windowRamDataInBus[56],windowRamDataInBus[55],
                          windowRamDataInBus[54],windowRamDataInBus[53],
                          windowRamDataInBus[52],windowRamDataInBus[51],
                          windowRamDataInBus[50],windowRamDataInBus[49],
                          windowRamDataInBus[48],windowRamDataInBus[47],
                          windowRamDataInBus[46],windowRamDataInBus[45],
                          windowRamDataInBus[44],windowRamDataInBus[43],
                          windowRamDataInBus[42],windowRamDataInBus[41],
                          windowRamDataInBus[40],windowRamDataInBus[39],
                          windowRamDataInBus[38],windowRamDataInBus[37],
                          windowRamDataInBus[36],windowRamDataInBus[35],
                          windowRamDataInBus[34],windowRamDataInBus[33],
                          windowRamDataInBus[32],windowRamDataInBus[31],
                          windowRamDataInBus[30],windowRamDataInBus[29],
                          windowRamDataInBus[28],windowRamDataInBus[27],
                          windowRamDataInBus[26],windowRamDataInBus[25],
                          windowRamDataInBus[24],windowRamDataInBus[23],
                          windowRamDataInBus[22],windowRamDataInBus[21],
                          windowRamDataInBus[20],windowRamDataInBus[19],
                          windowRamDataInBus[18],windowRamDataInBus[17],
                          windowRamDataInBus[16],windowRamDataInBus[15],
                          windowRamDataInBus[14],windowRamDataInBus[13],
                          windowRamDataInBus[12],windowRamDataInBus[11],
                          windowRamDataInBus[10],windowRamDataInBus[9],
                          windowRamDataInBus[8],windowRamDataInBus[7],
                          windowRamDataInBus[6],windowRamDataInBus[5],
                          windowRamDataInBus[4],windowRamDataInBus[3],
                          windowRamDataInBus[2],windowRamDataInBus[1],
                          windowRamDataInBus[0]}), .ramRead (windowRamRead), .ramAddress (
                          {windowRamAddressRead[12],windowRamAddressRead[11],
                          windowRamAddressRead[10],windowRamAddressRead[9],
                          windowRamAddressRead[8],windowRamAddressRead[7],
                          windowRamAddressRead[6],windowRamAddressRead[5],
                          windowRamAddressRead[4],windowRamAddressRead[3],
                          windowRamAddressRead[2],windowRamAddressRead[1],
                          windowRamAddressRead[0]}), .MFC (MFCWindowRam), .inputSize (
                          {inputSize[12],inputSize[11],inputSize[10],
                          inputSize[9],inputSize[8],inputSize[7],inputSize[6],
                          inputSize[5],inputSize[4],inputSize[3],inputSize[2],
                          inputSize[1],inputSize[0]}), .filterSize ({resetLogics
                          ,resetLogics,resetLogics,resetLogics,resetLogics,
                          resetLogics,resetLogics,resetLogics,resetLogics,
                          resetLogics,weightsSizeType,
                          NOT_weightsSizeType_dup_606,weightsSizeForWindow_0}), 
                          .isFilter (resetLogics), .loadNextWordList (
                          loadNextWindow), .loadWord (loadNextRow), .finishSlice (
                          sliceFinished), .readOne (windowReadOne), .readFinal (
                          windowReadFinal), .aluNumber ({windowAluNumber[2],
                          windowAluNumber[1],windowAluNumber[0]})) ;
    ReadLogic_12_40_true filterReadLogicEnt (.clk (clk), .resetState (
                         resetLogics), .switchRam (reset), .ramBasedAddress ({
                         filterRamBaseAddress[11],filterRamBaseAddress[10],
                         filterRamBaseAddress[9],filterRamBaseAddress[8],
                         filterRamBaseAddress[7],filterRamBaseAddress[6],
                         filterRamBaseAddress[5],filterRamBaseAddress[4],
                         filterRamBaseAddress[3],filterRamBaseAddress[2],
                         filterRamBaseAddress[1],filterRamBaseAddress[0]}), .internalBus (
                         {weightsInternalBus[39],weightsInternalBus[38],
                         weightsInternalBus[37],weightsInternalBus[36],
                         weightsInternalBus[35],weightsInternalBus[34],
                         weightsInternalBus[33],weightsInternalBus[32],
                         weightsInternalBus[31],weightsInternalBus[30],
                         weightsInternalBus[29],weightsInternalBus[28],
                         weightsInternalBus[27],weightsInternalBus[26],
                         weightsInternalBus[25],weightsInternalBus[24],
                         weightsInternalBus[23],weightsInternalBus[22],
                         weightsInternalBus[21],weightsInternalBus[20],
                         weightsInternalBus[19],weightsInternalBus[18],
                         weightsInternalBus[17],weightsInternalBus[16],
                         weightsInternalBus[15],weightsInternalBus[14],
                         weightsInternalBus[13],weightsInternalBus[12],
                         weightsInternalBus[11],weightsInternalBus[10],
                         weightsInternalBus[9],weightsInternalBus[8],
                         weightsInternalBus[7],weightsInternalBus[6],
                         weightsInternalBus[5],weightsInternalBus[4],
                         weightsInternalBus[3],weightsInternalBus[2],
                         weightsInternalBus[1],weightsInternalBus[0]}), .ramDataInBus (
                         {weightsRamDataInBus[39],weightsRamDataInBus[38],
                         weightsRamDataInBus[37],weightsRamDataInBus[36],
                         weightsRamDataInBus[35],weightsRamDataInBus[34],
                         weightsRamDataInBus[33],weightsRamDataInBus[32],
                         weightsRamDataInBus[31],weightsRamDataInBus[30],
                         weightsRamDataInBus[29],weightsRamDataInBus[28],
                         weightsRamDataInBus[27],weightsRamDataInBus[26],
                         weightsRamDataInBus[25],weightsRamDataInBus[24],
                         weightsRamDataInBus[23],weightsRamDataInBus[22],
                         weightsRamDataInBus[21],weightsRamDataInBus[20],
                         weightsRamDataInBus[19],weightsRamDataInBus[18],
                         weightsRamDataInBus[17],weightsRamDataInBus[16],
                         weightsRamDataInBus[15],weightsRamDataInBus[14],
                         weightsRamDataInBus[13],weightsRamDataInBus[12],
                         weightsRamDataInBus[11],weightsRamDataInBus[10],
                         weightsRamDataInBus[9],weightsRamDataInBus[8],
                         weightsRamDataInBus[7],weightsRamDataInBus[6],
                         weightsRamDataInBus[5],weightsRamDataInBus[4],
                         weightsRamDataInBus[3],weightsRamDataInBus[2],
                         weightsRamDataInBus[1],weightsRamDataInBus[0]}), .ramRead (
                         weightsRamRead), .ramAddress ({weightsRamAddress[11],
                         weightsRamAddress[10],weightsRamAddress[9],
                         weightsRamAddress[8],weightsRamAddress[7],
                         weightsRamAddress[6],weightsRamAddress[5],
                         weightsRamAddress[4],weightsRamAddress[3],
                         weightsRamAddress[2],weightsRamAddress[1],
                         weightsRamAddress[0]}), .MFC (MFCWeightsRam), .inputSize (
                         {resetLogics,resetLogics,resetLogics,resetLogics,
                         resetLogics,resetLogics,resetLogics,resetLogics,
                         resetLogics,filterStep_2,filterStep_1,
                         weightsSizeForWindow_0}), .filterSize ({resetLogics,
                         resetLogics,resetLogics,resetLogics,resetLogics,
                         resetLogics,resetLogics,resetLogics,resetLogics,
                         weightsSizeType,NOT_weightsSizeType_dup_606,
                         weightsSizeForWindow_0}), .isFilter (
                         weightsSizeForWindow_0), .loadNextWordList (
                         loadNextFilter), .loadWord (loadWord), .finishSlice (
                         resetLogics), .readOne (weightsReadOne), .readFinal (
                         weightsReadFinal), .aluNumber ({filterAluNumber[2],
                         filterAluNumber[1],filterAluNumber[0]})) ;
    WriteLogic_13_16 writeLogicEnt (.clk (clk), .resetState (resetLogics), .switchRam (
                     switchRam), .ramBasedAddress ({
                     currentWriteRamBaseAddress_12,currentWriteRamBaseAddress_11
                     ,currentWriteRamBaseAddress_10,currentWriteRamBaseAddress_9
                     ,currentWriteRamBaseAddress_8,currentWriteRamBaseAddress_7,
                     currentWriteRamBaseAddress_6,currentWriteRamBaseAddress_5,
                     currentWriteRamBaseAddress_4,currentWriteRamBaseAddress_3,
                     currentWriteRamBaseAddress_2,currentWriteRamBaseAddress_1,
                     currentWriteRamBaseAddress_0}), .internalBus ({
                     windowRamDataOutBus[15],windowRamDataOutBus[14],
                     windowRamDataOutBus[13],windowRamDataOutBus[12],
                     windowRamDataOutBus[11],windowRamDataOutBus[10],
                     windowRamDataOutBus[9],windowRamDataOutBus[8],
                     windowRamDataOutBus[7],windowRamDataOutBus[6],
                     windowRamDataOutBus[5],windowRamDataOutBus[4],
                     windowRamDataOutBus[3],windowRamDataOutBus[2],
                     windowRamDataOutBus[1],windowRamDataOutBus[0]}), .ramWrite (
                     windowRamWrite), .ramDataOutBus ({\$dummy [0],\$dummy [1],
                     \$dummy [2],\$dummy [3],\$dummy [4],\$dummy [5],\$dummy [6]
                     ,\$dummy [7],\$dummy [8],\$dummy [9],\$dummy [10],
                     \$dummy [11],\$dummy [12],\$dummy [13],\$dummy [14],
                     \$dummy [15]}), .ramAddress ({windowRamAddressWrite[12],
                     windowRamAddressWrite[11],windowRamAddressWrite[10],
                     windowRamAddressWrite[9],windowRamAddressWrite[8],
                     windowRamAddressWrite[7],windowRamAddressWrite[6],
                     windowRamAddressWrite[5],windowRamAddressWrite[4],
                     windowRamAddressWrite[3],windowRamAddressWrite[2],
                     windowRamAddressWrite[1],windowRamAddressWrite[0]}), .MFC (
                     MFCWrite), .outputSize ({outputSize[12],outputSize[11],
                     outputSize[10],outputSize[9],outputSize[8],outputSize[7],
                     outputSize[6],outputSize[5],outputSize[4],outputSize[3],
                     outputSize[2],outputSize[1],outputSize[0]}), .write (write)
                     , .finishFilter (writeFinishFilter), .writeDone (
                     writeDoneAll), .writeDoneOne (writeDoneOne)) ;
    inv01 ix608 (.Y (NOT_weightsSizeType_dup_606), .A (weightsSizeType)) ;
    fake_vcc ix596 (.Y (weightsSizeForWindow_0)) ;
    fake_gnd ix594 (.Y (resetLogics)) ;
    or02 ix9 (.Y (loadWord), .A0 (loadOneWord), .A1 (loadThreeWord)) ;
    ao21 ix29 (.Y (writeFinishFilter), .A0 (sliceFinished), .A1 (layerType), .B0 (
         filterFinished)) ;
    aoi21 ix7 (.Y (filterStep_1), .A0 (weightsSizeType), .A1 (nx614), .B0 (
          loadOneWord)) ;
    inv01 ix615 (.Y (nx614), .A (loadThreeWord)) ;
    nor02ii ix13 (.Y (filterStep_2), .A0 (loadWord), .A1 (weightsSizeType)) ;
    or02 ix23 (.Y (windowRLSwitchRam), .A0 (switchRam), .A1 (filterFinished)) ;
    or02 ix21 (.Y (switchRam), .A0 (reset), .A1 (layerFinished)) ;
    dffr reg_ramBaseAddressSelector (.Q (ramBaseAddressSelector), .QB (NOT__4681
         ), .D (NOT__4681), .CLK (layerFinished), .R (reset)) ;
endmodule


module WriteLogic_13_16 ( clk, resetState, switchRam, ramBasedAddress, 
                          internalBus, ramWrite, ramDataOutBus, ramAddress, MFC, 
                          outputSize, write, finishFilter, writeDone, 
                          writeDoneOne ) ;

    input clk ;
    input resetState ;
    input switchRam ;
    input [12:0]ramBasedAddress ;
    input [15:0]internalBus ;
    output ramWrite ;
    output [15:0]ramDataOutBus ;
    output [12:0]ramAddress ;
    input MFC ;
    input [12:0]outputSize ;
    input write ;
    input finishFilter ;
    output writeDone ;
    output writeDoneOne ;

    wire currentState_2, addressRegOut_12, addressRegOut_11, addressRegOut_10, 
         addressRegOut_9, addressRegOut_8, addressRegOut_7, addressRegOut_6, 
         addressRegOut_5, addressRegOut_4, addressRegOut_3, addressRegOut_2, 
         addressRegOut_1, addressRegOut_0, addressRegInFinal_12, 
         addressRegInFinal_11, addressRegInFinal_10, addressRegInFinal_9, 
         addressRegInFinal_8, addressRegInFinal_7, addressRegInFinal_6, 
         addressRegInFinal_5, addressRegInFinal_4, addressRegInFinal_3, 
         addressRegInFinal_2, addressRegInFinal_1, addressRegInFinal_0, 
         resetAddressReg, baseAddressCounterClk, ramAddressKeeperOut_12, 
         ramAddressKeeperOut_11, ramAddressKeeperOut_10, ramAddressKeeperOut_9, 
         ramAddressKeeperOut_8, ramAddressKeeperOut_7, ramAddressKeeperOut_6, 
         ramAddressKeeperOut_5, ramAddressKeeperOut_4, ramAddressKeeperOut_3, 
         ramAddressKeeperOut_2, ramAddressKeeperOut_1, ramAddressKeeperOut_0, 
         ramAddressKeeperOutPlus1_12, ramAddressKeeperOutPlus1_11, 
         ramAddressKeeperOutPlus1_10, ramAddressKeeperOutPlus1_9, 
         ramAddressKeeperOutPlus1_8, ramAddressKeeperOutPlus1_7, 
         ramAddressKeeperOutPlus1_6, ramAddressKeeperOutPlus1_5, 
         ramAddressKeeperOutPlus1_4, ramAddressKeeperOutPlus1_3, 
         ramAddressKeeperOutPlus1_2, ramAddressKeeperOutPlus1_1, 
         ramAddressKeeperOutPlus1_0, addressRegIn_12, addressRegIn_11, 
         addressRegIn_10, addressRegIn_9, addressRegIn_8, addressRegIn_7, 
         addressRegIn_6, addressRegIn_5, addressRegIn_4, addressRegIn_3, 
         addressRegIn_2, addressRegIn_1, addressRegIn_0, dmaCountIn_4, 
         dmaCountIn_3, dmaCountIn_2, dmaCountIn_1, dmaCountIn_0, nextState_1, 
         PWR, currentState_4, currentState_0, nx391, NOT_clk, nx10, 
         currentState_3, nx34, nx42, nx50, nx398, nx408, nx418, nx428, nx438, 
         nx458, nx463, nx467, nx469, nx471, nx473, nx501, nx503, nx513, nx515, 
         nx517, nx519, nx521;
    wire [20:0] \$dummy ;




    assign ramDataOutBus[15] = internalBus[15] ;
    assign ramDataOutBus[14] = internalBus[14] ;
    assign ramDataOutBus[13] = internalBus[13] ;
    assign ramDataOutBus[12] = internalBus[12] ;
    assign ramDataOutBus[11] = internalBus[11] ;
    assign ramDataOutBus[10] = internalBus[10] ;
    assign ramDataOutBus[9] = internalBus[9] ;
    assign ramDataOutBus[8] = internalBus[8] ;
    assign ramDataOutBus[7] = internalBus[7] ;
    assign ramDataOutBus[6] = internalBus[6] ;
    assign ramDataOutBus[5] = internalBus[5] ;
    assign ramDataOutBus[4] = internalBus[4] ;
    assign ramDataOutBus[3] = internalBus[3] ;
    assign ramDataOutBus[2] = internalBus[2] ;
    assign ramDataOutBus[1] = internalBus[1] ;
    assign ramDataOutBus[0] = internalBus[0] ;
    Reg_13 ramAddressKeeper (.D ({ramAddress[12],ramAddress[11],ramAddress[10],
           ramAddress[9],ramAddress[8],ramAddress[7],ramAddress[6],ramAddress[5]
           ,ramAddress[4],ramAddress[3],ramAddress[2],ramAddress[1],
           ramAddress[0]}), .en (ramWrite), .clk (clk), .rst (nextState_1), .Q (
           {ramAddressKeeperOut_12,ramAddressKeeperOut_11,ramAddressKeeperOut_10
           ,ramAddressKeeperOut_9,ramAddressKeeperOut_8,ramAddressKeeperOut_7,
           ramAddressKeeperOut_6,ramAddressKeeperOut_5,ramAddressKeeperOut_4,
           ramAddressKeeperOut_3,ramAddressKeeperOut_2,ramAddressKeeperOut_1,
           ramAddressKeeperOut_0})) ;
    WriteDMA_13_16 dma (.clk (clk), .writeBaseAddress ({addressRegOut_12,
                   addressRegOut_11,addressRegOut_10,addressRegOut_9,
                   addressRegOut_8,addressRegOut_7,addressRegOut_6,
                   addressRegOut_5,addressRegOut_4,addressRegOut_3,
                   addressRegOut_2,addressRegOut_1,addressRegOut_0}), .writeStep (
                   {outputSize[12],outputSize[11],outputSize[10],outputSize[9],
                   outputSize[8],outputSize[7],outputSize[6],outputSize[5],
                   outputSize[4],outputSize[3],outputSize[2],outputSize[1],
                   outputSize[0]}), .writeToRam (ramWrite), .counter ({
                   dmaCountIn_4,dmaCountIn_3,dmaCountIn_2,dmaCountIn_1,
                   dmaCountIn_0}), .initCounter (nx501), .initAddress (nx501), .internalBus (
                   {internalBus[15],internalBus[14],internalBus[13],
                   internalBus[12],internalBus[11],internalBus[10],
                   internalBus[9],internalBus[8],internalBus[7],internalBus[6],
                   internalBus[5],internalBus[4],internalBus[3],internalBus[2],
                   internalBus[1],internalBus[0]}), .ramWrite (\$dummy [0]), .ramDataOutBus (
                   {\$dummy [1],\$dummy [2],\$dummy [3],\$dummy [4],\$dummy [5],
                   \$dummy [6],\$dummy [7],\$dummy [8],\$dummy [9],\$dummy [10],
                   \$dummy [11],\$dummy [12],\$dummy [13],\$dummy [14],
                   \$dummy [15],\$dummy [16]}), .ramWriteAddress ({
                   ramAddress[12],ramAddress[11],ramAddress[10],ramAddress[9],
                   ramAddress[8],ramAddress[7],ramAddress[6],ramAddress[5],
                   ramAddress[4],ramAddress[3],ramAddress[2],ramAddress[1],
                   ramAddress[0]}), .MFC (MFC), .writeComplete (writeDone), .writeCompleteOneOut (
                   writeDoneOne)) ;
    NBitAdder_13 ramAddressIncrement (.a ({ramAddressKeeperOut_12,
                 ramAddressKeeperOut_11,ramAddressKeeperOut_10,
                 ramAddressKeeperOut_9,ramAddressKeeperOut_8,
                 ramAddressKeeperOut_7,ramAddressKeeperOut_6,
                 ramAddressKeeperOut_5,ramAddressKeeperOut_4,
                 ramAddressKeeperOut_3,ramAddressKeeperOut_2,
                 ramAddressKeeperOut_1,ramAddressKeeperOut_0}), .b ({nextState_1
                 ,nextState_1,nextState_1,nextState_1,nextState_1,nextState_1,
                 nextState_1,nextState_1,nextState_1,nextState_1,nextState_1,
                 nextState_1,nextState_1}), .carryIn (PWR), .sum ({
                 ramAddressKeeperOutPlus1_12,ramAddressKeeperOutPlus1_11,
                 ramAddressKeeperOutPlus1_10,ramAddressKeeperOutPlus1_9,
                 ramAddressKeeperOutPlus1_8,ramAddressKeeperOutPlus1_7,
                 ramAddressKeeperOutPlus1_6,ramAddressKeeperOutPlus1_5,
                 ramAddressKeeperOutPlus1_4,ramAddressKeeperOutPlus1_3,
                 ramAddressKeeperOutPlus1_2,ramAddressKeeperOutPlus1_1,
                 ramAddressKeeperOutPlus1_0}), .carryOut (\$dummy [17])) ;
    Mux2_13 baseAddressLoadMux (.A ({addressRegIn_12,addressRegIn_11,
            addressRegIn_10,addressRegIn_9,addressRegIn_8,addressRegIn_7,
            addressRegIn_6,addressRegIn_5,addressRegIn_4,addressRegIn_3,
            addressRegIn_2,addressRegIn_1,addressRegIn_0}), .B ({
            ramAddressKeeperOutPlus1_12,ramAddressKeeperOutPlus1_11,
            ramAddressKeeperOutPlus1_10,ramAddressKeeperOutPlus1_9,
            ramAddressKeeperOutPlus1_8,ramAddressKeeperOutPlus1_7,
            ramAddressKeeperOutPlus1_6,ramAddressKeeperOutPlus1_5,
            ramAddressKeeperOutPlus1_4,ramAddressKeeperOutPlus1_3,
            ramAddressKeeperOutPlus1_2,ramAddressKeeperOutPlus1_1,
            ramAddressKeeperOutPlus1_0}), .S (finishFilter), .C ({
            addressRegInFinal_12,addressRegInFinal_11,addressRegInFinal_10,
            addressRegInFinal_9,addressRegInFinal_8,addressRegInFinal_7,
            addressRegInFinal_6,addressRegInFinal_5,addressRegInFinal_4,
            addressRegInFinal_3,addressRegInFinal_2,addressRegInFinal_1,
            addressRegInFinal_0})) ;
    Counter2_13 baseAddressCounter (.load ({addressRegInFinal_12,
                addressRegInFinal_11,addressRegInFinal_10,addressRegInFinal_9,
                addressRegInFinal_8,addressRegInFinal_7,addressRegInFinal_6,
                addressRegInFinal_5,addressRegInFinal_4,addressRegInFinal_3,
                addressRegInFinal_2,addressRegInFinal_1,addressRegInFinal_0}), .reset (
                nextState_1), .clk (baseAddressCounterClk), .isLoad (
                resetAddressReg), .count ({addressRegOut_12,addressRegOut_11,
                addressRegOut_10,addressRegOut_9,addressRegOut_8,addressRegOut_7
                ,addressRegOut_6,addressRegOut_5,addressRegOut_4,addressRegOut_3
                ,addressRegOut_2,addressRegOut_1,addressRegOut_0})) ;
    fake_vcc ix365 (.Y (PWR)) ;
    fake_gnd ix363 (.Y (nextState_1)) ;
    mux21_ni ix439 (.Y (nx438), .A0 (currentState_4), .A1 (nx50), .S0 (nx391)) ;
    mux21_ni ix429 (.Y (nx428), .A0 (currentState_3), .A1 (nx42), .S0 (nx391)) ;
    dffr reg_currentState_3 (.Q (currentState_3), .QB (\$dummy [18]), .D (nx428)
         , .CLK (NOT_clk), .R (resetState)) ;
    inv01 ix453 (.Y (NOT_clk), .A (clk)) ;
    nor02ii ix43 (.Y (nx42), .A0 (switchRam), .A1 (nx503)) ;
    dffr reg_currentState_2 (.Q (currentState_2), .QB (\$dummy [19]), .D (nx418)
         , .CLK (NOT_clk), .R (resetState)) ;
    mux21_ni ix419 (.Y (nx418), .A0 (nx501), .A1 (nx34), .S0 (nx391)) ;
    mux21_ni ix409 (.Y (nx408), .A0 (currentState_0), .A1 (nx10), .S0 (nx391)) ;
    dffs_ni reg_currentState_0 (.Q (currentState_0), .QB (nx458), .D (nx408), .CLK (
            NOT_clk), .S (resetState)) ;
    aoi21 ix11 (.Y (nx10), .A0 (nx517), .A1 (nx471), .B0 (switchRam)) ;
    dffr reg_currentState_1 (.Q (\$dummy [20]), .QB (nx463), .D (nx398), .CLK (
         NOT_clk), .R (resetState)) ;
    oai21 ix399 (.Y (nx398), .A0 (nx517), .A1 (nx391), .B0 (nx473)) ;
    nand02 ix31 (.Y (nx391), .A0 (nx467), .A1 (nx469)) ;
    aoi21 ix468 (.Y (nx467), .A0 (writeDone), .A1 (currentState_4), .B0 (
          switchRam)) ;
    dffr reg_currentState_4 (.Q (currentState_4), .QB (nx471), .D (nx438), .CLK (
         NOT_clk), .R (resetState)) ;
    inv01 ix474 (.Y (nx473), .A (switchRam)) ;
    and02 ix59 (.Y (dmaCountIn_0), .A0 (outputSize[0]), .A1 (nx503)) ;
    and02 ix61 (.Y (dmaCountIn_1), .A0 (outputSize[1]), .A1 (nx503)) ;
    and02 ix63 (.Y (dmaCountIn_2), .A0 (outputSize[2]), .A1 (nx503)) ;
    and02 ix65 (.Y (dmaCountIn_3), .A0 (outputSize[3]), .A1 (nx503)) ;
    and02 ix67 (.Y (dmaCountIn_4), .A0 (outputSize[4]), .A1 (nx503)) ;
    mux21_ni ix103 (.Y (baseAddressCounterClk), .A0 (resetAddressReg), .A1 (
             currentState_3), .S0 (clk)) ;
    buf02 ix500 (.Y (nx501), .A (currentState_2)) ;
    buf02 ix502 (.Y (nx503), .A (currentState_2)) ;
    nor02ii ix57 (.Y (ramWrite), .A0 (nx471), .A1 (write)) ;
    nor02ii ix51 (.Y (nx50), .A0 (switchRam), .A1 (currentState_3)) ;
    nor02ii ix35 (.Y (nx34), .A0 (switchRam), .A1 (currentState_0)) ;
    mux21 ix470 (.Y (nx469), .A0 (write), .A1 (nx471), .S0 (nx458)) ;
    nor02ii ix69 (.Y (addressRegIn_0), .A0 (nx517), .A1 (ramBasedAddress[0])) ;
    nor02ii ix71 (.Y (addressRegIn_1), .A0 (nx517), .A1 (ramBasedAddress[1])) ;
    nor02ii ix73 (.Y (addressRegIn_2), .A0 (nx517), .A1 (ramBasedAddress[2])) ;
    nor02ii ix75 (.Y (addressRegIn_3), .A0 (nx517), .A1 (ramBasedAddress[3])) ;
    nor02ii ix77 (.Y (addressRegIn_4), .A0 (nx517), .A1 (ramBasedAddress[4])) ;
    nor02ii ix79 (.Y (addressRegIn_5), .A0 (nx519), .A1 (ramBasedAddress[5])) ;
    nor02ii ix81 (.Y (addressRegIn_6), .A0 (nx519), .A1 (ramBasedAddress[6])) ;
    nor02ii ix83 (.Y (addressRegIn_7), .A0 (nx519), .A1 (ramBasedAddress[7])) ;
    nor02ii ix85 (.Y (addressRegIn_8), .A0 (nx519), .A1 (ramBasedAddress[8])) ;
    nor02ii ix87 (.Y (addressRegIn_9), .A0 (nx519), .A1 (ramBasedAddress[9])) ;
    nor02ii ix89 (.Y (addressRegIn_10), .A0 (nx519), .A1 (ramBasedAddress[10])
            ) ;
    nor02ii ix91 (.Y (addressRegIn_11), .A0 (nx519), .A1 (ramBasedAddress[11])
            ) ;
    nor02ii ix93 (.Y (addressRegIn_12), .A0 (nx521), .A1 (ramBasedAddress[12])
            ) ;
    nand02 ix95 (.Y (resetAddressReg), .A0 (nx521), .A1 (nx513)) ;
    inv01 ix512 (.Y (nx513), .A (finishFilter)) ;
    inv01 ix514 (.Y (nx515), .A (nx463)) ;
    inv01 ix516 (.Y (nx517), .A (nx515)) ;
    inv01 ix518 (.Y (nx519), .A (nx515)) ;
    inv01 ix520 (.Y (nx521), .A (nx515)) ;
endmodule


module WriteDMA_13_16 ( clk, writeBaseAddress, writeStep, writeToRam, counter, 
                        initCounter, initAddress, internalBus, ramWrite, 
                        ramDataOutBus, ramWriteAddress, MFC, writeComplete, 
                        writeCompleteOneOut ) ;

    input clk ;
    input [12:0]writeBaseAddress ;
    input [12:0]writeStep ;
    input writeToRam ;
    input [4:0]counter ;
    input initCounter ;
    input initAddress ;
    input [15:0]internalBus ;
    output ramWrite ;
    output [15:0]ramDataOutBus ;
    output [12:0]ramWriteAddress ;
    input MFC ;
    output writeComplete ;
    output writeCompleteOneOut ;

    wire toBeAdded_12, toBeAdded_11, toBeAdded_10, toBeAdded_9, toBeAdded_8, 
         toBeAdded_7, toBeAdded_6, toBeAdded_5, toBeAdded_4, toBeAdded_3, 
         toBeAdded_2, toBeAdded_1, toBeAdded_0, currentCount_4, currentCount_3, 
         currentCount_2, currentCount_1, currentCount_0, enableCounter, GND, PWR, 
         NOT_MFC, nx26, nx101, nx103, nx105, nx1, nx5;



    assign ramWrite = writeToRam ;
    assign ramDataOutBus[15] = internalBus[15] ;
    assign ramDataOutBus[14] = internalBus[14] ;
    assign ramDataOutBus[13] = internalBus[13] ;
    assign ramDataOutBus[12] = internalBus[12] ;
    assign ramDataOutBus[11] = internalBus[11] ;
    assign ramDataOutBus[10] = internalBus[10] ;
    assign ramDataOutBus[9] = internalBus[9] ;
    assign ramDataOutBus[8] = internalBus[8] ;
    assign ramDataOutBus[7] = internalBus[7] ;
    assign ramDataOutBus[6] = internalBus[6] ;
    assign ramDataOutBus[5] = internalBus[5] ;
    assign ramDataOutBus[4] = internalBus[4] ;
    assign ramDataOutBus[3] = internalBus[3] ;
    assign ramDataOutBus[2] = internalBus[2] ;
    assign ramDataOutBus[1] = internalBus[1] ;
    assign ramDataOutBus[0] = internalBus[0] ;
    Reg_13 writeStepRegister (.D ({writeStep[12],writeStep[11],writeStep[10],
           writeStep[9],writeStep[8],writeStep[7],writeStep[6],writeStep[5],
           writeStep[4],writeStep[3],writeStep[2],writeStep[1],writeStep[0]}), .en (
           PWR), .clk (initCounter), .rst (GND), .Q ({toBeAdded_12,toBeAdded_11,
           toBeAdded_10,toBeAdded_9,toBeAdded_8,toBeAdded_7,toBeAdded_6,
           toBeAdded_5,toBeAdded_4,toBeAdded_3,toBeAdded_2,toBeAdded_1,
           toBeAdded_0})) ;
    MultiStepCounter_13 writeAddressRegister (.load ({writeBaseAddress[12],
                        writeBaseAddress[11],writeBaseAddress[10],
                        writeBaseAddress[9],writeBaseAddress[8],
                        writeBaseAddress[7],writeBaseAddress[6],
                        writeBaseAddress[5],writeBaseAddress[4],
                        writeBaseAddress[3],writeBaseAddress[2],
                        writeBaseAddress[1],writeBaseAddress[0]}), .toBeAdded ({
                        toBeAdded_12,toBeAdded_11,toBeAdded_10,toBeAdded_9,
                        toBeAdded_8,toBeAdded_7,toBeAdded_6,toBeAdded_5,
                        toBeAdded_4,toBeAdded_3,toBeAdded_2,toBeAdded_1,
                        toBeAdded_0}), .reset (GND), .clk (clk), .isLoad (
                        initAddress), .MFC (writeCompleteOneOut), .count ({
                        ramWriteAddress[12],ramWriteAddress[11],
                        ramWriteAddress[10],ramWriteAddress[9],
                        ramWriteAddress[8],ramWriteAddress[7],ramWriteAddress[6]
                        ,ramWriteAddress[5],ramWriteAddress[4],
                        ramWriteAddress[3],ramWriteAddress[2],ramWriteAddress[1]
                        ,ramWriteAddress[0]})) ;
    DownCounter_5 writecounter (.load ({counter[4],counter[3],counter[2],
                  counter[1],counter[0]}), .enable (enableCounter), .clk (clk), 
                  .isLoad (initCounter), .currentCount ({currentCount_4,
                  currentCount_3,currentCount_2,currentCount_1,currentCount_0})
                  ) ;
    fake_vcc ix82 (.Y (PWR)) ;
    fake_gnd ix80 (.Y (GND)) ;
    or02 ix33 (.Y (enableCounter), .A0 (writeCompleteOneOut), .A1 (initCounter)
         ) ;
    inv16 ix99 (.Y (NOT_MFC), .A (MFC)) ;
    nor04 ix27 (.Y (nx26), .A0 (nx101), .A1 (nx105), .A2 (currentCount_1), .A3 (
          clk)) ;
    or04 ix102 (.Y (nx101), .A0 (nx103), .A1 (currentCount_4), .A2 (
         currentCount_3), .A3 (currentCount_2)) ;
    inv01 ix104 (.Y (nx103), .A (currentCount_0)) ;
    nand02 ix106 (.Y (nx105), .A0 (writeToRam), .A1 (MFC)) ;
    inv01 ix17 (.Y (writeCompleteOneOut), .A (nx105)) ;
    latchs_ni lat_internalWriteComplete_u1 (.QB (nx5), .D (GND), .CLK (NOT_MFC)
              , .S (nx26)) ;
    inv02 lat_internalWriteComplete_u2 (.Y (writeComplete), .A (nx5)) ;
    buf02 lat_internalWriteComplete_u3 (.Y (nx1), .A (nx5)) ;
endmodule


module DownCounter_5 ( load, enable, clk, isLoad, currentCount ) ;

    input [4:0]load ;
    input enable ;
    input clk ;
    input isLoad ;
    inout [4:0]currentCount ;

    wire counterInput_4, counterInput_3, counterInput_2, counterInput_1, 
         counterInput_0, subtractorOutput_4, subtractorOutput_3, 
         subtractorOutput_2, subtractorOutput_1, subtractorOutput_0, PWR, 
         zerosSignal_4;
    wire [0:0] \$dummy ;




    Reg_5 counterReg (.D ({counterInput_4,counterInput_3,counterInput_2,
          counterInput_1,counterInput_0}), .en (enable), .clk (clk), .rst (
          zerosSignal_4), .Q ({currentCount[4],currentCount[3],currentCount[2],
          currentCount[1],currentCount[0]})) ;
    NBitSubtractor_5 nextCount (.x ({currentCount[4],currentCount[3],
                     currentCount[2],currentCount[1],currentCount[0]}), .y ({
                     zerosSignal_4,zerosSignal_4,zerosSignal_4,zerosSignal_4,
                     zerosSignal_4}), .bin (PWR), .difference ({
                     subtractorOutput_4,subtractorOutput_3,subtractorOutput_2,
                     subtractorOutput_1,subtractorOutput_0}), .borrowOut (
                     \$dummy [0])) ;
    Mux2_5 muxloadOrCurrent (.A ({subtractorOutput_4,subtractorOutput_3,
           subtractorOutput_2,subtractorOutput_1,subtractorOutput_0}), .B ({
           load[4],load[3],load[2],load[1],load[0]}), .S (isLoad), .C ({
           counterInput_4,counterInput_3,counterInput_2,counterInput_1,
           counterInput_0})) ;
    fake_gnd ix24 (.Y (zerosSignal_4)) ;
    fake_vcc ix22 (.Y (PWR)) ;
endmodule


module Mux2_5 ( A, B, S, C ) ;

    input [4:0]A ;
    input [4:0]B ;
    input S ;
    output [4:0]C ;

    wire nx96;



    mux21_ni ix7 (.Y (C[0]), .A0 (A[0]), .A1 (B[0]), .S0 (nx96)) ;
    mux21_ni ix15 (.Y (C[1]), .A0 (A[1]), .A1 (B[1]), .S0 (nx96)) ;
    mux21_ni ix23 (.Y (C[2]), .A0 (A[2]), .A1 (B[2]), .S0 (nx96)) ;
    mux21_ni ix31 (.Y (C[3]), .A0 (A[3]), .A1 (B[3]), .S0 (nx96)) ;
    mux21_ni ix39 (.Y (C[4]), .A0 (A[4]), .A1 (B[4]), .S0 (nx96)) ;
    buf02 ix95 (.Y (nx96), .A (S)) ;
endmodule


module NBitSubtractor_5 ( x, y, bin, difference, borrowOut ) ;

    input [4:0]x ;
    input [4:0]y ;
    input bin ;
    output [4:0]difference ;
    output borrowOut ;

    wire temp_3, temp_2, temp_1, temp_0;



    FullSubtractor f0 (.x (x[0]), .y (y[0]), .bin (bin), .difference (
                   difference[0]), .bout (temp_0)) ;
    FullSubtractor loop1_1_fx (.x (x[1]), .y (y[1]), .bin (temp_0), .difference (
                   difference[1]), .bout (temp_1)) ;
    FullSubtractor loop1_2_fx (.x (x[2]), .y (y[2]), .bin (temp_1), .difference (
                   difference[2]), .bout (temp_2)) ;
    FullSubtractor loop1_3_fx (.x (x[3]), .y (y[3]), .bin (temp_2), .difference (
                   difference[3]), .bout (temp_3)) ;
    FullSubtractor loop1_4_fx (.x (x[4]), .y (y[4]), .bin (temp_3), .difference (
                   difference[4]), .bout (borrowOut)) ;
endmodule


module ReadLogic_12_40_true ( clk, resetState, switchRam, ramBasedAddress, 
                              internalBus, ramDataInBus, ramRead, ramAddress, 
                              MFC, inputSize, filterSize, isFilter, 
                              loadNextWordList, loadWord, finishSlice, readOne, 
                              readFinal, aluNumber ) ;

    input clk ;
    input resetState ;
    input switchRam ;
    input [11:0]ramBasedAddress ;
    output [39:0]internalBus ;
    input [39:0]ramDataInBus ;
    output ramRead ;
    output [11:0]ramAddress ;
    input MFC ;
    input [11:0]inputSize ;
    input [11:0]filterSize ;
    input isFilter ;
    input loadNextWordList ;
    input loadWord ;
    input finishSlice ;
    output readOne ;
    output readFinal ;
    output [2:0]aluNumber ;

    wire aluNumberCounterClk, notClk, aluCounterOut_2, aluCounterOut_1, 
         aluCounterOut_0, dmaReadBaseAddress_11, dmaReadBaseAddress_10, 
         dmaReadBaseAddress_9, dmaReadBaseAddress_8, dmaReadBaseAddress_7, 
         dmaReadBaseAddress_6, dmaReadBaseAddress_5, dmaReadBaseAddress_4, 
         dmaReadBaseAddress_3, dmaReadBaseAddress_2, dmaReadBaseAddress_1, 
         dmaReadBaseAddress_0, dmaInitRamBaseAddress, dmaCountIn_2, dmaCountIn_1, 
         dmaCountIn_0, dmaInitCounter, PWR, addressRegOut_11, currentState_0, 
         nx387, nx12, nx16, NOT__4272, nx395, nx405, nx414, nx419, nx424, nx427, 
         nx432, nx434, nx437, nx440, nx444, nx451;
    wire [0:0] \$dummy ;




    Mux2_12 dmaReadBaseAddressMux (.A ({addressRegOut_11,addressRegOut_11,
            addressRegOut_11,addressRegOut_11,addressRegOut_11,addressRegOut_11,
            addressRegOut_11,addressRegOut_11,addressRegOut_11,addressRegOut_11,
            addressRegOut_11,addressRegOut_11}), .B ({ramBasedAddress[11],
            ramBasedAddress[10],ramBasedAddress[9],ramBasedAddress[8],
            ramBasedAddress[7],ramBasedAddress[6],ramBasedAddress[5],
            ramBasedAddress[4],ramBasedAddress[3],ramBasedAddress[2],
            ramBasedAddress[1],ramBasedAddress[0]}), .S (dmaInitRamBaseAddress)
            , .C ({dmaReadBaseAddress_11,dmaReadBaseAddress_10,
            dmaReadBaseAddress_9,dmaReadBaseAddress_8,dmaReadBaseAddress_7,
            dmaReadBaseAddress_6,dmaReadBaseAddress_5,dmaReadBaseAddress_4,
            dmaReadBaseAddress_3,dmaReadBaseAddress_2,dmaReadBaseAddress_1,
            dmaReadBaseAddress_0})) ;
    DMA_12_40 dma (.initialCount ({dmaCountIn_2,dmaCountIn_1,dmaCountIn_0}), .readBaseAddress (
              {dmaReadBaseAddress_11,dmaReadBaseAddress_10,dmaReadBaseAddress_9,
              dmaReadBaseAddress_8,dmaReadBaseAddress_7,dmaReadBaseAddress_6,
              dmaReadBaseAddress_5,dmaReadBaseAddress_4,dmaReadBaseAddress_3,
              dmaReadBaseAddress_2,dmaReadBaseAddress_1,dmaReadBaseAddress_0}), 
              .readStep ({inputSize[11],inputSize[10],inputSize[9],inputSize[8],
              inputSize[7],inputSize[6],inputSize[5],inputSize[4],inputSize[3],
              inputSize[2],inputSize[1],inputSize[0]}), .initAddress (
              dmaInitRamBaseAddress), .initCounter (nx451), .load (ramRead), .internalBus (
              {internalBus[39],internalBus[38],internalBus[37],internalBus[36],
              internalBus[35],internalBus[34],internalBus[33],internalBus[32],
              internalBus[31],internalBus[30],internalBus[29],internalBus[28],
              internalBus[27],internalBus[26],internalBus[25],internalBus[24],
              internalBus[23],internalBus[22],internalBus[21],internalBus[20],
              internalBus[19],internalBus[18],internalBus[17],internalBus[16],
              internalBus[15],internalBus[14],internalBus[13],internalBus[12],
              internalBus[11],internalBus[10],internalBus[9],internalBus[8],
              internalBus[7],internalBus[6],internalBus[5],internalBus[4],
              internalBus[3],internalBus[2],internalBus[1],internalBus[0]}), .finishedOneReadOut (
              readOne), .finishedReading (readFinal), .clk (clk), .ramDataInBus (
              {ramDataInBus[39],ramDataInBus[38],ramDataInBus[37],
              ramDataInBus[36],ramDataInBus[35],ramDataInBus[34],
              ramDataInBus[33],ramDataInBus[32],ramDataInBus[31],
              ramDataInBus[30],ramDataInBus[29],ramDataInBus[28],
              ramDataInBus[27],ramDataInBus[26],ramDataInBus[25],
              ramDataInBus[24],ramDataInBus[23],ramDataInBus[22],
              ramDataInBus[21],ramDataInBus[20],ramDataInBus[19],
              ramDataInBus[18],ramDataInBus[17],ramDataInBus[16],
              ramDataInBus[15],ramDataInBus[14],ramDataInBus[13],
              ramDataInBus[12],ramDataInBus[11],ramDataInBus[10],ramDataInBus[9]
              ,ramDataInBus[8],ramDataInBus[7],ramDataInBus[6],ramDataInBus[5],
              ramDataInBus[4],ramDataInBus[3],ramDataInBus[2],ramDataInBus[1],
              ramDataInBus[0]}), .ramRead (\$dummy [0]), .ramReadAddress ({
              ramAddress[11],ramAddress[10],ramAddress[9],ramAddress[8],
              ramAddress[7],ramAddress[6],ramAddress[5],ramAddress[4],
              ramAddress[3],ramAddress[2],ramAddress[1],ramAddress[0]}), .MFC (
              MFC)) ;
    Counter2_3 aluNumberCounter (.load ({addressRegOut_11,addressRegOut_11,
               addressRegOut_11}), .reset (NOT__4272), .clk (aluNumberCounterClk
               ), .isLoad (addressRegOut_11), .count ({aluCounterOut_2,
               aluCounterOut_1,aluCounterOut_0})) ;
    Reg_3 regCounterOut (.D ({aluCounterOut_2,aluCounterOut_1,aluCounterOut_0})
          , .en (PWR), .clk (notClk), .rst (addressRegOut_11), .Q ({aluNumber[2]
          ,aluNumber[1],aluNumber[0]})) ;
    oai32 ix406 (.Y (nx405), .A0 (switchRam), .A1 (currentState_0), .A2 (nx427)
          , .B0 (NOT__4272), .B1 (nx387)) ;
    oai21 ix396 (.Y (nx395), .A0 (nx414), .A1 (nx387), .B0 (nx424)) ;
    dffr reg_currentState_0 (.Q (currentState_0), .QB (nx414), .D (nx395), .CLK (
         notClk), .R (resetState)) ;
    inv01 ix417 (.Y (notClk), .A (clk)) ;
    nand02 ix23 (.Y (nx387), .A0 (nx419), .A1 (nx424)) ;
    aoi21 ix420 (.Y (nx419), .A0 (readFinal), .A1 (nx16), .B0 (
          dmaInitRamBaseAddress)) ;
    dffr reg_currentState_1 (.Q (ramRead), .QB (NOT__4272), .D (nx405), .CLK (
         notClk), .R (resetState)) ;
    nor02_2x ix425 (.Y (nx424), .A0 (nx12), .A1 (switchRam)) ;
    nor03_2x ix428 (.Y (nx427), .A0 (loadNextWordList), .A1 (loadWord), .A2 (
             ramRead)) ;
    fake_gnd ix375 (.Y (addressRegOut_11)) ;
    fake_vcc ix373 (.Y (PWR)) ;
    aoi21 ix41 (.Y (dmaInitCounter), .A0 (nx432), .A1 (nx434), .B0 (nx16)) ;
    inv01 ix433 (.Y (nx432), .A (loadNextWordList)) ;
    inv01 ix435 (.Y (nx434), .A (loadWord)) ;
    inv01 ix47 (.Y (dmaCountIn_0), .A (nx437)) ;
    oai21 ix438 (.Y (nx437), .A0 (nx432), .A1 (filterSize[0]), .B0 (nx451)) ;
    and03 ix53 (.Y (dmaCountIn_1), .A0 (nx440), .A1 (filterSize[1]), .A2 (
          loadNextWordList)) ;
    and03 ix59 (.Y (dmaCountIn_2), .A0 (nx440), .A1 (filterSize[2]), .A2 (
          loadNextWordList)) ;
    aoi21 ix67 (.Y (aluNumberCounterClk), .A0 (nx444), .A1 (ramRead), .B0 (
          notClk)) ;
    nand02 ix445 (.Y (nx444), .A0 (loadNextWordList), .A1 (readOne)) ;
    inv01 ix17 (.Y (nx16), .A (nx440)) ;
    buf02 ix450 (.Y (nx451), .A (dmaInitCounter)) ;
    and02 ix35 (.Y (dmaInitRamBaseAddress), .A0 (NOT__4272), .A1 (currentState_0
          )) ;
    nor02ii ix13 (.Y (nx12), .A0 (nx427), .A1 (nx414)) ;
    and02 ix441 (.Y (nx440), .A0 (nx414), .A1 (NOT__4272)) ;
endmodule


module DMA_12_40 ( initialCount, readBaseAddress, readStep, initAddress, 
                   initCounter, load, internalBus, finishedOneReadOut, 
                   finishedReading, clk, ramDataInBus, ramRead, ramReadAddress, 
                   MFC ) ;

    input [2:0]initialCount ;
    input [11:0]readBaseAddress ;
    input [11:0]readStep ;
    input initAddress ;
    input initCounter ;
    input load ;
    output [39:0]internalBus ;
    output finishedOneReadOut ;
    output finishedReading ;
    input clk ;
    input [39:0]ramDataInBus ;
    output ramRead ;
    output [11:0]ramReadAddress ;
    input MFC ;

    wire currentCount_2, currentCount_1, currentCount_0, tobeAdded_11, 
         tobeAdded_10, tobeAdded_9, tobeAdded_8, tobeAdded_7, tobeAdded_6, 
         tobeAdded_5, tobeAdded_4, tobeAdded_3, tobeAdded_2, tobeAdded_1, 
         tobeAdded_0, enableCount, PWR, GND, NOT_MFC, nx18, nx133, nx135, nx137, 
         nx1, nx5;



    assign ramRead = load ;
    MultiStepCounter_12 addressRegister (.load ({readBaseAddress[11],
                        readBaseAddress[10],readBaseAddress[9],
                        readBaseAddress[8],readBaseAddress[7],readBaseAddress[6]
                        ,readBaseAddress[5],readBaseAddress[4],
                        readBaseAddress[3],readBaseAddress[2],readBaseAddress[1]
                        ,readBaseAddress[0]}), .toBeAdded ({tobeAdded_11,
                        tobeAdded_10,tobeAdded_9,tobeAdded_8,tobeAdded_7,
                        tobeAdded_6,tobeAdded_5,tobeAdded_4,tobeAdded_3,
                        tobeAdded_2,tobeAdded_1,tobeAdded_0}), .reset (GND), .clk (
                        clk), .isLoad (initAddress), .MFC (finishedOneReadOut), 
                        .count ({ramReadAddress[11],ramReadAddress[10],
                        ramReadAddress[9],ramReadAddress[8],ramReadAddress[7],
                        ramReadAddress[6],ramReadAddress[5],ramReadAddress[4],
                        ramReadAddress[3],ramReadAddress[2],ramReadAddress[1],
                        ramReadAddress[0]})) ;
    DownCounter_3 counter (.load ({initialCount[2],initialCount[1],
                  initialCount[0]}), .enable (enableCount), .clk (clk), .isLoad (
                  initCounter), .currentCount ({currentCount_2,currentCount_1,
                  currentCount_0})) ;
    Reg_12 readStepRegister (.D ({readStep[11],readStep[10],readStep[9],
           readStep[8],readStep[7],readStep[6],readStep[5],readStep[4],
           readStep[3],readStep[2],readStep[1],readStep[0]}), .en (PWR), .clk (
           clk), .rst (GND), .Q ({tobeAdded_11,tobeAdded_10,tobeAdded_9,
           tobeAdded_8,tobeAdded_7,tobeAdded_6,tobeAdded_5,tobeAdded_4,
           tobeAdded_3,tobeAdded_2,tobeAdded_1,tobeAdded_0})) ;
    Tristate_40 tristateLabel (.\input  ({ramDataInBus[39],ramDataInBus[38],
                ramDataInBus[37],ramDataInBus[36],ramDataInBus[35],
                ramDataInBus[34],ramDataInBus[33],ramDataInBus[32],
                ramDataInBus[31],ramDataInBus[30],ramDataInBus[29],
                ramDataInBus[28],ramDataInBus[27],ramDataInBus[26],
                ramDataInBus[25],ramDataInBus[24],ramDataInBus[23],
                ramDataInBus[22],ramDataInBus[21],ramDataInBus[20],
                ramDataInBus[19],ramDataInBus[18],ramDataInBus[17],
                ramDataInBus[16],ramDataInBus[15],ramDataInBus[14],
                ramDataInBus[13],ramDataInBus[12],ramDataInBus[11],
                ramDataInBus[10],ramDataInBus[9],ramDataInBus[8],ramDataInBus[7]
                ,ramDataInBus[6],ramDataInBus[5],ramDataInBus[4],ramDataInBus[3]
                ,ramDataInBus[2],ramDataInBus[1],ramDataInBus[0]}), .en (
                finishedOneReadOut), .\output  ({internalBus[39],internalBus[38]
                ,internalBus[37],internalBus[36],internalBus[35],internalBus[34]
                ,internalBus[33],internalBus[32],internalBus[31],internalBus[30]
                ,internalBus[29],internalBus[28],internalBus[27],internalBus[26]
                ,internalBus[25],internalBus[24],internalBus[23],internalBus[22]
                ,internalBus[21],internalBus[20],internalBus[19],internalBus[18]
                ,internalBus[17],internalBus[16],internalBus[15],internalBus[14]
                ,internalBus[13],internalBus[12],internalBus[11],internalBus[10]
                ,internalBus[9],internalBus[8],internalBus[7],internalBus[6],
                internalBus[5],internalBus[4],internalBus[3],internalBus[2],
                internalBus[1],internalBus[0]})) ;
    fake_gnd ix116 (.Y (GND)) ;
    fake_vcc ix114 (.Y (PWR)) ;
    and02 ix13 (.Y (finishedOneReadOut), .A0 (load), .A1 (MFC)) ;
    or02 ix25 (.Y (enableCount), .A0 (MFC), .A1 (initCounter)) ;
    inv16 ix131 (.Y (NOT_MFC), .A (MFC)) ;
    nor04 ix19 (.Y (nx18), .A0 (currentCount_1), .A1 (nx133), .A2 (
          currentCount_2), .A3 (nx135)) ;
    inv01 ix134 (.Y (nx133), .A (currentCount_0)) ;
    nand02 ix136 (.Y (nx135), .A0 (nx137), .A1 (finishedOneReadOut)) ;
    inv01 ix138 (.Y (nx137), .A (clk)) ;
    latchs_ni lat_internalFinishedReading_u1 (.QB (nx5), .D (GND), .CLK (NOT_MFC
              ), .S (nx18)) ;
    inv02 lat_internalFinishedReading_u2 (.Y (finishedReading), .A (nx5)) ;
    buf02 lat_internalFinishedReading_u3 (.Y (nx1), .A (nx5)) ;
endmodule


module Tristate_40 ( \input , en, \output  ) ;

    input [39:0]\input  ;
    input en ;
    output [39:0]\output  ;

    wire nx375, nx378, nx381, nx384, nx387, nx390, nx393, nx396, nx399, nx402, 
         nx405, nx408, nx411, nx414, nx417, nx420, nx423, nx426, nx429, nx432, 
         nx435, nx438, nx441, nx444, nx447, nx450, nx453, nx456, nx459, nx462, 
         nx465, nx468, nx471, nx474, nx477, nx480, nx483, nx486, nx489, nx492, 
         nx499, nx501, nx503, nx505, nx507, nx509, nx511;



    tri01 tri_output_0 (.Y (\output [0]), .A (nx375), .E (nx501)) ;
    inv01 ix376 (.Y (nx375), .A (\input [0])) ;
    tri01 tri_output_1 (.Y (\output [1]), .A (nx378), .E (nx501)) ;
    inv01 ix379 (.Y (nx378), .A (\input [1])) ;
    tri01 tri_output_2 (.Y (\output [2]), .A (nx381), .E (nx501)) ;
    inv01 ix382 (.Y (nx381), .A (\input [2])) ;
    tri01 tri_output_3 (.Y (\output [3]), .A (nx384), .E (nx501)) ;
    inv01 ix385 (.Y (nx384), .A (\input [3])) ;
    tri01 tri_output_4 (.Y (\output [4]), .A (nx387), .E (nx501)) ;
    inv01 ix388 (.Y (nx387), .A (\input [4])) ;
    tri01 tri_output_5 (.Y (\output [5]), .A (nx390), .E (nx501)) ;
    inv01 ix391 (.Y (nx390), .A (\input [5])) ;
    tri01 tri_output_6 (.Y (\output [6]), .A (nx393), .E (nx501)) ;
    inv01 ix394 (.Y (nx393), .A (\input [6])) ;
    tri01 tri_output_7 (.Y (\output [7]), .A (nx396), .E (nx503)) ;
    inv01 ix397 (.Y (nx396), .A (\input [7])) ;
    tri01 tri_output_8 (.Y (\output [8]), .A (nx399), .E (nx503)) ;
    inv01 ix400 (.Y (nx399), .A (\input [8])) ;
    tri01 tri_output_9 (.Y (\output [9]), .A (nx402), .E (nx503)) ;
    inv01 ix403 (.Y (nx402), .A (\input [9])) ;
    tri01 tri_output_10 (.Y (\output [10]), .A (nx405), .E (nx503)) ;
    inv01 ix406 (.Y (nx405), .A (\input [10])) ;
    tri01 tri_output_11 (.Y (\output [11]), .A (nx408), .E (nx503)) ;
    inv01 ix409 (.Y (nx408), .A (\input [11])) ;
    tri01 tri_output_12 (.Y (\output [12]), .A (nx411), .E (nx503)) ;
    inv01 ix412 (.Y (nx411), .A (\input [12])) ;
    tri01 tri_output_13 (.Y (\output [13]), .A (nx414), .E (nx503)) ;
    inv01 ix415 (.Y (nx414), .A (\input [13])) ;
    tri01 tri_output_14 (.Y (\output [14]), .A (nx417), .E (nx505)) ;
    inv01 ix418 (.Y (nx417), .A (\input [14])) ;
    tri01 tri_output_15 (.Y (\output [15]), .A (nx420), .E (nx505)) ;
    inv01 ix421 (.Y (nx420), .A (\input [15])) ;
    tri01 tri_output_16 (.Y (\output [16]), .A (nx423), .E (nx505)) ;
    inv01 ix424 (.Y (nx423), .A (\input [16])) ;
    tri01 tri_output_17 (.Y (\output [17]), .A (nx426), .E (nx505)) ;
    inv01 ix427 (.Y (nx426), .A (\input [17])) ;
    tri01 tri_output_18 (.Y (\output [18]), .A (nx429), .E (nx505)) ;
    inv01 ix430 (.Y (nx429), .A (\input [18])) ;
    tri01 tri_output_19 (.Y (\output [19]), .A (nx432), .E (nx505)) ;
    inv01 ix433 (.Y (nx432), .A (\input [19])) ;
    tri01 tri_output_20 (.Y (\output [20]), .A (nx435), .E (nx505)) ;
    inv01 ix436 (.Y (nx435), .A (\input [20])) ;
    tri01 tri_output_21 (.Y (\output [21]), .A (nx438), .E (nx507)) ;
    inv01 ix439 (.Y (nx438), .A (\input [21])) ;
    tri01 tri_output_22 (.Y (\output [22]), .A (nx441), .E (nx507)) ;
    inv01 ix442 (.Y (nx441), .A (\input [22])) ;
    tri01 tri_output_23 (.Y (\output [23]), .A (nx444), .E (nx507)) ;
    inv01 ix445 (.Y (nx444), .A (\input [23])) ;
    tri01 tri_output_24 (.Y (\output [24]), .A (nx447), .E (nx507)) ;
    inv01 ix448 (.Y (nx447), .A (\input [24])) ;
    tri01 tri_output_25 (.Y (\output [25]), .A (nx450), .E (nx507)) ;
    inv01 ix451 (.Y (nx450), .A (\input [25])) ;
    tri01 tri_output_26 (.Y (\output [26]), .A (nx453), .E (nx507)) ;
    inv01 ix454 (.Y (nx453), .A (\input [26])) ;
    tri01 tri_output_27 (.Y (\output [27]), .A (nx456), .E (nx507)) ;
    inv01 ix457 (.Y (nx456), .A (\input [27])) ;
    tri01 tri_output_28 (.Y (\output [28]), .A (nx459), .E (nx509)) ;
    inv01 ix460 (.Y (nx459), .A (\input [28])) ;
    tri01 tri_output_29 (.Y (\output [29]), .A (nx462), .E (nx509)) ;
    inv01 ix463 (.Y (nx462), .A (\input [29])) ;
    tri01 tri_output_30 (.Y (\output [30]), .A (nx465), .E (nx509)) ;
    inv01 ix466 (.Y (nx465), .A (\input [30])) ;
    tri01 tri_output_31 (.Y (\output [31]), .A (nx468), .E (nx509)) ;
    inv01 ix469 (.Y (nx468), .A (\input [31])) ;
    tri01 tri_output_32 (.Y (\output [32]), .A (nx471), .E (nx509)) ;
    inv01 ix472 (.Y (nx471), .A (\input [32])) ;
    tri01 tri_output_33 (.Y (\output [33]), .A (nx474), .E (nx509)) ;
    inv01 ix475 (.Y (nx474), .A (\input [33])) ;
    tri01 tri_output_34 (.Y (\output [34]), .A (nx477), .E (nx509)) ;
    inv01 ix478 (.Y (nx477), .A (\input [34])) ;
    tri01 tri_output_35 (.Y (\output [35]), .A (nx480), .E (nx511)) ;
    inv01 ix481 (.Y (nx480), .A (\input [35])) ;
    tri01 tri_output_36 (.Y (\output [36]), .A (nx483), .E (nx511)) ;
    inv01 ix484 (.Y (nx483), .A (\input [36])) ;
    tri01 tri_output_37 (.Y (\output [37]), .A (nx486), .E (nx511)) ;
    inv01 ix487 (.Y (nx486), .A (\input [37])) ;
    tri01 tri_output_38 (.Y (\output [38]), .A (nx489), .E (nx511)) ;
    inv01 ix490 (.Y (nx489), .A (\input [38])) ;
    tri01 tri_output_39 (.Y (\output [39]), .A (nx492), .E (nx511)) ;
    inv01 ix493 (.Y (nx492), .A (\input [39])) ;
    inv01 ix498 (.Y (nx499), .A (en)) ;
    inv01 ix500 (.Y (nx501), .A (nx499)) ;
    inv01 ix502 (.Y (nx503), .A (nx499)) ;
    inv01 ix504 (.Y (nx505), .A (nx499)) ;
    inv01 ix506 (.Y (nx507), .A (nx499)) ;
    inv01 ix508 (.Y (nx509), .A (nx499)) ;
    inv01 ix510 (.Y (nx511), .A (nx499)) ;
endmodule


module MultiStepCounter_12 ( load, toBeAdded, reset, clk, isLoad, MFC, count ) ;

    input [11:0]load ;
    input [11:0]toBeAdded ;
    input reset ;
    input clk ;
    input isLoad ;
    input MFC ;
    output [11:0]count ;

    wire loadOrCurrent_11, loadOrCurrent_10, loadOrCurrent_9, loadOrCurrent_8, 
         loadOrCurrent_7, loadOrCurrent_6, loadOrCurrent_5, loadOrCurrent_4, 
         loadOrCurrent_3, loadOrCurrent_2, loadOrCurrent_1, loadOrCurrent_0, 
         counterInput_11, counterInput_10, counterInput_9, counterInput_8, 
         counterInput_7, counterInput_6, counterInput_5, counterInput_4, 
         counterInput_3, counterInput_2, counterInput_1, counterInput_0, 
         countAdded_11, countAdded_10, countAdded_9, countAdded_8, countAdded_7, 
         countAdded_6, countAdded_5, countAdded_4, countAdded_3, countAdded_2, 
         countAdded_1, countAdded_0, GND, PWR;
    wire [0:0] \$dummy ;




    Reg_12 counterReg (.D ({counterInput_11,counterInput_10,counterInput_9,
           counterInput_8,counterInput_7,counterInput_6,counterInput_5,
           counterInput_4,counterInput_3,counterInput_2,counterInput_1,
           counterInput_0}), .en (PWR), .clk (clk), .rst (reset), .Q ({count[11]
           ,count[10],count[9],count[8],count[7],count[6],count[5],count[4],
           count[3],count[2],count[1],count[0]})) ;
    NBitAdder_12 nextCount (.a ({count[11],count[10],count[9],count[8],count[7],
                 count[6],count[5],count[4],count[3],count[2],count[1],count[0]}
                 ), .b ({toBeAdded[11],toBeAdded[10],toBeAdded[9],toBeAdded[8],
                 toBeAdded[7],toBeAdded[6],toBeAdded[5],toBeAdded[4],
                 toBeAdded[3],toBeAdded[2],toBeAdded[1],toBeAdded[0]}), .carryIn (
                 GND), .sum ({countAdded_11,countAdded_10,countAdded_9,
                 countAdded_8,countAdded_7,countAdded_6,countAdded_5,
                 countAdded_4,countAdded_3,countAdded_2,countAdded_1,
                 countAdded_0}), .carryOut (\$dummy [0])) ;
    Mux2_12 muxloadOrCurrent (.A ({count[11],count[10],count[9],count[8],
            count[7],count[6],count[5],count[4],count[3],count[2],count[1],
            count[0]}), .B ({load[11],load[10],load[9],load[8],load[7],load[6],
            load[5],load[4],load[3],load[2],load[1],load[0]}), .S (isLoad), .C (
            {loadOrCurrent_11,loadOrCurrent_10,loadOrCurrent_9,loadOrCurrent_8,
            loadOrCurrent_7,loadOrCurrent_6,loadOrCurrent_5,loadOrCurrent_4,
            loadOrCurrent_3,loadOrCurrent_2,loadOrCurrent_1,loadOrCurrent_0})) ;
    Mux2_12 muxInput (.A ({loadOrCurrent_11,loadOrCurrent_10,loadOrCurrent_9,
            loadOrCurrent_8,loadOrCurrent_7,loadOrCurrent_6,loadOrCurrent_5,
            loadOrCurrent_4,loadOrCurrent_3,loadOrCurrent_2,loadOrCurrent_1,
            loadOrCurrent_0}), .B ({countAdded_11,countAdded_10,countAdded_9,
            countAdded_8,countAdded_7,countAdded_6,countAdded_5,countAdded_4,
            countAdded_3,countAdded_2,countAdded_1,countAdded_0}), .S (MFC), .C (
            {counterInput_11,counterInput_10,counterInput_9,counterInput_8,
            counterInput_7,counterInput_6,counterInput_5,counterInput_4,
            counterInput_3,counterInput_2,counterInput_1,counterInput_0})) ;
    fake_vcc ix69 (.Y (PWR)) ;
    fake_gnd ix67 (.Y (GND)) ;
endmodule


module NBitAdder_12 ( a, b, carryIn, sum, carryOut ) ;

    input [11:0]a ;
    input [11:0]b ;
    input carryIn ;
    output [11:0]sum ;
    output carryOut ;

    wire temp_10, temp_9, temp_8, temp_7, temp_6, temp_5, temp_4, temp_3, temp_2, 
         temp_1, temp_0;



    FullAdder f0 (.a (a[0]), .b (b[0]), .cin (carryIn), .s (sum[0]), .cout (
              temp_0)) ;
    FullAdder loop1_1_fx (.a (a[1]), .b (b[1]), .cin (temp_0), .s (sum[1]), .cout (
              temp_1)) ;
    FullAdder loop1_2_fx (.a (a[2]), .b (b[2]), .cin (temp_1), .s (sum[2]), .cout (
              temp_2)) ;
    FullAdder loop1_3_fx (.a (a[3]), .b (b[3]), .cin (temp_2), .s (sum[3]), .cout (
              temp_3)) ;
    FullAdder loop1_4_fx (.a (a[4]), .b (b[4]), .cin (temp_3), .s (sum[4]), .cout (
              temp_4)) ;
    FullAdder loop1_5_fx (.a (a[5]), .b (b[5]), .cin (temp_4), .s (sum[5]), .cout (
              temp_5)) ;
    FullAdder loop1_6_fx (.a (a[6]), .b (b[6]), .cin (temp_5), .s (sum[6]), .cout (
              temp_6)) ;
    FullAdder loop1_7_fx (.a (a[7]), .b (b[7]), .cin (temp_6), .s (sum[7]), .cout (
              temp_7)) ;
    FullAdder loop1_8_fx (.a (a[8]), .b (b[8]), .cin (temp_7), .s (sum[8]), .cout (
              temp_8)) ;
    FullAdder loop1_9_fx (.a (a[9]), .b (b[9]), .cin (temp_8), .s (sum[9]), .cout (
              temp_9)) ;
    FullAdder loop1_10_fx (.a (a[10]), .b (b[10]), .cin (temp_9), .s (sum[10]), 
              .cout (temp_10)) ;
    FullAdder loop1_11_fx (.a (a[11]), .b (b[11]), .cin (temp_10), .s (sum[11])
              , .cout (carryOut)) ;
endmodule


module Reg_12 ( D, en, clk, rst, Q ) ;

    input [11:0]D ;
    input en ;
    input clk ;
    input rst ;
    output [11:0]Q ;

    wire nx180, nx190, nx200, nx210, nx220, nx230, nx240, nx250, nx260, nx270, 
         nx280, nx290;
    wire [11:0] \$dummy ;




    dffr reg_Q_0 (.Q (Q[0]), .QB (\$dummy [0]), .D (nx180), .CLK (clk), .R (rst)
         ) ;
    mux21_ni ix181 (.Y (nx180), .A0 (Q[0]), .A1 (D[0]), .S0 (en)) ;
    dffr reg_Q_1 (.Q (Q[1]), .QB (\$dummy [1]), .D (nx190), .CLK (clk), .R (rst)
         ) ;
    mux21_ni ix191 (.Y (nx190), .A0 (Q[1]), .A1 (D[1]), .S0 (en)) ;
    dffr reg_Q_2 (.Q (Q[2]), .QB (\$dummy [2]), .D (nx200), .CLK (clk), .R (rst)
         ) ;
    mux21_ni ix201 (.Y (nx200), .A0 (Q[2]), .A1 (D[2]), .S0 (en)) ;
    dffr reg_Q_3 (.Q (Q[3]), .QB (\$dummy [3]), .D (nx210), .CLK (clk), .R (rst)
         ) ;
    mux21_ni ix211 (.Y (nx210), .A0 (Q[3]), .A1 (D[3]), .S0 (en)) ;
    dffr reg_Q_4 (.Q (Q[4]), .QB (\$dummy [4]), .D (nx220), .CLK (clk), .R (rst)
         ) ;
    mux21_ni ix221 (.Y (nx220), .A0 (Q[4]), .A1 (D[4]), .S0 (en)) ;
    dffr reg_Q_5 (.Q (Q[5]), .QB (\$dummy [5]), .D (nx230), .CLK (clk), .R (rst)
         ) ;
    mux21_ni ix231 (.Y (nx230), .A0 (Q[5]), .A1 (D[5]), .S0 (en)) ;
    dffr reg_Q_6 (.Q (Q[6]), .QB (\$dummy [6]), .D (nx240), .CLK (clk), .R (rst)
         ) ;
    mux21_ni ix241 (.Y (nx240), .A0 (Q[6]), .A1 (D[6]), .S0 (en)) ;
    dffr reg_Q_7 (.Q (Q[7]), .QB (\$dummy [7]), .D (nx250), .CLK (clk), .R (rst)
         ) ;
    mux21_ni ix251 (.Y (nx250), .A0 (Q[7]), .A1 (D[7]), .S0 (en)) ;
    dffr reg_Q_8 (.Q (Q[8]), .QB (\$dummy [8]), .D (nx260), .CLK (clk), .R (rst)
         ) ;
    mux21_ni ix261 (.Y (nx260), .A0 (Q[8]), .A1 (D[8]), .S0 (en)) ;
    dffr reg_Q_9 (.Q (Q[9]), .QB (\$dummy [9]), .D (nx270), .CLK (clk), .R (rst)
         ) ;
    mux21_ni ix271 (.Y (nx270), .A0 (Q[9]), .A1 (D[9]), .S0 (en)) ;
    dffr reg_Q_10 (.Q (Q[10]), .QB (\$dummy [10]), .D (nx280), .CLK (clk), .R (
         rst)) ;
    mux21_ni ix281 (.Y (nx280), .A0 (Q[10]), .A1 (D[10]), .S0 (en)) ;
    dffr reg_Q_11 (.Q (Q[11]), .QB (\$dummy [11]), .D (nx290), .CLK (clk), .R (
         rst)) ;
    mux21_ni ix291 (.Y (nx290), .A0 (Q[11]), .A1 (D[11]), .S0 (en)) ;
endmodule


module Mux2_12 ( A, B, S, C ) ;

    input [11:0]A ;
    input [11:0]B ;
    input S ;
    output [11:0]C ;

    wire nx145, nx147;



    mux21_ni ix7 (.Y (C[0]), .A0 (A[0]), .A1 (B[0]), .S0 (nx145)) ;
    mux21_ni ix15 (.Y (C[1]), .A0 (A[1]), .A1 (B[1]), .S0 (nx145)) ;
    mux21_ni ix23 (.Y (C[2]), .A0 (A[2]), .A1 (B[2]), .S0 (nx145)) ;
    mux21_ni ix31 (.Y (C[3]), .A0 (A[3]), .A1 (B[3]), .S0 (nx145)) ;
    mux21_ni ix39 (.Y (C[4]), .A0 (A[4]), .A1 (B[4]), .S0 (nx145)) ;
    mux21_ni ix47 (.Y (C[5]), .A0 (A[5]), .A1 (B[5]), .S0 (nx145)) ;
    mux21_ni ix55 (.Y (C[6]), .A0 (A[6]), .A1 (B[6]), .S0 (nx145)) ;
    mux21_ni ix63 (.Y (C[7]), .A0 (A[7]), .A1 (B[7]), .S0 (nx147)) ;
    mux21_ni ix71 (.Y (C[8]), .A0 (A[8]), .A1 (B[8]), .S0 (nx147)) ;
    mux21_ni ix79 (.Y (C[9]), .A0 (A[9]), .A1 (B[9]), .S0 (nx147)) ;
    mux21_ni ix87 (.Y (C[10]), .A0 (A[10]), .A1 (B[10]), .S0 (nx147)) ;
    mux21_ni ix95 (.Y (C[11]), .A0 (A[11]), .A1 (B[11]), .S0 (nx147)) ;
    buf02 ix144 (.Y (nx145), .A (S)) ;
    buf02 ix146 (.Y (nx147), .A (S)) ;
endmodule


module ReadLogic_13_80_false ( clk, resetState, switchRam, ramBasedAddress, 
                               internalBus, ramDataInBus, ramRead, ramAddress, 
                               MFC, inputSize, filterSize, isFilter, 
                               loadNextWordList, loadWord, finishSlice, readOne, 
                               readFinal, aluNumber ) ;

    input clk ;
    input resetState ;
    input switchRam ;
    input [12:0]ramBasedAddress ;
    output [79:0]internalBus ;
    input [79:0]ramDataInBus ;
    output ramRead ;
    output [12:0]ramAddress ;
    input MFC ;
    input [12:0]inputSize ;
    input [12:0]filterSize ;
    input isFilter ;
    input loadNextWordList ;
    input loadWord ;
    input finishSlice ;
    output readOne ;
    output readFinal ;
    output [2:0]aluNumber ;

    wire addressRegOut_12, addressRegOut_11, addressRegOut_10, addressRegOut_9, 
         addressRegOut_8, addressRegOut_7, addressRegOut_6, addressRegOut_5, 
         addressRegOut_4, addressRegOut_3, addressRegOut_2, addressRegOut_1, 
         addressRegOut_0, addressRegInFinal_12, addressRegInFinal_11, 
         addressRegInFinal_10, addressRegInFinal_9, addressRegInFinal_8, 
         addressRegInFinal_7, addressRegInFinal_6, addressRegInFinal_5, 
         addressRegInFinal_4, addressRegInFinal_3, addressRegInFinal_2, 
         addressRegInFinal_1, addressRegInFinal_0, dmaInitAddress, 
         resetAddressReg, baseAddressCounterClk, aluNumberCounterClk, notClk, 
         aluCounterOut_2, aluCounterOut_1, aluCounterOut_0, 
         dmaReadBaseAddress_12, dmaReadBaseAddress_11, dmaReadBaseAddress_10, 
         dmaReadBaseAddress_9, dmaReadBaseAddress_8, dmaReadBaseAddress_7, 
         dmaReadBaseAddress_6, dmaReadBaseAddress_5, dmaReadBaseAddress_4, 
         dmaReadBaseAddress_3, dmaReadBaseAddress_2, dmaReadBaseAddress_1, 
         dmaReadBaseAddress_0, ramAddressKeeperOut_12, ramAddressKeeperOut_11, 
         ramAddressKeeperOut_10, ramAddressKeeperOut_9, ramAddressKeeperOut_8, 
         ramAddressKeeperOut_7, ramAddressKeeperOut_6, ramAddressKeeperOut_5, 
         ramAddressKeeperOut_4, ramAddressKeeperOut_3, ramAddressKeeperOut_2, 
         ramAddressKeeperOut_1, ramAddressKeeperOut_0, 
         ramAddressKeeperOutPlusFS_12, ramAddressKeeperOutPlusFS_11, 
         ramAddressKeeperOutPlusFS_10, ramAddressKeeperOutPlusFS_9, 
         ramAddressKeeperOutPlusFS_8, ramAddressKeeperOutPlusFS_7, 
         ramAddressKeeperOutPlusFS_6, ramAddressKeeperOutPlusFS_5, 
         ramAddressKeeperOutPlusFS_4, ramAddressKeeperOutPlusFS_3, 
         ramAddressKeeperOutPlusFS_2, ramAddressKeeperOutPlusFS_1, 
         ramAddressKeeperOutPlusFS_0, addressRegIn_12, addressRegIn_11, 
         addressRegIn_10, addressRegIn_9, addressRegIn_8, addressRegIn_7, 
         addressRegIn_6, addressRegIn_5, addressRegIn_4, addressRegIn_3, 
         addressRegIn_2, addressRegIn_1, addressRegIn_0, dmaCountIn_2, 
         dmaCountIn_1, dmaCountIn_0, dmaInitCounter, PWR, dmaInitRamBaseAddress, 
         currentState_0, nx4, nx16, nx30, nx32, nx598, nx608, nx618, nx621, 
         nx623, nx626, nx628, nx630, nx633, nx635, nx640, nx644, nx662, nx673, 
         nx675, nx677, nx679, nx681, nx687, nx689;
    wire [2:0] \$dummy ;




    Mux2_13 dmaReadBaseAddressMux (.A ({addressRegOut_12,addressRegOut_11,
            addressRegOut_10,addressRegOut_9,addressRegOut_8,addressRegOut_7,
            addressRegOut_6,addressRegOut_5,addressRegOut_4,addressRegOut_3,
            addressRegOut_2,addressRegOut_1,addressRegOut_0}), .B ({
            ramBasedAddress[12],ramBasedAddress[11],ramBasedAddress[10],
            ramBasedAddress[9],ramBasedAddress[8],ramBasedAddress[7],
            ramBasedAddress[6],ramBasedAddress[5],ramBasedAddress[4],
            ramBasedAddress[3],ramBasedAddress[2],ramBasedAddress[1],
            ramBasedAddress[0]}), .S (dmaInitRamBaseAddress), .C ({
            dmaReadBaseAddress_12,dmaReadBaseAddress_11,dmaReadBaseAddress_10,
            dmaReadBaseAddress_9,dmaReadBaseAddress_8,dmaReadBaseAddress_7,
            dmaReadBaseAddress_6,dmaReadBaseAddress_5,dmaReadBaseAddress_4,
            dmaReadBaseAddress_3,dmaReadBaseAddress_2,dmaReadBaseAddress_1,
            dmaReadBaseAddress_0})) ;
    DMA_13_80 dma (.initialCount ({dmaCountIn_2,dmaCountIn_1,dmaCountIn_0}), .readBaseAddress (
              {dmaReadBaseAddress_12,dmaReadBaseAddress_11,dmaReadBaseAddress_10
              ,dmaReadBaseAddress_9,dmaReadBaseAddress_8,dmaReadBaseAddress_7,
              dmaReadBaseAddress_6,dmaReadBaseAddress_5,dmaReadBaseAddress_4,
              dmaReadBaseAddress_3,dmaReadBaseAddress_2,dmaReadBaseAddress_1,
              dmaReadBaseAddress_0}), .readStep ({inputSize[12],inputSize[11],
              inputSize[10],inputSize[9],inputSize[8],inputSize[7],inputSize[6],
              inputSize[5],inputSize[4],inputSize[3],inputSize[2],inputSize[1],
              inputSize[0]}), .initAddress (dmaInitAddress), .initCounter (nx677
              ), .load (nx673), .internalBus ({internalBus[79],internalBus[78],
              internalBus[77],internalBus[76],internalBus[75],internalBus[74],
              internalBus[73],internalBus[72],internalBus[71],internalBus[70],
              internalBus[69],internalBus[68],internalBus[67],internalBus[66],
              internalBus[65],internalBus[64],internalBus[63],internalBus[62],
              internalBus[61],internalBus[60],internalBus[59],internalBus[58],
              internalBus[57],internalBus[56],internalBus[55],internalBus[54],
              internalBus[53],internalBus[52],internalBus[51],internalBus[50],
              internalBus[49],internalBus[48],internalBus[47],internalBus[46],
              internalBus[45],internalBus[44],internalBus[43],internalBus[42],
              internalBus[41],internalBus[40],internalBus[39],internalBus[38],
              internalBus[37],internalBus[36],internalBus[35],internalBus[34],
              internalBus[33],internalBus[32],internalBus[31],internalBus[30],
              internalBus[29],internalBus[28],internalBus[27],internalBus[26],
              internalBus[25],internalBus[24],internalBus[23],internalBus[22],
              internalBus[21],internalBus[20],internalBus[19],internalBus[18],
              internalBus[17],internalBus[16],internalBus[15],internalBus[14],
              internalBus[13],internalBus[12],internalBus[11],internalBus[10],
              internalBus[9],internalBus[8],internalBus[7],internalBus[6],
              internalBus[5],internalBus[4],internalBus[3],internalBus[2],
              internalBus[1],internalBus[0]}), .finishedOneReadOut (readOne), .finishedReading (
              readFinal), .clk (clk), .ramDataInBus ({ramDataInBus[79],
              ramDataInBus[78],ramDataInBus[77],ramDataInBus[76],
              ramDataInBus[75],ramDataInBus[74],ramDataInBus[73],
              ramDataInBus[72],ramDataInBus[71],ramDataInBus[70],
              ramDataInBus[69],ramDataInBus[68],ramDataInBus[67],
              ramDataInBus[66],ramDataInBus[65],ramDataInBus[64],
              ramDataInBus[63],ramDataInBus[62],ramDataInBus[61],
              ramDataInBus[60],ramDataInBus[59],ramDataInBus[58],
              ramDataInBus[57],ramDataInBus[56],ramDataInBus[55],
              ramDataInBus[54],ramDataInBus[53],ramDataInBus[52],
              ramDataInBus[51],ramDataInBus[50],ramDataInBus[49],
              ramDataInBus[48],ramDataInBus[47],ramDataInBus[46],
              ramDataInBus[45],ramDataInBus[44],ramDataInBus[43],
              ramDataInBus[42],ramDataInBus[41],ramDataInBus[40],
              ramDataInBus[39],ramDataInBus[38],ramDataInBus[37],
              ramDataInBus[36],ramDataInBus[35],ramDataInBus[34],
              ramDataInBus[33],ramDataInBus[32],ramDataInBus[31],
              ramDataInBus[30],ramDataInBus[29],ramDataInBus[28],
              ramDataInBus[27],ramDataInBus[26],ramDataInBus[25],
              ramDataInBus[24],ramDataInBus[23],ramDataInBus[22],
              ramDataInBus[21],ramDataInBus[20],ramDataInBus[19],
              ramDataInBus[18],ramDataInBus[17],ramDataInBus[16],
              ramDataInBus[15],ramDataInBus[14],ramDataInBus[13],
              ramDataInBus[12],ramDataInBus[11],ramDataInBus[10],ramDataInBus[9]
              ,ramDataInBus[8],ramDataInBus[7],ramDataInBus[6],ramDataInBus[5],
              ramDataInBus[4],ramDataInBus[3],ramDataInBus[2],ramDataInBus[1],
              ramDataInBus[0]}), .ramRead (\$dummy [0]), .ramReadAddress ({
              ramAddress[12],ramAddress[11],ramAddress[10],ramAddress[9],
              ramAddress[8],ramAddress[7],ramAddress[6],ramAddress[5],
              ramAddress[4],ramAddress[3],ramAddress[2],ramAddress[1],
              ramAddress[0]}), .MFC (MFC)) ;
    NBitAdder_13 window_g_ramAddressIncrement (.a ({ramAddressKeeperOut_12,
                 ramAddressKeeperOut_11,ramAddressKeeperOut_10,
                 ramAddressKeeperOut_9,ramAddressKeeperOut_8,
                 ramAddressKeeperOut_7,ramAddressKeeperOut_6,
                 ramAddressKeeperOut_5,ramAddressKeeperOut_4,
                 ramAddressKeeperOut_3,ramAddressKeeperOut_2,
                 ramAddressKeeperOut_1,ramAddressKeeperOut_0}), .b ({
                 filterSize[12],filterSize[11],filterSize[10],filterSize[9],
                 filterSize[8],filterSize[7],filterSize[6],filterSize[5],
                 filterSize[4],filterSize[3],filterSize[2],filterSize[1],
                 filterSize[0]}), .carryIn (dmaInitRamBaseAddress), .sum ({
                 ramAddressKeeperOutPlusFS_12,ramAddressKeeperOutPlusFS_11,
                 ramAddressKeeperOutPlusFS_10,ramAddressKeeperOutPlusFS_9,
                 ramAddressKeeperOutPlusFS_8,ramAddressKeeperOutPlusFS_7,
                 ramAddressKeeperOutPlusFS_6,ramAddressKeeperOutPlusFS_5,
                 ramAddressKeeperOutPlusFS_4,ramAddressKeeperOutPlusFS_3,
                 ramAddressKeeperOutPlusFS_2,ramAddressKeeperOutPlusFS_1,
                 ramAddressKeeperOutPlusFS_0}), .carryOut (\$dummy [1])) ;
    Mux2_13 window_g_baseAddressLoadMux (.A ({addressRegIn_12,addressRegIn_11,
            addressRegIn_10,addressRegIn_9,addressRegIn_8,addressRegIn_7,
            addressRegIn_6,addressRegIn_5,addressRegIn_4,addressRegIn_3,
            addressRegIn_2,addressRegIn_1,addressRegIn_0}), .B ({
            ramAddressKeeperOutPlusFS_12,ramAddressKeeperOutPlusFS_11,
            ramAddressKeeperOutPlusFS_10,ramAddressKeeperOutPlusFS_9,
            ramAddressKeeperOutPlusFS_8,ramAddressKeeperOutPlusFS_7,
            ramAddressKeeperOutPlusFS_6,ramAddressKeeperOutPlusFS_5,
            ramAddressKeeperOutPlusFS_4,ramAddressKeeperOutPlusFS_3,
            ramAddressKeeperOutPlusFS_2,ramAddressKeeperOutPlusFS_1,
            ramAddressKeeperOutPlusFS_0}), .S (finishSlice), .C ({
            addressRegInFinal_12,addressRegInFinal_11,addressRegInFinal_10,
            addressRegInFinal_9,addressRegInFinal_8,addressRegInFinal_7,
            addressRegInFinal_6,addressRegInFinal_5,addressRegInFinal_4,
            addressRegInFinal_3,addressRegInFinal_2,addressRegInFinal_1,
            addressRegInFinal_0})) ;
    Counter2_13 window_g_baseAddressCounter (.load ({addressRegInFinal_12,
                addressRegInFinal_11,addressRegInFinal_10,addressRegInFinal_9,
                addressRegInFinal_8,addressRegInFinal_7,addressRegInFinal_6,
                addressRegInFinal_5,addressRegInFinal_4,addressRegInFinal_3,
                addressRegInFinal_2,addressRegInFinal_1,addressRegInFinal_0}), .reset (
                dmaInitRamBaseAddress), .clk (baseAddressCounterClk), .isLoad (
                resetAddressReg), .count ({addressRegOut_12,addressRegOut_11,
                addressRegOut_10,addressRegOut_9,addressRegOut_8,addressRegOut_7
                ,addressRegOut_6,addressRegOut_5,addressRegOut_4,addressRegOut_3
                ,addressRegOut_2,addressRegOut_1,addressRegOut_0})) ;
    Reg_13 window_g_ramAddressKeeper (.D ({ramAddress[12],ramAddress[11],
           ramAddress[10],ramAddress[9],ramAddress[8],ramAddress[7],
           ramAddress[6],ramAddress[5],ramAddress[4],ramAddress[3],ramAddress[2]
           ,ramAddress[1],ramAddress[0]}), .en (nx673), .clk (clk), .rst (
           dmaInitRamBaseAddress), .Q ({ramAddressKeeperOut_12,
           ramAddressKeeperOut_11,ramAddressKeeperOut_10,ramAddressKeeperOut_9,
           ramAddressKeeperOut_8,ramAddressKeeperOut_7,ramAddressKeeperOut_6,
           ramAddressKeeperOut_5,ramAddressKeeperOut_4,ramAddressKeeperOut_3,
           ramAddressKeeperOut_2,ramAddressKeeperOut_1,ramAddressKeeperOut_0})
           ) ;
    Counter2_3 aluNumberCounter (.load ({dmaInitRamBaseAddress,
               dmaInitRamBaseAddress,dmaInitRamBaseAddress}), .reset (nx687), .clk (
               aluNumberCounterClk), .isLoad (dmaInitRamBaseAddress), .count ({
               aluCounterOut_2,aluCounterOut_1,aluCounterOut_0})) ;
    Reg_3 regCounterOut (.D ({aluCounterOut_2,aluCounterOut_1,aluCounterOut_0})
          , .en (PWR), .clk (notClk), .rst (dmaInitRamBaseAddress), .Q ({
          aluNumber[2],aluNumber[1],aluNumber[0]})) ;
    ao21 ix609 (.Y (nx608), .A0 (nx673), .A1 (nx618), .B0 (nx16)) ;
    dffr reg_currentState_1 (.Q (ramRead), .QB (\$dummy [2]), .D (nx608), .CLK (
         notClk), .R (resetState)) ;
    inv01 ix617 (.Y (notClk), .A (clk)) ;
    nor04 ix619 (.Y (nx618), .A0 (nx16), .A1 (switchRam), .A2 (nx32), .A3 (nx679
          )) ;
    aoi21 ix17 (.Y (nx16), .A0 (nx621), .A1 (nx630), .B0 (switchRam)) ;
    oai21 ix622 (.Y (nx621), .A0 (loadNextWordList), .A1 (loadWord), .B0 (nx623)
          ) ;
    dffr reg_currentState_0 (.Q (currentState_0), .QB (nx623), .D (nx598), .CLK (
         notClk), .R (resetState)) ;
    mux21 ix599 (.Y (nx598), .A0 (nx626), .A1 (nx623), .S0 (nx618)) ;
    aoi221 ix627 (.Y (nx626), .A0 (nx673), .A1 (nx623), .B0 (nx628), .B1 (nx16)
           , .C0 (switchRam)) ;
    inv01 ix629 (.Y (nx628), .A (loadNextWordList)) ;
    nor02ii ix33 (.Y (nx32), .A0 (nx633), .A1 (readFinal)) ;
    fake_gnd ix564 (.Y (dmaInitRamBaseAddress)) ;
    fake_vcc ix562 (.Y (PWR)) ;
    aoi21 ix63 (.Y (dmaInitCounter), .A0 (nx628), .A1 (nx640), .B0 (nx30)) ;
    inv01 ix641 (.Y (nx640), .A (loadWord)) ;
    inv01 ix69 (.Y (dmaCountIn_0), .A (nx644)) ;
    oai21 ix645 (.Y (nx644), .A0 (nx628), .A1 (filterSize[0]), .B0 (nx677)) ;
    and03 ix75 (.Y (dmaCountIn_1), .A0 (nx633), .A1 (filterSize[1]), .A2 (
          loadNextWordList)) ;
    and03 ix81 (.Y (dmaCountIn_2), .A0 (nx633), .A1 (filterSize[2]), .A2 (
          loadNextWordList)) ;
    and02 ix85 (.Y (addressRegIn_0), .A0 (ramBasedAddress[0]), .A1 (nx679)) ;
    and02 ix89 (.Y (addressRegIn_1), .A0 (ramBasedAddress[1]), .A1 (nx679)) ;
    and02 ix93 (.Y (addressRegIn_2), .A0 (ramBasedAddress[2]), .A1 (nx679)) ;
    and02 ix97 (.Y (addressRegIn_3), .A0 (ramBasedAddress[3]), .A1 (nx679)) ;
    and02 ix101 (.Y (addressRegIn_4), .A0 (ramBasedAddress[4]), .A1 (nx679)) ;
    and02 ix105 (.Y (addressRegIn_5), .A0 (ramBasedAddress[5]), .A1 (nx679)) ;
    and02 ix109 (.Y (addressRegIn_6), .A0 (ramBasedAddress[6]), .A1 (nx681)) ;
    and02 ix113 (.Y (addressRegIn_7), .A0 (ramBasedAddress[7]), .A1 (nx681)) ;
    and02 ix117 (.Y (addressRegIn_8), .A0 (ramBasedAddress[8]), .A1 (nx681)) ;
    and02 ix121 (.Y (addressRegIn_9), .A0 (ramBasedAddress[9]), .A1 (nx681)) ;
    and02 ix125 (.Y (addressRegIn_10), .A0 (ramBasedAddress[10]), .A1 (nx681)) ;
    and02 ix129 (.Y (addressRegIn_11), .A0 (ramBasedAddress[11]), .A1 (nx681)) ;
    and02 ix133 (.Y (addressRegIn_12), .A0 (ramBasedAddress[12]), .A1 (nx681)) ;
    aoi21 ix141 (.Y (aluNumberCounterClk), .A0 (nx662), .A1 (nx675), .B0 (notClk
          )) ;
    nand02 ix663 (.Y (nx662), .A0 (loadNextWordList), .A1 (readOne)) ;
    mux21_ni ix155 (.Y (baseAddressCounterClk), .A0 (resetAddressReg), .A1 (nx4)
             , .S0 (clk)) ;
    or02 ix149 (.Y (resetAddressReg), .A0 (nx635), .A1 (finishSlice)) ;
    aoi21 ix57 (.Y (dmaInitAddress), .A0 (nx628), .A1 (nx623), .B0 (nx675)) ;
    inv01 ix31 (.Y (nx30), .A (nx633)) ;
    inv01 ix5 (.Y (nx4), .A (nx630)) ;
    inv02 ix672 (.Y (nx673), .A (nx687)) ;
    inv02 ix674 (.Y (nx675), .A (nx687)) ;
    buf02 ix676 (.Y (nx677), .A (dmaInitCounter)) ;
    or02 ix631 (.Y (nx630), .A0 (nx687), .A1 (currentState_0)) ;
    and02 ix634 (.Y (nx633), .A0 (nx623), .A1 (nx687)) ;
    and02 ix636 (.Y (nx635), .A0 (currentState_0), .A1 (nx689)) ;
    and02 ix678 (.Y (nx679), .A0 (currentState_0), .A1 (nx689)) ;
    and02 ix680 (.Y (nx681), .A0 (currentState_0), .A1 (nx689)) ;
    inv02 ix686 (.Y (nx687), .A (ramRead)) ;
    inv02 ix688 (.Y (nx689), .A (ramRead)) ;
endmodule


module Counter2_3 ( load, reset, clk, isLoad, count ) ;

    input [2:0]load ;
    input reset ;
    input clk ;
    input isLoad ;
    output [2:0]count ;

    wire counterInput_2, counterInput_1, counterInput_0, countAdded_2, 
         countAdded_1, countAdded_0, resetOrCurrent_2, resetOrCurrent_1, 
         resetOrCurrent_0, zerosSignal_2, PWR;
    wire [0:0] \$dummy ;




    Reg_3 counterReg (.D ({counterInput_2,counterInput_1,counterInput_0}), .en (
          PWR), .clk (clk), .rst (zerosSignal_2), .Q ({count[2],count[1],
          count[0]})) ;
    NBitAdder_3 nextCount (.a ({count[2],count[1],count[0]}), .b ({zerosSignal_2
                ,zerosSignal_2,zerosSignal_2}), .carryIn (PWR), .sum ({
                countAdded_2,countAdded_1,countAdded_0}), .carryOut (\$dummy [0]
                )) ;
    Mux2_3 muxloadOrCurrent (.A ({resetOrCurrent_2,resetOrCurrent_1,
           resetOrCurrent_0}), .B ({load[2],load[1],load[0]}), .S (isLoad), .C (
           {counterInput_2,counterInput_1,counterInput_0})) ;
    Mux2_3 muxInput (.A ({countAdded_2,countAdded_1,countAdded_0}), .B ({
           zerosSignal_2,zerosSignal_2,zerosSignal_2}), .S (reset), .C ({
           resetOrCurrent_2,resetOrCurrent_1,resetOrCurrent_0})) ;
    fake_vcc ix24 (.Y (PWR)) ;
    fake_gnd ix22 (.Y (zerosSignal_2)) ;
endmodule


module Counter2_13 ( load, reset, clk, isLoad, count ) ;

    input [12:0]load ;
    input reset ;
    input clk ;
    input isLoad ;
    output [12:0]count ;

    wire counterInput_12, counterInput_11, counterInput_10, counterInput_9, 
         counterInput_8, counterInput_7, counterInput_6, counterInput_5, 
         counterInput_4, counterInput_3, counterInput_2, counterInput_1, 
         counterInput_0, countAdded_12, countAdded_11, countAdded_10, 
         countAdded_9, countAdded_8, countAdded_7, countAdded_6, countAdded_5, 
         countAdded_4, countAdded_3, countAdded_2, countAdded_1, countAdded_0, 
         resetOrCurrent_12, resetOrCurrent_11, resetOrCurrent_10, 
         resetOrCurrent_9, resetOrCurrent_8, resetOrCurrent_7, resetOrCurrent_6, 
         resetOrCurrent_5, resetOrCurrent_4, resetOrCurrent_3, resetOrCurrent_2, 
         resetOrCurrent_1, resetOrCurrent_0, zerosSignal_12, PWR;
    wire [0:0] \$dummy ;




    Reg_13 counterReg (.D ({counterInput_12,counterInput_11,counterInput_10,
           counterInput_9,counterInput_8,counterInput_7,counterInput_6,
           counterInput_5,counterInput_4,counterInput_3,counterInput_2,
           counterInput_1,counterInput_0}), .en (PWR), .clk (clk), .rst (
           zerosSignal_12), .Q ({count[12],count[11],count[10],count[9],count[8]
           ,count[7],count[6],count[5],count[4],count[3],count[2],count[1],
           count[0]})) ;
    NBitAdder_13 nextCount (.a ({count[12],count[11],count[10],count[9],count[8]
                 ,count[7],count[6],count[5],count[4],count[3],count[2],count[1]
                 ,count[0]}), .b ({zerosSignal_12,zerosSignal_12,zerosSignal_12,
                 zerosSignal_12,zerosSignal_12,zerosSignal_12,zerosSignal_12,
                 zerosSignal_12,zerosSignal_12,zerosSignal_12,zerosSignal_12,
                 zerosSignal_12,zerosSignal_12}), .carryIn (PWR), .sum ({
                 countAdded_12,countAdded_11,countAdded_10,countAdded_9,
                 countAdded_8,countAdded_7,countAdded_6,countAdded_5,
                 countAdded_4,countAdded_3,countAdded_2,countAdded_1,
                 countAdded_0}), .carryOut (\$dummy [0])) ;
    Mux2_13 muxloadOrCurrent (.A ({resetOrCurrent_12,resetOrCurrent_11,
            resetOrCurrent_10,resetOrCurrent_9,resetOrCurrent_8,resetOrCurrent_7
            ,resetOrCurrent_6,resetOrCurrent_5,resetOrCurrent_4,resetOrCurrent_3
            ,resetOrCurrent_2,resetOrCurrent_1,resetOrCurrent_0}), .B ({load[12]
            ,load[11],load[10],load[9],load[8],load[7],load[6],load[5],load[4],
            load[3],load[2],load[1],load[0]}), .S (isLoad), .C ({counterInput_12
            ,counterInput_11,counterInput_10,counterInput_9,counterInput_8,
            counterInput_7,counterInput_6,counterInput_5,counterInput_4,
            counterInput_3,counterInput_2,counterInput_1,counterInput_0})) ;
    Mux2_13 muxInput (.A ({countAdded_12,countAdded_11,countAdded_10,
            countAdded_9,countAdded_8,countAdded_7,countAdded_6,countAdded_5,
            countAdded_4,countAdded_3,countAdded_2,countAdded_1,countAdded_0}), 
            .B ({zerosSignal_12,zerosSignal_12,zerosSignal_12,zerosSignal_12,
            zerosSignal_12,zerosSignal_12,zerosSignal_12,zerosSignal_12,
            zerosSignal_12,zerosSignal_12,zerosSignal_12,zerosSignal_12,
            zerosSignal_12}), .S (reset), .C ({resetOrCurrent_12,
            resetOrCurrent_11,resetOrCurrent_10,resetOrCurrent_9,
            resetOrCurrent_8,resetOrCurrent_7,resetOrCurrent_6,resetOrCurrent_5,
            resetOrCurrent_4,resetOrCurrent_3,resetOrCurrent_2,resetOrCurrent_1,
            resetOrCurrent_0})) ;
    fake_vcc ix74 (.Y (PWR)) ;
    fake_gnd ix72 (.Y (zerosSignal_12)) ;
endmodule


module DMA_13_80 ( initialCount, readBaseAddress, readStep, initAddress, 
                   initCounter, load, internalBus, finishedOneReadOut, 
                   finishedReading, clk, ramDataInBus, ramRead, ramReadAddress, 
                   MFC ) ;

    input [2:0]initialCount ;
    input [12:0]readBaseAddress ;
    input [12:0]readStep ;
    input initAddress ;
    input initCounter ;
    input load ;
    output [79:0]internalBus ;
    output finishedOneReadOut ;
    output finishedReading ;
    input clk ;
    input [79:0]ramDataInBus ;
    output ramRead ;
    output [12:0]ramReadAddress ;
    input MFC ;

    wire currentCount_2, currentCount_1, currentCount_0, tobeAdded_12, 
         tobeAdded_11, tobeAdded_10, tobeAdded_9, tobeAdded_8, tobeAdded_7, 
         tobeAdded_6, tobeAdded_5, tobeAdded_4, tobeAdded_3, tobeAdded_2, 
         tobeAdded_1, tobeAdded_0, enableCount, PWR, GND, NOT_MFC, nx18, nx175, 
         nx177, nx179, nx1, nx5;



    assign ramRead = load ;
    MultiStepCounter_13 addressRegister (.load ({readBaseAddress[12],
                        readBaseAddress[11],readBaseAddress[10],
                        readBaseAddress[9],readBaseAddress[8],readBaseAddress[7]
                        ,readBaseAddress[6],readBaseAddress[5],
                        readBaseAddress[4],readBaseAddress[3],readBaseAddress[2]
                        ,readBaseAddress[1],readBaseAddress[0]}), .toBeAdded ({
                        tobeAdded_12,tobeAdded_11,tobeAdded_10,tobeAdded_9,
                        tobeAdded_8,tobeAdded_7,tobeAdded_6,tobeAdded_5,
                        tobeAdded_4,tobeAdded_3,tobeAdded_2,tobeAdded_1,
                        tobeAdded_0}), .reset (GND), .clk (clk), .isLoad (
                        initAddress), .MFC (finishedOneReadOut), .count ({
                        ramReadAddress[12],ramReadAddress[11],ramReadAddress[10]
                        ,ramReadAddress[9],ramReadAddress[8],ramReadAddress[7],
                        ramReadAddress[6],ramReadAddress[5],ramReadAddress[4],
                        ramReadAddress[3],ramReadAddress[2],ramReadAddress[1],
                        ramReadAddress[0]})) ;
    DownCounter_3 counter (.load ({initialCount[2],initialCount[1],
                  initialCount[0]}), .enable (enableCount), .clk (clk), .isLoad (
                  initCounter), .currentCount ({currentCount_2,currentCount_1,
                  currentCount_0})) ;
    Reg_13 readStepRegister (.D ({readStep[12],readStep[11],readStep[10],
           readStep[9],readStep[8],readStep[7],readStep[6],readStep[5],
           readStep[4],readStep[3],readStep[2],readStep[1],readStep[0]}), .en (
           PWR), .clk (clk), .rst (GND), .Q ({tobeAdded_12,tobeAdded_11,
           tobeAdded_10,tobeAdded_9,tobeAdded_8,tobeAdded_7,tobeAdded_6,
           tobeAdded_5,tobeAdded_4,tobeAdded_3,tobeAdded_2,tobeAdded_1,
           tobeAdded_0})) ;
    Tristate_80 tristateLabel (.\input  ({ramDataInBus[79],ramDataInBus[78],
                ramDataInBus[77],ramDataInBus[76],ramDataInBus[75],
                ramDataInBus[74],ramDataInBus[73],ramDataInBus[72],
                ramDataInBus[71],ramDataInBus[70],ramDataInBus[69],
                ramDataInBus[68],ramDataInBus[67],ramDataInBus[66],
                ramDataInBus[65],ramDataInBus[64],ramDataInBus[63],
                ramDataInBus[62],ramDataInBus[61],ramDataInBus[60],
                ramDataInBus[59],ramDataInBus[58],ramDataInBus[57],
                ramDataInBus[56],ramDataInBus[55],ramDataInBus[54],
                ramDataInBus[53],ramDataInBus[52],ramDataInBus[51],
                ramDataInBus[50],ramDataInBus[49],ramDataInBus[48],
                ramDataInBus[47],ramDataInBus[46],ramDataInBus[45],
                ramDataInBus[44],ramDataInBus[43],ramDataInBus[42],
                ramDataInBus[41],ramDataInBus[40],ramDataInBus[39],
                ramDataInBus[38],ramDataInBus[37],ramDataInBus[36],
                ramDataInBus[35],ramDataInBus[34],ramDataInBus[33],
                ramDataInBus[32],ramDataInBus[31],ramDataInBus[30],
                ramDataInBus[29],ramDataInBus[28],ramDataInBus[27],
                ramDataInBus[26],ramDataInBus[25],ramDataInBus[24],
                ramDataInBus[23],ramDataInBus[22],ramDataInBus[21],
                ramDataInBus[20],ramDataInBus[19],ramDataInBus[18],
                ramDataInBus[17],ramDataInBus[16],ramDataInBus[15],
                ramDataInBus[14],ramDataInBus[13],ramDataInBus[12],
                ramDataInBus[11],ramDataInBus[10],ramDataInBus[9],
                ramDataInBus[8],ramDataInBus[7],ramDataInBus[6],ramDataInBus[5],
                ramDataInBus[4],ramDataInBus[3],ramDataInBus[2],ramDataInBus[1],
                ramDataInBus[0]}), .en (finishedOneReadOut), .\output  ({
                internalBus[79],internalBus[78],internalBus[77],internalBus[76],
                internalBus[75],internalBus[74],internalBus[73],internalBus[72],
                internalBus[71],internalBus[70],internalBus[69],internalBus[68],
                internalBus[67],internalBus[66],internalBus[65],internalBus[64],
                internalBus[63],internalBus[62],internalBus[61],internalBus[60],
                internalBus[59],internalBus[58],internalBus[57],internalBus[56],
                internalBus[55],internalBus[54],internalBus[53],internalBus[52],
                internalBus[51],internalBus[50],internalBus[49],internalBus[48],
                internalBus[47],internalBus[46],internalBus[45],internalBus[44],
                internalBus[43],internalBus[42],internalBus[41],internalBus[40],
                internalBus[39],internalBus[38],internalBus[37],internalBus[36],
                internalBus[35],internalBus[34],internalBus[33],internalBus[32],
                internalBus[31],internalBus[30],internalBus[29],internalBus[28],
                internalBus[27],internalBus[26],internalBus[25],internalBus[24],
                internalBus[23],internalBus[22],internalBus[21],internalBus[20],
                internalBus[19],internalBus[18],internalBus[17],internalBus[16],
                internalBus[15],internalBus[14],internalBus[13],internalBus[12],
                internalBus[11],internalBus[10],internalBus[9],internalBus[8],
                internalBus[7],internalBus[6],internalBus[5],internalBus[4],
                internalBus[3],internalBus[2],internalBus[1],internalBus[0]})) ;
    fake_gnd ix158 (.Y (GND)) ;
    fake_vcc ix156 (.Y (PWR)) ;
    and02 ix13 (.Y (finishedOneReadOut), .A0 (load), .A1 (MFC)) ;
    or02 ix25 (.Y (enableCount), .A0 (MFC), .A1 (initCounter)) ;
    inv16 ix173 (.Y (NOT_MFC), .A (MFC)) ;
    nor04 ix19 (.Y (nx18), .A0 (currentCount_1), .A1 (nx175), .A2 (
          currentCount_2), .A3 (nx177)) ;
    inv01 ix176 (.Y (nx175), .A (currentCount_0)) ;
    nand02 ix178 (.Y (nx177), .A0 (nx179), .A1 (finishedOneReadOut)) ;
    inv01 ix180 (.Y (nx179), .A (clk)) ;
    latchs_ni lat_internalFinishedReading_u1 (.QB (nx5), .D (GND), .CLK (NOT_MFC
              ), .S (nx18)) ;
    inv02 lat_internalFinishedReading_u2 (.Y (finishedReading), .A (nx5)) ;
    buf02 lat_internalFinishedReading_u3 (.Y (nx1), .A (nx5)) ;
endmodule


module DownCounter_3 ( load, enable, clk, isLoad, currentCount ) ;

    input [2:0]load ;
    input enable ;
    input clk ;
    input isLoad ;
    inout [2:0]currentCount ;

    wire counterInput_2, counterInput_1, counterInput_0, subtractorOutput_2, 
         subtractorOutput_1, subtractorOutput_0, PWR, zerosSignal_2;
    wire [0:0] \$dummy ;




    Reg_3 counterReg (.D ({counterInput_2,counterInput_1,counterInput_0}), .en (
          enable), .clk (clk), .rst (zerosSignal_2), .Q ({currentCount[2],
          currentCount[1],currentCount[0]})) ;
    NBitSubtractor_3 nextCount (.x ({currentCount[2],currentCount[1],
                     currentCount[0]}), .y ({zerosSignal_2,zerosSignal_2,
                     zerosSignal_2}), .bin (PWR), .difference ({
                     subtractorOutput_2,subtractorOutput_1,subtractorOutput_0})
                     , .borrowOut (\$dummy [0])) ;
    Mux2_3 muxloadOrCurrent (.A ({subtractorOutput_2,subtractorOutput_1,
           subtractorOutput_0}), .B ({load[2],load[1],load[0]}), .S (isLoad), .C (
           {counterInput_2,counterInput_1,counterInput_0})) ;
    fake_gnd ix18 (.Y (zerosSignal_2)) ;
    fake_vcc ix16 (.Y (PWR)) ;
endmodule


module Mux2_3 ( A, B, S, C ) ;

    input [2:0]A ;
    input [2:0]B ;
    input S ;
    output [2:0]C ;




    mux21_ni ix7 (.Y (C[0]), .A0 (A[0]), .A1 (B[0]), .S0 (S)) ;
    mux21_ni ix15 (.Y (C[1]), .A0 (A[1]), .A1 (B[1]), .S0 (S)) ;
    mux21_ni ix23 (.Y (C[2]), .A0 (A[2]), .A1 (B[2]), .S0 (S)) ;
endmodule


module NBitSubtractor_3 ( x, y, bin, difference, borrowOut ) ;

    input [2:0]x ;
    input [2:0]y ;
    input bin ;
    output [2:0]difference ;
    output borrowOut ;

    wire temp_1, temp_0;



    FullSubtractor f0 (.x (x[0]), .y (y[0]), .bin (bin), .difference (
                   difference[0]), .bout (temp_0)) ;
    FullSubtractor loop1_1_fx (.x (x[1]), .y (y[1]), .bin (temp_0), .difference (
                   difference[1]), .bout (temp_1)) ;
    FullSubtractor loop1_2_fx (.x (x[2]), .y (y[2]), .bin (temp_1), .difference (
                   difference[2]), .bout (borrowOut)) ;
endmodule


module FullSubtractor ( x, y, bin, difference, bout ) ;

    input x ;
    input y ;
    input bin ;
    output difference ;
    output bout ;

    wire nx71, nx73;



    mux21_ni ix11 (.Y (bout), .A0 (nx71), .A1 (bin), .S0 (nx73)) ;
    inv01 ix72 (.Y (nx71), .A (x)) ;
    xnor2 ix74 (.Y (nx73), .A0 (x), .A1 (y)) ;
    xnor2 ix13 (.Y (difference), .A0 (nx73), .A1 (bin)) ;
endmodule


module MultiStepCounter_13 ( load, toBeAdded, reset, clk, isLoad, MFC, count ) ;

    input [12:0]load ;
    input [12:0]toBeAdded ;
    input reset ;
    input clk ;
    input isLoad ;
    input MFC ;
    output [12:0]count ;

    wire loadOrCurrent_12, loadOrCurrent_11, loadOrCurrent_10, loadOrCurrent_9, 
         loadOrCurrent_8, loadOrCurrent_7, loadOrCurrent_6, loadOrCurrent_5, 
         loadOrCurrent_4, loadOrCurrent_3, loadOrCurrent_2, loadOrCurrent_1, 
         loadOrCurrent_0, counterInput_12, counterInput_11, counterInput_10, 
         counterInput_9, counterInput_8, counterInput_7, counterInput_6, 
         counterInput_5, counterInput_4, counterInput_3, counterInput_2, 
         counterInput_1, counterInput_0, countAdded_12, countAdded_11, 
         countAdded_10, countAdded_9, countAdded_8, countAdded_7, countAdded_6, 
         countAdded_5, countAdded_4, countAdded_3, countAdded_2, countAdded_1, 
         countAdded_0, GND, PWR;
    wire [0:0] \$dummy ;




    Reg_13 counterReg (.D ({counterInput_12,counterInput_11,counterInput_10,
           counterInput_9,counterInput_8,counterInput_7,counterInput_6,
           counterInput_5,counterInput_4,counterInput_3,counterInput_2,
           counterInput_1,counterInput_0}), .en (PWR), .clk (clk), .rst (reset)
           , .Q ({count[12],count[11],count[10],count[9],count[8],count[7],
           count[6],count[5],count[4],count[3],count[2],count[1],count[0]})) ;
    NBitAdder_13 nextCount (.a ({count[12],count[11],count[10],count[9],count[8]
                 ,count[7],count[6],count[5],count[4],count[3],count[2],count[1]
                 ,count[0]}), .b ({toBeAdded[12],toBeAdded[11],toBeAdded[10],
                 toBeAdded[9],toBeAdded[8],toBeAdded[7],toBeAdded[6],
                 toBeAdded[5],toBeAdded[4],toBeAdded[3],toBeAdded[2],
                 toBeAdded[1],toBeAdded[0]}), .carryIn (GND), .sum ({
                 countAdded_12,countAdded_11,countAdded_10,countAdded_9,
                 countAdded_8,countAdded_7,countAdded_6,countAdded_5,
                 countAdded_4,countAdded_3,countAdded_2,countAdded_1,
                 countAdded_0}), .carryOut (\$dummy [0])) ;
    Mux2_13 muxloadOrCurrent (.A ({count[12],count[11],count[10],count[9],
            count[8],count[7],count[6],count[5],count[4],count[3],count[2],
            count[1],count[0]}), .B ({load[12],load[11],load[10],load[9],load[8]
            ,load[7],load[6],load[5],load[4],load[3],load[2],load[1],load[0]}), 
            .S (isLoad), .C ({loadOrCurrent_12,loadOrCurrent_11,loadOrCurrent_10
            ,loadOrCurrent_9,loadOrCurrent_8,loadOrCurrent_7,loadOrCurrent_6,
            loadOrCurrent_5,loadOrCurrent_4,loadOrCurrent_3,loadOrCurrent_2,
            loadOrCurrent_1,loadOrCurrent_0})) ;
    Mux2_13 muxInput (.A ({loadOrCurrent_12,loadOrCurrent_11,loadOrCurrent_10,
            loadOrCurrent_9,loadOrCurrent_8,loadOrCurrent_7,loadOrCurrent_6,
            loadOrCurrent_5,loadOrCurrent_4,loadOrCurrent_3,loadOrCurrent_2,
            loadOrCurrent_1,loadOrCurrent_0}), .B ({countAdded_12,countAdded_11,
            countAdded_10,countAdded_9,countAdded_8,countAdded_7,countAdded_6,
            countAdded_5,countAdded_4,countAdded_3,countAdded_2,countAdded_1,
            countAdded_0}), .S (MFC), .C ({counterInput_12,counterInput_11,
            counterInput_10,counterInput_9,counterInput_8,counterInput_7,
            counterInput_6,counterInput_5,counterInput_4,counterInput_3,
            counterInput_2,counterInput_1,counterInput_0})) ;
    fake_vcc ix74 (.Y (PWR)) ;
    fake_gnd ix72 (.Y (GND)) ;
endmodule


module Reg_13 ( D, en, clk, rst, Q ) ;

    input [12:0]D ;
    input en ;
    input clk ;
    input rst ;
    output [12:0]Q ;

    wire nx192, nx202, nx212, nx222, nx232, nx242, nx252, nx262, nx272, nx282, 
         nx292, nx302, nx312, nx366, nx368, nx370, nx372;
    wire [12:0] \$dummy ;




    dffr reg_Q_0 (.Q (Q[0]), .QB (\$dummy [0]), .D (nx192), .CLK (nx370), .R (
         rst)) ;
    mux21_ni ix193 (.Y (nx192), .A0 (Q[0]), .A1 (D[0]), .S0 (nx366)) ;
    dffr reg_Q_1 (.Q (Q[1]), .QB (\$dummy [1]), .D (nx202), .CLK (nx370), .R (
         rst)) ;
    mux21_ni ix203 (.Y (nx202), .A0 (Q[1]), .A1 (D[1]), .S0 (nx366)) ;
    dffr reg_Q_2 (.Q (Q[2]), .QB (\$dummy [2]), .D (nx212), .CLK (nx370), .R (
         rst)) ;
    mux21_ni ix213 (.Y (nx212), .A0 (Q[2]), .A1 (D[2]), .S0 (nx366)) ;
    dffr reg_Q_3 (.Q (Q[3]), .QB (\$dummy [3]), .D (nx222), .CLK (nx370), .R (
         rst)) ;
    mux21_ni ix223 (.Y (nx222), .A0 (Q[3]), .A1 (D[3]), .S0 (nx366)) ;
    dffr reg_Q_4 (.Q (Q[4]), .QB (\$dummy [4]), .D (nx232), .CLK (nx370), .R (
         rst)) ;
    mux21_ni ix233 (.Y (nx232), .A0 (Q[4]), .A1 (D[4]), .S0 (nx366)) ;
    dffr reg_Q_5 (.Q (Q[5]), .QB (\$dummy [5]), .D (nx242), .CLK (nx370), .R (
         rst)) ;
    mux21_ni ix243 (.Y (nx242), .A0 (Q[5]), .A1 (D[5]), .S0 (nx366)) ;
    dffr reg_Q_6 (.Q (Q[6]), .QB (\$dummy [6]), .D (nx252), .CLK (nx370), .R (
         rst)) ;
    mux21_ni ix253 (.Y (nx252), .A0 (Q[6]), .A1 (D[6]), .S0 (nx366)) ;
    dffr reg_Q_7 (.Q (Q[7]), .QB (\$dummy [7]), .D (nx262), .CLK (nx372), .R (
         rst)) ;
    mux21_ni ix263 (.Y (nx262), .A0 (Q[7]), .A1 (D[7]), .S0 (nx368)) ;
    dffr reg_Q_8 (.Q (Q[8]), .QB (\$dummy [8]), .D (nx272), .CLK (nx372), .R (
         rst)) ;
    mux21_ni ix273 (.Y (nx272), .A0 (Q[8]), .A1 (D[8]), .S0 (nx368)) ;
    dffr reg_Q_9 (.Q (Q[9]), .QB (\$dummy [9]), .D (nx282), .CLK (nx372), .R (
         rst)) ;
    mux21_ni ix283 (.Y (nx282), .A0 (Q[9]), .A1 (D[9]), .S0 (nx368)) ;
    dffr reg_Q_10 (.Q (Q[10]), .QB (\$dummy [10]), .D (nx292), .CLK (nx372), .R (
         rst)) ;
    mux21_ni ix293 (.Y (nx292), .A0 (Q[10]), .A1 (D[10]), .S0 (nx368)) ;
    dffr reg_Q_11 (.Q (Q[11]), .QB (\$dummy [11]), .D (nx302), .CLK (nx372), .R (
         rst)) ;
    mux21_ni ix303 (.Y (nx302), .A0 (Q[11]), .A1 (D[11]), .S0 (nx368)) ;
    dffr reg_Q_12 (.Q (Q[12]), .QB (\$dummy [12]), .D (nx312), .CLK (nx372), .R (
         rst)) ;
    mux21_ni ix313 (.Y (nx312), .A0 (Q[12]), .A1 (D[12]), .S0 (nx368)) ;
    buf02 ix365 (.Y (nx366), .A (en)) ;
    buf02 ix367 (.Y (nx368), .A (en)) ;
    buf02 ix369 (.Y (nx370), .A (clk)) ;
    buf02 ix371 (.Y (nx372), .A (clk)) ;
endmodule


module Tristate_16 ( \input , en, \output  ) ;

    input [15:0]\input  ;
    input en ;
    output [15:0]\output  ;

    wire nx183, nx186, nx189, nx192, nx195, nx198, nx201, nx204, nx207, nx210, 
         nx213, nx216, nx219, nx222, nx225, nx228, nx235, nx237, nx239, nx241;



    tri01 tri_output_0 (.Y (\output [0]), .A (nx183), .E (nx237)) ;
    inv01 ix184 (.Y (nx183), .A (\input [0])) ;
    tri01 tri_output_1 (.Y (\output [1]), .A (nx186), .E (nx237)) ;
    inv01 ix187 (.Y (nx186), .A (\input [1])) ;
    tri01 tri_output_2 (.Y (\output [2]), .A (nx189), .E (nx237)) ;
    inv01 ix190 (.Y (nx189), .A (\input [2])) ;
    tri01 tri_output_3 (.Y (\output [3]), .A (nx192), .E (nx237)) ;
    inv01 ix193 (.Y (nx192), .A (\input [3])) ;
    tri01 tri_output_4 (.Y (\output [4]), .A (nx195), .E (nx237)) ;
    inv01 ix196 (.Y (nx195), .A (\input [4])) ;
    tri01 tri_output_5 (.Y (\output [5]), .A (nx198), .E (nx237)) ;
    inv01 ix199 (.Y (nx198), .A (\input [5])) ;
    tri01 tri_output_6 (.Y (\output [6]), .A (nx201), .E (nx237)) ;
    inv01 ix202 (.Y (nx201), .A (\input [6])) ;
    tri01 tri_output_7 (.Y (\output [7]), .A (nx204), .E (nx239)) ;
    inv01 ix205 (.Y (nx204), .A (\input [7])) ;
    tri01 tri_output_8 (.Y (\output [8]), .A (nx207), .E (nx239)) ;
    inv01 ix208 (.Y (nx207), .A (\input [8])) ;
    tri01 tri_output_9 (.Y (\output [9]), .A (nx210), .E (nx239)) ;
    inv01 ix211 (.Y (nx210), .A (\input [9])) ;
    tri01 tri_output_10 (.Y (\output [10]), .A (nx213), .E (nx239)) ;
    inv01 ix214 (.Y (nx213), .A (\input [10])) ;
    tri01 tri_output_11 (.Y (\output [11]), .A (nx216), .E (nx239)) ;
    inv01 ix217 (.Y (nx216), .A (\input [11])) ;
    tri01 tri_output_12 (.Y (\output [12]), .A (nx219), .E (nx239)) ;
    inv01 ix220 (.Y (nx219), .A (\input [12])) ;
    tri01 tri_output_13 (.Y (\output [13]), .A (nx222), .E (nx239)) ;
    inv01 ix223 (.Y (nx222), .A (\input [13])) ;
    tri01 tri_output_14 (.Y (\output [14]), .A (nx225), .E (nx241)) ;
    inv01 ix226 (.Y (nx225), .A (\input [14])) ;
    tri01 tri_output_15 (.Y (\output [15]), .A (nx228), .E (nx241)) ;
    inv01 ix229 (.Y (nx228), .A (\input [15])) ;
    inv01 ix234 (.Y (nx235), .A (en)) ;
    inv01 ix236 (.Y (nx237), .A (nx235)) ;
    inv01 ix238 (.Y (nx239), .A (nx235)) ;
    inv01 ix240 (.Y (nx241), .A (nx235)) ;
endmodule


module Tristate_80 ( \input , en, \output  ) ;

    input [79:0]\input  ;
    input en ;
    output [79:0]\output  ;

    wire nx695, nx698, nx701, nx704, nx707, nx710, nx713, nx716, nx719, nx722, 
         nx725, nx728, nx731, nx734, nx737, nx740, nx743, nx746, nx749, nx752, 
         nx755, nx758, nx761, nx764, nx767, nx770, nx773, nx776, nx779, nx782, 
         nx785, nx788, nx791, nx794, nx797, nx800, nx803, nx806, nx809, nx812, 
         nx815, nx818, nx821, nx824, nx827, nx830, nx833, nx836, nx839, nx842, 
         nx845, nx848, nx851, nx854, nx857, nx860, nx863, nx866, nx869, nx872, 
         nx875, nx878, nx881, nx884, nx887, nx890, nx893, nx896, nx899, nx902, 
         nx905, nx908, nx911, nx914, nx917, nx920, nx923, nx926, nx929, nx932, 
         nx939, nx941, nx943, nx945, nx947, nx949, nx951, nx953, nx955, nx957, 
         nx959, nx961, nx963, nx965;



    tri01 tri_output_0 (.Y (\output [0]), .A (nx695), .E (nx941)) ;
    inv01 ix696 (.Y (nx695), .A (\input [0])) ;
    tri01 tri_output_1 (.Y (\output [1]), .A (nx698), .E (nx941)) ;
    inv01 ix699 (.Y (nx698), .A (\input [1])) ;
    tri01 tri_output_2 (.Y (\output [2]), .A (nx701), .E (nx941)) ;
    inv01 ix702 (.Y (nx701), .A (\input [2])) ;
    tri01 tri_output_3 (.Y (\output [3]), .A (nx704), .E (nx941)) ;
    inv01 ix705 (.Y (nx704), .A (\input [3])) ;
    tri01 tri_output_4 (.Y (\output [4]), .A (nx707), .E (nx941)) ;
    inv01 ix708 (.Y (nx707), .A (\input [4])) ;
    tri01 tri_output_5 (.Y (\output [5]), .A (nx710), .E (nx941)) ;
    inv01 ix711 (.Y (nx710), .A (\input [5])) ;
    tri01 tri_output_6 (.Y (\output [6]), .A (nx713), .E (nx941)) ;
    inv01 ix714 (.Y (nx713), .A (\input [6])) ;
    tri01 tri_output_7 (.Y (\output [7]), .A (nx716), .E (nx943)) ;
    inv01 ix717 (.Y (nx716), .A (\input [7])) ;
    tri01 tri_output_8 (.Y (\output [8]), .A (nx719), .E (nx943)) ;
    inv01 ix720 (.Y (nx719), .A (\input [8])) ;
    tri01 tri_output_9 (.Y (\output [9]), .A (nx722), .E (nx943)) ;
    inv01 ix723 (.Y (nx722), .A (\input [9])) ;
    tri01 tri_output_10 (.Y (\output [10]), .A (nx725), .E (nx943)) ;
    inv01 ix726 (.Y (nx725), .A (\input [10])) ;
    tri01 tri_output_11 (.Y (\output [11]), .A (nx728), .E (nx943)) ;
    inv01 ix729 (.Y (nx728), .A (\input [11])) ;
    tri01 tri_output_12 (.Y (\output [12]), .A (nx731), .E (nx943)) ;
    inv01 ix732 (.Y (nx731), .A (\input [12])) ;
    tri01 tri_output_13 (.Y (\output [13]), .A (nx734), .E (nx943)) ;
    inv01 ix735 (.Y (nx734), .A (\input [13])) ;
    tri01 tri_output_14 (.Y (\output [14]), .A (nx737), .E (nx945)) ;
    inv01 ix738 (.Y (nx737), .A (\input [14])) ;
    tri01 tri_output_15 (.Y (\output [15]), .A (nx740), .E (nx945)) ;
    inv01 ix741 (.Y (nx740), .A (\input [15])) ;
    tri01 tri_output_16 (.Y (\output [16]), .A (nx743), .E (nx945)) ;
    inv01 ix744 (.Y (nx743), .A (\input [16])) ;
    tri01 tri_output_17 (.Y (\output [17]), .A (nx746), .E (nx945)) ;
    inv01 ix747 (.Y (nx746), .A (\input [17])) ;
    tri01 tri_output_18 (.Y (\output [18]), .A (nx749), .E (nx945)) ;
    inv01 ix750 (.Y (nx749), .A (\input [18])) ;
    tri01 tri_output_19 (.Y (\output [19]), .A (nx752), .E (nx945)) ;
    inv01 ix753 (.Y (nx752), .A (\input [19])) ;
    tri01 tri_output_20 (.Y (\output [20]), .A (nx755), .E (nx945)) ;
    inv01 ix756 (.Y (nx755), .A (\input [20])) ;
    tri01 tri_output_21 (.Y (\output [21]), .A (nx758), .E (nx947)) ;
    inv01 ix759 (.Y (nx758), .A (\input [21])) ;
    tri01 tri_output_22 (.Y (\output [22]), .A (nx761), .E (nx947)) ;
    inv01 ix762 (.Y (nx761), .A (\input [22])) ;
    tri01 tri_output_23 (.Y (\output [23]), .A (nx764), .E (nx947)) ;
    inv01 ix765 (.Y (nx764), .A (\input [23])) ;
    tri01 tri_output_24 (.Y (\output [24]), .A (nx767), .E (nx947)) ;
    inv01 ix768 (.Y (nx767), .A (\input [24])) ;
    tri01 tri_output_25 (.Y (\output [25]), .A (nx770), .E (nx947)) ;
    inv01 ix771 (.Y (nx770), .A (\input [25])) ;
    tri01 tri_output_26 (.Y (\output [26]), .A (nx773), .E (nx947)) ;
    inv01 ix774 (.Y (nx773), .A (\input [26])) ;
    tri01 tri_output_27 (.Y (\output [27]), .A (nx776), .E (nx947)) ;
    inv01 ix777 (.Y (nx776), .A (\input [27])) ;
    tri01 tri_output_28 (.Y (\output [28]), .A (nx779), .E (nx949)) ;
    inv01 ix780 (.Y (nx779), .A (\input [28])) ;
    tri01 tri_output_29 (.Y (\output [29]), .A (nx782), .E (nx949)) ;
    inv01 ix783 (.Y (nx782), .A (\input [29])) ;
    tri01 tri_output_30 (.Y (\output [30]), .A (nx785), .E (nx949)) ;
    inv01 ix786 (.Y (nx785), .A (\input [30])) ;
    tri01 tri_output_31 (.Y (\output [31]), .A (nx788), .E (nx949)) ;
    inv01 ix789 (.Y (nx788), .A (\input [31])) ;
    tri01 tri_output_32 (.Y (\output [32]), .A (nx791), .E (nx949)) ;
    inv01 ix792 (.Y (nx791), .A (\input [32])) ;
    tri01 tri_output_33 (.Y (\output [33]), .A (nx794), .E (nx949)) ;
    inv01 ix795 (.Y (nx794), .A (\input [33])) ;
    tri01 tri_output_34 (.Y (\output [34]), .A (nx797), .E (nx949)) ;
    inv01 ix798 (.Y (nx797), .A (\input [34])) ;
    tri01 tri_output_35 (.Y (\output [35]), .A (nx800), .E (nx951)) ;
    inv01 ix801 (.Y (nx800), .A (\input [35])) ;
    tri01 tri_output_36 (.Y (\output [36]), .A (nx803), .E (nx951)) ;
    inv01 ix804 (.Y (nx803), .A (\input [36])) ;
    tri01 tri_output_37 (.Y (\output [37]), .A (nx806), .E (nx951)) ;
    inv01 ix807 (.Y (nx806), .A (\input [37])) ;
    tri01 tri_output_38 (.Y (\output [38]), .A (nx809), .E (nx951)) ;
    inv01 ix810 (.Y (nx809), .A (\input [38])) ;
    tri01 tri_output_39 (.Y (\output [39]), .A (nx812), .E (nx951)) ;
    inv01 ix813 (.Y (nx812), .A (\input [39])) ;
    tri01 tri_output_40 (.Y (\output [40]), .A (nx815), .E (nx951)) ;
    inv01 ix816 (.Y (nx815), .A (\input [40])) ;
    tri01 tri_output_41 (.Y (\output [41]), .A (nx818), .E (nx951)) ;
    inv01 ix819 (.Y (nx818), .A (\input [41])) ;
    tri01 tri_output_42 (.Y (\output [42]), .A (nx821), .E (nx953)) ;
    inv01 ix822 (.Y (nx821), .A (\input [42])) ;
    tri01 tri_output_43 (.Y (\output [43]), .A (nx824), .E (nx953)) ;
    inv01 ix825 (.Y (nx824), .A (\input [43])) ;
    tri01 tri_output_44 (.Y (\output [44]), .A (nx827), .E (nx953)) ;
    inv01 ix828 (.Y (nx827), .A (\input [44])) ;
    tri01 tri_output_45 (.Y (\output [45]), .A (nx830), .E (nx953)) ;
    inv01 ix831 (.Y (nx830), .A (\input [45])) ;
    tri01 tri_output_46 (.Y (\output [46]), .A (nx833), .E (nx953)) ;
    inv01 ix834 (.Y (nx833), .A (\input [46])) ;
    tri01 tri_output_47 (.Y (\output [47]), .A (nx836), .E (nx953)) ;
    inv01 ix837 (.Y (nx836), .A (\input [47])) ;
    tri01 tri_output_48 (.Y (\output [48]), .A (nx839), .E (nx953)) ;
    inv01 ix840 (.Y (nx839), .A (\input [48])) ;
    tri01 tri_output_49 (.Y (\output [49]), .A (nx842), .E (nx955)) ;
    inv01 ix843 (.Y (nx842), .A (\input [49])) ;
    tri01 tri_output_50 (.Y (\output [50]), .A (nx845), .E (nx955)) ;
    inv01 ix846 (.Y (nx845), .A (\input [50])) ;
    tri01 tri_output_51 (.Y (\output [51]), .A (nx848), .E (nx955)) ;
    inv01 ix849 (.Y (nx848), .A (\input [51])) ;
    tri01 tri_output_52 (.Y (\output [52]), .A (nx851), .E (nx955)) ;
    inv01 ix852 (.Y (nx851), .A (\input [52])) ;
    tri01 tri_output_53 (.Y (\output [53]), .A (nx854), .E (nx955)) ;
    inv01 ix855 (.Y (nx854), .A (\input [53])) ;
    tri01 tri_output_54 (.Y (\output [54]), .A (nx857), .E (nx955)) ;
    inv01 ix858 (.Y (nx857), .A (\input [54])) ;
    tri01 tri_output_55 (.Y (\output [55]), .A (nx860), .E (nx955)) ;
    inv01 ix861 (.Y (nx860), .A (\input [55])) ;
    tri01 tri_output_56 (.Y (\output [56]), .A (nx863), .E (nx957)) ;
    inv01 ix864 (.Y (nx863), .A (\input [56])) ;
    tri01 tri_output_57 (.Y (\output [57]), .A (nx866), .E (nx957)) ;
    inv01 ix867 (.Y (nx866), .A (\input [57])) ;
    tri01 tri_output_58 (.Y (\output [58]), .A (nx869), .E (nx957)) ;
    inv01 ix870 (.Y (nx869), .A (\input [58])) ;
    tri01 tri_output_59 (.Y (\output [59]), .A (nx872), .E (nx957)) ;
    inv01 ix873 (.Y (nx872), .A (\input [59])) ;
    tri01 tri_output_60 (.Y (\output [60]), .A (nx875), .E (nx957)) ;
    inv01 ix876 (.Y (nx875), .A (\input [60])) ;
    tri01 tri_output_61 (.Y (\output [61]), .A (nx878), .E (nx957)) ;
    inv01 ix879 (.Y (nx878), .A (\input [61])) ;
    tri01 tri_output_62 (.Y (\output [62]), .A (nx881), .E (nx957)) ;
    inv01 ix882 (.Y (nx881), .A (\input [62])) ;
    tri01 tri_output_63 (.Y (\output [63]), .A (nx884), .E (nx959)) ;
    inv01 ix885 (.Y (nx884), .A (\input [63])) ;
    tri01 tri_output_64 (.Y (\output [64]), .A (nx887), .E (nx959)) ;
    inv01 ix888 (.Y (nx887), .A (\input [64])) ;
    tri01 tri_output_65 (.Y (\output [65]), .A (nx890), .E (nx959)) ;
    inv01 ix891 (.Y (nx890), .A (\input [65])) ;
    tri01 tri_output_66 (.Y (\output [66]), .A (nx893), .E (nx959)) ;
    inv01 ix894 (.Y (nx893), .A (\input [66])) ;
    tri01 tri_output_67 (.Y (\output [67]), .A (nx896), .E (nx959)) ;
    inv01 ix897 (.Y (nx896), .A (\input [67])) ;
    tri01 tri_output_68 (.Y (\output [68]), .A (nx899), .E (nx959)) ;
    inv01 ix900 (.Y (nx899), .A (\input [68])) ;
    tri01 tri_output_69 (.Y (\output [69]), .A (nx902), .E (nx959)) ;
    inv01 ix903 (.Y (nx902), .A (\input [69])) ;
    tri01 tri_output_70 (.Y (\output [70]), .A (nx905), .E (nx961)) ;
    inv01 ix906 (.Y (nx905), .A (\input [70])) ;
    tri01 tri_output_71 (.Y (\output [71]), .A (nx908), .E (nx961)) ;
    inv01 ix909 (.Y (nx908), .A (\input [71])) ;
    tri01 tri_output_72 (.Y (\output [72]), .A (nx911), .E (nx961)) ;
    inv01 ix912 (.Y (nx911), .A (\input [72])) ;
    tri01 tri_output_73 (.Y (\output [73]), .A (nx914), .E (nx961)) ;
    inv01 ix915 (.Y (nx914), .A (\input [73])) ;
    tri01 tri_output_74 (.Y (\output [74]), .A (nx917), .E (nx961)) ;
    inv01 ix918 (.Y (nx917), .A (\input [74])) ;
    tri01 tri_output_75 (.Y (\output [75]), .A (nx920), .E (nx961)) ;
    inv01 ix921 (.Y (nx920), .A (\input [75])) ;
    tri01 tri_output_76 (.Y (\output [76]), .A (nx923), .E (nx961)) ;
    inv01 ix924 (.Y (nx923), .A (\input [76])) ;
    tri01 tri_output_77 (.Y (\output [77]), .A (nx926), .E (nx963)) ;
    inv01 ix927 (.Y (nx926), .A (\input [77])) ;
    tri01 tri_output_78 (.Y (\output [78]), .A (nx929), .E (nx963)) ;
    inv01 ix930 (.Y (nx929), .A (\input [78])) ;
    tri01 tri_output_79 (.Y (\output [79]), .A (nx932), .E (nx963)) ;
    inv01 ix933 (.Y (nx932), .A (\input [79])) ;
    inv01 ix938 (.Y (nx939), .A (en)) ;
    inv01 ix940 (.Y (nx941), .A (nx965)) ;
    inv01 ix942 (.Y (nx943), .A (nx965)) ;
    inv01 ix944 (.Y (nx945), .A (nx965)) ;
    inv01 ix946 (.Y (nx947), .A (nx965)) ;
    inv01 ix948 (.Y (nx949), .A (nx965)) ;
    inv01 ix950 (.Y (nx951), .A (nx965)) ;
    inv01 ix952 (.Y (nx953), .A (nx965)) ;
    inv01 ix954 (.Y (nx955), .A (nx939)) ;
    inv01 ix956 (.Y (nx957), .A (nx939)) ;
    inv01 ix958 (.Y (nx959), .A (nx939)) ;
    inv01 ix960 (.Y (nx961), .A (nx939)) ;
    inv01 ix962 (.Y (nx963), .A (nx939)) ;
    inv01 ix964 (.Y (nx965), .A (en)) ;
endmodule


module Mux2_13 ( A, B, S, C ) ;

    input [12:0]A ;
    input [12:0]B ;
    input S ;
    output [12:0]C ;

    wire nx152, nx154;



    mux21_ni ix7 (.Y (C[0]), .A0 (A[0]), .A1 (B[0]), .S0 (nx152)) ;
    mux21_ni ix15 (.Y (C[1]), .A0 (A[1]), .A1 (B[1]), .S0 (nx152)) ;
    mux21_ni ix23 (.Y (C[2]), .A0 (A[2]), .A1 (B[2]), .S0 (nx152)) ;
    mux21_ni ix31 (.Y (C[3]), .A0 (A[3]), .A1 (B[3]), .S0 (nx152)) ;
    mux21_ni ix39 (.Y (C[4]), .A0 (A[4]), .A1 (B[4]), .S0 (nx152)) ;
    mux21_ni ix47 (.Y (C[5]), .A0 (A[5]), .A1 (B[5]), .S0 (nx152)) ;
    mux21_ni ix55 (.Y (C[6]), .A0 (A[6]), .A1 (B[6]), .S0 (nx152)) ;
    mux21_ni ix63 (.Y (C[7]), .A0 (A[7]), .A1 (B[7]), .S0 (nx154)) ;
    mux21_ni ix71 (.Y (C[8]), .A0 (A[8]), .A1 (B[8]), .S0 (nx154)) ;
    mux21_ni ix79 (.Y (C[9]), .A0 (A[9]), .A1 (B[9]), .S0 (nx154)) ;
    mux21_ni ix87 (.Y (C[10]), .A0 (A[10]), .A1 (B[10]), .S0 (nx154)) ;
    mux21_ni ix95 (.Y (C[11]), .A0 (A[11]), .A1 (B[11]), .S0 (nx154)) ;
    mux21_ni ix103 (.Y (C[12]), .A0 (A[12]), .A1 (B[12]), .S0 (nx154)) ;
    buf02 ix151 (.Y (nx152), .A (S)) ;
    buf02 ix153 (.Y (nx154), .A (S)) ;
endmodule


module NBitAdder_13 ( a, b, carryIn, sum, carryOut ) ;

    input [12:0]a ;
    input [12:0]b ;
    input carryIn ;
    output [12:0]sum ;
    output carryOut ;

    wire temp_11, temp_10, temp_9, temp_8, temp_7, temp_6, temp_5, temp_4, 
         temp_3, temp_2, temp_1, temp_0;



    FullAdder f0 (.a (a[0]), .b (b[0]), .cin (carryIn), .s (sum[0]), .cout (
              temp_0)) ;
    FullAdder loop1_1_fx (.a (a[1]), .b (b[1]), .cin (temp_0), .s (sum[1]), .cout (
              temp_1)) ;
    FullAdder loop1_2_fx (.a (a[2]), .b (b[2]), .cin (temp_1), .s (sum[2]), .cout (
              temp_2)) ;
    FullAdder loop1_3_fx (.a (a[3]), .b (b[3]), .cin (temp_2), .s (sum[3]), .cout (
              temp_3)) ;
    FullAdder loop1_4_fx (.a (a[4]), .b (b[4]), .cin (temp_3), .s (sum[4]), .cout (
              temp_4)) ;
    FullAdder loop1_5_fx (.a (a[5]), .b (b[5]), .cin (temp_4), .s (sum[5]), .cout (
              temp_5)) ;
    FullAdder loop1_6_fx (.a (a[6]), .b (b[6]), .cin (temp_5), .s (sum[6]), .cout (
              temp_6)) ;
    FullAdder loop1_7_fx (.a (a[7]), .b (b[7]), .cin (temp_6), .s (sum[7]), .cout (
              temp_7)) ;
    FullAdder loop1_8_fx (.a (a[8]), .b (b[8]), .cin (temp_7), .s (sum[8]), .cout (
              temp_8)) ;
    FullAdder loop1_9_fx (.a (a[9]), .b (b[9]), .cin (temp_8), .s (sum[9]), .cout (
              temp_9)) ;
    FullAdder loop1_10_fx (.a (a[10]), .b (b[10]), .cin (temp_9), .s (sum[10]), 
              .cout (temp_10)) ;
    FullAdder loop1_11_fx (.a (a[11]), .b (b[11]), .cin (temp_10), .s (sum[11])
              , .cout (temp_11)) ;
    FullAdder loop1_12_fx (.a (a[12]), .b (b[12]), .cin (temp_11), .s (sum[12])
              , .cout (carryOut)) ;
endmodule


module ControlUnit ( clk, layersNumber, filtersNumber, filterDepth, 
                     filterOutputSize, startNetwork, layerType, convFinish, 
                     dmaAFinish, dmaBFinish, dmaCFinish, resetNetwork, 
                     loadLayerConfig, loadNetworkConfig, loadFilterConfig, 
                     loadWindow, loadFilter, conv, pool, shift12, shift21, 
                     readNextCol, addToOutputBuffer, outputBufferEn, saveToRAM, 
                     currentPage, finishCurrentSlice, finishFilter, 
                     finishOneLayer, finishNetwork ) ;

    input clk ;
    input [1:0]layersNumber ;
    input [2:0]filtersNumber ;
    input [2:0]filterDepth ;
    input [4:0]filterOutputSize ;
    input startNetwork ;
    input layerType ;
    input convFinish ;
    input dmaAFinish ;
    input dmaBFinish ;
    input dmaCFinish ;
    input resetNetwork ;
    output loadLayerConfig ;
    output loadNetworkConfig ;
    output loadFilterConfig ;
    output loadWindow ;
    output loadFilter ;
    output conv ;
    output pool ;
    output shift12 ;
    output shift21 ;
    output readNextCol ;
    output addToOutputBuffer ;
    output outputBufferEn ;
    output saveToRAM ;
    output [0:0]currentPage ;
    output finishCurrentSlice ;
    output finishFilter ;
    output finishOneLayer ;
    output finishNetwork ;

    wire startOneLayer, startFilter, filterLastLayer, startSlice, nx94, nx96;



    NetworkController_2 networkMap (.start (startNetwork), .dmaFinish (
                        dmaAFinish), .oneLayerFinish (finishOneLayer), .resetState (
                        resetNetwork), .clk (clk), .layersNumber ({
                        layersNumber[1],layersNumber[0]}), .loadConfig (
                        loadNetworkConfig), .startOneLayer (startOneLayer), .finish (
                        finishNetwork)) ;
    LayerController_3 oneLayerMap (.start (startOneLayer), .dmaFinish (
                      dmaAFinish), .filterFinish (finishFilter), .resetState (
                      resetNetwork), .clk (clk), .filtersNumber ({
                      filtersNumber[2],filtersNumber[1],filtersNumber[0]}), .loadConfig (
                      loadLayerConfig), .startFilterConv (startFilter), .finish (
                      finishOneLayer)) ;
    FilterController_3 filterMap (.start (startFilter), .layerType (nx94), .dmaFinish (
                       dmaAFinish), .oneConvFinish (finishCurrentSlice), .resetState (
                       resetNetwork), .clk (clk), .depth ({filterDepth[2],
                       filterDepth[1],filterDepth[0]}), .startOneConv (
                       startSlice), .loadConfig (loadFilterConfig), .filterLastLayer (
                       filterLastLayer), .finish (finishFilter)) ;
    SliceFilterController_5 sliceFilterMap (.start (startSlice), .layerType (
                            nx96), .filterLastLayer (filterLastLayer), .finishConv (
                            convFinish), .dmaAFinish (dmaAFinish), .dmaBFinish (
                            dmaBFinish), .dmaCFinish (dmaCFinish), .resetState (
                            resetNetwork), .clk (clk), .outputSize ({
                            filterOutputSize[4],filterOutputSize[3],
                            filterOutputSize[2],filterOutputSize[1],
                            filterOutputSize[0]}), .pageTurn ({currentPage[0]})
                            , .loadFilter (loadFilter), .loadWindow (loadWindow)
                            , .conv (conv), .pool (pool), .shift12 (shift12), .shift21 (
                            shift21), .readNextCol (readNextCol), .addToOutputBuffer (
                            addToOutputBuffer), .outputBufferEn (outputBufferEn)
                            , .saveToRAM (saveToRAM), .finish (
                            finishCurrentSlice)) ;
    buf02 ix93 (.Y (nx94), .A (layerType)) ;
    buf02 ix95 (.Y (nx96), .A (layerType)) ;
endmodule


module SliceFilterController_5 ( start, layerType, filterLastLayer, finishConv, 
                                 dmaAFinish, dmaBFinish, dmaCFinish, resetState, 
                                 clk, outputSize, pageTurn, loadFilter, 
                                 loadWindow, conv, pool, shift12, shift21, 
                                 readNextCol, addToOutputBuffer, outputBufferEn, 
                                 saveToRAM, finish ) ;

    input start ;
    input layerType ;
    input filterLastLayer ;
    input finishConv ;
    input dmaAFinish ;
    input dmaBFinish ;
    input dmaCFinish ;
    input resetState ;
    input clk ;
    input [4:0]outputSize ;
    output [0:0]pageTurn ;
    output loadFilter ;
    output loadWindow ;
    output conv ;
    output pool ;
    output shift12 ;
    output shift21 ;
    output readNextCol ;
    output addToOutputBuffer ;
    output outputBufferEn ;
    output saveToRAM ;
    output finish ;

    wire currentState_0, outerCounterEn, altInnerCounterOut_4, 
         altInnerCounterOut_3, altInnerCounterOut_2, altInnerCounterOut_1, 
         altInnerCounterOut_0, altOuterCounterOut_4, altOuterCounterOut_3, 
         altOuterCounterOut_2, altOuterCounterOut_1, altOuterCounterOut_0, 
         innerCounterEn, currentState_1, currentState_3, nx603, NOT_clk, 
         currentState_2, outerCounterOut_1, outerCounterOut_4, outerCounterOut_0, 
         outerCounterOut_2, outerCounterOut_3, nx64, innerCounterOut_1, 
         innerCounterOut_4, innerCounterOut_0, innerCounterOut_2, 
         innerCounterOut_3, nx112, nx118, currentState_6, nx150, nx164, nx208, 
         nx212, NOT_pageTurn_0, nx608, nx618, nx628, nx640, nx650, nx660, nx670, 
         nx680, nx690, nx701, nx704, nx708, nx712, nx717, nx722, nx725, nx733, 
         nx735, nx739, nx743, nx747, nx751, nx756, nx758, nx762, nx766, nx770, 
         nx774, nx778, nx780, nx782, nx784, nx791, nx794, nx798, nx800, nx802, 
         nx805, nx807, nx809, nx811, nx813, nx816, nx824, nx830, nx835, nx837, 
         nx845, nx847;
    wire [15:0] \$dummy ;




    Counter_5 innerCounterMap (.en (innerCounterEn), .reset (outerCounterEn), .clk (
              clk), .count ({altInnerCounterOut_4,altInnerCounterOut_3,
              altInnerCounterOut_2,altInnerCounterOut_1,altInnerCounterOut_0})
              ) ;
    Counter_5 outerCounterMap (.en (outerCounterEn), .reset (nx845), .clk (clk)
              , .count ({altOuterCounterOut_4,altOuterCounterOut_3,
              altOuterCounterOut_2,altOuterCounterOut_1,altOuterCounterOut_0})
              ) ;
    Reg_1 pageRegMap (.D ({NOT_pageTurn_0}), .en (innerCounterEn), .clk (clk), .rst (
          nx845), .Q ({pageTurn[0]})) ;
    inv01 ix698 (.Y (NOT_pageTurn_0), .A (pageTurn[0])) ;
    aoi21 ix273 (.Y (conv), .A0 (nx701), .A1 (nx712), .B0 (layerType)) ;
    aoi21 ix705 (.Y (nx704), .A0 (outputBufferEn), .A1 (nx811), .B0 (
          currentState_1)) ;
    dffr reg_currentState_5 (.Q (outputBufferEn), .QB (\$dummy [0]), .D (nx618)
         , .CLK (NOT_clk), .R (resetState)) ;
    aoi21 ix709 (.Y (nx708), .A0 (layerType), .A1 (currentState_3), .B0 (
          addToOutputBuffer)) ;
    oai21 ix641 (.Y (nx640), .A0 (nx712), .A1 (nx603), .B0 (nx701)) ;
    dffr reg_currentState_3 (.Q (currentState_3), .QB (nx712), .D (nx640), .CLK (
         NOT_clk), .R (resetState)) ;
    inv02 ix715 (.Y (NOT_clk), .A (clk)) ;
    nand04 ix237 (.Y (nx603), .A0 (nx717), .A1 (nx725), .A2 (nx780), .A3 (nx784)
           ) ;
    nor03_2x ix718 (.Y (nx717), .A0 (currentState_2), .A1 (addToOutputBuffer), .A2 (
             outputBufferEn)) ;
    dffr reg_currentState_2 (.Q (currentState_2), .QB (nx701), .D (nx628), .CLK (
         NOT_clk), .R (resetState)) ;
    dffr reg_currentState_4 (.Q (addToOutputBuffer), .QB (\$dummy [1]), .D (
         nx608), .CLK (NOT_clk), .R (resetState)) ;
    nor03_2x ix609 (.Y (nx608), .A0 (layerType), .A1 (nx712), .A2 (nx722)) ;
    nand02 ix726 (.Y (nx725), .A0 (start), .A1 (nx845)) ;
    dffs_ni reg_currentState_0 (.Q (currentState_0), .QB (\$dummy [2]), .D (
            nx660), .CLK (NOT_clk), .S (resetState)) ;
    mux21_ni ix661 (.Y (nx660), .A0 (nx845), .A1 (currentState_6), .S0 (nx603)
             ) ;
    dffr reg_currentState_6 (.Q (currentState_6), .QB (nx778), .D (nx650), .CLK (
         NOT_clk), .R (resetState)) ;
    ao22 ix651 (.Y (nx650), .A0 (outputBufferEn), .A1 (nx118), .B0 (
         currentState_6), .B1 (nx722)) ;
    nor02_2x ix119 (.Y (nx118), .A0 (nx64), .A1 (nx112)) ;
    nand04 ix65 (.Y (nx64), .A0 (nx733), .A1 (nx743), .A2 (nx747), .A3 (nx751)
           ) ;
    and02 ix734 (.Y (nx733), .A0 (nx735), .A1 (nx739)) ;
    xnor2 ix736 (.Y (nx735), .A0 (outerCounterOut_3), .A1 (outputSize[3])) ;
    dff reg_outerCounterOut_3 (.Q (outerCounterOut_3), .QB (\$dummy [3]), .D (
        altOuterCounterOut_3), .CLK (clk)) ;
    xnor2 ix740 (.Y (nx739), .A0 (outerCounterOut_2), .A1 (outputSize[2])) ;
    dff reg_outerCounterOut_2 (.Q (outerCounterOut_2), .QB (\$dummy [4]), .D (
        altOuterCounterOut_2), .CLK (clk)) ;
    xnor2 ix744 (.Y (nx743), .A0 (outerCounterOut_0), .A1 (outputSize[0])) ;
    dff reg_outerCounterOut_0 (.Q (outerCounterOut_0), .QB (\$dummy [5]), .D (
        altOuterCounterOut_0), .CLK (clk)) ;
    xnor2 ix748 (.Y (nx747), .A0 (outerCounterOut_4), .A1 (outputSize[4])) ;
    dff reg_outerCounterOut_4 (.Q (outerCounterOut_4), .QB (\$dummy [6]), .D (
        altOuterCounterOut_4), .CLK (clk)) ;
    xnor2 ix752 (.Y (nx751), .A0 (outerCounterOut_1), .A1 (outputSize[1])) ;
    dff reg_outerCounterOut_1 (.Q (outerCounterOut_1), .QB (\$dummy [7]), .D (
        altOuterCounterOut_1), .CLK (clk)) ;
    nand04 ix113 (.Y (nx112), .A0 (nx756), .A1 (nx766), .A2 (nx770), .A3 (nx774)
           ) ;
    and02 ix757 (.Y (nx756), .A0 (nx758), .A1 (nx762)) ;
    xnor2 ix759 (.Y (nx758), .A0 (innerCounterOut_3), .A1 (outputSize[3])) ;
    dff reg_innerCounterOut_3 (.Q (innerCounterOut_3), .QB (\$dummy [8]), .D (
        altInnerCounterOut_3), .CLK (clk)) ;
    xnor2 ix763 (.Y (nx762), .A0 (innerCounterOut_2), .A1 (outputSize[2])) ;
    dff reg_innerCounterOut_2 (.Q (innerCounterOut_2), .QB (\$dummy [9]), .D (
        altInnerCounterOut_2), .CLK (clk)) ;
    xnor2 ix767 (.Y (nx766), .A0 (innerCounterOut_0), .A1 (outputSize[0])) ;
    dff reg_innerCounterOut_0 (.Q (innerCounterOut_0), .QB (\$dummy [10]), .D (
        altInnerCounterOut_0), .CLK (clk)) ;
    xnor2 ix771 (.Y (nx770), .A0 (innerCounterOut_4), .A1 (outputSize[4])) ;
    dff reg_innerCounterOut_4 (.Q (innerCounterOut_4), .QB (\$dummy [11]), .D (
        altInnerCounterOut_4), .CLK (clk)) ;
    xnor2 ix775 (.Y (nx774), .A0 (innerCounterOut_1), .A1 (outputSize[1])) ;
    dff reg_innerCounterOut_1 (.Q (innerCounterOut_1), .QB (\$dummy [12]), .D (
        altInnerCounterOut_1), .CLK (clk)) ;
    oai21 ix781 (.Y (nx780), .A0 (nx782), .A1 (dmaCFinish), .B0 (currentState_6)
          ) ;
    inv01 ix783 (.Y (nx782), .A (filterLastLayer)) ;
    aoi33 ix785 (.Y (nx784), .A0 (nx212), .A1 (dmaBFinish), .A2 (currentState_1)
          , .B0 (finishConv), .B1 (currentState_3), .B2 (nx208)) ;
    or02 ix213 (.Y (nx212), .A0 (layerType), .A1 (dmaAFinish)) ;
    dffr reg_currentState_1 (.Q (currentState_1), .QB (\$dummy [13]), .D (nx690)
         , .CLK (NOT_clk), .R (resetState)) ;
    mux21_ni ix691 (.Y (nx690), .A0 (currentState_1), .A1 (nx845), .S0 (nx603)
             ) ;
    aoi32 ix209 (.Y (nx208), .A0 (nx791), .A1 (filterLastLayer), .A2 (saveToRAM)
          , .B0 (nx811), .B1 (nx813)) ;
    dffr reg_finalDMACFinish (.Q (\$dummy [14]), .QB (nx791), .D (nx670), .CLK (
         clk), .R (nx164)) ;
    nand02 ix671 (.Y (nx670), .A0 (nx791), .A1 (nx794)) ;
    oai21 ix795 (.Y (nx794), .A0 (nx164), .A1 (currentState_3), .B0 (dmaCFinish)
          ) ;
    or02 ix165 (.Y (nx164), .A0 (nx845), .A1 (addToOutputBuffer)) ;
    aoi22 ix189 (.Y (saveToRAM), .A0 (nx798), .A1 (nx782), .B0 (nx800), .B1 (
          nx778)) ;
    inv01 ix799 (.Y (nx798), .A (layerType)) ;
    ao32 ix801 (.Y (nx800), .A0 (nx802), .A1 (nx805), .A2 (nx807), .B0 (nx809), 
         .B1 (nx701)) ;
    nor04 ix803 (.Y (nx802), .A0 (outerCounterOut_0), .A1 (outerCounterOut_1), .A2 (
          nx150), .A3 (outerCounterOut_2)) ;
    or02 ix151 (.Y (nx150), .A0 (outerCounterOut_3), .A1 (outerCounterOut_4)) ;
    nor02_2x ix806 (.Y (nx805), .A0 (innerCounterOut_0), .A1 (innerCounterOut_1)
             ) ;
    nor03_2x ix808 (.Y (nx807), .A0 (innerCounterOut_3), .A1 (innerCounterOut_4)
             , .A2 (innerCounterOut_2)) ;
    nand02 ix810 (.Y (nx809), .A0 (nx791), .A1 (currentState_3)) ;
    dffr reg_finalDMABFinish (.Q (\$dummy [15]), .QB (nx813), .D (nx680), .CLK (
         clk), .R (nx164)) ;
    nand02 ix681 (.Y (nx680), .A0 (nx813), .A1 (nx816)) ;
    oai21 ix817 (.Y (nx816), .A0 (nx164), .A1 (currentState_3), .B0 (dmaBFinish)
          ) ;
    aoi21 ix277 (.Y (pool), .A0 (nx701), .A1 (nx712), .B0 (nx798)) ;
    aoi21 ix831 (.Y (nx830), .A0 (nx782), .A1 (nx798), .B0 (dmaCFinish)) ;
    or02 ix301 (.Y (innerCounterEn), .A0 (nx845), .A1 (outputBufferEn)) ;
    ao21 ix255 (.Y (outerCounterEn), .A0 (outputBufferEn), .A1 (nx824), .B0 (
         nx847)) ;
    nand02 ix267 (.Y (loadWindow), .A0 (nx835), .A1 (nx837)) ;
    nand04 ix836 (.Y (nx835), .A0 (nx813), .A1 (currentState_3), .A2 (nx64), .A3 (
           nx824)) ;
    aoi21 ix838 (.Y (nx837), .A0 (start), .A1 (nx847), .B0 (currentState_1)) ;
    nor02_2x ix249 (.Y (loadFilter), .A0 (layerType), .A1 (nx837)) ;
    inv01 ix812 (.Y (nx811), .A (nx118)) ;
    inv01 ix825 (.Y (nx824), .A (nx112)) ;
    inv01 ix723 (.Y (nx722), .A (nx603)) ;
    buf02 ix844 (.Y (nx845), .A (currentState_0)) ;
    buf02 ix846 (.Y (nx847), .A (currentState_0)) ;
    nor02ii ix629 (.Y (nx628), .A0 (nx704), .A1 (nx603)) ;
    nor02ii ix619 (.Y (nx618), .A0 (nx708), .A1 (nx603)) ;
    nor02ii ix281 (.Y (shift12), .A0 (pageTurn[0]), .A1 (currentState_2)) ;
    nor02ii ix283 (.Y (shift21), .A0 (nx701), .A1 (pageTurn[0])) ;
    and03 ix289 (.Y (readNextCol), .A0 (nx112), .A1 (nx813), .A2 (currentState_3
          )) ;
    nor02ii ix299 (.Y (finish), .A0 (nx830), .A1 (currentState_6)) ;
endmodule


module Counter_5 ( en, reset, clk, count ) ;

    input en ;
    input reset ;
    input clk ;
    output [4:0]count ;

    wire addedOne_4, addedOne_3, addedOne_2, addedOne_1, addedOne_0, finalReset, 
         oneSignal_4, PWR;
    wire [0:0] \$dummy ;




    Reg_5 counterReg (.D ({addedOne_4,addedOne_3,addedOne_2,addedOne_1,
          addedOne_0}), .en (en), .clk (clk), .rst (finalReset), .Q ({count[4],
          count[3],count[2],count[1],count[0]})) ;
    NBitAdder_5 nextCount (.a ({count[4],count[3],count[2],count[1],count[0]}), 
                .b ({oneSignal_4,oneSignal_4,oneSignal_4,oneSignal_4,oneSignal_4
                }), .carryIn (PWR), .sum ({addedOne_4,addedOne_3,addedOne_2,
                addedOne_1,addedOne_0}), .carryOut (\$dummy [0])) ;
    fake_vcc ix21 (.Y (PWR)) ;
    fake_gnd ix19 (.Y (oneSignal_4)) ;
    and02 ix1 (.Y (finalReset), .A0 (reset), .A1 (clk)) ;
endmodule


module NBitAdder_5 ( a, b, carryIn, sum, carryOut ) ;

    input [4:0]a ;
    input [4:0]b ;
    input carryIn ;
    output [4:0]sum ;
    output carryOut ;

    wire temp_3, temp_2, temp_1, temp_0;



    FullAdder f0 (.a (a[0]), .b (b[0]), .cin (carryIn), .s (sum[0]), .cout (
              temp_0)) ;
    FullAdder loop1_1_fx (.a (a[1]), .b (b[1]), .cin (temp_0), .s (sum[1]), .cout (
              temp_1)) ;
    FullAdder loop1_2_fx (.a (a[2]), .b (b[2]), .cin (temp_1), .s (sum[2]), .cout (
              temp_2)) ;
    FullAdder loop1_3_fx (.a (a[3]), .b (b[3]), .cin (temp_2), .s (sum[3]), .cout (
              temp_3)) ;
    FullAdder loop1_4_fx (.a (a[4]), .b (b[4]), .cin (temp_3), .s (sum[4]), .cout (
              carryOut)) ;
endmodule


module Reg_5 ( D, en, clk, rst, Q ) ;

    input [4:0]D ;
    input en ;
    input clk ;
    input rst ;
    output [4:0]Q ;

    wire nx96, nx106, nx116, nx126, nx136, nx166;
    wire [4:0] \$dummy ;




    dffr reg_Q_0 (.Q (Q[0]), .QB (\$dummy [0]), .D (nx96), .CLK (clk), .R (rst)
         ) ;
    mux21_ni ix97 (.Y (nx96), .A0 (Q[0]), .A1 (D[0]), .S0 (nx166)) ;
    dffr reg_Q_1 (.Q (Q[1]), .QB (\$dummy [1]), .D (nx106), .CLK (clk), .R (rst)
         ) ;
    mux21_ni ix107 (.Y (nx106), .A0 (Q[1]), .A1 (D[1]), .S0 (nx166)) ;
    dffr reg_Q_2 (.Q (Q[2]), .QB (\$dummy [2]), .D (nx116), .CLK (clk), .R (rst)
         ) ;
    mux21_ni ix117 (.Y (nx116), .A0 (Q[2]), .A1 (D[2]), .S0 (nx166)) ;
    dffr reg_Q_3 (.Q (Q[3]), .QB (\$dummy [3]), .D (nx126), .CLK (clk), .R (rst)
         ) ;
    mux21_ni ix127 (.Y (nx126), .A0 (Q[3]), .A1 (D[3]), .S0 (nx166)) ;
    dffr reg_Q_4 (.Q (Q[4]), .QB (\$dummy [4]), .D (nx136), .CLK (clk), .R (rst)
         ) ;
    mux21_ni ix137 (.Y (nx136), .A0 (Q[4]), .A1 (D[4]), .S0 (nx166)) ;
    buf02 ix165 (.Y (nx166), .A (en)) ;
endmodule


module FilterController_3 ( start, layerType, dmaFinish, oneConvFinish, 
                            resetState, clk, depth, startOneConv, loadConfig, 
                            filterLastLayer, finish ) ;

    input start ;
    input layerType ;
    input dmaFinish ;
    input oneConvFinish ;
    input resetState ;
    input clk ;
    input [2:0]depth ;
    output startOneConv ;
    output loadConfig ;
    output filterLastLayer ;
    output finish ;

    wire counterEn, altCounterOut_2, altCounterOut_1, altCounterOut_0, 
         resetCounter, currentState_1, currentState_0, NOT_clk, nx12, 
         counterOut_2, counterOut_0, counterOut_1, nx76, nx86, nx161, nx171, 
         nx182, nx186, nx190, nx195, nx202, nx209, nx214, nx216, nx223;
    wire [2:0] \$dummy ;




    Counter_3 counterMap (.en (counterEn), .reset (resetCounter), .clk (clk), .count (
              {altCounterOut_2,altCounterOut_1,altCounterOut_0})) ;
    and04 ix65 (.Y (filterLastLayer), .A0 (nx182), .A1 (nx186), .A2 (nx190), .A3 (
          startOneConv)) ;
    xnor2 ix183 (.Y (nx182), .A0 (counterOut_2), .A1 (depth[2])) ;
    dff reg_counterOut_2 (.Q (counterOut_2), .QB (\$dummy [0]), .D (
        altCounterOut_2), .CLK (clk)) ;
    xnor2 ix187 (.Y (nx186), .A0 (counterOut_0), .A1 (depth[0])) ;
    dff reg_counterOut_0 (.Q (counterOut_0), .QB (\$dummy [1]), .D (
        altCounterOut_0), .CLK (clk)) ;
    xnor2 ix191 (.Y (nx190), .A0 (counterOut_1), .A1 (depth[1])) ;
    dff reg_counterOut_1 (.Q (counterOut_1), .QB (\$dummy [2]), .D (
        altCounterOut_1), .CLK (clk)) ;
    mux21_ni ix172 (.Y (nx171), .A0 (nx86), .A1 (currentState_1), .S0 (nx223)) ;
    oai22 ix87 (.Y (nx86), .A0 (nx12), .A1 (finish), .B0 (nx195), .B1 (
          currentState_0)) ;
    aoi21 ix13 (.Y (nx12), .A0 (layerType), .A1 (nx195), .B0 (currentState_0)) ;
    mux21_ni ix162 (.Y (nx161), .A0 (nx12), .A1 (currentState_0), .S0 (nx223)) ;
    aoi221 ix203 (.Y (nx202), .A0 (start), .A1 (resetCounter), .B0 (counterEn), 
           .B1 (filterLastLayer), .C0 (nx76)) ;
    dffr reg_currentState_1 (.Q (currentState_1), .QB (nx195), .D (nx171), .CLK (
         NOT_clk), .R (resetState)) ;
    inv01 ix207 (.Y (NOT_clk), .A (clk)) ;
    ao21 ix29 (.Y (counterEn), .A0 (oneConvFinish), .A1 (nx209), .B0 (
         resetCounter)) ;
    dffr reg_currentState_0 (.Q (currentState_0), .QB (nx209), .D (nx161), .CLK (
         NOT_clk), .R (resetState)) ;
    ao21 ix77 (.Y (nx76), .A0 (dmaFinish), .A1 (currentState_0), .B0 (finish)) ;
    aoi21 ix215 (.Y (nx214), .A0 (start), .A1 (nx216), .B0 (currentState_0)) ;
    inv01 ix217 (.Y (nx216), .A (layerType)) ;
    buf02 ix222 (.Y (nx223), .A (nx202)) ;
    and02 ix5 (.Y (startOneConv), .A0 (currentState_1), .A1 (nx209)) ;
    and02 ix23 (.Y (resetCounter), .A0 (nx195), .A1 (nx209)) ;
    and02 ix73 (.Y (finish), .A0 (currentState_1), .A1 (currentState_0)) ;
    nor02ii ix101 (.Y (loadConfig), .A0 (nx214), .A1 (nx195)) ;
endmodule


module LayerController_3 ( start, dmaFinish, filterFinish, resetState, clk, 
                           filtersNumber, loadConfig, startFilterConv, finish
                            ) ;

    input start ;
    input dmaFinish ;
    input filterFinish ;
    input resetState ;
    input clk ;
    input [2:0]filtersNumber ;
    output loadConfig ;
    output startFilterConv ;
    output finish ;

    wire counterEn, altCounterOut_2, altCounterOut_1, altCounterOut_0, 
         resetCounter, currentState_1, currentState_0, nx123, NOT_clk, 
         counterOut_2, counterOut_0, counterOut_1, nx58, nx78, nx130, nx140, 
         nx151, nx163, nx165, nx168, nx172, nx176, nx182, nx185;
    wire [2:0] \$dummy ;




    Counter_3 counterMap (.en (counterEn), .reset (resetCounter), .clk (clk), .count (
              {altCounterOut_2,altCounterOut_1,altCounterOut_0})) ;
    mux21_ni ix141 (.Y (nx140), .A0 (currentState_1), .A1 (nx78), .S0 (nx123)) ;
    dffr reg_currentState_1 (.Q (currentState_1), .QB (nx151), .D (nx140), .CLK (
         NOT_clk), .R (resetState)) ;
    inv01 ix156 (.Y (NOT_clk), .A (clk)) ;
    nor02_2x ix79 (.Y (nx78), .A0 (finish), .A1 (resetCounter)) ;
    oai21 ix164 (.Y (nx163), .A0 (currentState_1), .A1 (dmaFinish), .B0 (
          currentState_0)) ;
    oai21 ix166 (.Y (nx165), .A0 (nx58), .A1 (loadConfig), .B0 (counterEn)) ;
    and04 ix59 (.Y (nx58), .A0 (nx168), .A1 (nx172), .A2 (nx176), .A3 (
          startFilterConv)) ;
    xnor2 ix169 (.Y (nx168), .A0 (counterOut_2), .A1 (filtersNumber[2])) ;
    dff reg_counterOut_2 (.Q (counterOut_2), .QB (\$dummy [0]), .D (
        altCounterOut_2), .CLK (clk)) ;
    xnor2 ix173 (.Y (nx172), .A0 (counterOut_0), .A1 (filtersNumber[0])) ;
    dff reg_counterOut_0 (.Q (counterOut_0), .QB (\$dummy [1]), .D (
        altCounterOut_0), .CLK (clk)) ;
    xnor2 ix177 (.Y (nx176), .A0 (counterOut_1), .A1 (filtersNumber[1])) ;
    dff reg_counterOut_1 (.Q (counterOut_1), .QB (\$dummy [2]), .D (
        altCounterOut_1), .CLK (clk)) ;
    ao21 ix19 (.Y (counterEn), .A0 (filterFinish), .A1 (nx185), .B0 (
         resetCounter)) ;
    dffr reg_currentState_0 (.Q (currentState_0), .QB (nx185), .D (nx130), .CLK (
         NOT_clk), .R (resetState)) ;
    nand02 ix71 (.Y (nx123), .A0 (nx163), .A1 (nx165)) ;
    and02 ix73 (.Y (finish), .A0 (currentState_1), .A1 (currentState_0)) ;
    and02 ix13 (.Y (resetCounter), .A0 (nx151), .A1 (nx185)) ;
    xnor2 ix131 (.Y (nx130), .A0 (nx185), .A1 (nx123)) ;
    and02 ix53 (.Y (startFilterConv), .A0 (currentState_1), .A1 (nx185)) ;
    nor02ii ix89 (.Y (loadConfig), .A0 (nx182), .A1 (nx151)) ;
    nor02ii ix183 (.Y (nx182), .A0 (start), .A1 (nx185)) ;
endmodule


module Counter_3 ( en, reset, clk, count ) ;

    input en ;
    input reset ;
    input clk ;
    output [2:0]count ;

    wire addedOne_2, addedOne_1, addedOne_0, finalReset, oneSignal_2, PWR;
    wire [0:0] \$dummy ;




    Reg_3 counterReg (.D ({addedOne_2,addedOne_1,addedOne_0}), .en (en), .clk (
          clk), .rst (finalReset), .Q ({count[2],count[1],count[0]})) ;
    NBitAdder_3 nextCount (.a ({count[2],count[1],count[0]}), .b ({oneSignal_2,
                oneSignal_2,oneSignal_2}), .carryIn (PWR), .sum ({addedOne_2,
                addedOne_1,addedOne_0}), .carryOut (\$dummy [0])) ;
    fake_vcc ix17 (.Y (PWR)) ;
    fake_gnd ix15 (.Y (oneSignal_2)) ;
    and02 ix1 (.Y (finalReset), .A0 (reset), .A1 (clk)) ;
endmodule


module NBitAdder_3 ( a, b, carryIn, sum, carryOut ) ;

    input [2:0]a ;
    input [2:0]b ;
    input carryIn ;
    output [2:0]sum ;
    output carryOut ;

    wire temp_1, temp_0;



    FullAdder f0 (.a (a[0]), .b (b[0]), .cin (carryIn), .s (sum[0]), .cout (
              temp_0)) ;
    FullAdder loop1_1_fx (.a (a[1]), .b (b[1]), .cin (temp_0), .s (sum[1]), .cout (
              temp_1)) ;
    FullAdder loop1_2_fx (.a (a[2]), .b (b[2]), .cin (temp_1), .s (sum[2]), .cout (
              carryOut)) ;
endmodule


module Reg_3 ( D, en, clk, rst, Q ) ;

    input [2:0]D ;
    input en ;
    input clk ;
    input rst ;
    output [2:0]Q ;

    wire nx72, nx82, nx92;
    wire [2:0] \$dummy ;




    dffr reg_Q_0 (.Q (Q[0]), .QB (\$dummy [0]), .D (nx72), .CLK (clk), .R (rst)
         ) ;
    mux21_ni ix73 (.Y (nx72), .A0 (Q[0]), .A1 (D[0]), .S0 (en)) ;
    dffr reg_Q_1 (.Q (Q[1]), .QB (\$dummy [1]), .D (nx82), .CLK (clk), .R (rst)
         ) ;
    mux21_ni ix83 (.Y (nx82), .A0 (Q[1]), .A1 (D[1]), .S0 (en)) ;
    dffr reg_Q_2 (.Q (Q[2]), .QB (\$dummy [2]), .D (nx92), .CLK (clk), .R (rst)
         ) ;
    mux21_ni ix93 (.Y (nx92), .A0 (Q[2]), .A1 (D[2]), .S0 (en)) ;
endmodule


module NetworkController_2 ( start, dmaFinish, oneLayerFinish, resetState, clk, 
                             layersNumber, loadConfig, startOneLayer, finish ) ;

    input start ;
    input dmaFinish ;
    input oneLayerFinish ;
    input resetState ;
    input clk ;
    input [1:0]layersNumber ;
    output loadConfig ;
    output startOneLayer ;
    output finish ;

    wire counterEn, altCounterOut_1, altCounterOut_0, resetCounter, 
         currentState_1, currentState_0, nx119, NOT_clk, counterOut_0, 
         counterOut_1, nx46, nx66, nx126, nx136, nx147, nx159, nx161, nx165, 
         nx169, nx174, nx177;
    wire [1:0] \$dummy ;




    Counter_2 counterMap (.en (counterEn), .reset (resetCounter), .clk (clk), .count (
              {altCounterOut_1,altCounterOut_0})) ;
    mux21_ni ix137 (.Y (nx136), .A0 (currentState_1), .A1 (nx66), .S0 (nx119)) ;
    dffr reg_currentState_1 (.Q (currentState_1), .QB (nx147), .D (nx136), .CLK (
         NOT_clk), .R (resetState)) ;
    inv01 ix152 (.Y (NOT_clk), .A (clk)) ;
    nor02_2x ix67 (.Y (nx66), .A0 (finish), .A1 (resetCounter)) ;
    oai21 ix160 (.Y (nx159), .A0 (currentState_1), .A1 (dmaFinish), .B0 (
          currentState_0)) ;
    oai21 ix162 (.Y (nx161), .A0 (nx46), .A1 (loadConfig), .B0 (counterEn)) ;
    and03 ix47 (.Y (nx46), .A0 (startOneLayer), .A1 (nx165), .A2 (nx169)) ;
    xnor2 ix166 (.Y (nx165), .A0 (counterOut_0), .A1 (layersNumber[0])) ;
    dff reg_counterOut_0 (.Q (counterOut_0), .QB (\$dummy [0]), .D (
        altCounterOut_0), .CLK (clk)) ;
    xnor2 ix170 (.Y (nx169), .A0 (counterOut_1), .A1 (layersNumber[1])) ;
    dff reg_counterOut_1 (.Q (counterOut_1), .QB (\$dummy [1]), .D (
        altCounterOut_1), .CLK (clk)) ;
    ao21 ix19 (.Y (counterEn), .A0 (oneLayerFinish), .A1 (nx177), .B0 (
         resetCounter)) ;
    dffr reg_currentState_0 (.Q (currentState_0), .QB (nx177), .D (nx126), .CLK (
         NOT_clk), .R (resetState)) ;
    nand02 ix59 (.Y (nx119), .A0 (nx159), .A1 (nx161)) ;
    and02 ix61 (.Y (finish), .A0 (currentState_1), .A1 (currentState_0)) ;
    and02 ix13 (.Y (resetCounter), .A0 (nx147), .A1 (nx177)) ;
    xnor2 ix127 (.Y (nx126), .A0 (nx177), .A1 (nx119)) ;
    and02 ix23 (.Y (startOneLayer), .A0 (currentState_1), .A1 (nx177)) ;
    nor02ii ix77 (.Y (loadConfig), .A0 (nx174), .A1 (nx147)) ;
    nor02ii ix175 (.Y (nx174), .A0 (start), .A1 (nx177)) ;
endmodule


module Counter_2 ( en, reset, clk, count ) ;

    input en ;
    input reset ;
    input clk ;
    output [1:0]count ;

    wire addedOne_1, addedOne_0, finalReset, oneSignal_1, PWR;
    wire [0:0] \$dummy ;




    Reg_2 counterReg (.D ({addedOne_1,addedOne_0}), .en (en), .clk (clk), .rst (
          finalReset), .Q ({count[1],count[0]})) ;
    NBitAdder_2 nextCount (.a ({count[1],count[0]}), .b ({oneSignal_1,
                oneSignal_1}), .carryIn (PWR), .sum ({addedOne_1,addedOne_0}), .carryOut (
                \$dummy [0])) ;
    fake_vcc ix15 (.Y (PWR)) ;
    fake_gnd ix13 (.Y (oneSignal_1)) ;
    and02 ix1 (.Y (finalReset), .A0 (reset), .A1 (clk)) ;
endmodule


module NBitAdder_2 ( a, b, carryIn, sum, carryOut ) ;

    input [1:0]a ;
    input [1:0]b ;
    input carryIn ;
    output [1:0]sum ;
    output carryOut ;

    wire temp_0;



    FullAdder f0 (.a (a[0]), .b (b[0]), .cin (carryIn), .s (sum[0]), .cout (
              temp_0)) ;
    FullAdder loop1_1_fx (.a (a[1]), .b (b[1]), .cin (temp_0), .s (sum[1]), .cout (
              carryOut)) ;
endmodule


module Reg_2 ( D, en, clk, rst, Q ) ;

    input [1:0]D ;
    input en ;
    input clk ;
    input rst ;
    output [1:0]Q ;

    wire nx60, nx70;
    wire [1:0] \$dummy ;




    dffr reg_Q_0 (.Q (Q[0]), .QB (\$dummy [0]), .D (nx60), .CLK (clk), .R (rst)
         ) ;
    mux21_ni ix61 (.Y (nx60), .A0 (Q[0]), .A1 (D[0]), .S0 (en)) ;
    dffr reg_Q_1 (.Q (Q[1]), .QB (\$dummy [1]), .D (nx70), .CLK (clk), .R (rst)
         ) ;
    mux21_ni ix71 (.Y (nx70), .A0 (Q[1]), .A1 (D[1]), .S0 (en)) ;
endmodule


module CNNCores_8_16_5_5_3 ( filterBus, windowBus, decoderRow, clk, rst, 
                             writePage1, writePage2, writeFilter, shift2To1, 
                             shift1To2, pageTurn, start, layerType, filterType, 
                             doneCores, finalSumConv ) ;

    input [39:0]filterBus ;
    input [79:0]windowBus ;
    input [2:0]decoderRow ;
    input clk ;
    input rst ;
    input writePage1 ;
    input writePage2 ;
    input writeFilter ;
    input shift2To1 ;
    input shift1To2 ;
    input pageTurn ;
    input start ;
    input layerType ;
    input filterType ;
    output doneCores ;
    output [15:0]finalSumConv ;

    wire currentPage_0__15, currentPage_0__14, currentPage_0__13, 
         currentPage_0__12, currentPage_0__11, currentPage_0__10, 
         currentPage_0__9, currentPage_0__8, currentPage_0__7, currentPage_0__6, 
         currentPage_0__5, currentPage_0__4, currentPage_0__3, currentPage_0__2, 
         currentPage_0__1, currentPage_0__0, currentPage_1__15, 
         currentPage_1__14, currentPage_1__13, currentPage_1__12, 
         currentPage_1__11, currentPage_1__10, currentPage_1__9, 
         currentPage_1__8, currentPage_1__7, currentPage_1__6, currentPage_1__5, 
         currentPage_1__4, currentPage_1__3, currentPage_1__2, currentPage_1__1, 
         currentPage_1__0, currentPage_2__15, currentPage_2__14, 
         currentPage_2__13, currentPage_2__12, currentPage_2__11, 
         currentPage_2__10, currentPage_2__9, currentPage_2__8, currentPage_2__7, 
         currentPage_2__6, currentPage_2__5, currentPage_2__4, currentPage_2__3, 
         currentPage_2__2, currentPage_2__1, currentPage_2__0, currentPage_3__15, 
         currentPage_3__14, currentPage_3__13, currentPage_3__12, 
         currentPage_3__11, currentPage_3__10, currentPage_3__9, 
         currentPage_3__8, currentPage_3__7, currentPage_3__6, currentPage_3__5, 
         currentPage_3__4, currentPage_3__3, currentPage_3__2, currentPage_3__1, 
         currentPage_3__0, currentPage_4__15, currentPage_4__14, 
         currentPage_4__13, currentPage_4__12, currentPage_4__11, 
         currentPage_4__10, currentPage_4__9, currentPage_4__8, currentPage_4__7, 
         currentPage_4__6, currentPage_4__5, currentPage_4__4, currentPage_4__3, 
         currentPage_4__2, currentPage_4__1, currentPage_4__0, currentPage_5__15, 
         currentPage_5__14, currentPage_5__13, currentPage_5__12, 
         currentPage_5__11, currentPage_5__10, currentPage_5__9, 
         currentPage_5__8, currentPage_5__7, currentPage_5__6, currentPage_5__5, 
         currentPage_5__4, currentPage_5__3, currentPage_5__2, currentPage_5__1, 
         currentPage_5__0, currentPage_6__15, currentPage_6__14, 
         currentPage_6__13, currentPage_6__12, currentPage_6__11, 
         currentPage_6__10, currentPage_6__9, currentPage_6__8, currentPage_6__7, 
         currentPage_6__6, currentPage_6__5, currentPage_6__4, currentPage_6__3, 
         currentPage_6__2, currentPage_6__1, currentPage_6__0, currentPage_7__15, 
         currentPage_7__14, currentPage_7__13, currentPage_7__12, 
         currentPage_7__11, currentPage_7__10, currentPage_7__9, 
         currentPage_7__8, currentPage_7__7, currentPage_7__6, currentPage_7__5, 
         currentPage_7__4, currentPage_7__3, currentPage_7__2, currentPage_7__1, 
         currentPage_7__0, currentPage_8__15, currentPage_8__14, 
         currentPage_8__13, currentPage_8__12, currentPage_8__11, 
         currentPage_8__10, currentPage_8__9, currentPage_8__8, currentPage_8__7, 
         currentPage_8__6, currentPage_8__5, currentPage_8__4, currentPage_8__3, 
         currentPage_8__2, currentPage_8__1, currentPage_8__0, currentPage_9__15, 
         currentPage_9__14, currentPage_9__13, currentPage_9__12, 
         currentPage_9__11, currentPage_9__10, currentPage_9__9, 
         currentPage_9__8, currentPage_9__7, currentPage_9__6, currentPage_9__5, 
         currentPage_9__4, currentPage_9__3, currentPage_9__2, currentPage_9__1, 
         currentPage_9__0, currentPage_10__15, currentPage_10__14, 
         currentPage_10__13, currentPage_10__12, currentPage_10__11, 
         currentPage_10__10, currentPage_10__9, currentPage_10__8, 
         currentPage_10__7, currentPage_10__6, currentPage_10__5, 
         currentPage_10__4, currentPage_10__3, currentPage_10__2, 
         currentPage_10__1, currentPage_10__0, currentPage_11__15, 
         currentPage_11__14, currentPage_11__13, currentPage_11__12, 
         currentPage_11__11, currentPage_11__10, currentPage_11__9, 
         currentPage_11__8, currentPage_11__7, currentPage_11__6, 
         currentPage_11__5, currentPage_11__4, currentPage_11__3, 
         currentPage_11__2, currentPage_11__1, currentPage_11__0, 
         currentPage_12__15, currentPage_12__14, currentPage_12__13, 
         currentPage_12__12, currentPage_12__11, currentPage_12__10, 
         currentPage_12__9, currentPage_12__8, currentPage_12__7, 
         currentPage_12__6, currentPage_12__5, currentPage_12__4, 
         currentPage_12__3, currentPage_12__2, currentPage_12__1, 
         currentPage_12__0, currentPage_13__15, currentPage_13__14, 
         currentPage_13__13, currentPage_13__12, currentPage_13__11, 
         currentPage_13__10, currentPage_13__9, currentPage_13__8, 
         currentPage_13__7, currentPage_13__6, currentPage_13__5, 
         currentPage_13__4, currentPage_13__3, currentPage_13__2, 
         currentPage_13__1, currentPage_13__0, currentPage_14__15, 
         currentPage_14__14, currentPage_14__13, currentPage_14__12, 
         currentPage_14__11, currentPage_14__10, currentPage_14__9, 
         currentPage_14__8, currentPage_14__7, currentPage_14__6, 
         currentPage_14__5, currentPage_14__4, currentPage_14__3, 
         currentPage_14__2, currentPage_14__1, currentPage_14__0, 
         currentPage_15__15, currentPage_15__14, currentPage_15__13, 
         currentPage_15__12, currentPage_15__11, currentPage_15__10, 
         currentPage_15__9, currentPage_15__8, currentPage_15__7, 
         currentPage_15__6, currentPage_15__5, currentPage_15__4, 
         currentPage_15__3, currentPage_15__2, currentPage_15__1, 
         currentPage_15__0, currentPage_16__15, currentPage_16__14, 
         currentPage_16__13, currentPage_16__12, currentPage_16__11, 
         currentPage_16__10, currentPage_16__9, currentPage_16__8, 
         currentPage_16__7, currentPage_16__6, currentPage_16__5, 
         currentPage_16__4, currentPage_16__3, currentPage_16__2, 
         currentPage_16__1, currentPage_16__0, currentPage_17__15, 
         currentPage_17__14, currentPage_17__13, currentPage_17__12, 
         currentPage_17__11, currentPage_17__10, currentPage_17__9, 
         currentPage_17__8, currentPage_17__7, currentPage_17__6, 
         currentPage_17__5, currentPage_17__4, currentPage_17__3, 
         currentPage_17__2, currentPage_17__1, currentPage_17__0, 
         currentPage_18__15, currentPage_18__14, currentPage_18__13, 
         currentPage_18__12, currentPage_18__11, currentPage_18__10, 
         currentPage_18__9, currentPage_18__8, currentPage_18__7, 
         currentPage_18__6, currentPage_18__5, currentPage_18__4, 
         currentPage_18__3, currentPage_18__2, currentPage_18__1, 
         currentPage_18__0, currentPage_19__15, currentPage_19__14, 
         currentPage_19__13, currentPage_19__12, currentPage_19__11, 
         currentPage_19__10, currentPage_19__9, currentPage_19__8, 
         currentPage_19__7, currentPage_19__6, currentPage_19__5, 
         currentPage_19__4, currentPage_19__3, currentPage_19__2, 
         currentPage_19__1, currentPage_19__0, currentPage_20__15, 
         currentPage_20__14, currentPage_20__13, currentPage_20__12, 
         currentPage_20__11, currentPage_20__10, currentPage_20__9, 
         currentPage_20__8, currentPage_20__7, currentPage_20__6, 
         currentPage_20__5, currentPage_20__4, currentPage_20__3, 
         currentPage_20__2, currentPage_20__1, currentPage_20__0, 
         currentPage_21__15, currentPage_21__14, currentPage_21__13, 
         currentPage_21__12, currentPage_21__11, currentPage_21__10, 
         currentPage_21__9, currentPage_21__8, currentPage_21__7, 
         currentPage_21__6, currentPage_21__5, currentPage_21__4, 
         currentPage_21__3, currentPage_21__2, currentPage_21__1, 
         currentPage_21__0, currentPage_22__15, currentPage_22__14, 
         currentPage_22__13, currentPage_22__12, currentPage_22__11, 
         currentPage_22__10, currentPage_22__9, currentPage_22__8, 
         currentPage_22__7, currentPage_22__6, currentPage_22__5, 
         currentPage_22__4, currentPage_22__3, currentPage_22__2, 
         currentPage_22__1, currentPage_22__0, currentPage_23__15, 
         currentPage_23__14, currentPage_23__13, currentPage_23__12, 
         currentPage_23__11, currentPage_23__10, currentPage_23__9, 
         currentPage_23__8, currentPage_23__7, currentPage_23__6, 
         currentPage_23__5, currentPage_23__4, currentPage_23__3, 
         currentPage_23__2, currentPage_23__1, currentPage_23__0, 
         currentPage_24__15, currentPage_24__14, currentPage_24__13, 
         currentPage_24__12, currentPage_24__11, currentPage_24__10, 
         currentPage_24__9, currentPage_24__8, currentPage_24__7, 
         currentPage_24__6, currentPage_24__5, currentPage_24__4, 
         currentPage_24__3, currentPage_24__2, currentPage_24__1, 
         currentPage_24__0, outMuls_0__15, outMuls_0__14, outMuls_0__13, 
         outMuls_0__12, outMuls_0__11, outMuls_0__10, outMuls_0__9, outMuls_0__8, 
         outMuls_0__7, outMuls_0__6, outMuls_0__5, outMuls_0__4, outMuls_0__3, 
         outMuls_0__2, outMuls_0__1, outMuls_0__0, outMuls_1__15, outMuls_1__14, 
         outMuls_1__13, outMuls_1__12, outMuls_1__11, outMuls_1__10, 
         outMuls_1__9, outMuls_1__8, outMuls_1__7, outMuls_1__6, outMuls_1__5, 
         outMuls_1__4, outMuls_1__3, outMuls_1__2, outMuls_1__1, outMuls_1__0, 
         outMuls_2__15, outMuls_2__14, outMuls_2__13, outMuls_2__12, 
         outMuls_2__11, outMuls_2__10, outMuls_2__9, outMuls_2__8, outMuls_2__7, 
         outMuls_2__6, outMuls_2__5, outMuls_2__4, outMuls_2__3, outMuls_2__2, 
         outMuls_2__1, outMuls_2__0, outMuls_3__15, outMuls_3__14, outMuls_3__13, 
         outMuls_3__12, outMuls_3__11, outMuls_3__10, outMuls_3__9, outMuls_3__8, 
         outMuls_3__7, outMuls_3__6, outMuls_3__5, outMuls_3__4, outMuls_3__3, 
         outMuls_3__2, outMuls_3__1, outMuls_3__0, outMuls_4__15, outMuls_4__14, 
         outMuls_4__13, outMuls_4__12, outMuls_4__11, outMuls_4__10, 
         outMuls_4__9, outMuls_4__8, outMuls_4__7, outMuls_4__6, outMuls_4__5, 
         outMuls_4__4, outMuls_4__3, outMuls_4__2, outMuls_4__1, outMuls_4__0, 
         outMuls_5__15, outMuls_5__14, outMuls_5__13, outMuls_5__12, 
         outMuls_5__11, outMuls_5__10, outMuls_5__9, outMuls_5__8, outMuls_5__7, 
         outMuls_5__6, outMuls_5__5, outMuls_5__4, outMuls_5__3, outMuls_5__2, 
         outMuls_5__1, outMuls_5__0, outMuls_6__15, outMuls_6__14, outMuls_6__13, 
         outMuls_6__12, outMuls_6__11, outMuls_6__10, outMuls_6__9, outMuls_6__8, 
         outMuls_6__7, outMuls_6__6, outMuls_6__5, outMuls_6__4, outMuls_6__3, 
         outMuls_6__2, outMuls_6__1, outMuls_6__0, outMuls_7__15, outMuls_7__14, 
         outMuls_7__13, outMuls_7__12, outMuls_7__11, outMuls_7__10, 
         outMuls_7__9, outMuls_7__8, outMuls_7__7, outMuls_7__6, outMuls_7__5, 
         outMuls_7__4, outMuls_7__3, outMuls_7__2, outMuls_7__1, outMuls_7__0, 
         outMuls_8__15, outMuls_8__14, outMuls_8__13, outMuls_8__12, 
         outMuls_8__11, outMuls_8__10, outMuls_8__9, outMuls_8__8, outMuls_8__7, 
         outMuls_8__6, outMuls_8__5, outMuls_8__4, outMuls_8__3, outMuls_8__2, 
         outMuls_8__1, outMuls_8__0, outMuls_9__15, outMuls_9__14, outMuls_9__13, 
         outMuls_9__12, outMuls_9__11, outMuls_9__10, outMuls_9__9, outMuls_9__8, 
         outMuls_9__7, outMuls_9__6, outMuls_9__5, outMuls_9__4, outMuls_9__3, 
         outMuls_9__2, outMuls_9__1, outMuls_9__0, outMuls_10__15, 
         outMuls_10__14, outMuls_10__13, outMuls_10__12, outMuls_10__11, 
         outMuls_10__10, outMuls_10__9, outMuls_10__8, outMuls_10__7, 
         outMuls_10__6, outMuls_10__5, outMuls_10__4, outMuls_10__3, 
         outMuls_10__2, outMuls_10__1, outMuls_10__0, outMuls_11__15, 
         outMuls_11__14, outMuls_11__13, outMuls_11__12, outMuls_11__11, 
         outMuls_11__10, outMuls_11__9, outMuls_11__8, outMuls_11__7, 
         outMuls_11__6, outMuls_11__5, outMuls_11__4, outMuls_11__3, 
         outMuls_11__2, outMuls_11__1, outMuls_11__0, outMuls_12__15, 
         outMuls_12__14, outMuls_12__13, outMuls_12__12, outMuls_12__11, 
         outMuls_12__10, outMuls_12__9, outMuls_12__8, outMuls_12__7, 
         outMuls_12__6, outMuls_12__5, outMuls_12__4, outMuls_12__3, 
         outMuls_12__2, outMuls_12__1, outMuls_12__0, outMuls_13__15, 
         outMuls_13__14, outMuls_13__13, outMuls_13__12, outMuls_13__11, 
         outMuls_13__10, outMuls_13__9, outMuls_13__8, outMuls_13__7, 
         outMuls_13__6, outMuls_13__5, outMuls_13__4, outMuls_13__3, 
         outMuls_13__2, outMuls_13__1, outMuls_13__0, outMuls_14__15, 
         outMuls_14__14, outMuls_14__13, outMuls_14__12, outMuls_14__11, 
         outMuls_14__10, outMuls_14__9, outMuls_14__8, outMuls_14__7, 
         outMuls_14__6, outMuls_14__5, outMuls_14__4, outMuls_14__3, 
         outMuls_14__2, outMuls_14__1, outMuls_14__0, outMuls_15__15, 
         outMuls_15__14, outMuls_15__13, outMuls_15__12, outMuls_15__11, 
         outMuls_15__10, outMuls_15__9, outMuls_15__8, outMuls_15__7, 
         outMuls_15__6, outMuls_15__5, outMuls_15__4, outMuls_15__3, 
         outMuls_15__2, outMuls_15__1, outMuls_15__0, outMuls_16__15, 
         outMuls_16__14, outMuls_16__13, outMuls_16__12, outMuls_16__11, 
         outMuls_16__10, outMuls_16__9, outMuls_16__8, outMuls_16__7, 
         outMuls_16__6, outMuls_16__5, outMuls_16__4, outMuls_16__3, 
         outMuls_16__2, outMuls_16__1, outMuls_16__0, outMuls_17__15, 
         outMuls_17__14, outMuls_17__13, outMuls_17__12, outMuls_17__11, 
         outMuls_17__10, outMuls_17__9, outMuls_17__8, outMuls_17__7, 
         outMuls_17__6, outMuls_17__5, outMuls_17__4, outMuls_17__3, 
         outMuls_17__2, outMuls_17__1, outMuls_17__0, outMuls_18__15, 
         outMuls_18__14, outMuls_18__13, outMuls_18__12, outMuls_18__11, 
         outMuls_18__10, outMuls_18__9, outMuls_18__8, outMuls_18__7, 
         outMuls_18__6, outMuls_18__5, outMuls_18__4, outMuls_18__3, 
         outMuls_18__2, outMuls_18__1, outMuls_18__0, outMuls_19__15, 
         outMuls_19__14, outMuls_19__13, outMuls_19__12, outMuls_19__11, 
         outMuls_19__10, outMuls_19__9, outMuls_19__8, outMuls_19__7, 
         outMuls_19__6, outMuls_19__5, outMuls_19__4, outMuls_19__3, 
         outMuls_19__2, outMuls_19__1, outMuls_19__0, outMuls_20__15, 
         outMuls_20__14, outMuls_20__13, outMuls_20__12, outMuls_20__11, 
         outMuls_20__10, outMuls_20__9, outMuls_20__8, outMuls_20__7, 
         outMuls_20__6, outMuls_20__5, outMuls_20__4, outMuls_20__3, 
         outMuls_20__2, outMuls_20__1, outMuls_20__0, outMuls_21__15, 
         outMuls_21__14, outMuls_21__13, outMuls_21__12, outMuls_21__11, 
         outMuls_21__10, outMuls_21__9, outMuls_21__8, outMuls_21__7, 
         outMuls_21__6, outMuls_21__5, outMuls_21__4, outMuls_21__3, 
         outMuls_21__2, outMuls_21__1, outMuls_21__0, outMuls_22__15, 
         outMuls_22__14, outMuls_22__13, outMuls_22__12, outMuls_22__11, 
         outMuls_22__10, outMuls_22__9, outMuls_22__8, outMuls_22__7, 
         outMuls_22__6, outMuls_22__5, outMuls_22__4, outMuls_22__3, 
         outMuls_22__2, outMuls_22__1, outMuls_22__0, outMuls_23__15, 
         outMuls_23__14, outMuls_23__13, outMuls_23__12, outMuls_23__11, 
         outMuls_23__10, outMuls_23__9, outMuls_23__8, outMuls_23__7, 
         outMuls_23__6, outMuls_23__5, outMuls_23__4, outMuls_23__3, 
         outMuls_23__2, outMuls_23__1, outMuls_23__0, outMuls_24__15, 
         outMuls_24__14, outMuls_24__13, outMuls_24__12, outMuls_24__11, 
         outMuls_24__10, outMuls_24__9, outMuls_24__8, outMuls_24__7, 
         outMuls_24__6, outMuls_24__5, outMuls_24__4, outMuls_24__3, 
         outMuls_24__2, outMuls_24__1, outMuls_24__0, addersInputs_0__15, 
         addersInputs_0__14, addersInputs_0__13, addersInputs_0__12, 
         addersInputs_0__11, addersInputs_0__10, addersInputs_0__9, 
         addersInputs_0__8, addersInputs_0__7, addersInputs_0__6, 
         addersInputs_0__5, addersInputs_0__4, addersInputs_0__3, 
         addersInputs_0__2, addersInputs_0__1, addersInputs_0__0, 
         addersInputs_1__15, addersInputs_1__14, addersInputs_1__13, 
         addersInputs_1__12, addersInputs_1__11, addersInputs_1__10, 
         addersInputs_1__9, addersInputs_1__8, addersInputs_1__7, 
         addersInputs_1__6, addersInputs_1__5, addersInputs_1__4, 
         addersInputs_1__3, addersInputs_1__2, addersInputs_1__1, 
         addersInputs_1__0, addersInputs_2__15, addersInputs_2__14, 
         addersInputs_2__13, addersInputs_2__12, addersInputs_2__11, 
         addersInputs_2__10, addersInputs_2__9, addersInputs_2__8, 
         addersInputs_2__7, addersInputs_2__6, addersInputs_2__5, 
         addersInputs_2__4, addersInputs_2__3, addersInputs_2__2, 
         addersInputs_2__1, addersInputs_2__0, addersInputs_3__15, 
         addersInputs_3__14, addersInputs_3__13, addersInputs_3__12, 
         addersInputs_3__11, addersInputs_3__10, addersInputs_3__9, 
         addersInputs_3__8, addersInputs_3__7, addersInputs_3__6, 
         addersInputs_3__5, addersInputs_3__4, addersInputs_3__3, 
         addersInputs_3__2, addersInputs_3__1, addersInputs_3__0, 
         addersInputs_4__15, addersInputs_4__14, addersInputs_4__13, 
         addersInputs_4__12, addersInputs_4__11, addersInputs_4__10, 
         addersInputs_4__9, addersInputs_4__8, addersInputs_4__7, 
         addersInputs_4__6, addersInputs_4__5, addersInputs_4__4, 
         addersInputs_4__3, addersInputs_4__2, addersInputs_4__1, 
         addersInputs_4__0, addersInputs_5__15, addersInputs_5__14, 
         addersInputs_5__13, addersInputs_5__12, addersInputs_5__11, 
         addersInputs_5__10, addersInputs_5__9, addersInputs_5__8, 
         addersInputs_5__7, addersInputs_5__6, addersInputs_5__5, 
         addersInputs_5__4, addersInputs_5__3, addersInputs_5__2, 
         addersInputs_5__1, addersInputs_5__0, addersInputs_6__15, 
         addersInputs_6__14, addersInputs_6__13, addersInputs_6__12, 
         addersInputs_6__11, addersInputs_6__10, addersInputs_6__9, 
         addersInputs_6__8, addersInputs_6__7, addersInputs_6__6, 
         addersInputs_6__5, addersInputs_6__4, addersInputs_6__3, 
         addersInputs_6__2, addersInputs_6__1, addersInputs_6__0, 
         addersInputs_7__15, addersInputs_7__14, addersInputs_7__13, 
         addersInputs_7__12, addersInputs_7__11, addersInputs_7__10, 
         addersInputs_7__9, addersInputs_7__8, addersInputs_7__7, 
         addersInputs_7__6, addersInputs_7__5, addersInputs_7__4, 
         addersInputs_7__3, addersInputs_7__2, addersInputs_7__1, 
         addersInputs_7__0, addersInputs_8__15, addersInputs_8__14, 
         addersInputs_8__13, addersInputs_8__12, addersInputs_8__11, 
         addersInputs_8__10, addersInputs_8__9, addersInputs_8__8, 
         addersInputs_8__7, addersInputs_8__6, addersInputs_8__5, 
         addersInputs_8__4, addersInputs_8__3, addersInputs_8__2, 
         addersInputs_8__1, addersInputs_8__0, addersInputs_9__15, 
         addersInputs_9__14, addersInputs_9__13, addersInputs_9__12, 
         addersInputs_9__11, addersInputs_9__10, addersInputs_9__9, 
         addersInputs_9__8, addersInputs_9__7, addersInputs_9__6, 
         addersInputs_9__5, addersInputs_9__4, addersInputs_9__3, 
         addersInputs_9__2, addersInputs_9__1, addersInputs_9__0, 
         addersInputs_10__15, addersInputs_10__14, addersInputs_10__13, 
         addersInputs_10__12, addersInputs_10__11, addersInputs_10__10, 
         addersInputs_10__9, addersInputs_10__8, addersInputs_10__7, 
         addersInputs_10__6, addersInputs_10__5, addersInputs_10__4, 
         addersInputs_10__3, addersInputs_10__2, addersInputs_10__1, 
         addersInputs_10__0, addersInputs_11__15, addersInputs_11__14, 
         addersInputs_11__13, addersInputs_11__12, addersInputs_11__11, 
         addersInputs_11__10, addersInputs_11__9, addersInputs_11__8, 
         addersInputs_11__7, addersInputs_11__6, addersInputs_11__5, 
         addersInputs_11__4, addersInputs_11__3, addersInputs_11__2, 
         addersInputs_11__1, addersInputs_11__0, addersInputs_12__15, 
         addersInputs_12__14, addersInputs_12__13, addersInputs_12__12, 
         addersInputs_12__11, addersInputs_12__10, addersInputs_12__9, 
         addersInputs_12__8, addersInputs_12__7, addersInputs_12__6, 
         addersInputs_12__5, addersInputs_12__4, addersInputs_12__3, 
         addersInputs_12__2, addersInputs_12__1, addersInputs_12__0, 
         addersInputs_13__15, addersInputs_13__14, addersInputs_13__13, 
         addersInputs_13__12, addersInputs_13__11, addersInputs_13__10, 
         addersInputs_13__9, addersInputs_13__8, addersInputs_13__7, 
         addersInputs_13__6, addersInputs_13__5, addersInputs_13__4, 
         addersInputs_13__3, addersInputs_13__2, addersInputs_13__1, 
         addersInputs_13__0, addersInputs_14__15, addersInputs_14__14, 
         addersInputs_14__13, addersInputs_14__12, addersInputs_14__11, 
         addersInputs_14__10, addersInputs_14__9, addersInputs_14__8, 
         addersInputs_14__7, addersInputs_14__6, addersInputs_14__5, 
         addersInputs_14__4, addersInputs_14__3, addersInputs_14__2, 
         addersInputs_14__1, addersInputs_14__0, addersInputs_15__15, 
         addersInputs_15__14, addersInputs_15__13, addersInputs_15__12, 
         addersInputs_15__11, addersInputs_15__10, addersInputs_15__9, 
         addersInputs_15__8, addersInputs_15__7, addersInputs_15__6, 
         addersInputs_15__5, addersInputs_15__4, addersInputs_15__3, 
         addersInputs_15__2, addersInputs_15__1, addersInputs_15__0, 
         addersInputs_16__15, addersInputs_16__14, addersInputs_16__13, 
         addersInputs_16__12, addersInputs_16__11, addersInputs_16__10, 
         addersInputs_16__9, addersInputs_16__8, addersInputs_16__7, 
         addersInputs_16__6, addersInputs_16__5, addersInputs_16__4, 
         addersInputs_16__3, addersInputs_16__2, addersInputs_16__1, 
         addersInputs_16__0, addersInputs_17__15, addersInputs_17__14, 
         addersInputs_17__13, addersInputs_17__12, addersInputs_17__11, 
         addersInputs_17__10, addersInputs_17__9, addersInputs_17__8, 
         addersInputs_17__7, addersInputs_17__6, addersInputs_17__5, 
         addersInputs_17__4, addersInputs_17__3, addersInputs_17__2, 
         addersInputs_17__1, addersInputs_17__0, addersInputs_18__15, 
         addersInputs_18__14, addersInputs_18__13, addersInputs_18__12, 
         addersInputs_18__11, addersInputs_18__10, addersInputs_18__9, 
         addersInputs_18__8, addersInputs_18__7, addersInputs_18__6, 
         addersInputs_18__5, addersInputs_18__4, addersInputs_18__3, 
         addersInputs_18__2, addersInputs_18__1, addersInputs_18__0, 
         addersInputs_19__15, addersInputs_19__14, addersInputs_19__13, 
         addersInputs_19__12, addersInputs_19__11, addersInputs_19__10, 
         addersInputs_19__9, addersInputs_19__8, addersInputs_19__7, 
         addersInputs_19__6, addersInputs_19__5, addersInputs_19__4, 
         addersInputs_19__3, addersInputs_19__2, addersInputs_19__1, 
         addersInputs_19__0, addersInputs_20__15, addersInputs_20__14, 
         addersInputs_20__13, addersInputs_20__12, addersInputs_20__11, 
         addersInputs_20__10, addersInputs_20__9, addersInputs_20__8, 
         addersInputs_20__7, addersInputs_20__6, addersInputs_20__5, 
         addersInputs_20__4, addersInputs_20__3, addersInputs_20__2, 
         addersInputs_20__1, addersInputs_20__0, addersInputs_21__15, 
         addersInputs_21__14, addersInputs_21__13, addersInputs_21__12, 
         addersInputs_21__11, addersInputs_21__10, addersInputs_21__9, 
         addersInputs_21__8, addersInputs_21__7, addersInputs_21__6, 
         addersInputs_21__5, addersInputs_21__4, addersInputs_21__3, 
         addersInputs_21__2, addersInputs_21__1, addersInputs_21__0, 
         addersInputs_22__15, addersInputs_22__14, addersInputs_22__13, 
         addersInputs_22__12, addersInputs_22__11, addersInputs_22__10, 
         addersInputs_22__9, addersInputs_22__8, addersInputs_22__7, 
         addersInputs_22__6, addersInputs_22__5, addersInputs_22__4, 
         addersInputs_22__3, addersInputs_22__2, addersInputs_22__1, 
         addersInputs_22__0, addersInputs_23__15, addersInputs_23__14, 
         addersInputs_23__13, addersInputs_23__12, addersInputs_23__11, 
         addersInputs_23__10, addersInputs_23__9, addersInputs_23__8, 
         addersInputs_23__7, addersInputs_23__6, addersInputs_23__5, 
         addersInputs_23__4, addersInputs_23__3, addersInputs_23__2, 
         addersInputs_23__1, addersInputs_23__0, addersInputs_24__15, 
         addersInputs_24__14, addersInputs_24__13, addersInputs_24__12, 
         addersInputs_24__11, addersInputs_24__10, addersInputs_24__9, 
         addersInputs_24__8, addersInputs_24__7, addersInputs_24__6, 
         addersInputs_24__5, addersInputs_24__4, addersInputs_24__3, 
         addersInputs_24__2, addersInputs_24__1, addersInputs_24__0, filter_0__7, 
         filter_0__6, filter_0__5, filter_0__4, filter_0__3, filter_0__2, 
         filter_0__1, filter_0__0, filter_1__7, filter_1__6, filter_1__5, 
         filter_1__4, filter_1__3, filter_1__2, filter_1__1, filter_1__0, 
         filter_2__7, filter_2__6, filter_2__5, filter_2__4, filter_2__3, 
         filter_2__2, filter_2__1, filter_2__0, filter_3__7, filter_3__6, 
         filter_3__5, filter_3__4, filter_3__3, filter_3__2, filter_3__1, 
         filter_3__0, filter_4__7, filter_4__6, filter_4__5, filter_4__4, 
         filter_4__3, filter_4__2, filter_4__1, filter_4__0, filter_5__7, 
         filter_5__6, filter_5__5, filter_5__4, filter_5__3, filter_5__2, 
         filter_5__1, filter_5__0, filter_6__7, filter_6__6, filter_6__5, 
         filter_6__4, filter_6__3, filter_6__2, filter_6__1, filter_6__0, 
         filter_7__7, filter_7__6, filter_7__5, filter_7__4, filter_7__3, 
         filter_7__2, filter_7__1, filter_7__0, filter_8__7, filter_8__6, 
         filter_8__5, filter_8__4, filter_8__3, filter_8__2, filter_8__1, 
         filter_8__0, filter_9__7, filter_9__6, filter_9__5, filter_9__4, 
         filter_9__3, filter_9__2, filter_9__1, filter_9__0, filter_10__7, 
         filter_10__6, filter_10__5, filter_10__4, filter_10__3, filter_10__2, 
         filter_10__1, filter_10__0, filter_11__7, filter_11__6, filter_11__5, 
         filter_11__4, filter_11__3, filter_11__2, filter_11__1, filter_11__0, 
         filter_12__7, filter_12__6, filter_12__5, filter_12__4, filter_12__3, 
         filter_12__2, filter_12__1, filter_12__0, filter_13__7, filter_13__6, 
         filter_13__5, filter_13__4, filter_13__3, filter_13__2, filter_13__1, 
         filter_13__0, filter_14__7, filter_14__6, filter_14__5, filter_14__4, 
         filter_14__3, filter_14__2, filter_14__1, filter_14__0, filter_15__7, 
         filter_15__6, filter_15__5, filter_15__4, filter_15__3, filter_15__2, 
         filter_15__1, filter_15__0, filter_16__7, filter_16__6, filter_16__5, 
         filter_16__4, filter_16__3, filter_16__2, filter_16__1, filter_16__0, 
         filter_17__7, filter_17__6, filter_17__5, filter_17__4, filter_17__3, 
         filter_17__2, filter_17__1, filter_17__0, filter_18__7, filter_18__6, 
         filter_18__5, filter_18__4, filter_18__3, filter_18__2, filter_18__1, 
         filter_18__0, filter_19__7, filter_19__6, filter_19__5, filter_19__4, 
         filter_19__3, filter_19__2, filter_19__1, filter_19__0, filter_20__7, 
         filter_20__6, filter_20__5, filter_20__4, filter_20__3, filter_20__2, 
         filter_20__1, filter_20__0, filter_21__7, filter_21__6, filter_21__5, 
         filter_21__4, filter_21__3, filter_21__2, filter_21__1, filter_21__0, 
         filter_22__7, filter_22__6, filter_22__5, filter_22__4, filter_22__3, 
         filter_22__2, filter_22__1, filter_22__0, filter_23__7, filter_23__6, 
         filter_23__5, filter_23__4, filter_23__3, filter_23__2, filter_23__1, 
         filter_23__0, filter_24__7, filter_24__6, filter_24__5, filter_24__4, 
         filter_24__3, filter_24__2, filter_24__1, filter_24__0, doneMul, notClk, 
         outAdder_15, outAdder_14, outAdder_13, outAdder_12, outAdder_11, 
         outAdder_10, outAdder_9, outAdder_8, outAdder_7, outAdder_6, outAdder_5, 
         outAdder_4, outAdder_3, outAdder_2, outAdder_1, outAdder_0, 
         outShifter_11, outShifter_10, outShifter_9, outShifter_8, outShifter_7, 
         outShifter_6, outShifter_5, outShifter_4, outShifter_3, outShifter_2, 
         outShifter_1, outShifter_0, finalSum_15, finalSum_14, finalSum_13, 
         finalSum_12, finalSum_11, finalSum_10, finalSum_9, finalSum_8, 
         finalSum_7, finalSum_6, finalSum_5, finalSum_4, finalSum_3, finalSum_2, 
         finalSum_1, finalSum_0, nx1921, nx1944, nx1946, nx1948, nx1950, nx1952;
    wire [4:0] \$dummy ;




    RegFile_8_16_5_5_3_3 regFileMap (.filterBus ({filterBus[39],filterBus[38],
                         filterBus[37],filterBus[36],filterBus[35],filterBus[34]
                         ,filterBus[33],filterBus[32],filterBus[31],
                         filterBus[30],filterBus[29],filterBus[28],filterBus[27]
                         ,filterBus[26],filterBus[25],filterBus[24],
                         filterBus[23],filterBus[22],filterBus[21],filterBus[20]
                         ,filterBus[19],filterBus[18],filterBus[17],
                         filterBus[16],filterBus[15],filterBus[14],filterBus[13]
                         ,filterBus[12],filterBus[11],filterBus[10],filterBus[9]
                         ,filterBus[8],filterBus[7],filterBus[6],filterBus[5],
                         filterBus[4],filterBus[3],filterBus[2],filterBus[1],
                         filterBus[0]}), .windowBus ({windowBus[79],
                         windowBus[78],windowBus[77],windowBus[76],windowBus[75]
                         ,windowBus[74],windowBus[73],windowBus[72],
                         windowBus[71],windowBus[70],windowBus[69],windowBus[68]
                         ,windowBus[67],windowBus[66],windowBus[65],
                         windowBus[64],windowBus[63],windowBus[62],windowBus[61]
                         ,windowBus[60],windowBus[59],windowBus[58],
                         windowBus[57],windowBus[56],windowBus[55],windowBus[54]
                         ,windowBus[53],windowBus[52],windowBus[51],
                         windowBus[50],windowBus[49],windowBus[48],windowBus[47]
                         ,windowBus[46],windowBus[45],windowBus[44],
                         windowBus[43],windowBus[42],windowBus[41],windowBus[40]
                         ,windowBus[39],windowBus[38],windowBus[37],
                         windowBus[36],windowBus[35],windowBus[34],windowBus[33]
                         ,windowBus[32],windowBus[31],windowBus[30],
                         windowBus[29],windowBus[28],windowBus[27],windowBus[26]
                         ,windowBus[25],windowBus[24],windowBus[23],
                         windowBus[22],windowBus[21],windowBus[20],windowBus[19]
                         ,windowBus[18],windowBus[17],windowBus[16],
                         windowBus[15],windowBus[14],windowBus[13],windowBus[12]
                         ,windowBus[11],windowBus[10],windowBus[9],windowBus[8],
                         windowBus[7],windowBus[6],windowBus[5],windowBus[4],
                         windowBus[3],windowBus[2],windowBus[1],windowBus[0]}), 
                         .decoderRow ({decoderRow[2],decoderRow[1],decoderRow[0]
                         }), .clk (clk), .rst (rst), .enablePage1Read (
                         writePage1), .enablePage2Read (writePage2), .enableFilterRead (
                         writeFilter), .shift2To1 (shift2To1), .shift1To2 (
                         shift1To2), .pageTurn (pageTurn), .pagesOuts_0__15 (
                         currentPage_0__15), .pagesOuts_0__14 (currentPage_0__14
                         ), .pagesOuts_0__13 (currentPage_0__13), .pagesOuts_0__12 (
                         currentPage_0__12), .pagesOuts_0__11 (currentPage_0__11
                         ), .pagesOuts_0__10 (currentPage_0__10), .pagesOuts_0__9 (
                         currentPage_0__9), .pagesOuts_0__8 (currentPage_0__8), 
                         .pagesOuts_0__7 (currentPage_0__7), .pagesOuts_0__6 (
                         currentPage_0__6), .pagesOuts_0__5 (currentPage_0__5), 
                         .pagesOuts_0__4 (currentPage_0__4), .pagesOuts_0__3 (
                         currentPage_0__3), .pagesOuts_0__2 (currentPage_0__2), 
                         .pagesOuts_0__1 (currentPage_0__1), .pagesOuts_0__0 (
                         currentPage_0__0), .pagesOuts_1__15 (currentPage_1__15)
                         , .pagesOuts_1__14 (currentPage_1__14), .pagesOuts_1__13 (
                         currentPage_1__13), .pagesOuts_1__12 (currentPage_1__12
                         ), .pagesOuts_1__11 (currentPage_1__11), .pagesOuts_1__10 (
                         currentPage_1__10), .pagesOuts_1__9 (currentPage_1__9)
                         , .pagesOuts_1__8 (currentPage_1__8), .pagesOuts_1__7 (
                         currentPage_1__7), .pagesOuts_1__6 (currentPage_1__6), 
                         .pagesOuts_1__5 (currentPage_1__5), .pagesOuts_1__4 (
                         currentPage_1__4), .pagesOuts_1__3 (currentPage_1__3), 
                         .pagesOuts_1__2 (currentPage_1__2), .pagesOuts_1__1 (
                         currentPage_1__1), .pagesOuts_1__0 (currentPage_1__0), 
                         .pagesOuts_2__15 (currentPage_2__15), .pagesOuts_2__14 (
                         currentPage_2__14), .pagesOuts_2__13 (currentPage_2__13
                         ), .pagesOuts_2__12 (currentPage_2__12), .pagesOuts_2__11 (
                         currentPage_2__11), .pagesOuts_2__10 (currentPage_2__10
                         ), .pagesOuts_2__9 (currentPage_2__9), .pagesOuts_2__8 (
                         currentPage_2__8), .pagesOuts_2__7 (currentPage_2__7), 
                         .pagesOuts_2__6 (currentPage_2__6), .pagesOuts_2__5 (
                         currentPage_2__5), .pagesOuts_2__4 (currentPage_2__4), 
                         .pagesOuts_2__3 (currentPage_2__3), .pagesOuts_2__2 (
                         currentPage_2__2), .pagesOuts_2__1 (currentPage_2__1), 
                         .pagesOuts_2__0 (currentPage_2__0), .pagesOuts_3__15 (
                         currentPage_3__15), .pagesOuts_3__14 (currentPage_3__14
                         ), .pagesOuts_3__13 (currentPage_3__13), .pagesOuts_3__12 (
                         currentPage_3__12), .pagesOuts_3__11 (currentPage_3__11
                         ), .pagesOuts_3__10 (currentPage_3__10), .pagesOuts_3__9 (
                         currentPage_3__9), .pagesOuts_3__8 (currentPage_3__8), 
                         .pagesOuts_3__7 (currentPage_3__7), .pagesOuts_3__6 (
                         currentPage_3__6), .pagesOuts_3__5 (currentPage_3__5), 
                         .pagesOuts_3__4 (currentPage_3__4), .pagesOuts_3__3 (
                         currentPage_3__3), .pagesOuts_3__2 (currentPage_3__2), 
                         .pagesOuts_3__1 (currentPage_3__1), .pagesOuts_3__0 (
                         currentPage_3__0), .pagesOuts_4__15 (currentPage_4__15)
                         , .pagesOuts_4__14 (currentPage_4__14), .pagesOuts_4__13 (
                         currentPage_4__13), .pagesOuts_4__12 (currentPage_4__12
                         ), .pagesOuts_4__11 (currentPage_4__11), .pagesOuts_4__10 (
                         currentPage_4__10), .pagesOuts_4__9 (currentPage_4__9)
                         , .pagesOuts_4__8 (currentPage_4__8), .pagesOuts_4__7 (
                         currentPage_4__7), .pagesOuts_4__6 (currentPage_4__6), 
                         .pagesOuts_4__5 (currentPage_4__5), .pagesOuts_4__4 (
                         currentPage_4__4), .pagesOuts_4__3 (currentPage_4__3), 
                         .pagesOuts_4__2 (currentPage_4__2), .pagesOuts_4__1 (
                         currentPage_4__1), .pagesOuts_4__0 (currentPage_4__0), 
                         .pagesOuts_5__15 (currentPage_5__15), .pagesOuts_5__14 (
                         currentPage_5__14), .pagesOuts_5__13 (currentPage_5__13
                         ), .pagesOuts_5__12 (currentPage_5__12), .pagesOuts_5__11 (
                         currentPage_5__11), .pagesOuts_5__10 (currentPage_5__10
                         ), .pagesOuts_5__9 (currentPage_5__9), .pagesOuts_5__8 (
                         currentPage_5__8), .pagesOuts_5__7 (currentPage_5__7), 
                         .pagesOuts_5__6 (currentPage_5__6), .pagesOuts_5__5 (
                         currentPage_5__5), .pagesOuts_5__4 (currentPage_5__4), 
                         .pagesOuts_5__3 (currentPage_5__3), .pagesOuts_5__2 (
                         currentPage_5__2), .pagesOuts_5__1 (currentPage_5__1), 
                         .pagesOuts_5__0 (currentPage_5__0), .pagesOuts_6__15 (
                         currentPage_6__15), .pagesOuts_6__14 (currentPage_6__14
                         ), .pagesOuts_6__13 (currentPage_6__13), .pagesOuts_6__12 (
                         currentPage_6__12), .pagesOuts_6__11 (currentPage_6__11
                         ), .pagesOuts_6__10 (currentPage_6__10), .pagesOuts_6__9 (
                         currentPage_6__9), .pagesOuts_6__8 (currentPage_6__8), 
                         .pagesOuts_6__7 (currentPage_6__7), .pagesOuts_6__6 (
                         currentPage_6__6), .pagesOuts_6__5 (currentPage_6__5), 
                         .pagesOuts_6__4 (currentPage_6__4), .pagesOuts_6__3 (
                         currentPage_6__3), .pagesOuts_6__2 (currentPage_6__2), 
                         .pagesOuts_6__1 (currentPage_6__1), .pagesOuts_6__0 (
                         currentPage_6__0), .pagesOuts_7__15 (currentPage_7__15)
                         , .pagesOuts_7__14 (currentPage_7__14), .pagesOuts_7__13 (
                         currentPage_7__13), .pagesOuts_7__12 (currentPage_7__12
                         ), .pagesOuts_7__11 (currentPage_7__11), .pagesOuts_7__10 (
                         currentPage_7__10), .pagesOuts_7__9 (currentPage_7__9)
                         , .pagesOuts_7__8 (currentPage_7__8), .pagesOuts_7__7 (
                         currentPage_7__7), .pagesOuts_7__6 (currentPage_7__6), 
                         .pagesOuts_7__5 (currentPage_7__5), .pagesOuts_7__4 (
                         currentPage_7__4), .pagesOuts_7__3 (currentPage_7__3), 
                         .pagesOuts_7__2 (currentPage_7__2), .pagesOuts_7__1 (
                         currentPage_7__1), .pagesOuts_7__0 (currentPage_7__0), 
                         .pagesOuts_8__15 (currentPage_8__15), .pagesOuts_8__14 (
                         currentPage_8__14), .pagesOuts_8__13 (currentPage_8__13
                         ), .pagesOuts_8__12 (currentPage_8__12), .pagesOuts_8__11 (
                         currentPage_8__11), .pagesOuts_8__10 (currentPage_8__10
                         ), .pagesOuts_8__9 (currentPage_8__9), .pagesOuts_8__8 (
                         currentPage_8__8), .pagesOuts_8__7 (currentPage_8__7), 
                         .pagesOuts_8__6 (currentPage_8__6), .pagesOuts_8__5 (
                         currentPage_8__5), .pagesOuts_8__4 (currentPage_8__4), 
                         .pagesOuts_8__3 (currentPage_8__3), .pagesOuts_8__2 (
                         currentPage_8__2), .pagesOuts_8__1 (currentPage_8__1), 
                         .pagesOuts_8__0 (currentPage_8__0), .pagesOuts_9__15 (
                         currentPage_9__15), .pagesOuts_9__14 (currentPage_9__14
                         ), .pagesOuts_9__13 (currentPage_9__13), .pagesOuts_9__12 (
                         currentPage_9__12), .pagesOuts_9__11 (currentPage_9__11
                         ), .pagesOuts_9__10 (currentPage_9__10), .pagesOuts_9__9 (
                         currentPage_9__9), .pagesOuts_9__8 (currentPage_9__8), 
                         .pagesOuts_9__7 (currentPage_9__7), .pagesOuts_9__6 (
                         currentPage_9__6), .pagesOuts_9__5 (currentPage_9__5), 
                         .pagesOuts_9__4 (currentPage_9__4), .pagesOuts_9__3 (
                         currentPage_9__3), .pagesOuts_9__2 (currentPage_9__2), 
                         .pagesOuts_9__1 (currentPage_9__1), .pagesOuts_9__0 (
                         currentPage_9__0), .pagesOuts_10__15 (
                         currentPage_10__15), .pagesOuts_10__14 (
                         currentPage_10__14), .pagesOuts_10__13 (
                         currentPage_10__13), .pagesOuts_10__12 (
                         currentPage_10__12), .pagesOuts_10__11 (
                         currentPage_10__11), .pagesOuts_10__10 (
                         currentPage_10__10), .pagesOuts_10__9 (
                         currentPage_10__9), .pagesOuts_10__8 (currentPage_10__8
                         ), .pagesOuts_10__7 (currentPage_10__7), .pagesOuts_10__6 (
                         currentPage_10__6), .pagesOuts_10__5 (currentPage_10__5
                         ), .pagesOuts_10__4 (currentPage_10__4), .pagesOuts_10__3 (
                         currentPage_10__3), .pagesOuts_10__2 (currentPage_10__2
                         ), .pagesOuts_10__1 (currentPage_10__1), .pagesOuts_10__0 (
                         currentPage_10__0), .pagesOuts_11__15 (
                         currentPage_11__15), .pagesOuts_11__14 (
                         currentPage_11__14), .pagesOuts_11__13 (
                         currentPage_11__13), .pagesOuts_11__12 (
                         currentPage_11__12), .pagesOuts_11__11 (
                         currentPage_11__11), .pagesOuts_11__10 (
                         currentPage_11__10), .pagesOuts_11__9 (
                         currentPage_11__9), .pagesOuts_11__8 (currentPage_11__8
                         ), .pagesOuts_11__7 (currentPage_11__7), .pagesOuts_11__6 (
                         currentPage_11__6), .pagesOuts_11__5 (currentPage_11__5
                         ), .pagesOuts_11__4 (currentPage_11__4), .pagesOuts_11__3 (
                         currentPage_11__3), .pagesOuts_11__2 (currentPage_11__2
                         ), .pagesOuts_11__1 (currentPage_11__1), .pagesOuts_11__0 (
                         currentPage_11__0), .pagesOuts_12__15 (
                         currentPage_12__15), .pagesOuts_12__14 (
                         currentPage_12__14), .pagesOuts_12__13 (
                         currentPage_12__13), .pagesOuts_12__12 (
                         currentPage_12__12), .pagesOuts_12__11 (
                         currentPage_12__11), .pagesOuts_12__10 (
                         currentPage_12__10), .pagesOuts_12__9 (
                         currentPage_12__9), .pagesOuts_12__8 (currentPage_12__8
                         ), .pagesOuts_12__7 (currentPage_12__7), .pagesOuts_12__6 (
                         currentPage_12__6), .pagesOuts_12__5 (currentPage_12__5
                         ), .pagesOuts_12__4 (currentPage_12__4), .pagesOuts_12__3 (
                         currentPage_12__3), .pagesOuts_12__2 (currentPage_12__2
                         ), .pagesOuts_12__1 (currentPage_12__1), .pagesOuts_12__0 (
                         currentPage_12__0), .pagesOuts_13__15 (
                         currentPage_13__15), .pagesOuts_13__14 (
                         currentPage_13__14), .pagesOuts_13__13 (
                         currentPage_13__13), .pagesOuts_13__12 (
                         currentPage_13__12), .pagesOuts_13__11 (
                         currentPage_13__11), .pagesOuts_13__10 (
                         currentPage_13__10), .pagesOuts_13__9 (
                         currentPage_13__9), .pagesOuts_13__8 (currentPage_13__8
                         ), .pagesOuts_13__7 (currentPage_13__7), .pagesOuts_13__6 (
                         currentPage_13__6), .pagesOuts_13__5 (currentPage_13__5
                         ), .pagesOuts_13__4 (currentPage_13__4), .pagesOuts_13__3 (
                         currentPage_13__3), .pagesOuts_13__2 (currentPage_13__2
                         ), .pagesOuts_13__1 (currentPage_13__1), .pagesOuts_13__0 (
                         currentPage_13__0), .pagesOuts_14__15 (
                         currentPage_14__15), .pagesOuts_14__14 (
                         currentPage_14__14), .pagesOuts_14__13 (
                         currentPage_14__13), .pagesOuts_14__12 (
                         currentPage_14__12), .pagesOuts_14__11 (
                         currentPage_14__11), .pagesOuts_14__10 (
                         currentPage_14__10), .pagesOuts_14__9 (
                         currentPage_14__9), .pagesOuts_14__8 (currentPage_14__8
                         ), .pagesOuts_14__7 (currentPage_14__7), .pagesOuts_14__6 (
                         currentPage_14__6), .pagesOuts_14__5 (currentPage_14__5
                         ), .pagesOuts_14__4 (currentPage_14__4), .pagesOuts_14__3 (
                         currentPage_14__3), .pagesOuts_14__2 (currentPage_14__2
                         ), .pagesOuts_14__1 (currentPage_14__1), .pagesOuts_14__0 (
                         currentPage_14__0), .pagesOuts_15__15 (
                         currentPage_15__15), .pagesOuts_15__14 (
                         currentPage_15__14), .pagesOuts_15__13 (
                         currentPage_15__13), .pagesOuts_15__12 (
                         currentPage_15__12), .pagesOuts_15__11 (
                         currentPage_15__11), .pagesOuts_15__10 (
                         currentPage_15__10), .pagesOuts_15__9 (
                         currentPage_15__9), .pagesOuts_15__8 (currentPage_15__8
                         ), .pagesOuts_15__7 (currentPage_15__7), .pagesOuts_15__6 (
                         currentPage_15__6), .pagesOuts_15__5 (currentPage_15__5
                         ), .pagesOuts_15__4 (currentPage_15__4), .pagesOuts_15__3 (
                         currentPage_15__3), .pagesOuts_15__2 (currentPage_15__2
                         ), .pagesOuts_15__1 (currentPage_15__1), .pagesOuts_15__0 (
                         currentPage_15__0), .pagesOuts_16__15 (
                         currentPage_16__15), .pagesOuts_16__14 (
                         currentPage_16__14), .pagesOuts_16__13 (
                         currentPage_16__13), .pagesOuts_16__12 (
                         currentPage_16__12), .pagesOuts_16__11 (
                         currentPage_16__11), .pagesOuts_16__10 (
                         currentPage_16__10), .pagesOuts_16__9 (
                         currentPage_16__9), .pagesOuts_16__8 (currentPage_16__8
                         ), .pagesOuts_16__7 (currentPage_16__7), .pagesOuts_16__6 (
                         currentPage_16__6), .pagesOuts_16__5 (currentPage_16__5
                         ), .pagesOuts_16__4 (currentPage_16__4), .pagesOuts_16__3 (
                         currentPage_16__3), .pagesOuts_16__2 (currentPage_16__2
                         ), .pagesOuts_16__1 (currentPage_16__1), .pagesOuts_16__0 (
                         currentPage_16__0), .pagesOuts_17__15 (
                         currentPage_17__15), .pagesOuts_17__14 (
                         currentPage_17__14), .pagesOuts_17__13 (
                         currentPage_17__13), .pagesOuts_17__12 (
                         currentPage_17__12), .pagesOuts_17__11 (
                         currentPage_17__11), .pagesOuts_17__10 (
                         currentPage_17__10), .pagesOuts_17__9 (
                         currentPage_17__9), .pagesOuts_17__8 (currentPage_17__8
                         ), .pagesOuts_17__7 (currentPage_17__7), .pagesOuts_17__6 (
                         currentPage_17__6), .pagesOuts_17__5 (currentPage_17__5
                         ), .pagesOuts_17__4 (currentPage_17__4), .pagesOuts_17__3 (
                         currentPage_17__3), .pagesOuts_17__2 (currentPage_17__2
                         ), .pagesOuts_17__1 (currentPage_17__1), .pagesOuts_17__0 (
                         currentPage_17__0), .pagesOuts_18__15 (
                         currentPage_18__15), .pagesOuts_18__14 (
                         currentPage_18__14), .pagesOuts_18__13 (
                         currentPage_18__13), .pagesOuts_18__12 (
                         currentPage_18__12), .pagesOuts_18__11 (
                         currentPage_18__11), .pagesOuts_18__10 (
                         currentPage_18__10), .pagesOuts_18__9 (
                         currentPage_18__9), .pagesOuts_18__8 (currentPage_18__8
                         ), .pagesOuts_18__7 (currentPage_18__7), .pagesOuts_18__6 (
                         currentPage_18__6), .pagesOuts_18__5 (currentPage_18__5
                         ), .pagesOuts_18__4 (currentPage_18__4), .pagesOuts_18__3 (
                         currentPage_18__3), .pagesOuts_18__2 (currentPage_18__2
                         ), .pagesOuts_18__1 (currentPage_18__1), .pagesOuts_18__0 (
                         currentPage_18__0), .pagesOuts_19__15 (
                         currentPage_19__15), .pagesOuts_19__14 (
                         currentPage_19__14), .pagesOuts_19__13 (
                         currentPage_19__13), .pagesOuts_19__12 (
                         currentPage_19__12), .pagesOuts_19__11 (
                         currentPage_19__11), .pagesOuts_19__10 (
                         currentPage_19__10), .pagesOuts_19__9 (
                         currentPage_19__9), .pagesOuts_19__8 (currentPage_19__8
                         ), .pagesOuts_19__7 (currentPage_19__7), .pagesOuts_19__6 (
                         currentPage_19__6), .pagesOuts_19__5 (currentPage_19__5
                         ), .pagesOuts_19__4 (currentPage_19__4), .pagesOuts_19__3 (
                         currentPage_19__3), .pagesOuts_19__2 (currentPage_19__2
                         ), .pagesOuts_19__1 (currentPage_19__1), .pagesOuts_19__0 (
                         currentPage_19__0), .pagesOuts_20__15 (
                         currentPage_20__15), .pagesOuts_20__14 (
                         currentPage_20__14), .pagesOuts_20__13 (
                         currentPage_20__13), .pagesOuts_20__12 (
                         currentPage_20__12), .pagesOuts_20__11 (
                         currentPage_20__11), .pagesOuts_20__10 (
                         currentPage_20__10), .pagesOuts_20__9 (
                         currentPage_20__9), .pagesOuts_20__8 (currentPage_20__8
                         ), .pagesOuts_20__7 (currentPage_20__7), .pagesOuts_20__6 (
                         currentPage_20__6), .pagesOuts_20__5 (currentPage_20__5
                         ), .pagesOuts_20__4 (currentPage_20__4), .pagesOuts_20__3 (
                         currentPage_20__3), .pagesOuts_20__2 (currentPage_20__2
                         ), .pagesOuts_20__1 (currentPage_20__1), .pagesOuts_20__0 (
                         currentPage_20__0), .pagesOuts_21__15 (
                         currentPage_21__15), .pagesOuts_21__14 (
                         currentPage_21__14), .pagesOuts_21__13 (
                         currentPage_21__13), .pagesOuts_21__12 (
                         currentPage_21__12), .pagesOuts_21__11 (
                         currentPage_21__11), .pagesOuts_21__10 (
                         currentPage_21__10), .pagesOuts_21__9 (
                         currentPage_21__9), .pagesOuts_21__8 (currentPage_21__8
                         ), .pagesOuts_21__7 (currentPage_21__7), .pagesOuts_21__6 (
                         currentPage_21__6), .pagesOuts_21__5 (currentPage_21__5
                         ), .pagesOuts_21__4 (currentPage_21__4), .pagesOuts_21__3 (
                         currentPage_21__3), .pagesOuts_21__2 (currentPage_21__2
                         ), .pagesOuts_21__1 (currentPage_21__1), .pagesOuts_21__0 (
                         currentPage_21__0), .pagesOuts_22__15 (
                         currentPage_22__15), .pagesOuts_22__14 (
                         currentPage_22__14), .pagesOuts_22__13 (
                         currentPage_22__13), .pagesOuts_22__12 (
                         currentPage_22__12), .pagesOuts_22__11 (
                         currentPage_22__11), .pagesOuts_22__10 (
                         currentPage_22__10), .pagesOuts_22__9 (
                         currentPage_22__9), .pagesOuts_22__8 (currentPage_22__8
                         ), .pagesOuts_22__7 (currentPage_22__7), .pagesOuts_22__6 (
                         currentPage_22__6), .pagesOuts_22__5 (currentPage_22__5
                         ), .pagesOuts_22__4 (currentPage_22__4), .pagesOuts_22__3 (
                         currentPage_22__3), .pagesOuts_22__2 (currentPage_22__2
                         ), .pagesOuts_22__1 (currentPage_22__1), .pagesOuts_22__0 (
                         currentPage_22__0), .pagesOuts_23__15 (
                         currentPage_23__15), .pagesOuts_23__14 (
                         currentPage_23__14), .pagesOuts_23__13 (
                         currentPage_23__13), .pagesOuts_23__12 (
                         currentPage_23__12), .pagesOuts_23__11 (
                         currentPage_23__11), .pagesOuts_23__10 (
                         currentPage_23__10), .pagesOuts_23__9 (
                         currentPage_23__9), .pagesOuts_23__8 (currentPage_23__8
                         ), .pagesOuts_23__7 (currentPage_23__7), .pagesOuts_23__6 (
                         currentPage_23__6), .pagesOuts_23__5 (currentPage_23__5
                         ), .pagesOuts_23__4 (currentPage_23__4), .pagesOuts_23__3 (
                         currentPage_23__3), .pagesOuts_23__2 (currentPage_23__2
                         ), .pagesOuts_23__1 (currentPage_23__1), .pagesOuts_23__0 (
                         currentPage_23__0), .pagesOuts_24__15 (
                         currentPage_24__15), .pagesOuts_24__14 (
                         currentPage_24__14), .pagesOuts_24__13 (
                         currentPage_24__13), .pagesOuts_24__12 (
                         currentPage_24__12), .pagesOuts_24__11 (
                         currentPage_24__11), .pagesOuts_24__10 (
                         currentPage_24__10), .pagesOuts_24__9 (
                         currentPage_24__9), .pagesOuts_24__8 (currentPage_24__8
                         ), .pagesOuts_24__7 (currentPage_24__7), .pagesOuts_24__6 (
                         currentPage_24__6), .pagesOuts_24__5 (currentPage_24__5
                         ), .pagesOuts_24__4 (currentPage_24__4), .pagesOuts_24__3 (
                         currentPage_24__3), .pagesOuts_24__2 (currentPage_24__2
                         ), .pagesOuts_24__1 (currentPage_24__1), .pagesOuts_24__0 (
                         currentPage_24__0), .filtersOuts_0__7 (filter_0__7), .filtersOuts_0__6 (
                         filter_0__6), .filtersOuts_0__5 (filter_0__5), .filtersOuts_0__4 (
                         filter_0__4), .filtersOuts_0__3 (filter_0__3), .filtersOuts_0__2 (
                         filter_0__2), .filtersOuts_0__1 (filter_0__1), .filtersOuts_0__0 (
                         filter_0__0), .filtersOuts_1__7 (filter_1__7), .filtersOuts_1__6 (
                         filter_1__6), .filtersOuts_1__5 (filter_1__5), .filtersOuts_1__4 (
                         filter_1__4), .filtersOuts_1__3 (filter_1__3), .filtersOuts_1__2 (
                         filter_1__2), .filtersOuts_1__1 (filter_1__1), .filtersOuts_1__0 (
                         filter_1__0), .filtersOuts_2__7 (filter_2__7), .filtersOuts_2__6 (
                         filter_2__6), .filtersOuts_2__5 (filter_2__5), .filtersOuts_2__4 (
                         filter_2__4), .filtersOuts_2__3 (filter_2__3), .filtersOuts_2__2 (
                         filter_2__2), .filtersOuts_2__1 (filter_2__1), .filtersOuts_2__0 (
                         filter_2__0), .filtersOuts_3__7 (filter_3__7), .filtersOuts_3__6 (
                         filter_3__6), .filtersOuts_3__5 (filter_3__5), .filtersOuts_3__4 (
                         filter_3__4), .filtersOuts_3__3 (filter_3__3), .filtersOuts_3__2 (
                         filter_3__2), .filtersOuts_3__1 (filter_3__1), .filtersOuts_3__0 (
                         filter_3__0), .filtersOuts_4__7 (filter_4__7), .filtersOuts_4__6 (
                         filter_4__6), .filtersOuts_4__5 (filter_4__5), .filtersOuts_4__4 (
                         filter_4__4), .filtersOuts_4__3 (filter_4__3), .filtersOuts_4__2 (
                         filter_4__2), .filtersOuts_4__1 (filter_4__1), .filtersOuts_4__0 (
                         filter_4__0), .filtersOuts_5__7 (filter_5__7), .filtersOuts_5__6 (
                         filter_5__6), .filtersOuts_5__5 (filter_5__5), .filtersOuts_5__4 (
                         filter_5__4), .filtersOuts_5__3 (filter_5__3), .filtersOuts_5__2 (
                         filter_5__2), .filtersOuts_5__1 (filter_5__1), .filtersOuts_5__0 (
                         filter_5__0), .filtersOuts_6__7 (filter_6__7), .filtersOuts_6__6 (
                         filter_6__6), .filtersOuts_6__5 (filter_6__5), .filtersOuts_6__4 (
                         filter_6__4), .filtersOuts_6__3 (filter_6__3), .filtersOuts_6__2 (
                         filter_6__2), .filtersOuts_6__1 (filter_6__1), .filtersOuts_6__0 (
                         filter_6__0), .filtersOuts_7__7 (filter_7__7), .filtersOuts_7__6 (
                         filter_7__6), .filtersOuts_7__5 (filter_7__5), .filtersOuts_7__4 (
                         filter_7__4), .filtersOuts_7__3 (filter_7__3), .filtersOuts_7__2 (
                         filter_7__2), .filtersOuts_7__1 (filter_7__1), .filtersOuts_7__0 (
                         filter_7__0), .filtersOuts_8__7 (filter_8__7), .filtersOuts_8__6 (
                         filter_8__6), .filtersOuts_8__5 (filter_8__5), .filtersOuts_8__4 (
                         filter_8__4), .filtersOuts_8__3 (filter_8__3), .filtersOuts_8__2 (
                         filter_8__2), .filtersOuts_8__1 (filter_8__1), .filtersOuts_8__0 (
                         filter_8__0), .filtersOuts_9__7 (filter_9__7), .filtersOuts_9__6 (
                         filter_9__6), .filtersOuts_9__5 (filter_9__5), .filtersOuts_9__4 (
                         filter_9__4), .filtersOuts_9__3 (filter_9__3), .filtersOuts_9__2 (
                         filter_9__2), .filtersOuts_9__1 (filter_9__1), .filtersOuts_9__0 (
                         filter_9__0), .filtersOuts_10__7 (filter_10__7), .filtersOuts_10__6 (
                         filter_10__6), .filtersOuts_10__5 (filter_10__5), .filtersOuts_10__4 (
                         filter_10__4), .filtersOuts_10__3 (filter_10__3), .filtersOuts_10__2 (
                         filter_10__2), .filtersOuts_10__1 (filter_10__1), .filtersOuts_10__0 (
                         filter_10__0), .filtersOuts_11__7 (filter_11__7), .filtersOuts_11__6 (
                         filter_11__6), .filtersOuts_11__5 (filter_11__5), .filtersOuts_11__4 (
                         filter_11__4), .filtersOuts_11__3 (filter_11__3), .filtersOuts_11__2 (
                         filter_11__2), .filtersOuts_11__1 (filter_11__1), .filtersOuts_11__0 (
                         filter_11__0), .filtersOuts_12__7 (filter_12__7), .filtersOuts_12__6 (
                         filter_12__6), .filtersOuts_12__5 (filter_12__5), .filtersOuts_12__4 (
                         filter_12__4), .filtersOuts_12__3 (filter_12__3), .filtersOuts_12__2 (
                         filter_12__2), .filtersOuts_12__1 (filter_12__1), .filtersOuts_12__0 (
                         filter_12__0), .filtersOuts_13__7 (filter_13__7), .filtersOuts_13__6 (
                         filter_13__6), .filtersOuts_13__5 (filter_13__5), .filtersOuts_13__4 (
                         filter_13__4), .filtersOuts_13__3 (filter_13__3), .filtersOuts_13__2 (
                         filter_13__2), .filtersOuts_13__1 (filter_13__1), .filtersOuts_13__0 (
                         filter_13__0), .filtersOuts_14__7 (filter_14__7), .filtersOuts_14__6 (
                         filter_14__6), .filtersOuts_14__5 (filter_14__5), .filtersOuts_14__4 (
                         filter_14__4), .filtersOuts_14__3 (filter_14__3), .filtersOuts_14__2 (
                         filter_14__2), .filtersOuts_14__1 (filter_14__1), .filtersOuts_14__0 (
                         filter_14__0), .filtersOuts_15__7 (filter_15__7), .filtersOuts_15__6 (
                         filter_15__6), .filtersOuts_15__5 (filter_15__5), .filtersOuts_15__4 (
                         filter_15__4), .filtersOuts_15__3 (filter_15__3), .filtersOuts_15__2 (
                         filter_15__2), .filtersOuts_15__1 (filter_15__1), .filtersOuts_15__0 (
                         filter_15__0), .filtersOuts_16__7 (filter_16__7), .filtersOuts_16__6 (
                         filter_16__6), .filtersOuts_16__5 (filter_16__5), .filtersOuts_16__4 (
                         filter_16__4), .filtersOuts_16__3 (filter_16__3), .filtersOuts_16__2 (
                         filter_16__2), .filtersOuts_16__1 (filter_16__1), .filtersOuts_16__0 (
                         filter_16__0), .filtersOuts_17__7 (filter_17__7), .filtersOuts_17__6 (
                         filter_17__6), .filtersOuts_17__5 (filter_17__5), .filtersOuts_17__4 (
                         filter_17__4), .filtersOuts_17__3 (filter_17__3), .filtersOuts_17__2 (
                         filter_17__2), .filtersOuts_17__1 (filter_17__1), .filtersOuts_17__0 (
                         filter_17__0), .filtersOuts_18__7 (filter_18__7), .filtersOuts_18__6 (
                         filter_18__6), .filtersOuts_18__5 (filter_18__5), .filtersOuts_18__4 (
                         filter_18__4), .filtersOuts_18__3 (filter_18__3), .filtersOuts_18__2 (
                         filter_18__2), .filtersOuts_18__1 (filter_18__1), .filtersOuts_18__0 (
                         filter_18__0), .filtersOuts_19__7 (filter_19__7), .filtersOuts_19__6 (
                         filter_19__6), .filtersOuts_19__5 (filter_19__5), .filtersOuts_19__4 (
                         filter_19__4), .filtersOuts_19__3 (filter_19__3), .filtersOuts_19__2 (
                         filter_19__2), .filtersOuts_19__1 (filter_19__1), .filtersOuts_19__0 (
                         filter_19__0), .filtersOuts_20__7 (filter_20__7), .filtersOuts_20__6 (
                         filter_20__6), .filtersOuts_20__5 (filter_20__5), .filtersOuts_20__4 (
                         filter_20__4), .filtersOuts_20__3 (filter_20__3), .filtersOuts_20__2 (
                         filter_20__2), .filtersOuts_20__1 (filter_20__1), .filtersOuts_20__0 (
                         filter_20__0), .filtersOuts_21__7 (filter_21__7), .filtersOuts_21__6 (
                         filter_21__6), .filtersOuts_21__5 (filter_21__5), .filtersOuts_21__4 (
                         filter_21__4), .filtersOuts_21__3 (filter_21__3), .filtersOuts_21__2 (
                         filter_21__2), .filtersOuts_21__1 (filter_21__1), .filtersOuts_21__0 (
                         filter_21__0), .filtersOuts_22__7 (filter_22__7), .filtersOuts_22__6 (
                         filter_22__6), .filtersOuts_22__5 (filter_22__5), .filtersOuts_22__4 (
                         filter_22__4), .filtersOuts_22__3 (filter_22__3), .filtersOuts_22__2 (
                         filter_22__2), .filtersOuts_22__1 (filter_22__1), .filtersOuts_22__0 (
                         filter_22__0), .filtersOuts_23__7 (filter_23__7), .filtersOuts_23__6 (
                         filter_23__6), .filtersOuts_23__5 (filter_23__5), .filtersOuts_23__4 (
                         filter_23__4), .filtersOuts_23__3 (filter_23__3), .filtersOuts_23__2 (
                         filter_23__2), .filtersOuts_23__1 (filter_23__1), .filtersOuts_23__0 (
                         filter_23__0), .filtersOuts_24__7 (filter_24__7), .filtersOuts_24__6 (
                         filter_24__6), .filtersOuts_24__5 (filter_24__5), .filtersOuts_24__4 (
                         filter_24__4), .filtersOuts_24__3 (filter_24__3), .filtersOuts_24__2 (
                         filter_24__2), .filtersOuts_24__1 (filter_24__1), .filtersOuts_24__0 (
                         filter_24__0)) ;
    CNNMuls_25 mulsMap (.filter_24__7 (filter_0__7), .filter_24__6 (filter_0__6)
               , .filter_24__5 (filter_0__5), .filter_24__4 (filter_0__4), .filter_24__3 (
               filter_0__3), .filter_24__2 (filter_0__2), .filter_24__1 (
               filter_0__1), .filter_24__0 (filter_0__0), .filter_23__7 (
               filter_1__7), .filter_23__6 (filter_1__6), .filter_23__5 (
               filter_1__5), .filter_23__4 (filter_1__4), .filter_23__3 (
               filter_1__3), .filter_23__2 (filter_1__2), .filter_23__1 (
               filter_1__1), .filter_23__0 (filter_1__0), .filter_22__7 (
               filter_2__7), .filter_22__6 (filter_2__6), .filter_22__5 (
               filter_2__5), .filter_22__4 (filter_2__4), .filter_22__3 (
               filter_2__3), .filter_22__2 (filter_2__2), .filter_22__1 (
               filter_2__1), .filter_22__0 (filter_2__0), .filter_21__7 (
               filter_3__7), .filter_21__6 (filter_3__6), .filter_21__5 (
               filter_3__5), .filter_21__4 (filter_3__4), .filter_21__3 (
               filter_3__3), .filter_21__2 (filter_3__2), .filter_21__1 (
               filter_3__1), .filter_21__0 (filter_3__0), .filter_20__7 (
               filter_4__7), .filter_20__6 (filter_4__6), .filter_20__5 (
               filter_4__5), .filter_20__4 (filter_4__4), .filter_20__3 (
               filter_4__3), .filter_20__2 (filter_4__2), .filter_20__1 (
               filter_4__1), .filter_20__0 (filter_4__0), .filter_19__7 (
               filter_5__7), .filter_19__6 (filter_5__6), .filter_19__5 (
               filter_5__5), .filter_19__4 (filter_5__4), .filter_19__3 (
               filter_5__3), .filter_19__2 (filter_5__2), .filter_19__1 (
               filter_5__1), .filter_19__0 (filter_5__0), .filter_18__7 (
               filter_6__7), .filter_18__6 (filter_6__6), .filter_18__5 (
               filter_6__5), .filter_18__4 (filter_6__4), .filter_18__3 (
               filter_6__3), .filter_18__2 (filter_6__2), .filter_18__1 (
               filter_6__1), .filter_18__0 (filter_6__0), .filter_17__7 (
               filter_7__7), .filter_17__6 (filter_7__6), .filter_17__5 (
               filter_7__5), .filter_17__4 (filter_7__4), .filter_17__3 (
               filter_7__3), .filter_17__2 (filter_7__2), .filter_17__1 (
               filter_7__1), .filter_17__0 (filter_7__0), .filter_16__7 (
               filter_8__7), .filter_16__6 (filter_8__6), .filter_16__5 (
               filter_8__5), .filter_16__4 (filter_8__4), .filter_16__3 (
               filter_8__3), .filter_16__2 (filter_8__2), .filter_16__1 (
               filter_8__1), .filter_16__0 (filter_8__0), .filter_15__7 (
               filter_9__7), .filter_15__6 (filter_9__6), .filter_15__5 (
               filter_9__5), .filter_15__4 (filter_9__4), .filter_15__3 (
               filter_9__3), .filter_15__2 (filter_9__2), .filter_15__1 (
               filter_9__1), .filter_15__0 (filter_9__0), .filter_14__7 (
               filter_10__7), .filter_14__6 (filter_10__6), .filter_14__5 (
               filter_10__5), .filter_14__4 (filter_10__4), .filter_14__3 (
               filter_10__3), .filter_14__2 (filter_10__2), .filter_14__1 (
               filter_10__1), .filter_14__0 (filter_10__0), .filter_13__7 (
               filter_11__7), .filter_13__6 (filter_11__6), .filter_13__5 (
               filter_11__5), .filter_13__4 (filter_11__4), .filter_13__3 (
               filter_11__3), .filter_13__2 (filter_11__2), .filter_13__1 (
               filter_11__1), .filter_13__0 (filter_11__0), .filter_12__7 (
               filter_12__7), .filter_12__6 (filter_12__6), .filter_12__5 (
               filter_12__5), .filter_12__4 (filter_12__4), .filter_12__3 (
               filter_12__3), .filter_12__2 (filter_12__2), .filter_12__1 (
               filter_12__1), .filter_12__0 (filter_12__0), .filter_11__7 (
               filter_13__7), .filter_11__6 (filter_13__6), .filter_11__5 (
               filter_13__5), .filter_11__4 (filter_13__4), .filter_11__3 (
               filter_13__3), .filter_11__2 (filter_13__2), .filter_11__1 (
               filter_13__1), .filter_11__0 (filter_13__0), .filter_10__7 (
               filter_14__7), .filter_10__6 (filter_14__6), .filter_10__5 (
               filter_14__5), .filter_10__4 (filter_14__4), .filter_10__3 (
               filter_14__3), .filter_10__2 (filter_14__2), .filter_10__1 (
               filter_14__1), .filter_10__0 (filter_14__0), .filter_9__7 (
               filter_15__7), .filter_9__6 (filter_15__6), .filter_9__5 (
               filter_15__5), .filter_9__4 (filter_15__4), .filter_9__3 (
               filter_15__3), .filter_9__2 (filter_15__2), .filter_9__1 (
               filter_15__1), .filter_9__0 (filter_15__0), .filter_8__7 (
               filter_16__7), .filter_8__6 (filter_16__6), .filter_8__5 (
               filter_16__5), .filter_8__4 (filter_16__4), .filter_8__3 (
               filter_16__3), .filter_8__2 (filter_16__2), .filter_8__1 (
               filter_16__1), .filter_8__0 (filter_16__0), .filter_7__7 (
               filter_17__7), .filter_7__6 (filter_17__6), .filter_7__5 (
               filter_17__5), .filter_7__4 (filter_17__4), .filter_7__3 (
               filter_17__3), .filter_7__2 (filter_17__2), .filter_7__1 (
               filter_17__1), .filter_7__0 (filter_17__0), .filter_6__7 (
               filter_18__7), .filter_6__6 (filter_18__6), .filter_6__5 (
               filter_18__5), .filter_6__4 (filter_18__4), .filter_6__3 (
               filter_18__3), .filter_6__2 (filter_18__2), .filter_6__1 (
               filter_18__1), .filter_6__0 (filter_18__0), .filter_5__7 (
               filter_19__7), .filter_5__6 (filter_19__6), .filter_5__5 (
               filter_19__5), .filter_5__4 (filter_19__4), .filter_5__3 (
               filter_19__3), .filter_5__2 (filter_19__2), .filter_5__1 (
               filter_19__1), .filter_5__0 (filter_19__0), .filter_4__7 (
               filter_20__7), .filter_4__6 (filter_20__6), .filter_4__5 (
               filter_20__5), .filter_4__4 (filter_20__4), .filter_4__3 (
               filter_20__3), .filter_4__2 (filter_20__2), .filter_4__1 (
               filter_20__1), .filter_4__0 (filter_20__0), .filter_3__7 (
               filter_21__7), .filter_3__6 (filter_21__6), .filter_3__5 (
               filter_21__5), .filter_3__4 (filter_21__4), .filter_3__3 (
               filter_21__3), .filter_3__2 (filter_21__2), .filter_3__1 (
               filter_21__1), .filter_3__0 (filter_21__0), .filter_2__7 (
               filter_22__7), .filter_2__6 (filter_22__6), .filter_2__5 (
               filter_22__5), .filter_2__4 (filter_22__4), .filter_2__3 (
               filter_22__3), .filter_2__2 (filter_22__2), .filter_2__1 (
               filter_22__1), .filter_2__0 (filter_22__0), .filter_1__7 (
               filter_23__7), .filter_1__6 (filter_23__6), .filter_1__5 (
               filter_23__5), .filter_1__4 (filter_23__4), .filter_1__3 (
               filter_23__3), .filter_1__2 (filter_23__2), .filter_1__1 (
               filter_23__1), .filter_1__0 (filter_23__0), .filter_0__7 (
               filter_24__7), .filter_0__6 (filter_24__6), .filter_0__5 (
               filter_24__5), .filter_0__4 (filter_24__4), .filter_0__3 (
               filter_24__3), .filter_0__2 (filter_24__2), .filter_0__1 (
               filter_24__1), .filter_0__0 (filter_24__0), .window_24__15 (
               currentPage_0__15), .window_24__14 (currentPage_0__14), .window_24__13 (
               currentPage_0__13), .window_24__12 (currentPage_0__12), .window_24__11 (
               currentPage_0__11), .window_24__10 (currentPage_0__10), .window_24__9 (
               currentPage_0__9), .window_24__8 (currentPage_0__8), .window_24__7 (
               currentPage_0__7), .window_24__6 (currentPage_0__6), .window_24__5 (
               currentPage_0__5), .window_24__4 (currentPage_0__4), .window_24__3 (
               currentPage_0__3), .window_24__2 (currentPage_0__2), .window_24__1 (
               currentPage_0__1), .window_24__0 (currentPage_0__0), .window_23__15 (
               currentPage_1__15), .window_23__14 (currentPage_1__14), .window_23__13 (
               currentPage_1__13), .window_23__12 (currentPage_1__12), .window_23__11 (
               currentPage_1__11), .window_23__10 (currentPage_1__10), .window_23__9 (
               currentPage_1__9), .window_23__8 (currentPage_1__8), .window_23__7 (
               currentPage_1__7), .window_23__6 (currentPage_1__6), .window_23__5 (
               currentPage_1__5), .window_23__4 (currentPage_1__4), .window_23__3 (
               currentPage_1__3), .window_23__2 (currentPage_1__2), .window_23__1 (
               currentPage_1__1), .window_23__0 (currentPage_1__0), .window_22__15 (
               currentPage_2__15), .window_22__14 (currentPage_2__14), .window_22__13 (
               currentPage_2__13), .window_22__12 (currentPage_2__12), .window_22__11 (
               currentPage_2__11), .window_22__10 (currentPage_2__10), .window_22__9 (
               currentPage_2__9), .window_22__8 (currentPage_2__8), .window_22__7 (
               currentPage_2__7), .window_22__6 (currentPage_2__6), .window_22__5 (
               currentPage_2__5), .window_22__4 (currentPage_2__4), .window_22__3 (
               currentPage_2__3), .window_22__2 (currentPage_2__2), .window_22__1 (
               currentPage_2__1), .window_22__0 (currentPage_2__0), .window_21__15 (
               currentPage_3__15), .window_21__14 (currentPage_3__14), .window_21__13 (
               currentPage_3__13), .window_21__12 (currentPage_3__12), .window_21__11 (
               currentPage_3__11), .window_21__10 (currentPage_3__10), .window_21__9 (
               currentPage_3__9), .window_21__8 (currentPage_3__8), .window_21__7 (
               currentPage_3__7), .window_21__6 (currentPage_3__6), .window_21__5 (
               currentPage_3__5), .window_21__4 (currentPage_3__4), .window_21__3 (
               currentPage_3__3), .window_21__2 (currentPage_3__2), .window_21__1 (
               currentPage_3__1), .window_21__0 (currentPage_3__0), .window_20__15 (
               currentPage_4__15), .window_20__14 (currentPage_4__14), .window_20__13 (
               currentPage_4__13), .window_20__12 (currentPage_4__12), .window_20__11 (
               currentPage_4__11), .window_20__10 (currentPage_4__10), .window_20__9 (
               currentPage_4__9), .window_20__8 (currentPage_4__8), .window_20__7 (
               currentPage_4__7), .window_20__6 (currentPage_4__6), .window_20__5 (
               currentPage_4__5), .window_20__4 (currentPage_4__4), .window_20__3 (
               currentPage_4__3), .window_20__2 (currentPage_4__2), .window_20__1 (
               currentPage_4__1), .window_20__0 (currentPage_4__0), .window_19__15 (
               currentPage_5__15), .window_19__14 (currentPage_5__14), .window_19__13 (
               currentPage_5__13), .window_19__12 (currentPage_5__12), .window_19__11 (
               currentPage_5__11), .window_19__10 (currentPage_5__10), .window_19__9 (
               currentPage_5__9), .window_19__8 (currentPage_5__8), .window_19__7 (
               currentPage_5__7), .window_19__6 (currentPage_5__6), .window_19__5 (
               currentPage_5__5), .window_19__4 (currentPage_5__4), .window_19__3 (
               currentPage_5__3), .window_19__2 (currentPage_5__2), .window_19__1 (
               currentPage_5__1), .window_19__0 (currentPage_5__0), .window_18__15 (
               currentPage_6__15), .window_18__14 (currentPage_6__14), .window_18__13 (
               currentPage_6__13), .window_18__12 (currentPage_6__12), .window_18__11 (
               currentPage_6__11), .window_18__10 (currentPage_6__10), .window_18__9 (
               currentPage_6__9), .window_18__8 (currentPage_6__8), .window_18__7 (
               currentPage_6__7), .window_18__6 (currentPage_6__6), .window_18__5 (
               currentPage_6__5), .window_18__4 (currentPage_6__4), .window_18__3 (
               currentPage_6__3), .window_18__2 (currentPage_6__2), .window_18__1 (
               currentPage_6__1), .window_18__0 (currentPage_6__0), .window_17__15 (
               currentPage_7__15), .window_17__14 (currentPage_7__14), .window_17__13 (
               currentPage_7__13), .window_17__12 (currentPage_7__12), .window_17__11 (
               currentPage_7__11), .window_17__10 (currentPage_7__10), .window_17__9 (
               currentPage_7__9), .window_17__8 (currentPage_7__8), .window_17__7 (
               currentPage_7__7), .window_17__6 (currentPage_7__6), .window_17__5 (
               currentPage_7__5), .window_17__4 (currentPage_7__4), .window_17__3 (
               currentPage_7__3), .window_17__2 (currentPage_7__2), .window_17__1 (
               currentPage_7__1), .window_17__0 (currentPage_7__0), .window_16__15 (
               currentPage_8__15), .window_16__14 (currentPage_8__14), .window_16__13 (
               currentPage_8__13), .window_16__12 (currentPage_8__12), .window_16__11 (
               currentPage_8__11), .window_16__10 (currentPage_8__10), .window_16__9 (
               currentPage_8__9), .window_16__8 (currentPage_8__8), .window_16__7 (
               currentPage_8__7), .window_16__6 (currentPage_8__6), .window_16__5 (
               currentPage_8__5), .window_16__4 (currentPage_8__4), .window_16__3 (
               currentPage_8__3), .window_16__2 (currentPage_8__2), .window_16__1 (
               currentPage_8__1), .window_16__0 (currentPage_8__0), .window_15__15 (
               currentPage_9__15), .window_15__14 (currentPage_9__14), .window_15__13 (
               currentPage_9__13), .window_15__12 (currentPage_9__12), .window_15__11 (
               currentPage_9__11), .window_15__10 (currentPage_9__10), .window_15__9 (
               currentPage_9__9), .window_15__8 (currentPage_9__8), .window_15__7 (
               currentPage_9__7), .window_15__6 (currentPage_9__6), .window_15__5 (
               currentPage_9__5), .window_15__4 (currentPage_9__4), .window_15__3 (
               currentPage_9__3), .window_15__2 (currentPage_9__2), .window_15__1 (
               currentPage_9__1), .window_15__0 (currentPage_9__0), .window_14__15 (
               currentPage_10__15), .window_14__14 (currentPage_10__14), .window_14__13 (
               currentPage_10__13), .window_14__12 (currentPage_10__12), .window_14__11 (
               currentPage_10__11), .window_14__10 (currentPage_10__10), .window_14__9 (
               currentPage_10__9), .window_14__8 (currentPage_10__8), .window_14__7 (
               currentPage_10__7), .window_14__6 (currentPage_10__6), .window_14__5 (
               currentPage_10__5), .window_14__4 (currentPage_10__4), .window_14__3 (
               currentPage_10__3), .window_14__2 (currentPage_10__2), .window_14__1 (
               currentPage_10__1), .window_14__0 (currentPage_10__0), .window_13__15 (
               currentPage_11__15), .window_13__14 (currentPage_11__14), .window_13__13 (
               currentPage_11__13), .window_13__12 (currentPage_11__12), .window_13__11 (
               currentPage_11__11), .window_13__10 (currentPage_11__10), .window_13__9 (
               currentPage_11__9), .window_13__8 (currentPage_11__8), .window_13__7 (
               currentPage_11__7), .window_13__6 (currentPage_11__6), .window_13__5 (
               currentPage_11__5), .window_13__4 (currentPage_11__4), .window_13__3 (
               currentPage_11__3), .window_13__2 (currentPage_11__2), .window_13__1 (
               currentPage_11__1), .window_13__0 (currentPage_11__0), .window_12__15 (
               currentPage_12__15), .window_12__14 (currentPage_12__14), .window_12__13 (
               currentPage_12__13), .window_12__12 (currentPage_12__12), .window_12__11 (
               currentPage_12__11), .window_12__10 (currentPage_12__10), .window_12__9 (
               currentPage_12__9), .window_12__8 (currentPage_12__8), .window_12__7 (
               currentPage_12__7), .window_12__6 (currentPage_12__6), .window_12__5 (
               currentPage_12__5), .window_12__4 (currentPage_12__4), .window_12__3 (
               currentPage_12__3), .window_12__2 (currentPage_12__2), .window_12__1 (
               currentPage_12__1), .window_12__0 (currentPage_12__0), .window_11__15 (
               currentPage_13__15), .window_11__14 (currentPage_13__14), .window_11__13 (
               currentPage_13__13), .window_11__12 (currentPage_13__12), .window_11__11 (
               currentPage_13__11), .window_11__10 (currentPage_13__10), .window_11__9 (
               currentPage_13__9), .window_11__8 (currentPage_13__8), .window_11__7 (
               currentPage_13__7), .window_11__6 (currentPage_13__6), .window_11__5 (
               currentPage_13__5), .window_11__4 (currentPage_13__4), .window_11__3 (
               currentPage_13__3), .window_11__2 (currentPage_13__2), .window_11__1 (
               currentPage_13__1), .window_11__0 (currentPage_13__0), .window_10__15 (
               currentPage_14__15), .window_10__14 (currentPage_14__14), .window_10__13 (
               currentPage_14__13), .window_10__12 (currentPage_14__12), .window_10__11 (
               currentPage_14__11), .window_10__10 (currentPage_14__10), .window_10__9 (
               currentPage_14__9), .window_10__8 (currentPage_14__8), .window_10__7 (
               currentPage_14__7), .window_10__6 (currentPage_14__6), .window_10__5 (
               currentPage_14__5), .window_10__4 (currentPage_14__4), .window_10__3 (
               currentPage_14__3), .window_10__2 (currentPage_14__2), .window_10__1 (
               currentPage_14__1), .window_10__0 (currentPage_14__0), .window_9__15 (
               currentPage_15__15), .window_9__14 (currentPage_15__14), .window_9__13 (
               currentPage_15__13), .window_9__12 (currentPage_15__12), .window_9__11 (
               currentPage_15__11), .window_9__10 (currentPage_15__10), .window_9__9 (
               currentPage_15__9), .window_9__8 (currentPage_15__8), .window_9__7 (
               currentPage_15__7), .window_9__6 (currentPage_15__6), .window_9__5 (
               currentPage_15__5), .window_9__4 (currentPage_15__4), .window_9__3 (
               currentPage_15__3), .window_9__2 (currentPage_15__2), .window_9__1 (
               currentPage_15__1), .window_9__0 (currentPage_15__0), .window_8__15 (
               currentPage_16__15), .window_8__14 (currentPage_16__14), .window_8__13 (
               currentPage_16__13), .window_8__12 (currentPage_16__12), .window_8__11 (
               currentPage_16__11), .window_8__10 (currentPage_16__10), .window_8__9 (
               currentPage_16__9), .window_8__8 (currentPage_16__8), .window_8__7 (
               currentPage_16__7), .window_8__6 (currentPage_16__6), .window_8__5 (
               currentPage_16__5), .window_8__4 (currentPage_16__4), .window_8__3 (
               currentPage_16__3), .window_8__2 (currentPage_16__2), .window_8__1 (
               currentPage_16__1), .window_8__0 (currentPage_16__0), .window_7__15 (
               currentPage_17__15), .window_7__14 (currentPage_17__14), .window_7__13 (
               currentPage_17__13), .window_7__12 (currentPage_17__12), .window_7__11 (
               currentPage_17__11), .window_7__10 (currentPage_17__10), .window_7__9 (
               currentPage_17__9), .window_7__8 (currentPage_17__8), .window_7__7 (
               currentPage_17__7), .window_7__6 (currentPage_17__6), .window_7__5 (
               currentPage_17__5), .window_7__4 (currentPage_17__4), .window_7__3 (
               currentPage_17__3), .window_7__2 (currentPage_17__2), .window_7__1 (
               currentPage_17__1), .window_7__0 (currentPage_17__0), .window_6__15 (
               currentPage_18__15), .window_6__14 (currentPage_18__14), .window_6__13 (
               currentPage_18__13), .window_6__12 (currentPage_18__12), .window_6__11 (
               currentPage_18__11), .window_6__10 (currentPage_18__10), .window_6__9 (
               currentPage_18__9), .window_6__8 (currentPage_18__8), .window_6__7 (
               currentPage_18__7), .window_6__6 (currentPage_18__6), .window_6__5 (
               currentPage_18__5), .window_6__4 (currentPage_18__4), .window_6__3 (
               currentPage_18__3), .window_6__2 (currentPage_18__2), .window_6__1 (
               currentPage_18__1), .window_6__0 (currentPage_18__0), .window_5__15 (
               currentPage_19__15), .window_5__14 (currentPage_19__14), .window_5__13 (
               currentPage_19__13), .window_5__12 (currentPage_19__12), .window_5__11 (
               currentPage_19__11), .window_5__10 (currentPage_19__10), .window_5__9 (
               currentPage_19__9), .window_5__8 (currentPage_19__8), .window_5__7 (
               currentPage_19__7), .window_5__6 (currentPage_19__6), .window_5__5 (
               currentPage_19__5), .window_5__4 (currentPage_19__4), .window_5__3 (
               currentPage_19__3), .window_5__2 (currentPage_19__2), .window_5__1 (
               currentPage_19__1), .window_5__0 (currentPage_19__0), .window_4__15 (
               currentPage_20__15), .window_4__14 (currentPage_20__14), .window_4__13 (
               currentPage_20__13), .window_4__12 (currentPage_20__12), .window_4__11 (
               currentPage_20__11), .window_4__10 (currentPage_20__10), .window_4__9 (
               currentPage_20__9), .window_4__8 (currentPage_20__8), .window_4__7 (
               currentPage_20__7), .window_4__6 (currentPage_20__6), .window_4__5 (
               currentPage_20__5), .window_4__4 (currentPage_20__4), .window_4__3 (
               currentPage_20__3), .window_4__2 (currentPage_20__2), .window_4__1 (
               currentPage_20__1), .window_4__0 (currentPage_20__0), .window_3__15 (
               currentPage_21__15), .window_3__14 (currentPage_21__14), .window_3__13 (
               currentPage_21__13), .window_3__12 (currentPage_21__12), .window_3__11 (
               currentPage_21__11), .window_3__10 (currentPage_21__10), .window_3__9 (
               currentPage_21__9), .window_3__8 (currentPage_21__8), .window_3__7 (
               currentPage_21__7), .window_3__6 (currentPage_21__6), .window_3__5 (
               currentPage_21__5), .window_3__4 (currentPage_21__4), .window_3__3 (
               currentPage_21__3), .window_3__2 (currentPage_21__2), .window_3__1 (
               currentPage_21__1), .window_3__0 (currentPage_21__0), .window_2__15 (
               currentPage_22__15), .window_2__14 (currentPage_22__14), .window_2__13 (
               currentPage_22__13), .window_2__12 (currentPage_22__12), .window_2__11 (
               currentPage_22__11), .window_2__10 (currentPage_22__10), .window_2__9 (
               currentPage_22__9), .window_2__8 (currentPage_22__8), .window_2__7 (
               currentPage_22__7), .window_2__6 (currentPage_22__6), .window_2__5 (
               currentPage_22__5), .window_2__4 (currentPage_22__4), .window_2__3 (
               currentPage_22__3), .window_2__2 (currentPage_22__2), .window_2__1 (
               currentPage_22__1), .window_2__0 (currentPage_22__0), .window_1__15 (
               currentPage_23__15), .window_1__14 (currentPage_23__14), .window_1__13 (
               currentPage_23__13), .window_1__12 (currentPage_23__12), .window_1__11 (
               currentPage_23__11), .window_1__10 (currentPage_23__10), .window_1__9 (
               currentPage_23__9), .window_1__8 (currentPage_23__8), .window_1__7 (
               currentPage_23__7), .window_1__6 (currentPage_23__6), .window_1__5 (
               currentPage_23__5), .window_1__4 (currentPage_23__4), .window_1__3 (
               currentPage_23__3), .window_1__2 (currentPage_23__2), .window_1__1 (
               currentPage_23__1), .window_1__0 (currentPage_23__0), .window_0__15 (
               currentPage_24__15), .window_0__14 (currentPage_24__14), .window_0__13 (
               currentPage_24__13), .window_0__12 (currentPage_24__12), .window_0__11 (
               currentPage_24__11), .window_0__10 (currentPage_24__10), .window_0__9 (
               currentPage_24__9), .window_0__8 (currentPage_24__8), .window_0__7 (
               currentPage_24__7), .window_0__6 (currentPage_24__6), .window_0__5 (
               currentPage_24__5), .window_0__4 (currentPage_24__4), .window_0__3 (
               currentPage_24__3), .window_0__2 (currentPage_24__2), .window_0__1 (
               currentPage_24__1), .window_0__0 (currentPage_24__0), .outputs_24__15 (
               outMuls_0__15), .outputs_24__14 (outMuls_0__14), .outputs_24__13 (
               outMuls_0__13), .outputs_24__12 (outMuls_0__12), .outputs_24__11 (
               outMuls_0__11), .outputs_24__10 (outMuls_0__10), .outputs_24__9 (
               outMuls_0__9), .outputs_24__8 (outMuls_0__8), .outputs_24__7 (
               outMuls_0__7), .outputs_24__6 (outMuls_0__6), .outputs_24__5 (
               outMuls_0__5), .outputs_24__4 (outMuls_0__4), .outputs_24__3 (
               outMuls_0__3), .outputs_24__2 (outMuls_0__2), .outputs_24__1 (
               outMuls_0__1), .outputs_24__0 (outMuls_0__0), .outputs_23__15 (
               outMuls_1__15), .outputs_23__14 (outMuls_1__14), .outputs_23__13 (
               outMuls_1__13), .outputs_23__12 (outMuls_1__12), .outputs_23__11 (
               outMuls_1__11), .outputs_23__10 (outMuls_1__10), .outputs_23__9 (
               outMuls_1__9), .outputs_23__8 (outMuls_1__8), .outputs_23__7 (
               outMuls_1__7), .outputs_23__6 (outMuls_1__6), .outputs_23__5 (
               outMuls_1__5), .outputs_23__4 (outMuls_1__4), .outputs_23__3 (
               outMuls_1__3), .outputs_23__2 (outMuls_1__2), .outputs_23__1 (
               outMuls_1__1), .outputs_23__0 (outMuls_1__0), .outputs_22__15 (
               outMuls_2__15), .outputs_22__14 (outMuls_2__14), .outputs_22__13 (
               outMuls_2__13), .outputs_22__12 (outMuls_2__12), .outputs_22__11 (
               outMuls_2__11), .outputs_22__10 (outMuls_2__10), .outputs_22__9 (
               outMuls_2__9), .outputs_22__8 (outMuls_2__8), .outputs_22__7 (
               outMuls_2__7), .outputs_22__6 (outMuls_2__6), .outputs_22__5 (
               outMuls_2__5), .outputs_22__4 (outMuls_2__4), .outputs_22__3 (
               outMuls_2__3), .outputs_22__2 (outMuls_2__2), .outputs_22__1 (
               outMuls_2__1), .outputs_22__0 (outMuls_2__0), .outputs_21__15 (
               outMuls_3__15), .outputs_21__14 (outMuls_3__14), .outputs_21__13 (
               outMuls_3__13), .outputs_21__12 (outMuls_3__12), .outputs_21__11 (
               outMuls_3__11), .outputs_21__10 (outMuls_3__10), .outputs_21__9 (
               outMuls_3__9), .outputs_21__8 (outMuls_3__8), .outputs_21__7 (
               outMuls_3__7), .outputs_21__6 (outMuls_3__6), .outputs_21__5 (
               outMuls_3__5), .outputs_21__4 (outMuls_3__4), .outputs_21__3 (
               outMuls_3__3), .outputs_21__2 (outMuls_3__2), .outputs_21__1 (
               outMuls_3__1), .outputs_21__0 (outMuls_3__0), .outputs_20__15 (
               outMuls_4__15), .outputs_20__14 (outMuls_4__14), .outputs_20__13 (
               outMuls_4__13), .outputs_20__12 (outMuls_4__12), .outputs_20__11 (
               outMuls_4__11), .outputs_20__10 (outMuls_4__10), .outputs_20__9 (
               outMuls_4__9), .outputs_20__8 (outMuls_4__8), .outputs_20__7 (
               outMuls_4__7), .outputs_20__6 (outMuls_4__6), .outputs_20__5 (
               outMuls_4__5), .outputs_20__4 (outMuls_4__4), .outputs_20__3 (
               outMuls_4__3), .outputs_20__2 (outMuls_4__2), .outputs_20__1 (
               outMuls_4__1), .outputs_20__0 (outMuls_4__0), .outputs_19__15 (
               outMuls_5__15), .outputs_19__14 (outMuls_5__14), .outputs_19__13 (
               outMuls_5__13), .outputs_19__12 (outMuls_5__12), .outputs_19__11 (
               outMuls_5__11), .outputs_19__10 (outMuls_5__10), .outputs_19__9 (
               outMuls_5__9), .outputs_19__8 (outMuls_5__8), .outputs_19__7 (
               outMuls_5__7), .outputs_19__6 (outMuls_5__6), .outputs_19__5 (
               outMuls_5__5), .outputs_19__4 (outMuls_5__4), .outputs_19__3 (
               outMuls_5__3), .outputs_19__2 (outMuls_5__2), .outputs_19__1 (
               outMuls_5__1), .outputs_19__0 (outMuls_5__0), .outputs_18__15 (
               outMuls_6__15), .outputs_18__14 (outMuls_6__14), .outputs_18__13 (
               outMuls_6__13), .outputs_18__12 (outMuls_6__12), .outputs_18__11 (
               outMuls_6__11), .outputs_18__10 (outMuls_6__10), .outputs_18__9 (
               outMuls_6__9), .outputs_18__8 (outMuls_6__8), .outputs_18__7 (
               outMuls_6__7), .outputs_18__6 (outMuls_6__6), .outputs_18__5 (
               outMuls_6__5), .outputs_18__4 (outMuls_6__4), .outputs_18__3 (
               outMuls_6__3), .outputs_18__2 (outMuls_6__2), .outputs_18__1 (
               outMuls_6__1), .outputs_18__0 (outMuls_6__0), .outputs_17__15 (
               outMuls_7__15), .outputs_17__14 (outMuls_7__14), .outputs_17__13 (
               outMuls_7__13), .outputs_17__12 (outMuls_7__12), .outputs_17__11 (
               outMuls_7__11), .outputs_17__10 (outMuls_7__10), .outputs_17__9 (
               outMuls_7__9), .outputs_17__8 (outMuls_7__8), .outputs_17__7 (
               outMuls_7__7), .outputs_17__6 (outMuls_7__6), .outputs_17__5 (
               outMuls_7__5), .outputs_17__4 (outMuls_7__4), .outputs_17__3 (
               outMuls_7__3), .outputs_17__2 (outMuls_7__2), .outputs_17__1 (
               outMuls_7__1), .outputs_17__0 (outMuls_7__0), .outputs_16__15 (
               outMuls_8__15), .outputs_16__14 (outMuls_8__14), .outputs_16__13 (
               outMuls_8__13), .outputs_16__12 (outMuls_8__12), .outputs_16__11 (
               outMuls_8__11), .outputs_16__10 (outMuls_8__10), .outputs_16__9 (
               outMuls_8__9), .outputs_16__8 (outMuls_8__8), .outputs_16__7 (
               outMuls_8__7), .outputs_16__6 (outMuls_8__6), .outputs_16__5 (
               outMuls_8__5), .outputs_16__4 (outMuls_8__4), .outputs_16__3 (
               outMuls_8__3), .outputs_16__2 (outMuls_8__2), .outputs_16__1 (
               outMuls_8__1), .outputs_16__0 (outMuls_8__0), .outputs_15__15 (
               outMuls_9__15), .outputs_15__14 (outMuls_9__14), .outputs_15__13 (
               outMuls_9__13), .outputs_15__12 (outMuls_9__12), .outputs_15__11 (
               outMuls_9__11), .outputs_15__10 (outMuls_9__10), .outputs_15__9 (
               outMuls_9__9), .outputs_15__8 (outMuls_9__8), .outputs_15__7 (
               outMuls_9__7), .outputs_15__6 (outMuls_9__6), .outputs_15__5 (
               outMuls_9__5), .outputs_15__4 (outMuls_9__4), .outputs_15__3 (
               outMuls_9__3), .outputs_15__2 (outMuls_9__2), .outputs_15__1 (
               outMuls_9__1), .outputs_15__0 (outMuls_9__0), .outputs_14__15 (
               outMuls_10__15), .outputs_14__14 (outMuls_10__14), .outputs_14__13 (
               outMuls_10__13), .outputs_14__12 (outMuls_10__12), .outputs_14__11 (
               outMuls_10__11), .outputs_14__10 (outMuls_10__10), .outputs_14__9 (
               outMuls_10__9), .outputs_14__8 (outMuls_10__8), .outputs_14__7 (
               outMuls_10__7), .outputs_14__6 (outMuls_10__6), .outputs_14__5 (
               outMuls_10__5), .outputs_14__4 (outMuls_10__4), .outputs_14__3 (
               outMuls_10__3), .outputs_14__2 (outMuls_10__2), .outputs_14__1 (
               outMuls_10__1), .outputs_14__0 (outMuls_10__0), .outputs_13__15 (
               outMuls_11__15), .outputs_13__14 (outMuls_11__14), .outputs_13__13 (
               outMuls_11__13), .outputs_13__12 (outMuls_11__12), .outputs_13__11 (
               outMuls_11__11), .outputs_13__10 (outMuls_11__10), .outputs_13__9 (
               outMuls_11__9), .outputs_13__8 (outMuls_11__8), .outputs_13__7 (
               outMuls_11__7), .outputs_13__6 (outMuls_11__6), .outputs_13__5 (
               outMuls_11__5), .outputs_13__4 (outMuls_11__4), .outputs_13__3 (
               outMuls_11__3), .outputs_13__2 (outMuls_11__2), .outputs_13__1 (
               outMuls_11__1), .outputs_13__0 (outMuls_11__0), .outputs_12__15 (
               outMuls_12__15), .outputs_12__14 (outMuls_12__14), .outputs_12__13 (
               outMuls_12__13), .outputs_12__12 (outMuls_12__12), .outputs_12__11 (
               outMuls_12__11), .outputs_12__10 (outMuls_12__10), .outputs_12__9 (
               outMuls_12__9), .outputs_12__8 (outMuls_12__8), .outputs_12__7 (
               outMuls_12__7), .outputs_12__6 (outMuls_12__6), .outputs_12__5 (
               outMuls_12__5), .outputs_12__4 (outMuls_12__4), .outputs_12__3 (
               outMuls_12__3), .outputs_12__2 (outMuls_12__2), .outputs_12__1 (
               outMuls_12__1), .outputs_12__0 (outMuls_12__0), .outputs_11__15 (
               outMuls_13__15), .outputs_11__14 (outMuls_13__14), .outputs_11__13 (
               outMuls_13__13), .outputs_11__12 (outMuls_13__12), .outputs_11__11 (
               outMuls_13__11), .outputs_11__10 (outMuls_13__10), .outputs_11__9 (
               outMuls_13__9), .outputs_11__8 (outMuls_13__8), .outputs_11__7 (
               outMuls_13__7), .outputs_11__6 (outMuls_13__6), .outputs_11__5 (
               outMuls_13__5), .outputs_11__4 (outMuls_13__4), .outputs_11__3 (
               outMuls_13__3), .outputs_11__2 (outMuls_13__2), .outputs_11__1 (
               outMuls_13__1), .outputs_11__0 (outMuls_13__0), .outputs_10__15 (
               outMuls_14__15), .outputs_10__14 (outMuls_14__14), .outputs_10__13 (
               outMuls_14__13), .outputs_10__12 (outMuls_14__12), .outputs_10__11 (
               outMuls_14__11), .outputs_10__10 (outMuls_14__10), .outputs_10__9 (
               outMuls_14__9), .outputs_10__8 (outMuls_14__8), .outputs_10__7 (
               outMuls_14__7), .outputs_10__6 (outMuls_14__6), .outputs_10__5 (
               outMuls_14__5), .outputs_10__4 (outMuls_14__4), .outputs_10__3 (
               outMuls_14__3), .outputs_10__2 (outMuls_14__2), .outputs_10__1 (
               outMuls_14__1), .outputs_10__0 (outMuls_14__0), .outputs_9__15 (
               outMuls_15__15), .outputs_9__14 (outMuls_15__14), .outputs_9__13 (
               outMuls_15__13), .outputs_9__12 (outMuls_15__12), .outputs_9__11 (
               outMuls_15__11), .outputs_9__10 (outMuls_15__10), .outputs_9__9 (
               outMuls_15__9), .outputs_9__8 (outMuls_15__8), .outputs_9__7 (
               outMuls_15__7), .outputs_9__6 (outMuls_15__6), .outputs_9__5 (
               outMuls_15__5), .outputs_9__4 (outMuls_15__4), .outputs_9__3 (
               outMuls_15__3), .outputs_9__2 (outMuls_15__2), .outputs_9__1 (
               outMuls_15__1), .outputs_9__0 (outMuls_15__0), .outputs_8__15 (
               outMuls_16__15), .outputs_8__14 (outMuls_16__14), .outputs_8__13 (
               outMuls_16__13), .outputs_8__12 (outMuls_16__12), .outputs_8__11 (
               outMuls_16__11), .outputs_8__10 (outMuls_16__10), .outputs_8__9 (
               outMuls_16__9), .outputs_8__8 (outMuls_16__8), .outputs_8__7 (
               outMuls_16__7), .outputs_8__6 (outMuls_16__6), .outputs_8__5 (
               outMuls_16__5), .outputs_8__4 (outMuls_16__4), .outputs_8__3 (
               outMuls_16__3), .outputs_8__2 (outMuls_16__2), .outputs_8__1 (
               outMuls_16__1), .outputs_8__0 (outMuls_16__0), .outputs_7__15 (
               outMuls_17__15), .outputs_7__14 (outMuls_17__14), .outputs_7__13 (
               outMuls_17__13), .outputs_7__12 (outMuls_17__12), .outputs_7__11 (
               outMuls_17__11), .outputs_7__10 (outMuls_17__10), .outputs_7__9 (
               outMuls_17__9), .outputs_7__8 (outMuls_17__8), .outputs_7__7 (
               outMuls_17__7), .outputs_7__6 (outMuls_17__6), .outputs_7__5 (
               outMuls_17__5), .outputs_7__4 (outMuls_17__4), .outputs_7__3 (
               outMuls_17__3), .outputs_7__2 (outMuls_17__2), .outputs_7__1 (
               outMuls_17__1), .outputs_7__0 (outMuls_17__0), .outputs_6__15 (
               outMuls_18__15), .outputs_6__14 (outMuls_18__14), .outputs_6__13 (
               outMuls_18__13), .outputs_6__12 (outMuls_18__12), .outputs_6__11 (
               outMuls_18__11), .outputs_6__10 (outMuls_18__10), .outputs_6__9 (
               outMuls_18__9), .outputs_6__8 (outMuls_18__8), .outputs_6__7 (
               outMuls_18__7), .outputs_6__6 (outMuls_18__6), .outputs_6__5 (
               outMuls_18__5), .outputs_6__4 (outMuls_18__4), .outputs_6__3 (
               outMuls_18__3), .outputs_6__2 (outMuls_18__2), .outputs_6__1 (
               outMuls_18__1), .outputs_6__0 (outMuls_18__0), .outputs_5__15 (
               outMuls_19__15), .outputs_5__14 (outMuls_19__14), .outputs_5__13 (
               outMuls_19__13), .outputs_5__12 (outMuls_19__12), .outputs_5__11 (
               outMuls_19__11), .outputs_5__10 (outMuls_19__10), .outputs_5__9 (
               outMuls_19__9), .outputs_5__8 (outMuls_19__8), .outputs_5__7 (
               outMuls_19__7), .outputs_5__6 (outMuls_19__6), .outputs_5__5 (
               outMuls_19__5), .outputs_5__4 (outMuls_19__4), .outputs_5__3 (
               outMuls_19__3), .outputs_5__2 (outMuls_19__2), .outputs_5__1 (
               outMuls_19__1), .outputs_5__0 (outMuls_19__0), .outputs_4__15 (
               outMuls_20__15), .outputs_4__14 (outMuls_20__14), .outputs_4__13 (
               outMuls_20__13), .outputs_4__12 (outMuls_20__12), .outputs_4__11 (
               outMuls_20__11), .outputs_4__10 (outMuls_20__10), .outputs_4__9 (
               outMuls_20__9), .outputs_4__8 (outMuls_20__8), .outputs_4__7 (
               outMuls_20__7), .outputs_4__6 (outMuls_20__6), .outputs_4__5 (
               outMuls_20__5), .outputs_4__4 (outMuls_20__4), .outputs_4__3 (
               outMuls_20__3), .outputs_4__2 (outMuls_20__2), .outputs_4__1 (
               outMuls_20__1), .outputs_4__0 (outMuls_20__0), .outputs_3__15 (
               outMuls_21__15), .outputs_3__14 (outMuls_21__14), .outputs_3__13 (
               outMuls_21__13), .outputs_3__12 (outMuls_21__12), .outputs_3__11 (
               outMuls_21__11), .outputs_3__10 (outMuls_21__10), .outputs_3__9 (
               outMuls_21__9), .outputs_3__8 (outMuls_21__8), .outputs_3__7 (
               outMuls_21__7), .outputs_3__6 (outMuls_21__6), .outputs_3__5 (
               outMuls_21__5), .outputs_3__4 (outMuls_21__4), .outputs_3__3 (
               outMuls_21__3), .outputs_3__2 (outMuls_21__2), .outputs_3__1 (
               outMuls_21__1), .outputs_3__0 (outMuls_21__0), .outputs_2__15 (
               outMuls_22__15), .outputs_2__14 (outMuls_22__14), .outputs_2__13 (
               outMuls_22__13), .outputs_2__12 (outMuls_22__12), .outputs_2__11 (
               outMuls_22__11), .outputs_2__10 (outMuls_22__10), .outputs_2__9 (
               outMuls_22__9), .outputs_2__8 (outMuls_22__8), .outputs_2__7 (
               outMuls_22__7), .outputs_2__6 (outMuls_22__6), .outputs_2__5 (
               outMuls_22__5), .outputs_2__4 (outMuls_22__4), .outputs_2__3 (
               outMuls_22__3), .outputs_2__2 (outMuls_22__2), .outputs_2__1 (
               outMuls_22__1), .outputs_2__0 (outMuls_22__0), .outputs_1__15 (
               outMuls_23__15), .outputs_1__14 (outMuls_23__14), .outputs_1__13 (
               outMuls_23__13), .outputs_1__12 (outMuls_23__12), .outputs_1__11 (
               outMuls_23__11), .outputs_1__10 (outMuls_23__10), .outputs_1__9 (
               outMuls_23__9), .outputs_1__8 (outMuls_23__8), .outputs_1__7 (
               outMuls_23__7), .outputs_1__6 (outMuls_23__6), .outputs_1__5 (
               outMuls_23__5), .outputs_1__4 (outMuls_23__4), .outputs_1__3 (
               outMuls_23__3), .outputs_1__2 (outMuls_23__2), .outputs_1__1 (
               outMuls_23__1), .outputs_1__0 (outMuls_23__0), .outputs_0__15 (
               outMuls_24__15), .outputs_0__14 (outMuls_24__14), .outputs_0__13 (
               outMuls_24__13), .outputs_0__12 (outMuls_24__12), .outputs_0__11 (
               outMuls_24__11), .outputs_0__10 (outMuls_24__10), .outputs_0__9 (
               outMuls_24__9), .outputs_0__8 (outMuls_24__8), .outputs_0__7 (
               outMuls_24__7), .outputs_0__6 (outMuls_24__6), .outputs_0__5 (
               outMuls_24__5), .outputs_0__4 (outMuls_24__4), .outputs_0__3 (
               outMuls_24__3), .outputs_0__2 (outMuls_24__2), .outputs_0__1 (
               outMuls_24__1), .outputs_0__0 (outMuls_24__0), .clk (clk), .start (
               start), .rst (rst), .doneOut (doneMul), .workingOut (\$dummy [0])
               ) ;
    Mux2_16 loop1_0_inputAddersMap (.A ({outMuls_0__15,outMuls_0__14,
            outMuls_0__13,outMuls_0__12,outMuls_0__11,outMuls_0__10,outMuls_0__9
            ,outMuls_0__8,outMuls_0__7,outMuls_0__6,outMuls_0__5,outMuls_0__4,
            outMuls_0__3,outMuls_0__2,outMuls_0__1,outMuls_0__0}), .B ({
            currentPage_0__15,currentPage_0__14,currentPage_0__13,
            currentPage_0__12,currentPage_0__11,currentPage_0__10,
            currentPage_0__9,currentPage_0__8,currentPage_0__7,currentPage_0__6,
            currentPage_0__5,currentPage_0__4,currentPage_0__3,currentPage_0__2,
            currentPage_0__1,currentPage_0__0}), .S (nx1946), .C ({
            addersInputs_0__15,addersInputs_0__14,addersInputs_0__13,
            addersInputs_0__12,addersInputs_0__11,addersInputs_0__10,
            addersInputs_0__9,addersInputs_0__8,addersInputs_0__7,
            addersInputs_0__6,addersInputs_0__5,addersInputs_0__4,
            addersInputs_0__3,addersInputs_0__2,addersInputs_0__1,
            addersInputs_0__0})) ;
    Mux2_16 loop1_1_inputAddersMap (.A ({outMuls_1__15,outMuls_1__14,
            outMuls_1__13,outMuls_1__12,outMuls_1__11,outMuls_1__10,outMuls_1__9
            ,outMuls_1__8,outMuls_1__7,outMuls_1__6,outMuls_1__5,outMuls_1__4,
            outMuls_1__3,outMuls_1__2,outMuls_1__1,outMuls_1__0}), .B ({
            currentPage_1__15,currentPage_1__14,currentPage_1__13,
            currentPage_1__12,currentPage_1__11,currentPage_1__10,
            currentPage_1__9,currentPage_1__8,currentPage_1__7,currentPage_1__6,
            currentPage_1__5,currentPage_1__4,currentPage_1__3,currentPage_1__2,
            currentPage_1__1,currentPage_1__0}), .S (nx1946), .C ({
            addersInputs_1__15,addersInputs_1__14,addersInputs_1__13,
            addersInputs_1__12,addersInputs_1__11,addersInputs_1__10,
            addersInputs_1__9,addersInputs_1__8,addersInputs_1__7,
            addersInputs_1__6,addersInputs_1__5,addersInputs_1__4,
            addersInputs_1__3,addersInputs_1__2,addersInputs_1__1,
            addersInputs_1__0})) ;
    Mux2_16 loop1_2_inputAddersMap (.A ({outMuls_2__15,outMuls_2__14,
            outMuls_2__13,outMuls_2__12,outMuls_2__11,outMuls_2__10,outMuls_2__9
            ,outMuls_2__8,outMuls_2__7,outMuls_2__6,outMuls_2__5,outMuls_2__4,
            outMuls_2__3,outMuls_2__2,outMuls_2__1,outMuls_2__0}), .B ({
            currentPage_2__15,currentPage_2__14,currentPage_2__13,
            currentPage_2__12,currentPage_2__11,currentPage_2__10,
            currentPage_2__9,currentPage_2__8,currentPage_2__7,currentPage_2__6,
            currentPage_2__5,currentPage_2__4,currentPage_2__3,currentPage_2__2,
            currentPage_2__1,currentPage_2__0}), .S (nx1946), .C ({
            addersInputs_2__15,addersInputs_2__14,addersInputs_2__13,
            addersInputs_2__12,addersInputs_2__11,addersInputs_2__10,
            addersInputs_2__9,addersInputs_2__8,addersInputs_2__7,
            addersInputs_2__6,addersInputs_2__5,addersInputs_2__4,
            addersInputs_2__3,addersInputs_2__2,addersInputs_2__1,
            addersInputs_2__0})) ;
    Mux2_16 loop1_3_inputAddersMap (.A ({outMuls_3__15,outMuls_3__14,
            outMuls_3__13,outMuls_3__12,outMuls_3__11,outMuls_3__10,outMuls_3__9
            ,outMuls_3__8,outMuls_3__7,outMuls_3__6,outMuls_3__5,outMuls_3__4,
            outMuls_3__3,outMuls_3__2,outMuls_3__1,outMuls_3__0}), .B ({
            currentPage_3__15,currentPage_3__14,currentPage_3__13,
            currentPage_3__12,currentPage_3__11,currentPage_3__10,
            currentPage_3__9,currentPage_3__8,currentPage_3__7,currentPage_3__6,
            currentPage_3__5,currentPage_3__4,currentPage_3__3,currentPage_3__2,
            currentPage_3__1,currentPage_3__0}), .S (nx1946), .C ({
            addersInputs_3__15,addersInputs_3__14,addersInputs_3__13,
            addersInputs_3__12,addersInputs_3__11,addersInputs_3__10,
            addersInputs_3__9,addersInputs_3__8,addersInputs_3__7,
            addersInputs_3__6,addersInputs_3__5,addersInputs_3__4,
            addersInputs_3__3,addersInputs_3__2,addersInputs_3__1,
            addersInputs_3__0})) ;
    Mux2_16 loop1_4_inputAddersMap (.A ({outMuls_4__15,outMuls_4__14,
            outMuls_4__13,outMuls_4__12,outMuls_4__11,outMuls_4__10,outMuls_4__9
            ,outMuls_4__8,outMuls_4__7,outMuls_4__6,outMuls_4__5,outMuls_4__4,
            outMuls_4__3,outMuls_4__2,outMuls_4__1,outMuls_4__0}), .B ({
            currentPage_4__15,currentPage_4__14,currentPage_4__13,
            currentPage_4__12,currentPage_4__11,currentPage_4__10,
            currentPage_4__9,currentPage_4__8,currentPage_4__7,currentPage_4__6,
            currentPage_4__5,currentPage_4__4,currentPage_4__3,currentPage_4__2,
            currentPage_4__1,currentPage_4__0}), .S (nx1946), .C ({
            addersInputs_4__15,addersInputs_4__14,addersInputs_4__13,
            addersInputs_4__12,addersInputs_4__11,addersInputs_4__10,
            addersInputs_4__9,addersInputs_4__8,addersInputs_4__7,
            addersInputs_4__6,addersInputs_4__5,addersInputs_4__4,
            addersInputs_4__3,addersInputs_4__2,addersInputs_4__1,
            addersInputs_4__0})) ;
    Mux2_16 loop1_5_inputAddersMap (.A ({outMuls_5__15,outMuls_5__14,
            outMuls_5__13,outMuls_5__12,outMuls_5__11,outMuls_5__10,outMuls_5__9
            ,outMuls_5__8,outMuls_5__7,outMuls_5__6,outMuls_5__5,outMuls_5__4,
            outMuls_5__3,outMuls_5__2,outMuls_5__1,outMuls_5__0}), .B ({
            currentPage_5__15,currentPage_5__14,currentPage_5__13,
            currentPage_5__12,currentPage_5__11,currentPage_5__10,
            currentPage_5__9,currentPage_5__8,currentPage_5__7,currentPage_5__6,
            currentPage_5__5,currentPage_5__4,currentPage_5__3,currentPage_5__2,
            currentPage_5__1,currentPage_5__0}), .S (nx1946), .C ({
            addersInputs_5__15,addersInputs_5__14,addersInputs_5__13,
            addersInputs_5__12,addersInputs_5__11,addersInputs_5__10,
            addersInputs_5__9,addersInputs_5__8,addersInputs_5__7,
            addersInputs_5__6,addersInputs_5__5,addersInputs_5__4,
            addersInputs_5__3,addersInputs_5__2,addersInputs_5__1,
            addersInputs_5__0})) ;
    Mux2_16 loop1_6_inputAddersMap (.A ({outMuls_6__15,outMuls_6__14,
            outMuls_6__13,outMuls_6__12,outMuls_6__11,outMuls_6__10,outMuls_6__9
            ,outMuls_6__8,outMuls_6__7,outMuls_6__6,outMuls_6__5,outMuls_6__4,
            outMuls_6__3,outMuls_6__2,outMuls_6__1,outMuls_6__0}), .B ({
            currentPage_6__15,currentPage_6__14,currentPage_6__13,
            currentPage_6__12,currentPage_6__11,currentPage_6__10,
            currentPage_6__9,currentPage_6__8,currentPage_6__7,currentPage_6__6,
            currentPage_6__5,currentPage_6__4,currentPage_6__3,currentPage_6__2,
            currentPage_6__1,currentPage_6__0}), .S (nx1946), .C ({
            addersInputs_6__15,addersInputs_6__14,addersInputs_6__13,
            addersInputs_6__12,addersInputs_6__11,addersInputs_6__10,
            addersInputs_6__9,addersInputs_6__8,addersInputs_6__7,
            addersInputs_6__6,addersInputs_6__5,addersInputs_6__4,
            addersInputs_6__3,addersInputs_6__2,addersInputs_6__1,
            addersInputs_6__0})) ;
    Mux2_16 loop1_7_inputAddersMap (.A ({outMuls_7__15,outMuls_7__14,
            outMuls_7__13,outMuls_7__12,outMuls_7__11,outMuls_7__10,outMuls_7__9
            ,outMuls_7__8,outMuls_7__7,outMuls_7__6,outMuls_7__5,outMuls_7__4,
            outMuls_7__3,outMuls_7__2,outMuls_7__1,outMuls_7__0}), .B ({
            currentPage_7__15,currentPage_7__14,currentPage_7__13,
            currentPage_7__12,currentPage_7__11,currentPage_7__10,
            currentPage_7__9,currentPage_7__8,currentPage_7__7,currentPage_7__6,
            currentPage_7__5,currentPage_7__4,currentPage_7__3,currentPage_7__2,
            currentPage_7__1,currentPage_7__0}), .S (nx1948), .C ({
            addersInputs_7__15,addersInputs_7__14,addersInputs_7__13,
            addersInputs_7__12,addersInputs_7__11,addersInputs_7__10,
            addersInputs_7__9,addersInputs_7__8,addersInputs_7__7,
            addersInputs_7__6,addersInputs_7__5,addersInputs_7__4,
            addersInputs_7__3,addersInputs_7__2,addersInputs_7__1,
            addersInputs_7__0})) ;
    Mux2_16 loop1_8_inputAddersMap (.A ({outMuls_8__15,outMuls_8__14,
            outMuls_8__13,outMuls_8__12,outMuls_8__11,outMuls_8__10,outMuls_8__9
            ,outMuls_8__8,outMuls_8__7,outMuls_8__6,outMuls_8__5,outMuls_8__4,
            outMuls_8__3,outMuls_8__2,outMuls_8__1,outMuls_8__0}), .B ({
            currentPage_8__15,currentPage_8__14,currentPage_8__13,
            currentPage_8__12,currentPage_8__11,currentPage_8__10,
            currentPage_8__9,currentPage_8__8,currentPage_8__7,currentPage_8__6,
            currentPage_8__5,currentPage_8__4,currentPage_8__3,currentPage_8__2,
            currentPage_8__1,currentPage_8__0}), .S (nx1948), .C ({
            addersInputs_8__15,addersInputs_8__14,addersInputs_8__13,
            addersInputs_8__12,addersInputs_8__11,addersInputs_8__10,
            addersInputs_8__9,addersInputs_8__8,addersInputs_8__7,
            addersInputs_8__6,addersInputs_8__5,addersInputs_8__4,
            addersInputs_8__3,addersInputs_8__2,addersInputs_8__1,
            addersInputs_8__0})) ;
    Mux2_16 loop1_9_inputAddersMap (.A ({outMuls_9__15,outMuls_9__14,
            outMuls_9__13,outMuls_9__12,outMuls_9__11,outMuls_9__10,outMuls_9__9
            ,outMuls_9__8,outMuls_9__7,outMuls_9__6,outMuls_9__5,outMuls_9__4,
            outMuls_9__3,outMuls_9__2,outMuls_9__1,outMuls_9__0}), .B ({
            currentPage_9__15,currentPage_9__14,currentPage_9__13,
            currentPage_9__12,currentPage_9__11,currentPage_9__10,
            currentPage_9__9,currentPage_9__8,currentPage_9__7,currentPage_9__6,
            currentPage_9__5,currentPage_9__4,currentPage_9__3,currentPage_9__2,
            currentPage_9__1,currentPage_9__0}), .S (nx1948), .C ({
            addersInputs_9__15,addersInputs_9__14,addersInputs_9__13,
            addersInputs_9__12,addersInputs_9__11,addersInputs_9__10,
            addersInputs_9__9,addersInputs_9__8,addersInputs_9__7,
            addersInputs_9__6,addersInputs_9__5,addersInputs_9__4,
            addersInputs_9__3,addersInputs_9__2,addersInputs_9__1,
            addersInputs_9__0})) ;
    Mux2_16 loop1_10_inputAddersMap (.A ({outMuls_10__15,outMuls_10__14,
            outMuls_10__13,outMuls_10__12,outMuls_10__11,outMuls_10__10,
            outMuls_10__9,outMuls_10__8,outMuls_10__7,outMuls_10__6,
            outMuls_10__5,outMuls_10__4,outMuls_10__3,outMuls_10__2,
            outMuls_10__1,outMuls_10__0}), .B ({currentPage_10__15,
            currentPage_10__14,currentPage_10__13,currentPage_10__12,
            currentPage_10__11,currentPage_10__10,currentPage_10__9,
            currentPage_10__8,currentPage_10__7,currentPage_10__6,
            currentPage_10__5,currentPage_10__4,currentPage_10__3,
            currentPage_10__2,currentPage_10__1,currentPage_10__0}), .S (nx1948)
            , .C ({addersInputs_10__15,addersInputs_10__14,addersInputs_10__13,
            addersInputs_10__12,addersInputs_10__11,addersInputs_10__10,
            addersInputs_10__9,addersInputs_10__8,addersInputs_10__7,
            addersInputs_10__6,addersInputs_10__5,addersInputs_10__4,
            addersInputs_10__3,addersInputs_10__2,addersInputs_10__1,
            addersInputs_10__0})) ;
    Mux2_16 loop1_11_inputAddersMap (.A ({outMuls_11__15,outMuls_11__14,
            outMuls_11__13,outMuls_11__12,outMuls_11__11,outMuls_11__10,
            outMuls_11__9,outMuls_11__8,outMuls_11__7,outMuls_11__6,
            outMuls_11__5,outMuls_11__4,outMuls_11__3,outMuls_11__2,
            outMuls_11__1,outMuls_11__0}), .B ({currentPage_11__15,
            currentPage_11__14,currentPage_11__13,currentPage_11__12,
            currentPage_11__11,currentPage_11__10,currentPage_11__9,
            currentPage_11__8,currentPage_11__7,currentPage_11__6,
            currentPage_11__5,currentPage_11__4,currentPage_11__3,
            currentPage_11__2,currentPage_11__1,currentPage_11__0}), .S (nx1948)
            , .C ({addersInputs_11__15,addersInputs_11__14,addersInputs_11__13,
            addersInputs_11__12,addersInputs_11__11,addersInputs_11__10,
            addersInputs_11__9,addersInputs_11__8,addersInputs_11__7,
            addersInputs_11__6,addersInputs_11__5,addersInputs_11__4,
            addersInputs_11__3,addersInputs_11__2,addersInputs_11__1,
            addersInputs_11__0})) ;
    Mux2_16 loop1_12_inputAddersMap (.A ({outMuls_12__15,outMuls_12__14,
            outMuls_12__13,outMuls_12__12,outMuls_12__11,outMuls_12__10,
            outMuls_12__9,outMuls_12__8,outMuls_12__7,outMuls_12__6,
            outMuls_12__5,outMuls_12__4,outMuls_12__3,outMuls_12__2,
            outMuls_12__1,outMuls_12__0}), .B ({currentPage_12__15,
            currentPage_12__14,currentPage_12__13,currentPage_12__12,
            currentPage_12__11,currentPage_12__10,currentPage_12__9,
            currentPage_12__8,currentPage_12__7,currentPage_12__6,
            currentPage_12__5,currentPage_12__4,currentPage_12__3,
            currentPage_12__2,currentPage_12__1,currentPage_12__0}), .S (nx1948)
            , .C ({addersInputs_12__15,addersInputs_12__14,addersInputs_12__13,
            addersInputs_12__12,addersInputs_12__11,addersInputs_12__10,
            addersInputs_12__9,addersInputs_12__8,addersInputs_12__7,
            addersInputs_12__6,addersInputs_12__5,addersInputs_12__4,
            addersInputs_12__3,addersInputs_12__2,addersInputs_12__1,
            addersInputs_12__0})) ;
    Mux2_16 loop1_13_inputAddersMap (.A ({outMuls_13__15,outMuls_13__14,
            outMuls_13__13,outMuls_13__12,outMuls_13__11,outMuls_13__10,
            outMuls_13__9,outMuls_13__8,outMuls_13__7,outMuls_13__6,
            outMuls_13__5,outMuls_13__4,outMuls_13__3,outMuls_13__2,
            outMuls_13__1,outMuls_13__0}), .B ({currentPage_13__15,
            currentPage_13__14,currentPage_13__13,currentPage_13__12,
            currentPage_13__11,currentPage_13__10,currentPage_13__9,
            currentPage_13__8,currentPage_13__7,currentPage_13__6,
            currentPage_13__5,currentPage_13__4,currentPage_13__3,
            currentPage_13__2,currentPage_13__1,currentPage_13__0}), .S (nx1948)
            , .C ({addersInputs_13__15,addersInputs_13__14,addersInputs_13__13,
            addersInputs_13__12,addersInputs_13__11,addersInputs_13__10,
            addersInputs_13__9,addersInputs_13__8,addersInputs_13__7,
            addersInputs_13__6,addersInputs_13__5,addersInputs_13__4,
            addersInputs_13__3,addersInputs_13__2,addersInputs_13__1,
            addersInputs_13__0})) ;
    Mux2_16 loop1_14_inputAddersMap (.A ({outMuls_14__15,outMuls_14__14,
            outMuls_14__13,outMuls_14__12,outMuls_14__11,outMuls_14__10,
            outMuls_14__9,outMuls_14__8,outMuls_14__7,outMuls_14__6,
            outMuls_14__5,outMuls_14__4,outMuls_14__3,outMuls_14__2,
            outMuls_14__1,outMuls_14__0}), .B ({currentPage_14__15,
            currentPage_14__14,currentPage_14__13,currentPage_14__12,
            currentPage_14__11,currentPage_14__10,currentPage_14__9,
            currentPage_14__8,currentPage_14__7,currentPage_14__6,
            currentPage_14__5,currentPage_14__4,currentPage_14__3,
            currentPage_14__2,currentPage_14__1,currentPage_14__0}), .S (nx1950)
            , .C ({addersInputs_14__15,addersInputs_14__14,addersInputs_14__13,
            addersInputs_14__12,addersInputs_14__11,addersInputs_14__10,
            addersInputs_14__9,addersInputs_14__8,addersInputs_14__7,
            addersInputs_14__6,addersInputs_14__5,addersInputs_14__4,
            addersInputs_14__3,addersInputs_14__2,addersInputs_14__1,
            addersInputs_14__0})) ;
    Mux2_16 loop1_15_inputAddersMap (.A ({outMuls_15__15,outMuls_15__14,
            outMuls_15__13,outMuls_15__12,outMuls_15__11,outMuls_15__10,
            outMuls_15__9,outMuls_15__8,outMuls_15__7,outMuls_15__6,
            outMuls_15__5,outMuls_15__4,outMuls_15__3,outMuls_15__2,
            outMuls_15__1,outMuls_15__0}), .B ({currentPage_15__15,
            currentPage_15__14,currentPage_15__13,currentPage_15__12,
            currentPage_15__11,currentPage_15__10,currentPage_15__9,
            currentPage_15__8,currentPage_15__7,currentPage_15__6,
            currentPage_15__5,currentPage_15__4,currentPage_15__3,
            currentPage_15__2,currentPage_15__1,currentPage_15__0}), .S (nx1950)
            , .C ({addersInputs_15__15,addersInputs_15__14,addersInputs_15__13,
            addersInputs_15__12,addersInputs_15__11,addersInputs_15__10,
            addersInputs_15__9,addersInputs_15__8,addersInputs_15__7,
            addersInputs_15__6,addersInputs_15__5,addersInputs_15__4,
            addersInputs_15__3,addersInputs_15__2,addersInputs_15__1,
            addersInputs_15__0})) ;
    Mux2_16 loop1_16_inputAddersMap (.A ({outMuls_16__15,outMuls_16__14,
            outMuls_16__13,outMuls_16__12,outMuls_16__11,outMuls_16__10,
            outMuls_16__9,outMuls_16__8,outMuls_16__7,outMuls_16__6,
            outMuls_16__5,outMuls_16__4,outMuls_16__3,outMuls_16__2,
            outMuls_16__1,outMuls_16__0}), .B ({currentPage_16__15,
            currentPage_16__14,currentPage_16__13,currentPage_16__12,
            currentPage_16__11,currentPage_16__10,currentPage_16__9,
            currentPage_16__8,currentPage_16__7,currentPage_16__6,
            currentPage_16__5,currentPage_16__4,currentPage_16__3,
            currentPage_16__2,currentPage_16__1,currentPage_16__0}), .S (nx1950)
            , .C ({addersInputs_16__15,addersInputs_16__14,addersInputs_16__13,
            addersInputs_16__12,addersInputs_16__11,addersInputs_16__10,
            addersInputs_16__9,addersInputs_16__8,addersInputs_16__7,
            addersInputs_16__6,addersInputs_16__5,addersInputs_16__4,
            addersInputs_16__3,addersInputs_16__2,addersInputs_16__1,
            addersInputs_16__0})) ;
    Mux2_16 loop1_17_inputAddersMap (.A ({outMuls_17__15,outMuls_17__14,
            outMuls_17__13,outMuls_17__12,outMuls_17__11,outMuls_17__10,
            outMuls_17__9,outMuls_17__8,outMuls_17__7,outMuls_17__6,
            outMuls_17__5,outMuls_17__4,outMuls_17__3,outMuls_17__2,
            outMuls_17__1,outMuls_17__0}), .B ({currentPage_17__15,
            currentPage_17__14,currentPage_17__13,currentPage_17__12,
            currentPage_17__11,currentPage_17__10,currentPage_17__9,
            currentPage_17__8,currentPage_17__7,currentPage_17__6,
            currentPage_17__5,currentPage_17__4,currentPage_17__3,
            currentPage_17__2,currentPage_17__1,currentPage_17__0}), .S (nx1950)
            , .C ({addersInputs_17__15,addersInputs_17__14,addersInputs_17__13,
            addersInputs_17__12,addersInputs_17__11,addersInputs_17__10,
            addersInputs_17__9,addersInputs_17__8,addersInputs_17__7,
            addersInputs_17__6,addersInputs_17__5,addersInputs_17__4,
            addersInputs_17__3,addersInputs_17__2,addersInputs_17__1,
            addersInputs_17__0})) ;
    Mux2_16 loop1_18_inputAddersMap (.A ({outMuls_18__15,outMuls_18__14,
            outMuls_18__13,outMuls_18__12,outMuls_18__11,outMuls_18__10,
            outMuls_18__9,outMuls_18__8,outMuls_18__7,outMuls_18__6,
            outMuls_18__5,outMuls_18__4,outMuls_18__3,outMuls_18__2,
            outMuls_18__1,outMuls_18__0}), .B ({currentPage_18__15,
            currentPage_18__14,currentPage_18__13,currentPage_18__12,
            currentPage_18__11,currentPage_18__10,currentPage_18__9,
            currentPage_18__8,currentPage_18__7,currentPage_18__6,
            currentPage_18__5,currentPage_18__4,currentPage_18__3,
            currentPage_18__2,currentPage_18__1,currentPage_18__0}), .S (nx1950)
            , .C ({addersInputs_18__15,addersInputs_18__14,addersInputs_18__13,
            addersInputs_18__12,addersInputs_18__11,addersInputs_18__10,
            addersInputs_18__9,addersInputs_18__8,addersInputs_18__7,
            addersInputs_18__6,addersInputs_18__5,addersInputs_18__4,
            addersInputs_18__3,addersInputs_18__2,addersInputs_18__1,
            addersInputs_18__0})) ;
    Mux2_16 loop1_19_inputAddersMap (.A ({outMuls_19__15,outMuls_19__14,
            outMuls_19__13,outMuls_19__12,outMuls_19__11,outMuls_19__10,
            outMuls_19__9,outMuls_19__8,outMuls_19__7,outMuls_19__6,
            outMuls_19__5,outMuls_19__4,outMuls_19__3,outMuls_19__2,
            outMuls_19__1,outMuls_19__0}), .B ({currentPage_19__15,
            currentPage_19__14,currentPage_19__13,currentPage_19__12,
            currentPage_19__11,currentPage_19__10,currentPage_19__9,
            currentPage_19__8,currentPage_19__7,currentPage_19__6,
            currentPage_19__5,currentPage_19__4,currentPage_19__3,
            currentPage_19__2,currentPage_19__1,currentPage_19__0}), .S (nx1950)
            , .C ({addersInputs_19__15,addersInputs_19__14,addersInputs_19__13,
            addersInputs_19__12,addersInputs_19__11,addersInputs_19__10,
            addersInputs_19__9,addersInputs_19__8,addersInputs_19__7,
            addersInputs_19__6,addersInputs_19__5,addersInputs_19__4,
            addersInputs_19__3,addersInputs_19__2,addersInputs_19__1,
            addersInputs_19__0})) ;
    Mux2_16 loop1_20_inputAddersMap (.A ({outMuls_20__15,outMuls_20__14,
            outMuls_20__13,outMuls_20__12,outMuls_20__11,outMuls_20__10,
            outMuls_20__9,outMuls_20__8,outMuls_20__7,outMuls_20__6,
            outMuls_20__5,outMuls_20__4,outMuls_20__3,outMuls_20__2,
            outMuls_20__1,outMuls_20__0}), .B ({currentPage_20__15,
            currentPage_20__14,currentPage_20__13,currentPage_20__12,
            currentPage_20__11,currentPage_20__10,currentPage_20__9,
            currentPage_20__8,currentPage_20__7,currentPage_20__6,
            currentPage_20__5,currentPage_20__4,currentPage_20__3,
            currentPage_20__2,currentPage_20__1,currentPage_20__0}), .S (nx1950)
            , .C ({addersInputs_20__15,addersInputs_20__14,addersInputs_20__13,
            addersInputs_20__12,addersInputs_20__11,addersInputs_20__10,
            addersInputs_20__9,addersInputs_20__8,addersInputs_20__7,
            addersInputs_20__6,addersInputs_20__5,addersInputs_20__4,
            addersInputs_20__3,addersInputs_20__2,addersInputs_20__1,
            addersInputs_20__0})) ;
    Mux2_16 loop1_21_inputAddersMap (.A ({outMuls_21__15,outMuls_21__14,
            outMuls_21__13,outMuls_21__12,outMuls_21__11,outMuls_21__10,
            outMuls_21__9,outMuls_21__8,outMuls_21__7,outMuls_21__6,
            outMuls_21__5,outMuls_21__4,outMuls_21__3,outMuls_21__2,
            outMuls_21__1,outMuls_21__0}), .B ({currentPage_21__15,
            currentPage_21__14,currentPage_21__13,currentPage_21__12,
            currentPage_21__11,currentPage_21__10,currentPage_21__9,
            currentPage_21__8,currentPage_21__7,currentPage_21__6,
            currentPage_21__5,currentPage_21__4,currentPage_21__3,
            currentPage_21__2,currentPage_21__1,currentPage_21__0}), .S (nx1952)
            , .C ({addersInputs_21__15,addersInputs_21__14,addersInputs_21__13,
            addersInputs_21__12,addersInputs_21__11,addersInputs_21__10,
            addersInputs_21__9,addersInputs_21__8,addersInputs_21__7,
            addersInputs_21__6,addersInputs_21__5,addersInputs_21__4,
            addersInputs_21__3,addersInputs_21__2,addersInputs_21__1,
            addersInputs_21__0})) ;
    Mux2_16 loop1_22_inputAddersMap (.A ({outMuls_22__15,outMuls_22__14,
            outMuls_22__13,outMuls_22__12,outMuls_22__11,outMuls_22__10,
            outMuls_22__9,outMuls_22__8,outMuls_22__7,outMuls_22__6,
            outMuls_22__5,outMuls_22__4,outMuls_22__3,outMuls_22__2,
            outMuls_22__1,outMuls_22__0}), .B ({currentPage_22__15,
            currentPage_22__14,currentPage_22__13,currentPage_22__12,
            currentPage_22__11,currentPage_22__10,currentPage_22__9,
            currentPage_22__8,currentPage_22__7,currentPage_22__6,
            currentPage_22__5,currentPage_22__4,currentPage_22__3,
            currentPage_22__2,currentPage_22__1,currentPage_22__0}), .S (nx1952)
            , .C ({addersInputs_22__15,addersInputs_22__14,addersInputs_22__13,
            addersInputs_22__12,addersInputs_22__11,addersInputs_22__10,
            addersInputs_22__9,addersInputs_22__8,addersInputs_22__7,
            addersInputs_22__6,addersInputs_22__5,addersInputs_22__4,
            addersInputs_22__3,addersInputs_22__2,addersInputs_22__1,
            addersInputs_22__0})) ;
    Mux2_16 loop1_23_inputAddersMap (.A ({outMuls_23__15,outMuls_23__14,
            outMuls_23__13,outMuls_23__12,outMuls_23__11,outMuls_23__10,
            outMuls_23__9,outMuls_23__8,outMuls_23__7,outMuls_23__6,
            outMuls_23__5,outMuls_23__4,outMuls_23__3,outMuls_23__2,
            outMuls_23__1,outMuls_23__0}), .B ({currentPage_23__15,
            currentPage_23__14,currentPage_23__13,currentPage_23__12,
            currentPage_23__11,currentPage_23__10,currentPage_23__9,
            currentPage_23__8,currentPage_23__7,currentPage_23__6,
            currentPage_23__5,currentPage_23__4,currentPage_23__3,
            currentPage_23__2,currentPage_23__1,currentPage_23__0}), .S (nx1952)
            , .C ({addersInputs_23__15,addersInputs_23__14,addersInputs_23__13,
            addersInputs_23__12,addersInputs_23__11,addersInputs_23__10,
            addersInputs_23__9,addersInputs_23__8,addersInputs_23__7,
            addersInputs_23__6,addersInputs_23__5,addersInputs_23__4,
            addersInputs_23__3,addersInputs_23__2,addersInputs_23__1,
            addersInputs_23__0})) ;
    Mux2_16 loop1_24_inputAddersMap (.A ({outMuls_24__15,outMuls_24__14,
            outMuls_24__13,outMuls_24__12,outMuls_24__11,outMuls_24__10,
            outMuls_24__9,outMuls_24__8,outMuls_24__7,outMuls_24__6,
            outMuls_24__5,outMuls_24__4,outMuls_24__3,outMuls_24__2,
            outMuls_24__1,outMuls_24__0}), .B ({currentPage_24__15,
            currentPage_24__14,currentPage_24__13,currentPage_24__12,
            currentPage_24__11,currentPage_24__10,currentPage_24__9,
            currentPage_24__8,currentPage_24__7,currentPage_24__6,
            currentPage_24__5,currentPage_24__4,currentPage_24__3,
            currentPage_24__2,currentPage_24__1,currentPage_24__0}), .S (nx1952)
            , .C ({addersInputs_24__15,addersInputs_24__14,addersInputs_24__13,
            addersInputs_24__12,addersInputs_24__11,addersInputs_24__10,
            addersInputs_24__9,addersInputs_24__8,addersInputs_24__7,
            addersInputs_24__6,addersInputs_24__5,addersInputs_24__4,
            addersInputs_24__3,addersInputs_24__2,addersInputs_24__1,
            addersInputs_24__0})) ;
    CNNAdders_16 addersMap (.inputs_0__15 (addersInputs_0__15), .inputs_0__14 (
                 addersInputs_0__14), .inputs_0__13 (addersInputs_0__13), .inputs_0__12 (
                 addersInputs_0__12), .inputs_0__11 (addersInputs_0__11), .inputs_0__10 (
                 addersInputs_0__10), .inputs_0__9 (addersInputs_0__9), .inputs_0__8 (
                 addersInputs_0__8), .inputs_0__7 (addersInputs_0__7), .inputs_0__6 (
                 addersInputs_0__6), .inputs_0__5 (addersInputs_0__5), .inputs_0__4 (
                 addersInputs_0__4), .inputs_0__3 (addersInputs_0__3), .inputs_0__2 (
                 addersInputs_0__2), .inputs_0__1 (addersInputs_0__1), .inputs_0__0 (
                 addersInputs_0__0), .inputs_1__15 (addersInputs_1__15), .inputs_1__14 (
                 addersInputs_1__14), .inputs_1__13 (addersInputs_1__13), .inputs_1__12 (
                 addersInputs_1__12), .inputs_1__11 (addersInputs_1__11), .inputs_1__10 (
                 addersInputs_1__10), .inputs_1__9 (addersInputs_1__9), .inputs_1__8 (
                 addersInputs_1__8), .inputs_1__7 (addersInputs_1__7), .inputs_1__6 (
                 addersInputs_1__6), .inputs_1__5 (addersInputs_1__5), .inputs_1__4 (
                 addersInputs_1__4), .inputs_1__3 (addersInputs_1__3), .inputs_1__2 (
                 addersInputs_1__2), .inputs_1__1 (addersInputs_1__1), .inputs_1__0 (
                 addersInputs_1__0), .inputs_2__15 (addersInputs_2__15), .inputs_2__14 (
                 addersInputs_2__14), .inputs_2__13 (addersInputs_2__13), .inputs_2__12 (
                 addersInputs_2__12), .inputs_2__11 (addersInputs_2__11), .inputs_2__10 (
                 addersInputs_2__10), .inputs_2__9 (addersInputs_2__9), .inputs_2__8 (
                 addersInputs_2__8), .inputs_2__7 (addersInputs_2__7), .inputs_2__6 (
                 addersInputs_2__6), .inputs_2__5 (addersInputs_2__5), .inputs_2__4 (
                 addersInputs_2__4), .inputs_2__3 (addersInputs_2__3), .inputs_2__2 (
                 addersInputs_2__2), .inputs_2__1 (addersInputs_2__1), .inputs_2__0 (
                 addersInputs_2__0), .inputs_3__15 (addersInputs_3__15), .inputs_3__14 (
                 addersInputs_3__14), .inputs_3__13 (addersInputs_3__13), .inputs_3__12 (
                 addersInputs_3__12), .inputs_3__11 (addersInputs_3__11), .inputs_3__10 (
                 addersInputs_3__10), .inputs_3__9 (addersInputs_3__9), .inputs_3__8 (
                 addersInputs_3__8), .inputs_3__7 (addersInputs_3__7), .inputs_3__6 (
                 addersInputs_3__6), .inputs_3__5 (addersInputs_3__5), .inputs_3__4 (
                 addersInputs_3__4), .inputs_3__3 (addersInputs_3__3), .inputs_3__2 (
                 addersInputs_3__2), .inputs_3__1 (addersInputs_3__1), .inputs_3__0 (
                 addersInputs_3__0), .inputs_4__15 (addersInputs_4__15), .inputs_4__14 (
                 addersInputs_4__14), .inputs_4__13 (addersInputs_4__13), .inputs_4__12 (
                 addersInputs_4__12), .inputs_4__11 (addersInputs_4__11), .inputs_4__10 (
                 addersInputs_4__10), .inputs_4__9 (addersInputs_4__9), .inputs_4__8 (
                 addersInputs_4__8), .inputs_4__7 (addersInputs_4__7), .inputs_4__6 (
                 addersInputs_4__6), .inputs_4__5 (addersInputs_4__5), .inputs_4__4 (
                 addersInputs_4__4), .inputs_4__3 (addersInputs_4__3), .inputs_4__2 (
                 addersInputs_4__2), .inputs_4__1 (addersInputs_4__1), .inputs_4__0 (
                 addersInputs_4__0), .inputs_5__15 (addersInputs_5__15), .inputs_5__14 (
                 addersInputs_5__14), .inputs_5__13 (addersInputs_5__13), .inputs_5__12 (
                 addersInputs_5__12), .inputs_5__11 (addersInputs_5__11), .inputs_5__10 (
                 addersInputs_5__10), .inputs_5__9 (addersInputs_5__9), .inputs_5__8 (
                 addersInputs_5__8), .inputs_5__7 (addersInputs_5__7), .inputs_5__6 (
                 addersInputs_5__6), .inputs_5__5 (addersInputs_5__5), .inputs_5__4 (
                 addersInputs_5__4), .inputs_5__3 (addersInputs_5__3), .inputs_5__2 (
                 addersInputs_5__2), .inputs_5__1 (addersInputs_5__1), .inputs_5__0 (
                 addersInputs_5__0), .inputs_6__15 (addersInputs_6__15), .inputs_6__14 (
                 addersInputs_6__14), .inputs_6__13 (addersInputs_6__13), .inputs_6__12 (
                 addersInputs_6__12), .inputs_6__11 (addersInputs_6__11), .inputs_6__10 (
                 addersInputs_6__10), .inputs_6__9 (addersInputs_6__9), .inputs_6__8 (
                 addersInputs_6__8), .inputs_6__7 (addersInputs_6__7), .inputs_6__6 (
                 addersInputs_6__6), .inputs_6__5 (addersInputs_6__5), .inputs_6__4 (
                 addersInputs_6__4), .inputs_6__3 (addersInputs_6__3), .inputs_6__2 (
                 addersInputs_6__2), .inputs_6__1 (addersInputs_6__1), .inputs_6__0 (
                 addersInputs_6__0), .inputs_7__15 (addersInputs_7__15), .inputs_7__14 (
                 addersInputs_7__14), .inputs_7__13 (addersInputs_7__13), .inputs_7__12 (
                 addersInputs_7__12), .inputs_7__11 (addersInputs_7__11), .inputs_7__10 (
                 addersInputs_7__10), .inputs_7__9 (addersInputs_7__9), .inputs_7__8 (
                 addersInputs_7__8), .inputs_7__7 (addersInputs_7__7), .inputs_7__6 (
                 addersInputs_7__6), .inputs_7__5 (addersInputs_7__5), .inputs_7__4 (
                 addersInputs_7__4), .inputs_7__3 (addersInputs_7__3), .inputs_7__2 (
                 addersInputs_7__2), .inputs_7__1 (addersInputs_7__1), .inputs_7__0 (
                 addersInputs_7__0), .inputs_8__15 (addersInputs_8__15), .inputs_8__14 (
                 addersInputs_8__14), .inputs_8__13 (addersInputs_8__13), .inputs_8__12 (
                 addersInputs_8__12), .inputs_8__11 (addersInputs_8__11), .inputs_8__10 (
                 addersInputs_8__10), .inputs_8__9 (addersInputs_8__9), .inputs_8__8 (
                 addersInputs_8__8), .inputs_8__7 (addersInputs_8__7), .inputs_8__6 (
                 addersInputs_8__6), .inputs_8__5 (addersInputs_8__5), .inputs_8__4 (
                 addersInputs_8__4), .inputs_8__3 (addersInputs_8__3), .inputs_8__2 (
                 addersInputs_8__2), .inputs_8__1 (addersInputs_8__1), .inputs_8__0 (
                 addersInputs_8__0), .inputs_9__15 (addersInputs_9__15), .inputs_9__14 (
                 addersInputs_9__14), .inputs_9__13 (addersInputs_9__13), .inputs_9__12 (
                 addersInputs_9__12), .inputs_9__11 (addersInputs_9__11), .inputs_9__10 (
                 addersInputs_9__10), .inputs_9__9 (addersInputs_9__9), .inputs_9__8 (
                 addersInputs_9__8), .inputs_9__7 (addersInputs_9__7), .inputs_9__6 (
                 addersInputs_9__6), .inputs_9__5 (addersInputs_9__5), .inputs_9__4 (
                 addersInputs_9__4), .inputs_9__3 (addersInputs_9__3), .inputs_9__2 (
                 addersInputs_9__2), .inputs_9__1 (addersInputs_9__1), .inputs_9__0 (
                 addersInputs_9__0), .inputs_10__15 (addersInputs_10__15), .inputs_10__14 (
                 addersInputs_10__14), .inputs_10__13 (addersInputs_10__13), .inputs_10__12 (
                 addersInputs_10__12), .inputs_10__11 (addersInputs_10__11), .inputs_10__10 (
                 addersInputs_10__10), .inputs_10__9 (addersInputs_10__9), .inputs_10__8 (
                 addersInputs_10__8), .inputs_10__7 (addersInputs_10__7), .inputs_10__6 (
                 addersInputs_10__6), .inputs_10__5 (addersInputs_10__5), .inputs_10__4 (
                 addersInputs_10__4), .inputs_10__3 (addersInputs_10__3), .inputs_10__2 (
                 addersInputs_10__2), .inputs_10__1 (addersInputs_10__1), .inputs_10__0 (
                 addersInputs_10__0), .inputs_11__15 (addersInputs_11__15), .inputs_11__14 (
                 addersInputs_11__14), .inputs_11__13 (addersInputs_11__13), .inputs_11__12 (
                 addersInputs_11__12), .inputs_11__11 (addersInputs_11__11), .inputs_11__10 (
                 addersInputs_11__10), .inputs_11__9 (addersInputs_11__9), .inputs_11__8 (
                 addersInputs_11__8), .inputs_11__7 (addersInputs_11__7), .inputs_11__6 (
                 addersInputs_11__6), .inputs_11__5 (addersInputs_11__5), .inputs_11__4 (
                 addersInputs_11__4), .inputs_11__3 (addersInputs_11__3), .inputs_11__2 (
                 addersInputs_11__2), .inputs_11__1 (addersInputs_11__1), .inputs_11__0 (
                 addersInputs_11__0), .inputs_12__15 (addersInputs_12__15), .inputs_12__14 (
                 addersInputs_12__14), .inputs_12__13 (addersInputs_12__13), .inputs_12__12 (
                 addersInputs_12__12), .inputs_12__11 (addersInputs_12__11), .inputs_12__10 (
                 addersInputs_12__10), .inputs_12__9 (addersInputs_12__9), .inputs_12__8 (
                 addersInputs_12__8), .inputs_12__7 (addersInputs_12__7), .inputs_12__6 (
                 addersInputs_12__6), .inputs_12__5 (addersInputs_12__5), .inputs_12__4 (
                 addersInputs_12__4), .inputs_12__3 (addersInputs_12__3), .inputs_12__2 (
                 addersInputs_12__2), .inputs_12__1 (addersInputs_12__1), .inputs_12__0 (
                 addersInputs_12__0), .inputs_13__15 (addersInputs_13__15), .inputs_13__14 (
                 addersInputs_13__14), .inputs_13__13 (addersInputs_13__13), .inputs_13__12 (
                 addersInputs_13__12), .inputs_13__11 (addersInputs_13__11), .inputs_13__10 (
                 addersInputs_13__10), .inputs_13__9 (addersInputs_13__9), .inputs_13__8 (
                 addersInputs_13__8), .inputs_13__7 (addersInputs_13__7), .inputs_13__6 (
                 addersInputs_13__6), .inputs_13__5 (addersInputs_13__5), .inputs_13__4 (
                 addersInputs_13__4), .inputs_13__3 (addersInputs_13__3), .inputs_13__2 (
                 addersInputs_13__2), .inputs_13__1 (addersInputs_13__1), .inputs_13__0 (
                 addersInputs_13__0), .inputs_14__15 (addersInputs_14__15), .inputs_14__14 (
                 addersInputs_14__14), .inputs_14__13 (addersInputs_14__13), .inputs_14__12 (
                 addersInputs_14__12), .inputs_14__11 (addersInputs_14__11), .inputs_14__10 (
                 addersInputs_14__10), .inputs_14__9 (addersInputs_14__9), .inputs_14__8 (
                 addersInputs_14__8), .inputs_14__7 (addersInputs_14__7), .inputs_14__6 (
                 addersInputs_14__6), .inputs_14__5 (addersInputs_14__5), .inputs_14__4 (
                 addersInputs_14__4), .inputs_14__3 (addersInputs_14__3), .inputs_14__2 (
                 addersInputs_14__2), .inputs_14__1 (addersInputs_14__1), .inputs_14__0 (
                 addersInputs_14__0), .inputs_15__15 (addersInputs_15__15), .inputs_15__14 (
                 addersInputs_15__14), .inputs_15__13 (addersInputs_15__13), .inputs_15__12 (
                 addersInputs_15__12), .inputs_15__11 (addersInputs_15__11), .inputs_15__10 (
                 addersInputs_15__10), .inputs_15__9 (addersInputs_15__9), .inputs_15__8 (
                 addersInputs_15__8), .inputs_15__7 (addersInputs_15__7), .inputs_15__6 (
                 addersInputs_15__6), .inputs_15__5 (addersInputs_15__5), .inputs_15__4 (
                 addersInputs_15__4), .inputs_15__3 (addersInputs_15__3), .inputs_15__2 (
                 addersInputs_15__2), .inputs_15__1 (addersInputs_15__1), .inputs_15__0 (
                 addersInputs_15__0), .inputs_16__15 (addersInputs_16__15), .inputs_16__14 (
                 addersInputs_16__14), .inputs_16__13 (addersInputs_16__13), .inputs_16__12 (
                 addersInputs_16__12), .inputs_16__11 (addersInputs_16__11), .inputs_16__10 (
                 addersInputs_16__10), .inputs_16__9 (addersInputs_16__9), .inputs_16__8 (
                 addersInputs_16__8), .inputs_16__7 (addersInputs_16__7), .inputs_16__6 (
                 addersInputs_16__6), .inputs_16__5 (addersInputs_16__5), .inputs_16__4 (
                 addersInputs_16__4), .inputs_16__3 (addersInputs_16__3), .inputs_16__2 (
                 addersInputs_16__2), .inputs_16__1 (addersInputs_16__1), .inputs_16__0 (
                 addersInputs_16__0), .inputs_17__15 (addersInputs_17__15), .inputs_17__14 (
                 addersInputs_17__14), .inputs_17__13 (addersInputs_17__13), .inputs_17__12 (
                 addersInputs_17__12), .inputs_17__11 (addersInputs_17__11), .inputs_17__10 (
                 addersInputs_17__10), .inputs_17__9 (addersInputs_17__9), .inputs_17__8 (
                 addersInputs_17__8), .inputs_17__7 (addersInputs_17__7), .inputs_17__6 (
                 addersInputs_17__6), .inputs_17__5 (addersInputs_17__5), .inputs_17__4 (
                 addersInputs_17__4), .inputs_17__3 (addersInputs_17__3), .inputs_17__2 (
                 addersInputs_17__2), .inputs_17__1 (addersInputs_17__1), .inputs_17__0 (
                 addersInputs_17__0), .inputs_18__15 (addersInputs_18__15), .inputs_18__14 (
                 addersInputs_18__14), .inputs_18__13 (addersInputs_18__13), .inputs_18__12 (
                 addersInputs_18__12), .inputs_18__11 (addersInputs_18__11), .inputs_18__10 (
                 addersInputs_18__10), .inputs_18__9 (addersInputs_18__9), .inputs_18__8 (
                 addersInputs_18__8), .inputs_18__7 (addersInputs_18__7), .inputs_18__6 (
                 addersInputs_18__6), .inputs_18__5 (addersInputs_18__5), .inputs_18__4 (
                 addersInputs_18__4), .inputs_18__3 (addersInputs_18__3), .inputs_18__2 (
                 addersInputs_18__2), .inputs_18__1 (addersInputs_18__1), .inputs_18__0 (
                 addersInputs_18__0), .inputs_19__15 (addersInputs_19__15), .inputs_19__14 (
                 addersInputs_19__14), .inputs_19__13 (addersInputs_19__13), .inputs_19__12 (
                 addersInputs_19__12), .inputs_19__11 (addersInputs_19__11), .inputs_19__10 (
                 addersInputs_19__10), .inputs_19__9 (addersInputs_19__9), .inputs_19__8 (
                 addersInputs_19__8), .inputs_19__7 (addersInputs_19__7), .inputs_19__6 (
                 addersInputs_19__6), .inputs_19__5 (addersInputs_19__5), .inputs_19__4 (
                 addersInputs_19__4), .inputs_19__3 (addersInputs_19__3), .inputs_19__2 (
                 addersInputs_19__2), .inputs_19__1 (addersInputs_19__1), .inputs_19__0 (
                 addersInputs_19__0), .inputs_20__15 (addersInputs_20__15), .inputs_20__14 (
                 addersInputs_20__14), .inputs_20__13 (addersInputs_20__13), .inputs_20__12 (
                 addersInputs_20__12), .inputs_20__11 (addersInputs_20__11), .inputs_20__10 (
                 addersInputs_20__10), .inputs_20__9 (addersInputs_20__9), .inputs_20__8 (
                 addersInputs_20__8), .inputs_20__7 (addersInputs_20__7), .inputs_20__6 (
                 addersInputs_20__6), .inputs_20__5 (addersInputs_20__5), .inputs_20__4 (
                 addersInputs_20__4), .inputs_20__3 (addersInputs_20__3), .inputs_20__2 (
                 addersInputs_20__2), .inputs_20__1 (addersInputs_20__1), .inputs_20__0 (
                 addersInputs_20__0), .inputs_21__15 (addersInputs_21__15), .inputs_21__14 (
                 addersInputs_21__14), .inputs_21__13 (addersInputs_21__13), .inputs_21__12 (
                 addersInputs_21__12), .inputs_21__11 (addersInputs_21__11), .inputs_21__10 (
                 addersInputs_21__10), .inputs_21__9 (addersInputs_21__9), .inputs_21__8 (
                 addersInputs_21__8), .inputs_21__7 (addersInputs_21__7), .inputs_21__6 (
                 addersInputs_21__6), .inputs_21__5 (addersInputs_21__5), .inputs_21__4 (
                 addersInputs_21__4), .inputs_21__3 (addersInputs_21__3), .inputs_21__2 (
                 addersInputs_21__2), .inputs_21__1 (addersInputs_21__1), .inputs_21__0 (
                 addersInputs_21__0), .inputs_22__15 (addersInputs_22__15), .inputs_22__14 (
                 addersInputs_22__14), .inputs_22__13 (addersInputs_22__13), .inputs_22__12 (
                 addersInputs_22__12), .inputs_22__11 (addersInputs_22__11), .inputs_22__10 (
                 addersInputs_22__10), .inputs_22__9 (addersInputs_22__9), .inputs_22__8 (
                 addersInputs_22__8), .inputs_22__7 (addersInputs_22__7), .inputs_22__6 (
                 addersInputs_22__6), .inputs_22__5 (addersInputs_22__5), .inputs_22__4 (
                 addersInputs_22__4), .inputs_22__3 (addersInputs_22__3), .inputs_22__2 (
                 addersInputs_22__2), .inputs_22__1 (addersInputs_22__1), .inputs_22__0 (
                 addersInputs_22__0), .inputs_23__15 (addersInputs_23__15), .inputs_23__14 (
                 addersInputs_23__14), .inputs_23__13 (addersInputs_23__13), .inputs_23__12 (
                 addersInputs_23__12), .inputs_23__11 (addersInputs_23__11), .inputs_23__10 (
                 addersInputs_23__10), .inputs_23__9 (addersInputs_23__9), .inputs_23__8 (
                 addersInputs_23__8), .inputs_23__7 (addersInputs_23__7), .inputs_23__6 (
                 addersInputs_23__6), .inputs_23__5 (addersInputs_23__5), .inputs_23__4 (
                 addersInputs_23__4), .inputs_23__3 (addersInputs_23__3), .inputs_23__2 (
                 addersInputs_23__2), .inputs_23__1 (addersInputs_23__1), .inputs_23__0 (
                 addersInputs_23__0), .inputs_24__15 (addersInputs_24__15), .inputs_24__14 (
                 addersInputs_24__14), .inputs_24__13 (addersInputs_24__13), .inputs_24__12 (
                 addersInputs_24__12), .inputs_24__11 (addersInputs_24__11), .inputs_24__10 (
                 addersInputs_24__10), .inputs_24__9 (addersInputs_24__9), .inputs_24__8 (
                 addersInputs_24__8), .inputs_24__7 (addersInputs_24__7), .inputs_24__6 (
                 addersInputs_24__6), .inputs_24__5 (addersInputs_24__5), .inputs_24__4 (
                 addersInputs_24__4), .inputs_24__3 (addersInputs_24__3), .inputs_24__2 (
                 addersInputs_24__2), .inputs_24__1 (addersInputs_24__1), .inputs_24__0 (
                 addersInputs_24__0), .filterType (filterType), .finalSum ({
                 outAdder_15,outAdder_14,outAdder_13,outAdder_12,outAdder_11,
                 outAdder_10,outAdder_9,outAdder_8,outAdder_7,outAdder_6,
                 outAdder_5,outAdder_4,outAdder_3,outAdder_2,outAdder_1,
                 outAdder_0})) ;
    CNNShifter_16 shifterMap (.A ({outAdder_15,outAdder_14,outAdder_13,
                  outAdder_12,outAdder_11,outAdder_10,outAdder_9,outAdder_8,
                  outAdder_7,outAdder_6,outAdder_5,outAdder_4,outAdder_3,nx1921,
                  nx1921,nx1921}), .filterSize (filterType), .shiftedOut ({
                  \$dummy [1],\$dummy [2],\$dummy [3],\$dummy [4],outShifter_11,
                  outShifter_10,outShifter_9,outShifter_8,outShifter_7,
                  outShifter_6,outShifter_5,outShifter_4,outShifter_3,
                  outShifter_2,outShifter_1,outShifter_0})) ;
    Mux2_16 finalOutMap (.A ({outAdder_15,outAdder_14,outAdder_13,outAdder_12,
            outAdder_11,outAdder_10,outAdder_9,outAdder_8,outAdder_7,outAdder_6,
            outAdder_5,outAdder_4,outAdder_3,outAdder_2,outAdder_1,outAdder_0})
            , .B ({outAdder_15,outAdder_15,outAdder_15,outAdder_15,outShifter_11
            ,outShifter_10,outShifter_9,outShifter_8,outShifter_7,outShifter_6,
            outShifter_5,outShifter_4,outShifter_3,outShifter_2,outShifter_1,
            outShifter_0}), .S (nx1952), .C ({finalSum_15,finalSum_14,
            finalSum_13,finalSum_12,finalSum_11,finalSum_10,finalSum_9,
            finalSum_8,finalSum_7,finalSum_6,finalSum_5,finalSum_4,finalSum_3,
            finalSum_2,finalSum_1,finalSum_0})) ;
    Reg_16 captureReg (.D ({finalSum_15,finalSum_14,finalSum_13,finalSum_12,
           finalSum_11,finalSum_10,finalSum_9,finalSum_8,finalSum_7,finalSum_6,
           finalSum_5,finalSum_4,finalSum_3,finalSum_2,finalSum_1,finalSum_0}), 
           .en (doneCores), .clk (notClk), .rst (rst), .Q ({finalSumConv[15],
           finalSumConv[14],finalSumConv[13],finalSumConv[12],finalSumConv[11],
           finalSumConv[10],finalSumConv[9],finalSumConv[8],finalSumConv[7],
           finalSumConv[6],finalSumConv[5],finalSumConv[4],finalSumConv[3],
           finalSumConv[2],finalSumConv[1],finalSumConv[0]})) ;
    fake_gnd ix1922 (.Y (nx1921)) ;
    inv01 ix1933 (.Y (notClk), .A (clk)) ;
    or02 ix3 (.Y (doneCores), .A0 (nx1952), .A1 (doneMul)) ;
    inv01 ix1943 (.Y (nx1944), .A (layerType)) ;
    inv01 ix1945 (.Y (nx1946), .A (nx1944)) ;
    inv01 ix1947 (.Y (nx1948), .A (nx1944)) ;
    inv01 ix1949 (.Y (nx1950), .A (nx1944)) ;
    inv01 ix1951 (.Y (nx1952), .A (nx1944)) ;
endmodule


module CNNShifter_16 ( A, filterSize, shiftedOut ) ;

    input [15:0]A ;
    input filterSize ;
    output [15:0]shiftedOut ;

    wire nx134, nx136;



    assign shiftedOut[15] = A[15] ;
    assign shiftedOut[14] = A[15] ;
    assign shiftedOut[13] = A[15] ;
    assign shiftedOut[12] = A[15] ;
    mux21_ni ix7 (.Y (shiftedOut[0]), .A0 (A[3]), .A1 (A[5]), .S0 (nx134)) ;
    mux21_ni ix15 (.Y (shiftedOut[1]), .A0 (A[4]), .A1 (A[6]), .S0 (nx134)) ;
    mux21_ni ix23 (.Y (shiftedOut[2]), .A0 (A[5]), .A1 (A[7]), .S0 (nx134)) ;
    mux21_ni ix31 (.Y (shiftedOut[3]), .A0 (A[6]), .A1 (A[8]), .S0 (nx134)) ;
    mux21_ni ix39 (.Y (shiftedOut[4]), .A0 (A[7]), .A1 (A[9]), .S0 (nx134)) ;
    mux21_ni ix47 (.Y (shiftedOut[5]), .A0 (A[8]), .A1 (A[10]), .S0 (nx134)) ;
    mux21_ni ix55 (.Y (shiftedOut[6]), .A0 (A[9]), .A1 (A[11]), .S0 (nx134)) ;
    mux21_ni ix63 (.Y (shiftedOut[7]), .A0 (A[10]), .A1 (A[12]), .S0 (nx136)) ;
    mux21_ni ix71 (.Y (shiftedOut[8]), .A0 (A[11]), .A1 (A[13]), .S0 (nx136)) ;
    mux21_ni ix79 (.Y (shiftedOut[9]), .A0 (A[12]), .A1 (A[14]), .S0 (nx136)) ;
    mux21_ni ix87 (.Y (shiftedOut[10]), .A0 (A[13]), .A1 (A[15]), .S0 (nx136)) ;
    mux21_ni ix95 (.Y (shiftedOut[11]), .A0 (A[14]), .A1 (A[15]), .S0 (nx136)) ;
    buf02 ix133 (.Y (nx134), .A (filterSize)) ;
    buf02 ix135 (.Y (nx136), .A (filterSize)) ;
endmodule


module CNNAdders_16 ( inputs_0__15, inputs_0__14, inputs_0__13, inputs_0__12, 
                      inputs_0__11, inputs_0__10, inputs_0__9, inputs_0__8, 
                      inputs_0__7, inputs_0__6, inputs_0__5, inputs_0__4, 
                      inputs_0__3, inputs_0__2, inputs_0__1, inputs_0__0, 
                      inputs_1__15, inputs_1__14, inputs_1__13, inputs_1__12, 
                      inputs_1__11, inputs_1__10, inputs_1__9, inputs_1__8, 
                      inputs_1__7, inputs_1__6, inputs_1__5, inputs_1__4, 
                      inputs_1__3, inputs_1__2, inputs_1__1, inputs_1__0, 
                      inputs_2__15, inputs_2__14, inputs_2__13, inputs_2__12, 
                      inputs_2__11, inputs_2__10, inputs_2__9, inputs_2__8, 
                      inputs_2__7, inputs_2__6, inputs_2__5, inputs_2__4, 
                      inputs_2__3, inputs_2__2, inputs_2__1, inputs_2__0, 
                      inputs_3__15, inputs_3__14, inputs_3__13, inputs_3__12, 
                      inputs_3__11, inputs_3__10, inputs_3__9, inputs_3__8, 
                      inputs_3__7, inputs_3__6, inputs_3__5, inputs_3__4, 
                      inputs_3__3, inputs_3__2, inputs_3__1, inputs_3__0, 
                      inputs_4__15, inputs_4__14, inputs_4__13, inputs_4__12, 
                      inputs_4__11, inputs_4__10, inputs_4__9, inputs_4__8, 
                      inputs_4__7, inputs_4__6, inputs_4__5, inputs_4__4, 
                      inputs_4__3, inputs_4__2, inputs_4__1, inputs_4__0, 
                      inputs_5__15, inputs_5__14, inputs_5__13, inputs_5__12, 
                      inputs_5__11, inputs_5__10, inputs_5__9, inputs_5__8, 
                      inputs_5__7, inputs_5__6, inputs_5__5, inputs_5__4, 
                      inputs_5__3, inputs_5__2, inputs_5__1, inputs_5__0, 
                      inputs_6__15, inputs_6__14, inputs_6__13, inputs_6__12, 
                      inputs_6__11, inputs_6__10, inputs_6__9, inputs_6__8, 
                      inputs_6__7, inputs_6__6, inputs_6__5, inputs_6__4, 
                      inputs_6__3, inputs_6__2, inputs_6__1, inputs_6__0, 
                      inputs_7__15, inputs_7__14, inputs_7__13, inputs_7__12, 
                      inputs_7__11, inputs_7__10, inputs_7__9, inputs_7__8, 
                      inputs_7__7, inputs_7__6, inputs_7__5, inputs_7__4, 
                      inputs_7__3, inputs_7__2, inputs_7__1, inputs_7__0, 
                      inputs_8__15, inputs_8__14, inputs_8__13, inputs_8__12, 
                      inputs_8__11, inputs_8__10, inputs_8__9, inputs_8__8, 
                      inputs_8__7, inputs_8__6, inputs_8__5, inputs_8__4, 
                      inputs_8__3, inputs_8__2, inputs_8__1, inputs_8__0, 
                      inputs_9__15, inputs_9__14, inputs_9__13, inputs_9__12, 
                      inputs_9__11, inputs_9__10, inputs_9__9, inputs_9__8, 
                      inputs_9__7, inputs_9__6, inputs_9__5, inputs_9__4, 
                      inputs_9__3, inputs_9__2, inputs_9__1, inputs_9__0, 
                      inputs_10__15, inputs_10__14, inputs_10__13, inputs_10__12, 
                      inputs_10__11, inputs_10__10, inputs_10__9, inputs_10__8, 
                      inputs_10__7, inputs_10__6, inputs_10__5, inputs_10__4, 
                      inputs_10__3, inputs_10__2, inputs_10__1, inputs_10__0, 
                      inputs_11__15, inputs_11__14, inputs_11__13, inputs_11__12, 
                      inputs_11__11, inputs_11__10, inputs_11__9, inputs_11__8, 
                      inputs_11__7, inputs_11__6, inputs_11__5, inputs_11__4, 
                      inputs_11__3, inputs_11__2, inputs_11__1, inputs_11__0, 
                      inputs_12__15, inputs_12__14, inputs_12__13, inputs_12__12, 
                      inputs_12__11, inputs_12__10, inputs_12__9, inputs_12__8, 
                      inputs_12__7, inputs_12__6, inputs_12__5, inputs_12__4, 
                      inputs_12__3, inputs_12__2, inputs_12__1, inputs_12__0, 
                      inputs_13__15, inputs_13__14, inputs_13__13, inputs_13__12, 
                      inputs_13__11, inputs_13__10, inputs_13__9, inputs_13__8, 
                      inputs_13__7, inputs_13__6, inputs_13__5, inputs_13__4, 
                      inputs_13__3, inputs_13__2, inputs_13__1, inputs_13__0, 
                      inputs_14__15, inputs_14__14, inputs_14__13, inputs_14__12, 
                      inputs_14__11, inputs_14__10, inputs_14__9, inputs_14__8, 
                      inputs_14__7, inputs_14__6, inputs_14__5, inputs_14__4, 
                      inputs_14__3, inputs_14__2, inputs_14__1, inputs_14__0, 
                      inputs_15__15, inputs_15__14, inputs_15__13, inputs_15__12, 
                      inputs_15__11, inputs_15__10, inputs_15__9, inputs_15__8, 
                      inputs_15__7, inputs_15__6, inputs_15__5, inputs_15__4, 
                      inputs_15__3, inputs_15__2, inputs_15__1, inputs_15__0, 
                      inputs_16__15, inputs_16__14, inputs_16__13, inputs_16__12, 
                      inputs_16__11, inputs_16__10, inputs_16__9, inputs_16__8, 
                      inputs_16__7, inputs_16__6, inputs_16__5, inputs_16__4, 
                      inputs_16__3, inputs_16__2, inputs_16__1, inputs_16__0, 
                      inputs_17__15, inputs_17__14, inputs_17__13, inputs_17__12, 
                      inputs_17__11, inputs_17__10, inputs_17__9, inputs_17__8, 
                      inputs_17__7, inputs_17__6, inputs_17__5, inputs_17__4, 
                      inputs_17__3, inputs_17__2, inputs_17__1, inputs_17__0, 
                      inputs_18__15, inputs_18__14, inputs_18__13, inputs_18__12, 
                      inputs_18__11, inputs_18__10, inputs_18__9, inputs_18__8, 
                      inputs_18__7, inputs_18__6, inputs_18__5, inputs_18__4, 
                      inputs_18__3, inputs_18__2, inputs_18__1, inputs_18__0, 
                      inputs_19__15, inputs_19__14, inputs_19__13, inputs_19__12, 
                      inputs_19__11, inputs_19__10, inputs_19__9, inputs_19__8, 
                      inputs_19__7, inputs_19__6, inputs_19__5, inputs_19__4, 
                      inputs_19__3, inputs_19__2, inputs_19__1, inputs_19__0, 
                      inputs_20__15, inputs_20__14, inputs_20__13, inputs_20__12, 
                      inputs_20__11, inputs_20__10, inputs_20__9, inputs_20__8, 
                      inputs_20__7, inputs_20__6, inputs_20__5, inputs_20__4, 
                      inputs_20__3, inputs_20__2, inputs_20__1, inputs_20__0, 
                      inputs_21__15, inputs_21__14, inputs_21__13, inputs_21__12, 
                      inputs_21__11, inputs_21__10, inputs_21__9, inputs_21__8, 
                      inputs_21__7, inputs_21__6, inputs_21__5, inputs_21__4, 
                      inputs_21__3, inputs_21__2, inputs_21__1, inputs_21__0, 
                      inputs_22__15, inputs_22__14, inputs_22__13, inputs_22__12, 
                      inputs_22__11, inputs_22__10, inputs_22__9, inputs_22__8, 
                      inputs_22__7, inputs_22__6, inputs_22__5, inputs_22__4, 
                      inputs_22__3, inputs_22__2, inputs_22__1, inputs_22__0, 
                      inputs_23__15, inputs_23__14, inputs_23__13, inputs_23__12, 
                      inputs_23__11, inputs_23__10, inputs_23__9, inputs_23__8, 
                      inputs_23__7, inputs_23__6, inputs_23__5, inputs_23__4, 
                      inputs_23__3, inputs_23__2, inputs_23__1, inputs_23__0, 
                      inputs_24__15, inputs_24__14, inputs_24__13, inputs_24__12, 
                      inputs_24__11, inputs_24__10, inputs_24__9, inputs_24__8, 
                      inputs_24__7, inputs_24__6, inputs_24__5, inputs_24__4, 
                      inputs_24__3, inputs_24__2, inputs_24__1, inputs_24__0, 
                      filterType, finalSum ) ;

    input inputs_0__15 ;
    input inputs_0__14 ;
    input inputs_0__13 ;
    input inputs_0__12 ;
    input inputs_0__11 ;
    input inputs_0__10 ;
    input inputs_0__9 ;
    input inputs_0__8 ;
    input inputs_0__7 ;
    input inputs_0__6 ;
    input inputs_0__5 ;
    input inputs_0__4 ;
    input inputs_0__3 ;
    input inputs_0__2 ;
    input inputs_0__1 ;
    input inputs_0__0 ;
    input inputs_1__15 ;
    input inputs_1__14 ;
    input inputs_1__13 ;
    input inputs_1__12 ;
    input inputs_1__11 ;
    input inputs_1__10 ;
    input inputs_1__9 ;
    input inputs_1__8 ;
    input inputs_1__7 ;
    input inputs_1__6 ;
    input inputs_1__5 ;
    input inputs_1__4 ;
    input inputs_1__3 ;
    input inputs_1__2 ;
    input inputs_1__1 ;
    input inputs_1__0 ;
    input inputs_2__15 ;
    input inputs_2__14 ;
    input inputs_2__13 ;
    input inputs_2__12 ;
    input inputs_2__11 ;
    input inputs_2__10 ;
    input inputs_2__9 ;
    input inputs_2__8 ;
    input inputs_2__7 ;
    input inputs_2__6 ;
    input inputs_2__5 ;
    input inputs_2__4 ;
    input inputs_2__3 ;
    input inputs_2__2 ;
    input inputs_2__1 ;
    input inputs_2__0 ;
    input inputs_3__15 ;
    input inputs_3__14 ;
    input inputs_3__13 ;
    input inputs_3__12 ;
    input inputs_3__11 ;
    input inputs_3__10 ;
    input inputs_3__9 ;
    input inputs_3__8 ;
    input inputs_3__7 ;
    input inputs_3__6 ;
    input inputs_3__5 ;
    input inputs_3__4 ;
    input inputs_3__3 ;
    input inputs_3__2 ;
    input inputs_3__1 ;
    input inputs_3__0 ;
    input inputs_4__15 ;
    input inputs_4__14 ;
    input inputs_4__13 ;
    input inputs_4__12 ;
    input inputs_4__11 ;
    input inputs_4__10 ;
    input inputs_4__9 ;
    input inputs_4__8 ;
    input inputs_4__7 ;
    input inputs_4__6 ;
    input inputs_4__5 ;
    input inputs_4__4 ;
    input inputs_4__3 ;
    input inputs_4__2 ;
    input inputs_4__1 ;
    input inputs_4__0 ;
    input inputs_5__15 ;
    input inputs_5__14 ;
    input inputs_5__13 ;
    input inputs_5__12 ;
    input inputs_5__11 ;
    input inputs_5__10 ;
    input inputs_5__9 ;
    input inputs_5__8 ;
    input inputs_5__7 ;
    input inputs_5__6 ;
    input inputs_5__5 ;
    input inputs_5__4 ;
    input inputs_5__3 ;
    input inputs_5__2 ;
    input inputs_5__1 ;
    input inputs_5__0 ;
    input inputs_6__15 ;
    input inputs_6__14 ;
    input inputs_6__13 ;
    input inputs_6__12 ;
    input inputs_6__11 ;
    input inputs_6__10 ;
    input inputs_6__9 ;
    input inputs_6__8 ;
    input inputs_6__7 ;
    input inputs_6__6 ;
    input inputs_6__5 ;
    input inputs_6__4 ;
    input inputs_6__3 ;
    input inputs_6__2 ;
    input inputs_6__1 ;
    input inputs_6__0 ;
    input inputs_7__15 ;
    input inputs_7__14 ;
    input inputs_7__13 ;
    input inputs_7__12 ;
    input inputs_7__11 ;
    input inputs_7__10 ;
    input inputs_7__9 ;
    input inputs_7__8 ;
    input inputs_7__7 ;
    input inputs_7__6 ;
    input inputs_7__5 ;
    input inputs_7__4 ;
    input inputs_7__3 ;
    input inputs_7__2 ;
    input inputs_7__1 ;
    input inputs_7__0 ;
    input inputs_8__15 ;
    input inputs_8__14 ;
    input inputs_8__13 ;
    input inputs_8__12 ;
    input inputs_8__11 ;
    input inputs_8__10 ;
    input inputs_8__9 ;
    input inputs_8__8 ;
    input inputs_8__7 ;
    input inputs_8__6 ;
    input inputs_8__5 ;
    input inputs_8__4 ;
    input inputs_8__3 ;
    input inputs_8__2 ;
    input inputs_8__1 ;
    input inputs_8__0 ;
    input inputs_9__15 ;
    input inputs_9__14 ;
    input inputs_9__13 ;
    input inputs_9__12 ;
    input inputs_9__11 ;
    input inputs_9__10 ;
    input inputs_9__9 ;
    input inputs_9__8 ;
    input inputs_9__7 ;
    input inputs_9__6 ;
    input inputs_9__5 ;
    input inputs_9__4 ;
    input inputs_9__3 ;
    input inputs_9__2 ;
    input inputs_9__1 ;
    input inputs_9__0 ;
    input inputs_10__15 ;
    input inputs_10__14 ;
    input inputs_10__13 ;
    input inputs_10__12 ;
    input inputs_10__11 ;
    input inputs_10__10 ;
    input inputs_10__9 ;
    input inputs_10__8 ;
    input inputs_10__7 ;
    input inputs_10__6 ;
    input inputs_10__5 ;
    input inputs_10__4 ;
    input inputs_10__3 ;
    input inputs_10__2 ;
    input inputs_10__1 ;
    input inputs_10__0 ;
    input inputs_11__15 ;
    input inputs_11__14 ;
    input inputs_11__13 ;
    input inputs_11__12 ;
    input inputs_11__11 ;
    input inputs_11__10 ;
    input inputs_11__9 ;
    input inputs_11__8 ;
    input inputs_11__7 ;
    input inputs_11__6 ;
    input inputs_11__5 ;
    input inputs_11__4 ;
    input inputs_11__3 ;
    input inputs_11__2 ;
    input inputs_11__1 ;
    input inputs_11__0 ;
    input inputs_12__15 ;
    input inputs_12__14 ;
    input inputs_12__13 ;
    input inputs_12__12 ;
    input inputs_12__11 ;
    input inputs_12__10 ;
    input inputs_12__9 ;
    input inputs_12__8 ;
    input inputs_12__7 ;
    input inputs_12__6 ;
    input inputs_12__5 ;
    input inputs_12__4 ;
    input inputs_12__3 ;
    input inputs_12__2 ;
    input inputs_12__1 ;
    input inputs_12__0 ;
    input inputs_13__15 ;
    input inputs_13__14 ;
    input inputs_13__13 ;
    input inputs_13__12 ;
    input inputs_13__11 ;
    input inputs_13__10 ;
    input inputs_13__9 ;
    input inputs_13__8 ;
    input inputs_13__7 ;
    input inputs_13__6 ;
    input inputs_13__5 ;
    input inputs_13__4 ;
    input inputs_13__3 ;
    input inputs_13__2 ;
    input inputs_13__1 ;
    input inputs_13__0 ;
    input inputs_14__15 ;
    input inputs_14__14 ;
    input inputs_14__13 ;
    input inputs_14__12 ;
    input inputs_14__11 ;
    input inputs_14__10 ;
    input inputs_14__9 ;
    input inputs_14__8 ;
    input inputs_14__7 ;
    input inputs_14__6 ;
    input inputs_14__5 ;
    input inputs_14__4 ;
    input inputs_14__3 ;
    input inputs_14__2 ;
    input inputs_14__1 ;
    input inputs_14__0 ;
    input inputs_15__15 ;
    input inputs_15__14 ;
    input inputs_15__13 ;
    input inputs_15__12 ;
    input inputs_15__11 ;
    input inputs_15__10 ;
    input inputs_15__9 ;
    input inputs_15__8 ;
    input inputs_15__7 ;
    input inputs_15__6 ;
    input inputs_15__5 ;
    input inputs_15__4 ;
    input inputs_15__3 ;
    input inputs_15__2 ;
    input inputs_15__1 ;
    input inputs_15__0 ;
    input inputs_16__15 ;
    input inputs_16__14 ;
    input inputs_16__13 ;
    input inputs_16__12 ;
    input inputs_16__11 ;
    input inputs_16__10 ;
    input inputs_16__9 ;
    input inputs_16__8 ;
    input inputs_16__7 ;
    input inputs_16__6 ;
    input inputs_16__5 ;
    input inputs_16__4 ;
    input inputs_16__3 ;
    input inputs_16__2 ;
    input inputs_16__1 ;
    input inputs_16__0 ;
    input inputs_17__15 ;
    input inputs_17__14 ;
    input inputs_17__13 ;
    input inputs_17__12 ;
    input inputs_17__11 ;
    input inputs_17__10 ;
    input inputs_17__9 ;
    input inputs_17__8 ;
    input inputs_17__7 ;
    input inputs_17__6 ;
    input inputs_17__5 ;
    input inputs_17__4 ;
    input inputs_17__3 ;
    input inputs_17__2 ;
    input inputs_17__1 ;
    input inputs_17__0 ;
    input inputs_18__15 ;
    input inputs_18__14 ;
    input inputs_18__13 ;
    input inputs_18__12 ;
    input inputs_18__11 ;
    input inputs_18__10 ;
    input inputs_18__9 ;
    input inputs_18__8 ;
    input inputs_18__7 ;
    input inputs_18__6 ;
    input inputs_18__5 ;
    input inputs_18__4 ;
    input inputs_18__3 ;
    input inputs_18__2 ;
    input inputs_18__1 ;
    input inputs_18__0 ;
    input inputs_19__15 ;
    input inputs_19__14 ;
    input inputs_19__13 ;
    input inputs_19__12 ;
    input inputs_19__11 ;
    input inputs_19__10 ;
    input inputs_19__9 ;
    input inputs_19__8 ;
    input inputs_19__7 ;
    input inputs_19__6 ;
    input inputs_19__5 ;
    input inputs_19__4 ;
    input inputs_19__3 ;
    input inputs_19__2 ;
    input inputs_19__1 ;
    input inputs_19__0 ;
    input inputs_20__15 ;
    input inputs_20__14 ;
    input inputs_20__13 ;
    input inputs_20__12 ;
    input inputs_20__11 ;
    input inputs_20__10 ;
    input inputs_20__9 ;
    input inputs_20__8 ;
    input inputs_20__7 ;
    input inputs_20__6 ;
    input inputs_20__5 ;
    input inputs_20__4 ;
    input inputs_20__3 ;
    input inputs_20__2 ;
    input inputs_20__1 ;
    input inputs_20__0 ;
    input inputs_21__15 ;
    input inputs_21__14 ;
    input inputs_21__13 ;
    input inputs_21__12 ;
    input inputs_21__11 ;
    input inputs_21__10 ;
    input inputs_21__9 ;
    input inputs_21__8 ;
    input inputs_21__7 ;
    input inputs_21__6 ;
    input inputs_21__5 ;
    input inputs_21__4 ;
    input inputs_21__3 ;
    input inputs_21__2 ;
    input inputs_21__1 ;
    input inputs_21__0 ;
    input inputs_22__15 ;
    input inputs_22__14 ;
    input inputs_22__13 ;
    input inputs_22__12 ;
    input inputs_22__11 ;
    input inputs_22__10 ;
    input inputs_22__9 ;
    input inputs_22__8 ;
    input inputs_22__7 ;
    input inputs_22__6 ;
    input inputs_22__5 ;
    input inputs_22__4 ;
    input inputs_22__3 ;
    input inputs_22__2 ;
    input inputs_22__1 ;
    input inputs_22__0 ;
    input inputs_23__15 ;
    input inputs_23__14 ;
    input inputs_23__13 ;
    input inputs_23__12 ;
    input inputs_23__11 ;
    input inputs_23__10 ;
    input inputs_23__9 ;
    input inputs_23__8 ;
    input inputs_23__7 ;
    input inputs_23__6 ;
    input inputs_23__5 ;
    input inputs_23__4 ;
    input inputs_23__3 ;
    input inputs_23__2 ;
    input inputs_23__1 ;
    input inputs_23__0 ;
    input inputs_24__15 ;
    input inputs_24__14 ;
    input inputs_24__13 ;
    input inputs_24__12 ;
    input inputs_24__11 ;
    input inputs_24__10 ;
    input inputs_24__9 ;
    input inputs_24__8 ;
    input inputs_24__7 ;
    input inputs_24__6 ;
    input inputs_24__5 ;
    input inputs_24__4 ;
    input inputs_24__3 ;
    input inputs_24__2 ;
    input inputs_24__1 ;
    input inputs_24__0 ;
    input filterType ;
    output [15:0]finalSum ;

    wire sum1_15, sum1_14, sum1_13, sum1_12, sum1_11, sum1_10, sum1_9, sum1_8, 
         sum1_7, sum1_6, sum1_5, sum1_4, sum1_3, sum1_2, sum1_1, sum1_0, sum2_15, 
         sum2_14, sum2_13, sum2_12, sum2_11, sum2_10, sum2_9, sum2_8, sum2_7, 
         sum2_6, sum2_5, sum2_4, sum2_3, sum2_2, sum2_1, sum2_0, sum3_15, 
         sum3_14, sum3_13, sum3_12, sum3_11, sum3_10, sum3_9, sum3_8, sum3_7, 
         sum3_6, sum3_5, sum3_4, sum3_3, sum3_2, sum3_1, sum3_0, sum3Filter_15, 
         sum3Filter_14, sum3Filter_13, sum3Filter_12, sum3Filter_11, 
         sum3Filter_10, sum3Filter_9, sum3Filter_8, sum3Filter_7, sum3Filter_6, 
         sum3Filter_5, sum3Filter_4, sum3Filter_3, sum3Filter_2, sum3Filter_1, 
         sum3Filter_0, sum4_15, sum4_14, sum4_13, sum4_12, sum4_11, sum4_10, 
         sum4_9, sum4_8, sum4_7, sum4_6, sum4_5, sum4_4, sum4_3, sum4_2, sum4_1, 
         sum4_0, totalSum_15, totalSum_14, totalSum_13, totalSum_12, totalSum_11, 
         totalSum_10, totalSum_9, totalSum_8, totalSum_7, totalSum_6, totalSum_5, 
         totalSum_4, totalSum_3, totalSum_2, totalSum_1, totalSum_0, GND;
    wire [2:0] \$dummy ;




    Adder8Values_16 sum1Map (.inputs_0__15 (inputs_0__15), .inputs_0__14 (
                    inputs_0__14), .inputs_0__13 (inputs_0__13), .inputs_0__12 (
                    inputs_0__12), .inputs_0__11 (inputs_0__11), .inputs_0__10 (
                    inputs_0__10), .inputs_0__9 (inputs_0__9), .inputs_0__8 (
                    inputs_0__8), .inputs_0__7 (inputs_0__7), .inputs_0__6 (
                    inputs_0__6), .inputs_0__5 (inputs_0__5), .inputs_0__4 (
                    inputs_0__4), .inputs_0__3 (inputs_0__3), .inputs_0__2 (
                    inputs_0__2), .inputs_0__1 (inputs_0__1), .inputs_0__0 (
                    inputs_0__0), .inputs_1__15 (inputs_1__15), .inputs_1__14 (
                    inputs_1__14), .inputs_1__13 (inputs_1__13), .inputs_1__12 (
                    inputs_1__12), .inputs_1__11 (inputs_1__11), .inputs_1__10 (
                    inputs_1__10), .inputs_1__9 (inputs_1__9), .inputs_1__8 (
                    inputs_1__8), .inputs_1__7 (inputs_1__7), .inputs_1__6 (
                    inputs_1__6), .inputs_1__5 (inputs_1__5), .inputs_1__4 (
                    inputs_1__4), .inputs_1__3 (inputs_1__3), .inputs_1__2 (
                    inputs_1__2), .inputs_1__1 (inputs_1__1), .inputs_1__0 (
                    inputs_1__0), .inputs_2__15 (inputs_2__15), .inputs_2__14 (
                    inputs_2__14), .inputs_2__13 (inputs_2__13), .inputs_2__12 (
                    inputs_2__12), .inputs_2__11 (inputs_2__11), .inputs_2__10 (
                    inputs_2__10), .inputs_2__9 (inputs_2__9), .inputs_2__8 (
                    inputs_2__8), .inputs_2__7 (inputs_2__7), .inputs_2__6 (
                    inputs_2__6), .inputs_2__5 (inputs_2__5), .inputs_2__4 (
                    inputs_2__4), .inputs_2__3 (inputs_2__3), .inputs_2__2 (
                    inputs_2__2), .inputs_2__1 (inputs_2__1), .inputs_2__0 (
                    inputs_2__0), .inputs_3__15 (inputs_3__15), .inputs_3__14 (
                    inputs_3__14), .inputs_3__13 (inputs_3__13), .inputs_3__12 (
                    inputs_3__12), .inputs_3__11 (inputs_3__11), .inputs_3__10 (
                    inputs_3__10), .inputs_3__9 (inputs_3__9), .inputs_3__8 (
                    inputs_3__8), .inputs_3__7 (inputs_3__7), .inputs_3__6 (
                    inputs_3__6), .inputs_3__5 (inputs_3__5), .inputs_3__4 (
                    inputs_3__4), .inputs_3__3 (inputs_3__3), .inputs_3__2 (
                    inputs_3__2), .inputs_3__1 (inputs_3__1), .inputs_3__0 (
                    inputs_3__0), .inputs_4__15 (inputs_4__15), .inputs_4__14 (
                    inputs_4__14), .inputs_4__13 (inputs_4__13), .inputs_4__12 (
                    inputs_4__12), .inputs_4__11 (inputs_4__11), .inputs_4__10 (
                    inputs_4__10), .inputs_4__9 (inputs_4__9), .inputs_4__8 (
                    inputs_4__8), .inputs_4__7 (inputs_4__7), .inputs_4__6 (
                    inputs_4__6), .inputs_4__5 (inputs_4__5), .inputs_4__4 (
                    inputs_4__4), .inputs_4__3 (inputs_4__3), .inputs_4__2 (
                    inputs_4__2), .inputs_4__1 (inputs_4__1), .inputs_4__0 (
                    inputs_4__0), .inputs_5__15 (inputs_5__15), .inputs_5__14 (
                    inputs_5__14), .inputs_5__13 (inputs_5__13), .inputs_5__12 (
                    inputs_5__12), .inputs_5__11 (inputs_5__11), .inputs_5__10 (
                    inputs_5__10), .inputs_5__9 (inputs_5__9), .inputs_5__8 (
                    inputs_5__8), .inputs_5__7 (inputs_5__7), .inputs_5__6 (
                    inputs_5__6), .inputs_5__5 (inputs_5__5), .inputs_5__4 (
                    inputs_5__4), .inputs_5__3 (inputs_5__3), .inputs_5__2 (
                    inputs_5__2), .inputs_5__1 (inputs_5__1), .inputs_5__0 (
                    inputs_5__0), .inputs_6__15 (inputs_6__15), .inputs_6__14 (
                    inputs_6__14), .inputs_6__13 (inputs_6__13), .inputs_6__12 (
                    inputs_6__12), .inputs_6__11 (inputs_6__11), .inputs_6__10 (
                    inputs_6__10), .inputs_6__9 (inputs_6__9), .inputs_6__8 (
                    inputs_6__8), .inputs_6__7 (inputs_6__7), .inputs_6__6 (
                    inputs_6__6), .inputs_6__5 (inputs_6__5), .inputs_6__4 (
                    inputs_6__4), .inputs_6__3 (inputs_6__3), .inputs_6__2 (
                    inputs_6__2), .inputs_6__1 (inputs_6__1), .inputs_6__0 (
                    inputs_6__0), .inputs_7__15 (inputs_7__15), .inputs_7__14 (
                    inputs_7__14), .inputs_7__13 (inputs_7__13), .inputs_7__12 (
                    inputs_7__12), .inputs_7__11 (inputs_7__11), .inputs_7__10 (
                    inputs_7__10), .inputs_7__9 (inputs_7__9), .inputs_7__8 (
                    inputs_7__8), .inputs_7__7 (inputs_7__7), .inputs_7__6 (
                    inputs_7__6), .inputs_7__5 (inputs_7__5), .inputs_7__4 (
                    inputs_7__4), .inputs_7__3 (inputs_7__3), .inputs_7__2 (
                    inputs_7__2), .inputs_7__1 (inputs_7__1), .inputs_7__0 (
                    inputs_7__0), .sum ({sum1_15,sum1_14,sum1_13,sum1_12,sum1_11
                    ,sum1_10,sum1_9,sum1_8,sum1_7,sum1_6,sum1_5,sum1_4,sum1_3,
                    sum1_2,sum1_1,sum1_0})) ;
    Adder8Values_16 sum2Map (.inputs_0__15 (inputs_9__15), .inputs_0__14 (
                    inputs_9__14), .inputs_0__13 (inputs_9__13), .inputs_0__12 (
                    inputs_9__12), .inputs_0__11 (inputs_9__11), .inputs_0__10 (
                    inputs_9__10), .inputs_0__9 (inputs_9__9), .inputs_0__8 (
                    inputs_9__8), .inputs_0__7 (inputs_9__7), .inputs_0__6 (
                    inputs_9__6), .inputs_0__5 (inputs_9__5), .inputs_0__4 (
                    inputs_9__4), .inputs_0__3 (inputs_9__3), .inputs_0__2 (
                    inputs_9__2), .inputs_0__1 (inputs_9__1), .inputs_0__0 (
                    inputs_9__0), .inputs_1__15 (inputs_10__15), .inputs_1__14 (
                    inputs_10__14), .inputs_1__13 (inputs_10__13), .inputs_1__12 (
                    inputs_10__12), .inputs_1__11 (inputs_10__11), .inputs_1__10 (
                    inputs_10__10), .inputs_1__9 (inputs_10__9), .inputs_1__8 (
                    inputs_10__8), .inputs_1__7 (inputs_10__7), .inputs_1__6 (
                    inputs_10__6), .inputs_1__5 (inputs_10__5), .inputs_1__4 (
                    inputs_10__4), .inputs_1__3 (inputs_10__3), .inputs_1__2 (
                    inputs_10__2), .inputs_1__1 (inputs_10__1), .inputs_1__0 (
                    inputs_10__0), .inputs_2__15 (inputs_11__15), .inputs_2__14 (
                    inputs_11__14), .inputs_2__13 (inputs_11__13), .inputs_2__12 (
                    inputs_11__12), .inputs_2__11 (inputs_11__11), .inputs_2__10 (
                    inputs_11__10), .inputs_2__9 (inputs_11__9), .inputs_2__8 (
                    inputs_11__8), .inputs_2__7 (inputs_11__7), .inputs_2__6 (
                    inputs_11__6), .inputs_2__5 (inputs_11__5), .inputs_2__4 (
                    inputs_11__4), .inputs_2__3 (inputs_11__3), .inputs_2__2 (
                    inputs_11__2), .inputs_2__1 (inputs_11__1), .inputs_2__0 (
                    inputs_11__0), .inputs_3__15 (inputs_12__15), .inputs_3__14 (
                    inputs_12__14), .inputs_3__13 (inputs_12__13), .inputs_3__12 (
                    inputs_12__12), .inputs_3__11 (inputs_12__11), .inputs_3__10 (
                    inputs_12__10), .inputs_3__9 (inputs_12__9), .inputs_3__8 (
                    inputs_12__8), .inputs_3__7 (inputs_12__7), .inputs_3__6 (
                    inputs_12__6), .inputs_3__5 (inputs_12__5), .inputs_3__4 (
                    inputs_12__4), .inputs_3__3 (inputs_12__3), .inputs_3__2 (
                    inputs_12__2), .inputs_3__1 (inputs_12__1), .inputs_3__0 (
                    inputs_12__0), .inputs_4__15 (inputs_13__15), .inputs_4__14 (
                    inputs_13__14), .inputs_4__13 (inputs_13__13), .inputs_4__12 (
                    inputs_13__12), .inputs_4__11 (inputs_13__11), .inputs_4__10 (
                    inputs_13__10), .inputs_4__9 (inputs_13__9), .inputs_4__8 (
                    inputs_13__8), .inputs_4__7 (inputs_13__7), .inputs_4__6 (
                    inputs_13__6), .inputs_4__5 (inputs_13__5), .inputs_4__4 (
                    inputs_13__4), .inputs_4__3 (inputs_13__3), .inputs_4__2 (
                    inputs_13__2), .inputs_4__1 (inputs_13__1), .inputs_4__0 (
                    inputs_13__0), .inputs_5__15 (inputs_14__15), .inputs_5__14 (
                    inputs_14__14), .inputs_5__13 (inputs_14__13), .inputs_5__12 (
                    inputs_14__12), .inputs_5__11 (inputs_14__11), .inputs_5__10 (
                    inputs_14__10), .inputs_5__9 (inputs_14__9), .inputs_5__8 (
                    inputs_14__8), .inputs_5__7 (inputs_14__7), .inputs_5__6 (
                    inputs_14__6), .inputs_5__5 (inputs_14__5), .inputs_5__4 (
                    inputs_14__4), .inputs_5__3 (inputs_14__3), .inputs_5__2 (
                    inputs_14__2), .inputs_5__1 (inputs_14__1), .inputs_5__0 (
                    inputs_14__0), .inputs_6__15 (inputs_15__15), .inputs_6__14 (
                    inputs_15__14), .inputs_6__13 (inputs_15__13), .inputs_6__12 (
                    inputs_15__12), .inputs_6__11 (inputs_15__11), .inputs_6__10 (
                    inputs_15__10), .inputs_6__9 (inputs_15__9), .inputs_6__8 (
                    inputs_15__8), .inputs_6__7 (inputs_15__7), .inputs_6__6 (
                    inputs_15__6), .inputs_6__5 (inputs_15__5), .inputs_6__4 (
                    inputs_15__4), .inputs_6__3 (inputs_15__3), .inputs_6__2 (
                    inputs_15__2), .inputs_6__1 (inputs_15__1), .inputs_6__0 (
                    inputs_15__0), .inputs_7__15 (inputs_16__15), .inputs_7__14 (
                    inputs_16__14), .inputs_7__13 (inputs_16__13), .inputs_7__12 (
                    inputs_16__12), .inputs_7__11 (inputs_16__11), .inputs_7__10 (
                    inputs_16__10), .inputs_7__9 (inputs_16__9), .inputs_7__8 (
                    inputs_16__8), .inputs_7__7 (inputs_16__7), .inputs_7__6 (
                    inputs_16__6), .inputs_7__5 (inputs_16__5), .inputs_7__4 (
                    inputs_16__4), .inputs_7__3 (inputs_16__3), .inputs_7__2 (
                    inputs_16__2), .inputs_7__1 (inputs_16__1), .inputs_7__0 (
                    inputs_16__0), .sum ({sum2_15,sum2_14,sum2_13,sum2_12,
                    sum2_11,sum2_10,sum2_9,sum2_8,sum2_7,sum2_6,sum2_5,sum2_4,
                    sum2_3,sum2_2,sum2_1,sum2_0})) ;
    Adder8Values_16 sum3Map (.inputs_0__15 (inputs_17__15), .inputs_0__14 (
                    inputs_17__14), .inputs_0__13 (inputs_17__13), .inputs_0__12 (
                    inputs_17__12), .inputs_0__11 (inputs_17__11), .inputs_0__10 (
                    inputs_17__10), .inputs_0__9 (inputs_17__9), .inputs_0__8 (
                    inputs_17__8), .inputs_0__7 (inputs_17__7), .inputs_0__6 (
                    inputs_17__6), .inputs_0__5 (inputs_17__5), .inputs_0__4 (
                    inputs_17__4), .inputs_0__3 (inputs_17__3), .inputs_0__2 (
                    inputs_17__2), .inputs_0__1 (inputs_17__1), .inputs_0__0 (
                    inputs_17__0), .inputs_1__15 (inputs_18__15), .inputs_1__14 (
                    inputs_18__14), .inputs_1__13 (inputs_18__13), .inputs_1__12 (
                    inputs_18__12), .inputs_1__11 (inputs_18__11), .inputs_1__10 (
                    inputs_18__10), .inputs_1__9 (inputs_18__9), .inputs_1__8 (
                    inputs_18__8), .inputs_1__7 (inputs_18__7), .inputs_1__6 (
                    inputs_18__6), .inputs_1__5 (inputs_18__5), .inputs_1__4 (
                    inputs_18__4), .inputs_1__3 (inputs_18__3), .inputs_1__2 (
                    inputs_18__2), .inputs_1__1 (inputs_18__1), .inputs_1__0 (
                    inputs_18__0), .inputs_2__15 (inputs_19__15), .inputs_2__14 (
                    inputs_19__14), .inputs_2__13 (inputs_19__13), .inputs_2__12 (
                    inputs_19__12), .inputs_2__11 (inputs_19__11), .inputs_2__10 (
                    inputs_19__10), .inputs_2__9 (inputs_19__9), .inputs_2__8 (
                    inputs_19__8), .inputs_2__7 (inputs_19__7), .inputs_2__6 (
                    inputs_19__6), .inputs_2__5 (inputs_19__5), .inputs_2__4 (
                    inputs_19__4), .inputs_2__3 (inputs_19__3), .inputs_2__2 (
                    inputs_19__2), .inputs_2__1 (inputs_19__1), .inputs_2__0 (
                    inputs_19__0), .inputs_3__15 (inputs_20__15), .inputs_3__14 (
                    inputs_20__14), .inputs_3__13 (inputs_20__13), .inputs_3__12 (
                    inputs_20__12), .inputs_3__11 (inputs_20__11), .inputs_3__10 (
                    inputs_20__10), .inputs_3__9 (inputs_20__9), .inputs_3__8 (
                    inputs_20__8), .inputs_3__7 (inputs_20__7), .inputs_3__6 (
                    inputs_20__6), .inputs_3__5 (inputs_20__5), .inputs_3__4 (
                    inputs_20__4), .inputs_3__3 (inputs_20__3), .inputs_3__2 (
                    inputs_20__2), .inputs_3__1 (inputs_20__1), .inputs_3__0 (
                    inputs_20__0), .inputs_4__15 (inputs_21__15), .inputs_4__14 (
                    inputs_21__14), .inputs_4__13 (inputs_21__13), .inputs_4__12 (
                    inputs_21__12), .inputs_4__11 (inputs_21__11), .inputs_4__10 (
                    inputs_21__10), .inputs_4__9 (inputs_21__9), .inputs_4__8 (
                    inputs_21__8), .inputs_4__7 (inputs_21__7), .inputs_4__6 (
                    inputs_21__6), .inputs_4__5 (inputs_21__5), .inputs_4__4 (
                    inputs_21__4), .inputs_4__3 (inputs_21__3), .inputs_4__2 (
                    inputs_21__2), .inputs_4__1 (inputs_21__1), .inputs_4__0 (
                    inputs_21__0), .inputs_5__15 (inputs_22__15), .inputs_5__14 (
                    inputs_22__14), .inputs_5__13 (inputs_22__13), .inputs_5__12 (
                    inputs_22__12), .inputs_5__11 (inputs_22__11), .inputs_5__10 (
                    inputs_22__10), .inputs_5__9 (inputs_22__9), .inputs_5__8 (
                    inputs_22__8), .inputs_5__7 (inputs_22__7), .inputs_5__6 (
                    inputs_22__6), .inputs_5__5 (inputs_22__5), .inputs_5__4 (
                    inputs_22__4), .inputs_5__3 (inputs_22__3), .inputs_5__2 (
                    inputs_22__2), .inputs_5__1 (inputs_22__1), .inputs_5__0 (
                    inputs_22__0), .inputs_6__15 (inputs_23__15), .inputs_6__14 (
                    inputs_23__14), .inputs_6__13 (inputs_23__13), .inputs_6__12 (
                    inputs_23__12), .inputs_6__11 (inputs_23__11), .inputs_6__10 (
                    inputs_23__10), .inputs_6__9 (inputs_23__9), .inputs_6__8 (
                    inputs_23__8), .inputs_6__7 (inputs_23__7), .inputs_6__6 (
                    inputs_23__6), .inputs_6__5 (inputs_23__5), .inputs_6__4 (
                    inputs_23__4), .inputs_6__3 (inputs_23__3), .inputs_6__2 (
                    inputs_23__2), .inputs_6__1 (inputs_23__1), .inputs_6__0 (
                    inputs_23__0), .inputs_7__15 (inputs_24__15), .inputs_7__14 (
                    inputs_24__14), .inputs_7__13 (inputs_24__13), .inputs_7__12 (
                    inputs_24__12), .inputs_7__11 (inputs_24__11), .inputs_7__10 (
                    inputs_24__10), .inputs_7__9 (inputs_24__9), .inputs_7__8 (
                    inputs_24__8), .inputs_7__7 (inputs_24__7), .inputs_7__6 (
                    inputs_24__6), .inputs_7__5 (inputs_24__5), .inputs_7__4 (
                    inputs_24__4), .inputs_7__3 (inputs_24__3), .inputs_7__2 (
                    inputs_24__2), .inputs_7__1 (inputs_24__1), .inputs_7__0 (
                    inputs_24__0), .sum ({sum3_15,sum3_14,sum3_13,sum3_12,
                    sum3_11,sum3_10,sum3_9,sum3_8,sum3_7,sum3_6,sum3_5,sum3_4,
                    sum3_3,sum3_2,sum3_1,sum3_0})) ;
    NBitAdder_16 sum3FilterMap (.a ({sum1_15,sum1_14,sum1_13,sum1_12,sum1_11,
                 sum1_10,sum1_9,sum1_8,sum1_7,sum1_6,sum1_5,sum1_4,sum1_3,sum1_2
                 ,sum1_1,sum1_0}), .b ({inputs_8__15,inputs_8__14,inputs_8__13,
                 inputs_8__12,inputs_8__11,inputs_8__10,inputs_8__9,inputs_8__8,
                 inputs_8__7,inputs_8__6,inputs_8__5,inputs_8__4,inputs_8__3,
                 inputs_8__2,inputs_8__1,inputs_8__0}), .carryIn (GND), .sum ({
                 sum3Filter_15,sum3Filter_14,sum3Filter_13,sum3Filter_12,
                 sum3Filter_11,sum3Filter_10,sum3Filter_9,sum3Filter_8,
                 sum3Filter_7,sum3Filter_6,sum3Filter_5,sum3Filter_4,
                 sum3Filter_3,sum3Filter_2,sum3Filter_1,sum3Filter_0}), .carryOut (
                 \$dummy [0])) ;
    NBitAdder_16 sumRestMap (.a ({sum2_15,sum2_14,sum2_13,sum2_12,sum2_11,
                 sum2_10,sum2_9,sum2_8,sum2_7,sum2_6,sum2_5,sum2_4,sum2_3,sum2_2
                 ,sum2_1,sum2_0}), .b ({sum3_15,sum3_14,sum3_13,sum3_12,sum3_11,
                 sum3_10,sum3_9,sum3_8,sum3_7,sum3_6,sum3_5,sum3_4,sum3_3,sum3_2
                 ,sum3_1,sum3_0}), .carryIn (GND), .sum ({sum4_15,sum4_14,
                 sum4_13,sum4_12,sum4_11,sum4_10,sum4_9,sum4_8,sum4_7,sum4_6,
                 sum4_5,sum4_4,sum4_3,sum4_2,sum4_1,sum4_0}), .carryOut (
                 \$dummy [1])) ;
    NBitAdder_16 sumFinalMap (.a ({sum3Filter_15,sum3Filter_14,sum3Filter_13,
                 sum3Filter_12,sum3Filter_11,sum3Filter_10,sum3Filter_9,
                 sum3Filter_8,sum3Filter_7,sum3Filter_6,sum3Filter_5,
                 sum3Filter_4,sum3Filter_3,sum3Filter_2,sum3Filter_1,
                 sum3Filter_0}), .b ({sum4_15,sum4_14,sum4_13,sum4_12,sum4_11,
                 sum4_10,sum4_9,sum4_8,sum4_7,sum4_6,sum4_5,sum4_4,sum4_3,sum4_2
                 ,sum4_1,sum4_0}), .carryIn (GND), .sum ({totalSum_15,
                 totalSum_14,totalSum_13,totalSum_12,totalSum_11,totalSum_10,
                 totalSum_9,totalSum_8,totalSum_7,totalSum_6,totalSum_5,
                 totalSum_4,totalSum_3,totalSum_2,totalSum_1,totalSum_0}), .carryOut (
                 \$dummy [2])) ;
    Mux2_16 finalSumMap (.A ({sum3Filter_15,sum3Filter_14,sum3Filter_13,
            sum3Filter_12,sum3Filter_11,sum3Filter_10,sum3Filter_9,sum3Filter_8,
            sum3Filter_7,sum3Filter_6,sum3Filter_5,sum3Filter_4,sum3Filter_3,
            sum3Filter_2,sum3Filter_1,sum3Filter_0}), .B ({totalSum_15,
            totalSum_14,totalSum_13,totalSum_12,totalSum_11,totalSum_10,
            totalSum_9,totalSum_8,totalSum_7,totalSum_6,totalSum_5,totalSum_4,
            totalSum_3,totalSum_2,totalSum_1,totalSum_0}), .S (filterType), .C (
            {finalSum[15],finalSum[14],finalSum[13],finalSum[12],finalSum[11],
            finalSum[10],finalSum[9],finalSum[8],finalSum[7],finalSum[6],
            finalSum[5],finalSum[4],finalSum[3],finalSum[2],finalSum[1],
            finalSum[0]})) ;
    fake_gnd ix221 (.Y (GND)) ;
endmodule


module Adder8Values_16 ( inputs_0__15, inputs_0__14, inputs_0__13, inputs_0__12, 
                         inputs_0__11, inputs_0__10, inputs_0__9, inputs_0__8, 
                         inputs_0__7, inputs_0__6, inputs_0__5, inputs_0__4, 
                         inputs_0__3, inputs_0__2, inputs_0__1, inputs_0__0, 
                         inputs_1__15, inputs_1__14, inputs_1__13, inputs_1__12, 
                         inputs_1__11, inputs_1__10, inputs_1__9, inputs_1__8, 
                         inputs_1__7, inputs_1__6, inputs_1__5, inputs_1__4, 
                         inputs_1__3, inputs_1__2, inputs_1__1, inputs_1__0, 
                         inputs_2__15, inputs_2__14, inputs_2__13, inputs_2__12, 
                         inputs_2__11, inputs_2__10, inputs_2__9, inputs_2__8, 
                         inputs_2__7, inputs_2__6, inputs_2__5, inputs_2__4, 
                         inputs_2__3, inputs_2__2, inputs_2__1, inputs_2__0, 
                         inputs_3__15, inputs_3__14, inputs_3__13, inputs_3__12, 
                         inputs_3__11, inputs_3__10, inputs_3__9, inputs_3__8, 
                         inputs_3__7, inputs_3__6, inputs_3__5, inputs_3__4, 
                         inputs_3__3, inputs_3__2, inputs_3__1, inputs_3__0, 
                         inputs_4__15, inputs_4__14, inputs_4__13, inputs_4__12, 
                         inputs_4__11, inputs_4__10, inputs_4__9, inputs_4__8, 
                         inputs_4__7, inputs_4__6, inputs_4__5, inputs_4__4, 
                         inputs_4__3, inputs_4__2, inputs_4__1, inputs_4__0, 
                         inputs_5__15, inputs_5__14, inputs_5__13, inputs_5__12, 
                         inputs_5__11, inputs_5__10, inputs_5__9, inputs_5__8, 
                         inputs_5__7, inputs_5__6, inputs_5__5, inputs_5__4, 
                         inputs_5__3, inputs_5__2, inputs_5__1, inputs_5__0, 
                         inputs_6__15, inputs_6__14, inputs_6__13, inputs_6__12, 
                         inputs_6__11, inputs_6__10, inputs_6__9, inputs_6__8, 
                         inputs_6__7, inputs_6__6, inputs_6__5, inputs_6__4, 
                         inputs_6__3, inputs_6__2, inputs_6__1, inputs_6__0, 
                         inputs_7__15, inputs_7__14, inputs_7__13, inputs_7__12, 
                         inputs_7__11, inputs_7__10, inputs_7__9, inputs_7__8, 
                         inputs_7__7, inputs_7__6, inputs_7__5, inputs_7__4, 
                         inputs_7__3, inputs_7__2, inputs_7__1, inputs_7__0, sum
                          ) ;

    input inputs_0__15 ;
    input inputs_0__14 ;
    input inputs_0__13 ;
    input inputs_0__12 ;
    input inputs_0__11 ;
    input inputs_0__10 ;
    input inputs_0__9 ;
    input inputs_0__8 ;
    input inputs_0__7 ;
    input inputs_0__6 ;
    input inputs_0__5 ;
    input inputs_0__4 ;
    input inputs_0__3 ;
    input inputs_0__2 ;
    input inputs_0__1 ;
    input inputs_0__0 ;
    input inputs_1__15 ;
    input inputs_1__14 ;
    input inputs_1__13 ;
    input inputs_1__12 ;
    input inputs_1__11 ;
    input inputs_1__10 ;
    input inputs_1__9 ;
    input inputs_1__8 ;
    input inputs_1__7 ;
    input inputs_1__6 ;
    input inputs_1__5 ;
    input inputs_1__4 ;
    input inputs_1__3 ;
    input inputs_1__2 ;
    input inputs_1__1 ;
    input inputs_1__0 ;
    input inputs_2__15 ;
    input inputs_2__14 ;
    input inputs_2__13 ;
    input inputs_2__12 ;
    input inputs_2__11 ;
    input inputs_2__10 ;
    input inputs_2__9 ;
    input inputs_2__8 ;
    input inputs_2__7 ;
    input inputs_2__6 ;
    input inputs_2__5 ;
    input inputs_2__4 ;
    input inputs_2__3 ;
    input inputs_2__2 ;
    input inputs_2__1 ;
    input inputs_2__0 ;
    input inputs_3__15 ;
    input inputs_3__14 ;
    input inputs_3__13 ;
    input inputs_3__12 ;
    input inputs_3__11 ;
    input inputs_3__10 ;
    input inputs_3__9 ;
    input inputs_3__8 ;
    input inputs_3__7 ;
    input inputs_3__6 ;
    input inputs_3__5 ;
    input inputs_3__4 ;
    input inputs_3__3 ;
    input inputs_3__2 ;
    input inputs_3__1 ;
    input inputs_3__0 ;
    input inputs_4__15 ;
    input inputs_4__14 ;
    input inputs_4__13 ;
    input inputs_4__12 ;
    input inputs_4__11 ;
    input inputs_4__10 ;
    input inputs_4__9 ;
    input inputs_4__8 ;
    input inputs_4__7 ;
    input inputs_4__6 ;
    input inputs_4__5 ;
    input inputs_4__4 ;
    input inputs_4__3 ;
    input inputs_4__2 ;
    input inputs_4__1 ;
    input inputs_4__0 ;
    input inputs_5__15 ;
    input inputs_5__14 ;
    input inputs_5__13 ;
    input inputs_5__12 ;
    input inputs_5__11 ;
    input inputs_5__10 ;
    input inputs_5__9 ;
    input inputs_5__8 ;
    input inputs_5__7 ;
    input inputs_5__6 ;
    input inputs_5__5 ;
    input inputs_5__4 ;
    input inputs_5__3 ;
    input inputs_5__2 ;
    input inputs_5__1 ;
    input inputs_5__0 ;
    input inputs_6__15 ;
    input inputs_6__14 ;
    input inputs_6__13 ;
    input inputs_6__12 ;
    input inputs_6__11 ;
    input inputs_6__10 ;
    input inputs_6__9 ;
    input inputs_6__8 ;
    input inputs_6__7 ;
    input inputs_6__6 ;
    input inputs_6__5 ;
    input inputs_6__4 ;
    input inputs_6__3 ;
    input inputs_6__2 ;
    input inputs_6__1 ;
    input inputs_6__0 ;
    input inputs_7__15 ;
    input inputs_7__14 ;
    input inputs_7__13 ;
    input inputs_7__12 ;
    input inputs_7__11 ;
    input inputs_7__10 ;
    input inputs_7__9 ;
    input inputs_7__8 ;
    input inputs_7__7 ;
    input inputs_7__6 ;
    input inputs_7__5 ;
    input inputs_7__4 ;
    input inputs_7__3 ;
    input inputs_7__2 ;
    input inputs_7__1 ;
    input inputs_7__0 ;
    output [15:0]sum ;

    wire sum1_15, sum1_14, sum1_13, sum1_12, sum1_11, sum1_10, sum1_9, sum1_8, 
         sum1_7, sum1_6, sum1_5, sum1_4, sum1_3, sum1_2, sum1_1, sum1_0, sum2_15, 
         sum2_14, sum2_13, sum2_12, sum2_11, sum2_10, sum2_9, sum2_8, sum2_7, 
         sum2_6, sum2_5, sum2_4, sum2_3, sum2_2, sum2_1, sum2_0, GND;
    wire [0:0] \$dummy ;




    Adder4Values_16 sum1Map (.a ({inputs_0__15,inputs_0__14,inputs_0__13,
                    inputs_0__12,inputs_0__11,inputs_0__10,inputs_0__9,
                    inputs_0__8,inputs_0__7,inputs_0__6,inputs_0__5,inputs_0__4,
                    inputs_0__3,inputs_0__2,inputs_0__1,inputs_0__0}), .b ({
                    inputs_1__15,inputs_1__14,inputs_1__13,inputs_1__12,
                    inputs_1__11,inputs_1__10,inputs_1__9,inputs_1__8,
                    inputs_1__7,inputs_1__6,inputs_1__5,inputs_1__4,inputs_1__3,
                    inputs_1__2,inputs_1__1,inputs_1__0}), .c ({inputs_2__15,
                    inputs_2__14,inputs_2__13,inputs_2__12,inputs_2__11,
                    inputs_2__10,inputs_2__9,inputs_2__8,inputs_2__7,inputs_2__6
                    ,inputs_2__5,inputs_2__4,inputs_2__3,inputs_2__2,inputs_2__1
                    ,inputs_2__0}), .d ({inputs_3__15,inputs_3__14,inputs_3__13,
                    inputs_3__12,inputs_3__11,inputs_3__10,inputs_3__9,
                    inputs_3__8,inputs_3__7,inputs_3__6,inputs_3__5,inputs_3__4,
                    inputs_3__3,inputs_3__2,inputs_3__1,inputs_3__0}), .sum ({
                    sum1_15,sum1_14,sum1_13,sum1_12,sum1_11,sum1_10,sum1_9,
                    sum1_8,sum1_7,sum1_6,sum1_5,sum1_4,sum1_3,sum1_2,sum1_1,
                    sum1_0})) ;
    Adder4Values_16 sum2Map (.a ({inputs_4__15,inputs_4__14,inputs_4__13,
                    inputs_4__12,inputs_4__11,inputs_4__10,inputs_4__9,
                    inputs_4__8,inputs_4__7,inputs_4__6,inputs_4__5,inputs_4__4,
                    inputs_4__3,inputs_4__2,inputs_4__1,inputs_4__0}), .b ({
                    inputs_5__15,inputs_5__14,inputs_5__13,inputs_5__12,
                    inputs_5__11,inputs_5__10,inputs_5__9,inputs_5__8,
                    inputs_5__7,inputs_5__6,inputs_5__5,inputs_5__4,inputs_5__3,
                    inputs_5__2,inputs_5__1,inputs_5__0}), .c ({inputs_6__15,
                    inputs_6__14,inputs_6__13,inputs_6__12,inputs_6__11,
                    inputs_6__10,inputs_6__9,inputs_6__8,inputs_6__7,inputs_6__6
                    ,inputs_6__5,inputs_6__4,inputs_6__3,inputs_6__2,inputs_6__1
                    ,inputs_6__0}), .d ({inputs_7__15,inputs_7__14,inputs_7__13,
                    inputs_7__12,inputs_7__11,inputs_7__10,inputs_7__9,
                    inputs_7__8,inputs_7__7,inputs_7__6,inputs_7__5,inputs_7__4,
                    inputs_7__3,inputs_7__2,inputs_7__1,inputs_7__0}), .sum ({
                    sum2_15,sum2_14,sum2_13,sum2_12,sum2_11,sum2_10,sum2_9,
                    sum2_8,sum2_7,sum2_6,sum2_5,sum2_4,sum2_3,sum2_2,sum2_1,
                    sum2_0})) ;
    NBitAdder_16 sumFinalMap (.a ({sum1_15,sum1_14,sum1_13,sum1_12,sum1_11,
                 sum1_10,sum1_9,sum1_8,sum1_7,sum1_6,sum1_5,sum1_4,sum1_3,sum1_2
                 ,sum1_1,sum1_0}), .b ({sum2_15,sum2_14,sum2_13,sum2_12,sum2_11,
                 sum2_10,sum2_9,sum2_8,sum2_7,sum2_6,sum2_5,sum2_4,sum2_3,sum2_2
                 ,sum2_1,sum2_0}), .carryIn (GND), .sum ({sum[15],sum[14],
                 sum[13],sum[12],sum[11],sum[10],sum[9],sum[8],sum[7],sum[6],
                 sum[5],sum[4],sum[3],sum[2],sum[1],sum[0]}), .carryOut (
                 \$dummy [0])) ;
    fake_gnd ix121 (.Y (GND)) ;
endmodule


module Adder4Values_16 ( a, b, c, d, sum ) ;

    input [15:0]a ;
    input [15:0]b ;
    input [15:0]c ;
    input [15:0]d ;
    output [15:0]sum ;

    wire sum1_15, sum1_14, sum1_13, sum1_12, sum1_11, sum1_10, sum1_9, sum1_8, 
         sum1_7, sum1_6, sum1_5, sum1_4, sum1_3, sum1_2, sum1_1, sum1_0, sum2_15, 
         sum2_14, sum2_13, sum2_12, sum2_11, sum2_10, sum2_9, sum2_8, sum2_7, 
         sum2_6, sum2_5, sum2_4, sum2_3, sum2_2, sum2_1, sum2_0, GND;
    wire [2:0] \$dummy ;




    NBitAdder_16 sum1Map (.a ({a[15],a[14],a[13],a[12],a[11],a[10],a[9],a[8],
                 a[7],a[6],a[5],a[4],a[3],a[2],a[1],a[0]}), .b ({b[15],b[14],
                 b[13],b[12],b[11],b[10],b[9],b[8],b[7],b[6],b[5],b[4],b[3],b[2]
                 ,b[1],b[0]}), .carryIn (GND), .sum ({sum1_15,sum1_14,sum1_13,
                 sum1_12,sum1_11,sum1_10,sum1_9,sum1_8,sum1_7,sum1_6,sum1_5,
                 sum1_4,sum1_3,sum1_2,sum1_1,sum1_0}), .carryOut (\$dummy [0])
                 ) ;
    NBitAdder_16 sum2Map (.a ({c[15],c[14],c[13],c[12],c[11],c[10],c[9],c[8],
                 c[7],c[6],c[5],c[4],c[3],c[2],c[1],c[0]}), .b ({d[15],d[14],
                 d[13],d[12],d[11],d[10],d[9],d[8],d[7],d[6],d[5],d[4],d[3],d[2]
                 ,d[1],d[0]}), .carryIn (GND), .sum ({sum2_15,sum2_14,sum2_13,
                 sum2_12,sum2_11,sum2_10,sum2_9,sum2_8,sum2_7,sum2_6,sum2_5,
                 sum2_4,sum2_3,sum2_2,sum2_1,sum2_0}), .carryOut (\$dummy [1])
                 ) ;
    NBitAdder_16 sumFinalMap (.a ({sum1_15,sum1_14,sum1_13,sum1_12,sum1_11,
                 sum1_10,sum1_9,sum1_8,sum1_7,sum1_6,sum1_5,sum1_4,sum1_3,sum1_2
                 ,sum1_1,sum1_0}), .b ({sum2_15,sum2_14,sum2_13,sum2_12,sum2_11,
                 sum2_10,sum2_9,sum2_8,sum2_7,sum2_6,sum2_5,sum2_4,sum2_3,sum2_2
                 ,sum2_1,sum2_0}), .carryIn (GND), .sum ({sum[15],sum[14],
                 sum[13],sum[12],sum[11],sum[10],sum[9],sum[8],sum[7],sum[6],
                 sum[5],sum[4],sum[3],sum[2],sum[1],sum[0]}), .carryOut (
                 \$dummy [2])) ;
    fake_gnd ix125 (.Y (GND)) ;
endmodule


module NBitAdder_16 ( a, b, carryIn, sum, carryOut ) ;

    input [15:0]a ;
    input [15:0]b ;
    input carryIn ;
    output [15:0]sum ;
    output carryOut ;

    wire temp_14, temp_13, temp_12, temp_11, temp_10, temp_9, temp_8, temp_7, 
         temp_6, temp_5, temp_4, temp_3, temp_2, temp_1, temp_0;



    FullAdder f0 (.a (a[0]), .b (b[0]), .cin (carryIn), .s (sum[0]), .cout (
              temp_0)) ;
    FullAdder loop1_1_fx (.a (a[1]), .b (b[1]), .cin (temp_0), .s (sum[1]), .cout (
              temp_1)) ;
    FullAdder loop1_2_fx (.a (a[2]), .b (b[2]), .cin (temp_1), .s (sum[2]), .cout (
              temp_2)) ;
    FullAdder loop1_3_fx (.a (a[3]), .b (b[3]), .cin (temp_2), .s (sum[3]), .cout (
              temp_3)) ;
    FullAdder loop1_4_fx (.a (a[4]), .b (b[4]), .cin (temp_3), .s (sum[4]), .cout (
              temp_4)) ;
    FullAdder loop1_5_fx (.a (a[5]), .b (b[5]), .cin (temp_4), .s (sum[5]), .cout (
              temp_5)) ;
    FullAdder loop1_6_fx (.a (a[6]), .b (b[6]), .cin (temp_5), .s (sum[6]), .cout (
              temp_6)) ;
    FullAdder loop1_7_fx (.a (a[7]), .b (b[7]), .cin (temp_6), .s (sum[7]), .cout (
              temp_7)) ;
    FullAdder loop1_8_fx (.a (a[8]), .b (b[8]), .cin (temp_7), .s (sum[8]), .cout (
              temp_8)) ;
    FullAdder loop1_9_fx (.a (a[9]), .b (b[9]), .cin (temp_8), .s (sum[9]), .cout (
              temp_9)) ;
    FullAdder loop1_10_fx (.a (a[10]), .b (b[10]), .cin (temp_9), .s (sum[10]), 
              .cout (temp_10)) ;
    FullAdder loop1_11_fx (.a (a[11]), .b (b[11]), .cin (temp_10), .s (sum[11])
              , .cout (temp_11)) ;
    FullAdder loop1_12_fx (.a (a[12]), .b (b[12]), .cin (temp_11), .s (sum[12])
              , .cout (temp_12)) ;
    FullAdder loop1_13_fx (.a (a[13]), .b (b[13]), .cin (temp_12), .s (sum[13])
              , .cout (temp_13)) ;
    FullAdder loop1_14_fx (.a (a[14]), .b (b[14]), .cin (temp_13), .s (sum[14])
              , .cout (temp_14)) ;
    FullAdder loop1_15_fx (.a (a[15]), .b (b[15]), .cin (temp_14), .s (sum[15])
              , .cout (carryOut)) ;
endmodule


module CNNMuls_25 ( filter_24__7, filter_24__6, filter_24__5, filter_24__4, 
                    filter_24__3, filter_24__2, filter_24__1, filter_24__0, 
                    filter_23__7, filter_23__6, filter_23__5, filter_23__4, 
                    filter_23__3, filter_23__2, filter_23__1, filter_23__0, 
                    filter_22__7, filter_22__6, filter_22__5, filter_22__4, 
                    filter_22__3, filter_22__2, filter_22__1, filter_22__0, 
                    filter_21__7, filter_21__6, filter_21__5, filter_21__4, 
                    filter_21__3, filter_21__2, filter_21__1, filter_21__0, 
                    filter_20__7, filter_20__6, filter_20__5, filter_20__4, 
                    filter_20__3, filter_20__2, filter_20__1, filter_20__0, 
                    filter_19__7, filter_19__6, filter_19__5, filter_19__4, 
                    filter_19__3, filter_19__2, filter_19__1, filter_19__0, 
                    filter_18__7, filter_18__6, filter_18__5, filter_18__4, 
                    filter_18__3, filter_18__2, filter_18__1, filter_18__0, 
                    filter_17__7, filter_17__6, filter_17__5, filter_17__4, 
                    filter_17__3, filter_17__2, filter_17__1, filter_17__0, 
                    filter_16__7, filter_16__6, filter_16__5, filter_16__4, 
                    filter_16__3, filter_16__2, filter_16__1, filter_16__0, 
                    filter_15__7, filter_15__6, filter_15__5, filter_15__4, 
                    filter_15__3, filter_15__2, filter_15__1, filter_15__0, 
                    filter_14__7, filter_14__6, filter_14__5, filter_14__4, 
                    filter_14__3, filter_14__2, filter_14__1, filter_14__0, 
                    filter_13__7, filter_13__6, filter_13__5, filter_13__4, 
                    filter_13__3, filter_13__2, filter_13__1, filter_13__0, 
                    filter_12__7, filter_12__6, filter_12__5, filter_12__4, 
                    filter_12__3, filter_12__2, filter_12__1, filter_12__0, 
                    filter_11__7, filter_11__6, filter_11__5, filter_11__4, 
                    filter_11__3, filter_11__2, filter_11__1, filter_11__0, 
                    filter_10__7, filter_10__6, filter_10__5, filter_10__4, 
                    filter_10__3, filter_10__2, filter_10__1, filter_10__0, 
                    filter_9__7, filter_9__6, filter_9__5, filter_9__4, 
                    filter_9__3, filter_9__2, filter_9__1, filter_9__0, 
                    filter_8__7, filter_8__6, filter_8__5, filter_8__4, 
                    filter_8__3, filter_8__2, filter_8__1, filter_8__0, 
                    filter_7__7, filter_7__6, filter_7__5, filter_7__4, 
                    filter_7__3, filter_7__2, filter_7__1, filter_7__0, 
                    filter_6__7, filter_6__6, filter_6__5, filter_6__4, 
                    filter_6__3, filter_6__2, filter_6__1, filter_6__0, 
                    filter_5__7, filter_5__6, filter_5__5, filter_5__4, 
                    filter_5__3, filter_5__2, filter_5__1, filter_5__0, 
                    filter_4__7, filter_4__6, filter_4__5, filter_4__4, 
                    filter_4__3, filter_4__2, filter_4__1, filter_4__0, 
                    filter_3__7, filter_3__6, filter_3__5, filter_3__4, 
                    filter_3__3, filter_3__2, filter_3__1, filter_3__0, 
                    filter_2__7, filter_2__6, filter_2__5, filter_2__4, 
                    filter_2__3, filter_2__2, filter_2__1, filter_2__0, 
                    filter_1__7, filter_1__6, filter_1__5, filter_1__4, 
                    filter_1__3, filter_1__2, filter_1__1, filter_1__0, 
                    filter_0__7, filter_0__6, filter_0__5, filter_0__4, 
                    filter_0__3, filter_0__2, filter_0__1, filter_0__0, 
                    window_24__15, window_24__14, window_24__13, window_24__12, 
                    window_24__11, window_24__10, window_24__9, window_24__8, 
                    window_24__7, window_24__6, window_24__5, window_24__4, 
                    window_24__3, window_24__2, window_24__1, window_24__0, 
                    window_23__15, window_23__14, window_23__13, window_23__12, 
                    window_23__11, window_23__10, window_23__9, window_23__8, 
                    window_23__7, window_23__6, window_23__5, window_23__4, 
                    window_23__3, window_23__2, window_23__1, window_23__0, 
                    window_22__15, window_22__14, window_22__13, window_22__12, 
                    window_22__11, window_22__10, window_22__9, window_22__8, 
                    window_22__7, window_22__6, window_22__5, window_22__4, 
                    window_22__3, window_22__2, window_22__1, window_22__0, 
                    window_21__15, window_21__14, window_21__13, window_21__12, 
                    window_21__11, window_21__10, window_21__9, window_21__8, 
                    window_21__7, window_21__6, window_21__5, window_21__4, 
                    window_21__3, window_21__2, window_21__1, window_21__0, 
                    window_20__15, window_20__14, window_20__13, window_20__12, 
                    window_20__11, window_20__10, window_20__9, window_20__8, 
                    window_20__7, window_20__6, window_20__5, window_20__4, 
                    window_20__3, window_20__2, window_20__1, window_20__0, 
                    window_19__15, window_19__14, window_19__13, window_19__12, 
                    window_19__11, window_19__10, window_19__9, window_19__8, 
                    window_19__7, window_19__6, window_19__5, window_19__4, 
                    window_19__3, window_19__2, window_19__1, window_19__0, 
                    window_18__15, window_18__14, window_18__13, window_18__12, 
                    window_18__11, window_18__10, window_18__9, window_18__8, 
                    window_18__7, window_18__6, window_18__5, window_18__4, 
                    window_18__3, window_18__2, window_18__1, window_18__0, 
                    window_17__15, window_17__14, window_17__13, window_17__12, 
                    window_17__11, window_17__10, window_17__9, window_17__8, 
                    window_17__7, window_17__6, window_17__5, window_17__4, 
                    window_17__3, window_17__2, window_17__1, window_17__0, 
                    window_16__15, window_16__14, window_16__13, window_16__12, 
                    window_16__11, window_16__10, window_16__9, window_16__8, 
                    window_16__7, window_16__6, window_16__5, window_16__4, 
                    window_16__3, window_16__2, window_16__1, window_16__0, 
                    window_15__15, window_15__14, window_15__13, window_15__12, 
                    window_15__11, window_15__10, window_15__9, window_15__8, 
                    window_15__7, window_15__6, window_15__5, window_15__4, 
                    window_15__3, window_15__2, window_15__1, window_15__0, 
                    window_14__15, window_14__14, window_14__13, window_14__12, 
                    window_14__11, window_14__10, window_14__9, window_14__8, 
                    window_14__7, window_14__6, window_14__5, window_14__4, 
                    window_14__3, window_14__2, window_14__1, window_14__0, 
                    window_13__15, window_13__14, window_13__13, window_13__12, 
                    window_13__11, window_13__10, window_13__9, window_13__8, 
                    window_13__7, window_13__6, window_13__5, window_13__4, 
                    window_13__3, window_13__2, window_13__1, window_13__0, 
                    window_12__15, window_12__14, window_12__13, window_12__12, 
                    window_12__11, window_12__10, window_12__9, window_12__8, 
                    window_12__7, window_12__6, window_12__5, window_12__4, 
                    window_12__3, window_12__2, window_12__1, window_12__0, 
                    window_11__15, window_11__14, window_11__13, window_11__12, 
                    window_11__11, window_11__10, window_11__9, window_11__8, 
                    window_11__7, window_11__6, window_11__5, window_11__4, 
                    window_11__3, window_11__2, window_11__1, window_11__0, 
                    window_10__15, window_10__14, window_10__13, window_10__12, 
                    window_10__11, window_10__10, window_10__9, window_10__8, 
                    window_10__7, window_10__6, window_10__5, window_10__4, 
                    window_10__3, window_10__2, window_10__1, window_10__0, 
                    window_9__15, window_9__14, window_9__13, window_9__12, 
                    window_9__11, window_9__10, window_9__9, window_9__8, 
                    window_9__7, window_9__6, window_9__5, window_9__4, 
                    window_9__3, window_9__2, window_9__1, window_9__0, 
                    window_8__15, window_8__14, window_8__13, window_8__12, 
                    window_8__11, window_8__10, window_8__9, window_8__8, 
                    window_8__7, window_8__6, window_8__5, window_8__4, 
                    window_8__3, window_8__2, window_8__1, window_8__0, 
                    window_7__15, window_7__14, window_7__13, window_7__12, 
                    window_7__11, window_7__10, window_7__9, window_7__8, 
                    window_7__7, window_7__6, window_7__5, window_7__4, 
                    window_7__3, window_7__2, window_7__1, window_7__0, 
                    window_6__15, window_6__14, window_6__13, window_6__12, 
                    window_6__11, window_6__10, window_6__9, window_6__8, 
                    window_6__7, window_6__6, window_6__5, window_6__4, 
                    window_6__3, window_6__2, window_6__1, window_6__0, 
                    window_5__15, window_5__14, window_5__13, window_5__12, 
                    window_5__11, window_5__10, window_5__9, window_5__8, 
                    window_5__7, window_5__6, window_5__5, window_5__4, 
                    window_5__3, window_5__2, window_5__1, window_5__0, 
                    window_4__15, window_4__14, window_4__13, window_4__12, 
                    window_4__11, window_4__10, window_4__9, window_4__8, 
                    window_4__7, window_4__6, window_4__5, window_4__4, 
                    window_4__3, window_4__2, window_4__1, window_4__0, 
                    window_3__15, window_3__14, window_3__13, window_3__12, 
                    window_3__11, window_3__10, window_3__9, window_3__8, 
                    window_3__7, window_3__6, window_3__5, window_3__4, 
                    window_3__3, window_3__2, window_3__1, window_3__0, 
                    window_2__15, window_2__14, window_2__13, window_2__12, 
                    window_2__11, window_2__10, window_2__9, window_2__8, 
                    window_2__7, window_2__6, window_2__5, window_2__4, 
                    window_2__3, window_2__2, window_2__1, window_2__0, 
                    window_1__15, window_1__14, window_1__13, window_1__12, 
                    window_1__11, window_1__10, window_1__9, window_1__8, 
                    window_1__7, window_1__6, window_1__5, window_1__4, 
                    window_1__3, window_1__2, window_1__1, window_1__0, 
                    window_0__15, window_0__14, window_0__13, window_0__12, 
                    window_0__11, window_0__10, window_0__9, window_0__8, 
                    window_0__7, window_0__6, window_0__5, window_0__4, 
                    window_0__3, window_0__2, window_0__1, window_0__0, 
                    outputs_24__15, outputs_24__14, outputs_24__13, 
                    outputs_24__12, outputs_24__11, outputs_24__10, 
                    outputs_24__9, outputs_24__8, outputs_24__7, outputs_24__6, 
                    outputs_24__5, outputs_24__4, outputs_24__3, outputs_24__2, 
                    outputs_24__1, outputs_24__0, outputs_23__15, outputs_23__14, 
                    outputs_23__13, outputs_23__12, outputs_23__11, 
                    outputs_23__10, outputs_23__9, outputs_23__8, outputs_23__7, 
                    outputs_23__6, outputs_23__5, outputs_23__4, outputs_23__3, 
                    outputs_23__2, outputs_23__1, outputs_23__0, outputs_22__15, 
                    outputs_22__14, outputs_22__13, outputs_22__12, 
                    outputs_22__11, outputs_22__10, outputs_22__9, outputs_22__8, 
                    outputs_22__7, outputs_22__6, outputs_22__5, outputs_22__4, 
                    outputs_22__3, outputs_22__2, outputs_22__1, outputs_22__0, 
                    outputs_21__15, outputs_21__14, outputs_21__13, 
                    outputs_21__12, outputs_21__11, outputs_21__10, 
                    outputs_21__9, outputs_21__8, outputs_21__7, outputs_21__6, 
                    outputs_21__5, outputs_21__4, outputs_21__3, outputs_21__2, 
                    outputs_21__1, outputs_21__0, outputs_20__15, outputs_20__14, 
                    outputs_20__13, outputs_20__12, outputs_20__11, 
                    outputs_20__10, outputs_20__9, outputs_20__8, outputs_20__7, 
                    outputs_20__6, outputs_20__5, outputs_20__4, outputs_20__3, 
                    outputs_20__2, outputs_20__1, outputs_20__0, outputs_19__15, 
                    outputs_19__14, outputs_19__13, outputs_19__12, 
                    outputs_19__11, outputs_19__10, outputs_19__9, outputs_19__8, 
                    outputs_19__7, outputs_19__6, outputs_19__5, outputs_19__4, 
                    outputs_19__3, outputs_19__2, outputs_19__1, outputs_19__0, 
                    outputs_18__15, outputs_18__14, outputs_18__13, 
                    outputs_18__12, outputs_18__11, outputs_18__10, 
                    outputs_18__9, outputs_18__8, outputs_18__7, outputs_18__6, 
                    outputs_18__5, outputs_18__4, outputs_18__3, outputs_18__2, 
                    outputs_18__1, outputs_18__0, outputs_17__15, outputs_17__14, 
                    outputs_17__13, outputs_17__12, outputs_17__11, 
                    outputs_17__10, outputs_17__9, outputs_17__8, outputs_17__7, 
                    outputs_17__6, outputs_17__5, outputs_17__4, outputs_17__3, 
                    outputs_17__2, outputs_17__1, outputs_17__0, outputs_16__15, 
                    outputs_16__14, outputs_16__13, outputs_16__12, 
                    outputs_16__11, outputs_16__10, outputs_16__9, outputs_16__8, 
                    outputs_16__7, outputs_16__6, outputs_16__5, outputs_16__4, 
                    outputs_16__3, outputs_16__2, outputs_16__1, outputs_16__0, 
                    outputs_15__15, outputs_15__14, outputs_15__13, 
                    outputs_15__12, outputs_15__11, outputs_15__10, 
                    outputs_15__9, outputs_15__8, outputs_15__7, outputs_15__6, 
                    outputs_15__5, outputs_15__4, outputs_15__3, outputs_15__2, 
                    outputs_15__1, outputs_15__0, outputs_14__15, outputs_14__14, 
                    outputs_14__13, outputs_14__12, outputs_14__11, 
                    outputs_14__10, outputs_14__9, outputs_14__8, outputs_14__7, 
                    outputs_14__6, outputs_14__5, outputs_14__4, outputs_14__3, 
                    outputs_14__2, outputs_14__1, outputs_14__0, outputs_13__15, 
                    outputs_13__14, outputs_13__13, outputs_13__12, 
                    outputs_13__11, outputs_13__10, outputs_13__9, outputs_13__8, 
                    outputs_13__7, outputs_13__6, outputs_13__5, outputs_13__4, 
                    outputs_13__3, outputs_13__2, outputs_13__1, outputs_13__0, 
                    outputs_12__15, outputs_12__14, outputs_12__13, 
                    outputs_12__12, outputs_12__11, outputs_12__10, 
                    outputs_12__9, outputs_12__8, outputs_12__7, outputs_12__6, 
                    outputs_12__5, outputs_12__4, outputs_12__3, outputs_12__2, 
                    outputs_12__1, outputs_12__0, outputs_11__15, outputs_11__14, 
                    outputs_11__13, outputs_11__12, outputs_11__11, 
                    outputs_11__10, outputs_11__9, outputs_11__8, outputs_11__7, 
                    outputs_11__6, outputs_11__5, outputs_11__4, outputs_11__3, 
                    outputs_11__2, outputs_11__1, outputs_11__0, outputs_10__15, 
                    outputs_10__14, outputs_10__13, outputs_10__12, 
                    outputs_10__11, outputs_10__10, outputs_10__9, outputs_10__8, 
                    outputs_10__7, outputs_10__6, outputs_10__5, outputs_10__4, 
                    outputs_10__3, outputs_10__2, outputs_10__1, outputs_10__0, 
                    outputs_9__15, outputs_9__14, outputs_9__13, outputs_9__12, 
                    outputs_9__11, outputs_9__10, outputs_9__9, outputs_9__8, 
                    outputs_9__7, outputs_9__6, outputs_9__5, outputs_9__4, 
                    outputs_9__3, outputs_9__2, outputs_9__1, outputs_9__0, 
                    outputs_8__15, outputs_8__14, outputs_8__13, outputs_8__12, 
                    outputs_8__11, outputs_8__10, outputs_8__9, outputs_8__8, 
                    outputs_8__7, outputs_8__6, outputs_8__5, outputs_8__4, 
                    outputs_8__3, outputs_8__2, outputs_8__1, outputs_8__0, 
                    outputs_7__15, outputs_7__14, outputs_7__13, outputs_7__12, 
                    outputs_7__11, outputs_7__10, outputs_7__9, outputs_7__8, 
                    outputs_7__7, outputs_7__6, outputs_7__5, outputs_7__4, 
                    outputs_7__3, outputs_7__2, outputs_7__1, outputs_7__0, 
                    outputs_6__15, outputs_6__14, outputs_6__13, outputs_6__12, 
                    outputs_6__11, outputs_6__10, outputs_6__9, outputs_6__8, 
                    outputs_6__7, outputs_6__6, outputs_6__5, outputs_6__4, 
                    outputs_6__3, outputs_6__2, outputs_6__1, outputs_6__0, 
                    outputs_5__15, outputs_5__14, outputs_5__13, outputs_5__12, 
                    outputs_5__11, outputs_5__10, outputs_5__9, outputs_5__8, 
                    outputs_5__7, outputs_5__6, outputs_5__5, outputs_5__4, 
                    outputs_5__3, outputs_5__2, outputs_5__1, outputs_5__0, 
                    outputs_4__15, outputs_4__14, outputs_4__13, outputs_4__12, 
                    outputs_4__11, outputs_4__10, outputs_4__9, outputs_4__8, 
                    outputs_4__7, outputs_4__6, outputs_4__5, outputs_4__4, 
                    outputs_4__3, outputs_4__2, outputs_4__1, outputs_4__0, 
                    outputs_3__15, outputs_3__14, outputs_3__13, outputs_3__12, 
                    outputs_3__11, outputs_3__10, outputs_3__9, outputs_3__8, 
                    outputs_3__7, outputs_3__6, outputs_3__5, outputs_3__4, 
                    outputs_3__3, outputs_3__2, outputs_3__1, outputs_3__0, 
                    outputs_2__15, outputs_2__14, outputs_2__13, outputs_2__12, 
                    outputs_2__11, outputs_2__10, outputs_2__9, outputs_2__8, 
                    outputs_2__7, outputs_2__6, outputs_2__5, outputs_2__4, 
                    outputs_2__3, outputs_2__2, outputs_2__1, outputs_2__0, 
                    outputs_1__15, outputs_1__14, outputs_1__13, outputs_1__12, 
                    outputs_1__11, outputs_1__10, outputs_1__9, outputs_1__8, 
                    outputs_1__7, outputs_1__6, outputs_1__5, outputs_1__4, 
                    outputs_1__3, outputs_1__2, outputs_1__1, outputs_1__0, 
                    outputs_0__15, outputs_0__14, outputs_0__13, outputs_0__12, 
                    outputs_0__11, outputs_0__10, outputs_0__9, outputs_0__8, 
                    outputs_0__7, outputs_0__6, outputs_0__5, outputs_0__4, 
                    outputs_0__3, outputs_0__2, outputs_0__1, outputs_0__0, clk, 
                    start, rst, doneOut, workingOut ) ;

    input filter_24__7 ;
    input filter_24__6 ;
    input filter_24__5 ;
    input filter_24__4 ;
    input filter_24__3 ;
    input filter_24__2 ;
    input filter_24__1 ;
    input filter_24__0 ;
    input filter_23__7 ;
    input filter_23__6 ;
    input filter_23__5 ;
    input filter_23__4 ;
    input filter_23__3 ;
    input filter_23__2 ;
    input filter_23__1 ;
    input filter_23__0 ;
    input filter_22__7 ;
    input filter_22__6 ;
    input filter_22__5 ;
    input filter_22__4 ;
    input filter_22__3 ;
    input filter_22__2 ;
    input filter_22__1 ;
    input filter_22__0 ;
    input filter_21__7 ;
    input filter_21__6 ;
    input filter_21__5 ;
    input filter_21__4 ;
    input filter_21__3 ;
    input filter_21__2 ;
    input filter_21__1 ;
    input filter_21__0 ;
    input filter_20__7 ;
    input filter_20__6 ;
    input filter_20__5 ;
    input filter_20__4 ;
    input filter_20__3 ;
    input filter_20__2 ;
    input filter_20__1 ;
    input filter_20__0 ;
    input filter_19__7 ;
    input filter_19__6 ;
    input filter_19__5 ;
    input filter_19__4 ;
    input filter_19__3 ;
    input filter_19__2 ;
    input filter_19__1 ;
    input filter_19__0 ;
    input filter_18__7 ;
    input filter_18__6 ;
    input filter_18__5 ;
    input filter_18__4 ;
    input filter_18__3 ;
    input filter_18__2 ;
    input filter_18__1 ;
    input filter_18__0 ;
    input filter_17__7 ;
    input filter_17__6 ;
    input filter_17__5 ;
    input filter_17__4 ;
    input filter_17__3 ;
    input filter_17__2 ;
    input filter_17__1 ;
    input filter_17__0 ;
    input filter_16__7 ;
    input filter_16__6 ;
    input filter_16__5 ;
    input filter_16__4 ;
    input filter_16__3 ;
    input filter_16__2 ;
    input filter_16__1 ;
    input filter_16__0 ;
    input filter_15__7 ;
    input filter_15__6 ;
    input filter_15__5 ;
    input filter_15__4 ;
    input filter_15__3 ;
    input filter_15__2 ;
    input filter_15__1 ;
    input filter_15__0 ;
    input filter_14__7 ;
    input filter_14__6 ;
    input filter_14__5 ;
    input filter_14__4 ;
    input filter_14__3 ;
    input filter_14__2 ;
    input filter_14__1 ;
    input filter_14__0 ;
    input filter_13__7 ;
    input filter_13__6 ;
    input filter_13__5 ;
    input filter_13__4 ;
    input filter_13__3 ;
    input filter_13__2 ;
    input filter_13__1 ;
    input filter_13__0 ;
    input filter_12__7 ;
    input filter_12__6 ;
    input filter_12__5 ;
    input filter_12__4 ;
    input filter_12__3 ;
    input filter_12__2 ;
    input filter_12__1 ;
    input filter_12__0 ;
    input filter_11__7 ;
    input filter_11__6 ;
    input filter_11__5 ;
    input filter_11__4 ;
    input filter_11__3 ;
    input filter_11__2 ;
    input filter_11__1 ;
    input filter_11__0 ;
    input filter_10__7 ;
    input filter_10__6 ;
    input filter_10__5 ;
    input filter_10__4 ;
    input filter_10__3 ;
    input filter_10__2 ;
    input filter_10__1 ;
    input filter_10__0 ;
    input filter_9__7 ;
    input filter_9__6 ;
    input filter_9__5 ;
    input filter_9__4 ;
    input filter_9__3 ;
    input filter_9__2 ;
    input filter_9__1 ;
    input filter_9__0 ;
    input filter_8__7 ;
    input filter_8__6 ;
    input filter_8__5 ;
    input filter_8__4 ;
    input filter_8__3 ;
    input filter_8__2 ;
    input filter_8__1 ;
    input filter_8__0 ;
    input filter_7__7 ;
    input filter_7__6 ;
    input filter_7__5 ;
    input filter_7__4 ;
    input filter_7__3 ;
    input filter_7__2 ;
    input filter_7__1 ;
    input filter_7__0 ;
    input filter_6__7 ;
    input filter_6__6 ;
    input filter_6__5 ;
    input filter_6__4 ;
    input filter_6__3 ;
    input filter_6__2 ;
    input filter_6__1 ;
    input filter_6__0 ;
    input filter_5__7 ;
    input filter_5__6 ;
    input filter_5__5 ;
    input filter_5__4 ;
    input filter_5__3 ;
    input filter_5__2 ;
    input filter_5__1 ;
    input filter_5__0 ;
    input filter_4__7 ;
    input filter_4__6 ;
    input filter_4__5 ;
    input filter_4__4 ;
    input filter_4__3 ;
    input filter_4__2 ;
    input filter_4__1 ;
    input filter_4__0 ;
    input filter_3__7 ;
    input filter_3__6 ;
    input filter_3__5 ;
    input filter_3__4 ;
    input filter_3__3 ;
    input filter_3__2 ;
    input filter_3__1 ;
    input filter_3__0 ;
    input filter_2__7 ;
    input filter_2__6 ;
    input filter_2__5 ;
    input filter_2__4 ;
    input filter_2__3 ;
    input filter_2__2 ;
    input filter_2__1 ;
    input filter_2__0 ;
    input filter_1__7 ;
    input filter_1__6 ;
    input filter_1__5 ;
    input filter_1__4 ;
    input filter_1__3 ;
    input filter_1__2 ;
    input filter_1__1 ;
    input filter_1__0 ;
    input filter_0__7 ;
    input filter_0__6 ;
    input filter_0__5 ;
    input filter_0__4 ;
    input filter_0__3 ;
    input filter_0__2 ;
    input filter_0__1 ;
    input filter_0__0 ;
    input window_24__15 ;
    input window_24__14 ;
    input window_24__13 ;
    input window_24__12 ;
    input window_24__11 ;
    input window_24__10 ;
    input window_24__9 ;
    input window_24__8 ;
    input window_24__7 ;
    input window_24__6 ;
    input window_24__5 ;
    input window_24__4 ;
    input window_24__3 ;
    input window_24__2 ;
    input window_24__1 ;
    input window_24__0 ;
    input window_23__15 ;
    input window_23__14 ;
    input window_23__13 ;
    input window_23__12 ;
    input window_23__11 ;
    input window_23__10 ;
    input window_23__9 ;
    input window_23__8 ;
    input window_23__7 ;
    input window_23__6 ;
    input window_23__5 ;
    input window_23__4 ;
    input window_23__3 ;
    input window_23__2 ;
    input window_23__1 ;
    input window_23__0 ;
    input window_22__15 ;
    input window_22__14 ;
    input window_22__13 ;
    input window_22__12 ;
    input window_22__11 ;
    input window_22__10 ;
    input window_22__9 ;
    input window_22__8 ;
    input window_22__7 ;
    input window_22__6 ;
    input window_22__5 ;
    input window_22__4 ;
    input window_22__3 ;
    input window_22__2 ;
    input window_22__1 ;
    input window_22__0 ;
    input window_21__15 ;
    input window_21__14 ;
    input window_21__13 ;
    input window_21__12 ;
    input window_21__11 ;
    input window_21__10 ;
    input window_21__9 ;
    input window_21__8 ;
    input window_21__7 ;
    input window_21__6 ;
    input window_21__5 ;
    input window_21__4 ;
    input window_21__3 ;
    input window_21__2 ;
    input window_21__1 ;
    input window_21__0 ;
    input window_20__15 ;
    input window_20__14 ;
    input window_20__13 ;
    input window_20__12 ;
    input window_20__11 ;
    input window_20__10 ;
    input window_20__9 ;
    input window_20__8 ;
    input window_20__7 ;
    input window_20__6 ;
    input window_20__5 ;
    input window_20__4 ;
    input window_20__3 ;
    input window_20__2 ;
    input window_20__1 ;
    input window_20__0 ;
    input window_19__15 ;
    input window_19__14 ;
    input window_19__13 ;
    input window_19__12 ;
    input window_19__11 ;
    input window_19__10 ;
    input window_19__9 ;
    input window_19__8 ;
    input window_19__7 ;
    input window_19__6 ;
    input window_19__5 ;
    input window_19__4 ;
    input window_19__3 ;
    input window_19__2 ;
    input window_19__1 ;
    input window_19__0 ;
    input window_18__15 ;
    input window_18__14 ;
    input window_18__13 ;
    input window_18__12 ;
    input window_18__11 ;
    input window_18__10 ;
    input window_18__9 ;
    input window_18__8 ;
    input window_18__7 ;
    input window_18__6 ;
    input window_18__5 ;
    input window_18__4 ;
    input window_18__3 ;
    input window_18__2 ;
    input window_18__1 ;
    input window_18__0 ;
    input window_17__15 ;
    input window_17__14 ;
    input window_17__13 ;
    input window_17__12 ;
    input window_17__11 ;
    input window_17__10 ;
    input window_17__9 ;
    input window_17__8 ;
    input window_17__7 ;
    input window_17__6 ;
    input window_17__5 ;
    input window_17__4 ;
    input window_17__3 ;
    input window_17__2 ;
    input window_17__1 ;
    input window_17__0 ;
    input window_16__15 ;
    input window_16__14 ;
    input window_16__13 ;
    input window_16__12 ;
    input window_16__11 ;
    input window_16__10 ;
    input window_16__9 ;
    input window_16__8 ;
    input window_16__7 ;
    input window_16__6 ;
    input window_16__5 ;
    input window_16__4 ;
    input window_16__3 ;
    input window_16__2 ;
    input window_16__1 ;
    input window_16__0 ;
    input window_15__15 ;
    input window_15__14 ;
    input window_15__13 ;
    input window_15__12 ;
    input window_15__11 ;
    input window_15__10 ;
    input window_15__9 ;
    input window_15__8 ;
    input window_15__7 ;
    input window_15__6 ;
    input window_15__5 ;
    input window_15__4 ;
    input window_15__3 ;
    input window_15__2 ;
    input window_15__1 ;
    input window_15__0 ;
    input window_14__15 ;
    input window_14__14 ;
    input window_14__13 ;
    input window_14__12 ;
    input window_14__11 ;
    input window_14__10 ;
    input window_14__9 ;
    input window_14__8 ;
    input window_14__7 ;
    input window_14__6 ;
    input window_14__5 ;
    input window_14__4 ;
    input window_14__3 ;
    input window_14__2 ;
    input window_14__1 ;
    input window_14__0 ;
    input window_13__15 ;
    input window_13__14 ;
    input window_13__13 ;
    input window_13__12 ;
    input window_13__11 ;
    input window_13__10 ;
    input window_13__9 ;
    input window_13__8 ;
    input window_13__7 ;
    input window_13__6 ;
    input window_13__5 ;
    input window_13__4 ;
    input window_13__3 ;
    input window_13__2 ;
    input window_13__1 ;
    input window_13__0 ;
    input window_12__15 ;
    input window_12__14 ;
    input window_12__13 ;
    input window_12__12 ;
    input window_12__11 ;
    input window_12__10 ;
    input window_12__9 ;
    input window_12__8 ;
    input window_12__7 ;
    input window_12__6 ;
    input window_12__5 ;
    input window_12__4 ;
    input window_12__3 ;
    input window_12__2 ;
    input window_12__1 ;
    input window_12__0 ;
    input window_11__15 ;
    input window_11__14 ;
    input window_11__13 ;
    input window_11__12 ;
    input window_11__11 ;
    input window_11__10 ;
    input window_11__9 ;
    input window_11__8 ;
    input window_11__7 ;
    input window_11__6 ;
    input window_11__5 ;
    input window_11__4 ;
    input window_11__3 ;
    input window_11__2 ;
    input window_11__1 ;
    input window_11__0 ;
    input window_10__15 ;
    input window_10__14 ;
    input window_10__13 ;
    input window_10__12 ;
    input window_10__11 ;
    input window_10__10 ;
    input window_10__9 ;
    input window_10__8 ;
    input window_10__7 ;
    input window_10__6 ;
    input window_10__5 ;
    input window_10__4 ;
    input window_10__3 ;
    input window_10__2 ;
    input window_10__1 ;
    input window_10__0 ;
    input window_9__15 ;
    input window_9__14 ;
    input window_9__13 ;
    input window_9__12 ;
    input window_9__11 ;
    input window_9__10 ;
    input window_9__9 ;
    input window_9__8 ;
    input window_9__7 ;
    input window_9__6 ;
    input window_9__5 ;
    input window_9__4 ;
    input window_9__3 ;
    input window_9__2 ;
    input window_9__1 ;
    input window_9__0 ;
    input window_8__15 ;
    input window_8__14 ;
    input window_8__13 ;
    input window_8__12 ;
    input window_8__11 ;
    input window_8__10 ;
    input window_8__9 ;
    input window_8__8 ;
    input window_8__7 ;
    input window_8__6 ;
    input window_8__5 ;
    input window_8__4 ;
    input window_8__3 ;
    input window_8__2 ;
    input window_8__1 ;
    input window_8__0 ;
    input window_7__15 ;
    input window_7__14 ;
    input window_7__13 ;
    input window_7__12 ;
    input window_7__11 ;
    input window_7__10 ;
    input window_7__9 ;
    input window_7__8 ;
    input window_7__7 ;
    input window_7__6 ;
    input window_7__5 ;
    input window_7__4 ;
    input window_7__3 ;
    input window_7__2 ;
    input window_7__1 ;
    input window_7__0 ;
    input window_6__15 ;
    input window_6__14 ;
    input window_6__13 ;
    input window_6__12 ;
    input window_6__11 ;
    input window_6__10 ;
    input window_6__9 ;
    input window_6__8 ;
    input window_6__7 ;
    input window_6__6 ;
    input window_6__5 ;
    input window_6__4 ;
    input window_6__3 ;
    input window_6__2 ;
    input window_6__1 ;
    input window_6__0 ;
    input window_5__15 ;
    input window_5__14 ;
    input window_5__13 ;
    input window_5__12 ;
    input window_5__11 ;
    input window_5__10 ;
    input window_5__9 ;
    input window_5__8 ;
    input window_5__7 ;
    input window_5__6 ;
    input window_5__5 ;
    input window_5__4 ;
    input window_5__3 ;
    input window_5__2 ;
    input window_5__1 ;
    input window_5__0 ;
    input window_4__15 ;
    input window_4__14 ;
    input window_4__13 ;
    input window_4__12 ;
    input window_4__11 ;
    input window_4__10 ;
    input window_4__9 ;
    input window_4__8 ;
    input window_4__7 ;
    input window_4__6 ;
    input window_4__5 ;
    input window_4__4 ;
    input window_4__3 ;
    input window_4__2 ;
    input window_4__1 ;
    input window_4__0 ;
    input window_3__15 ;
    input window_3__14 ;
    input window_3__13 ;
    input window_3__12 ;
    input window_3__11 ;
    input window_3__10 ;
    input window_3__9 ;
    input window_3__8 ;
    input window_3__7 ;
    input window_3__6 ;
    input window_3__5 ;
    input window_3__4 ;
    input window_3__3 ;
    input window_3__2 ;
    input window_3__1 ;
    input window_3__0 ;
    input window_2__15 ;
    input window_2__14 ;
    input window_2__13 ;
    input window_2__12 ;
    input window_2__11 ;
    input window_2__10 ;
    input window_2__9 ;
    input window_2__8 ;
    input window_2__7 ;
    input window_2__6 ;
    input window_2__5 ;
    input window_2__4 ;
    input window_2__3 ;
    input window_2__2 ;
    input window_2__1 ;
    input window_2__0 ;
    input window_1__15 ;
    input window_1__14 ;
    input window_1__13 ;
    input window_1__12 ;
    input window_1__11 ;
    input window_1__10 ;
    input window_1__9 ;
    input window_1__8 ;
    input window_1__7 ;
    input window_1__6 ;
    input window_1__5 ;
    input window_1__4 ;
    input window_1__3 ;
    input window_1__2 ;
    input window_1__1 ;
    input window_1__0 ;
    input window_0__15 ;
    input window_0__14 ;
    input window_0__13 ;
    input window_0__12 ;
    input window_0__11 ;
    input window_0__10 ;
    input window_0__9 ;
    input window_0__8 ;
    input window_0__7 ;
    input window_0__6 ;
    input window_0__5 ;
    input window_0__4 ;
    input window_0__3 ;
    input window_0__2 ;
    input window_0__1 ;
    input window_0__0 ;
    output outputs_24__15 ;
    output outputs_24__14 ;
    output outputs_24__13 ;
    output outputs_24__12 ;
    output outputs_24__11 ;
    output outputs_24__10 ;
    output outputs_24__9 ;
    output outputs_24__8 ;
    output outputs_24__7 ;
    output outputs_24__6 ;
    output outputs_24__5 ;
    output outputs_24__4 ;
    output outputs_24__3 ;
    output outputs_24__2 ;
    output outputs_24__1 ;
    output outputs_24__0 ;
    output outputs_23__15 ;
    output outputs_23__14 ;
    output outputs_23__13 ;
    output outputs_23__12 ;
    output outputs_23__11 ;
    output outputs_23__10 ;
    output outputs_23__9 ;
    output outputs_23__8 ;
    output outputs_23__7 ;
    output outputs_23__6 ;
    output outputs_23__5 ;
    output outputs_23__4 ;
    output outputs_23__3 ;
    output outputs_23__2 ;
    output outputs_23__1 ;
    output outputs_23__0 ;
    output outputs_22__15 ;
    output outputs_22__14 ;
    output outputs_22__13 ;
    output outputs_22__12 ;
    output outputs_22__11 ;
    output outputs_22__10 ;
    output outputs_22__9 ;
    output outputs_22__8 ;
    output outputs_22__7 ;
    output outputs_22__6 ;
    output outputs_22__5 ;
    output outputs_22__4 ;
    output outputs_22__3 ;
    output outputs_22__2 ;
    output outputs_22__1 ;
    output outputs_22__0 ;
    output outputs_21__15 ;
    output outputs_21__14 ;
    output outputs_21__13 ;
    output outputs_21__12 ;
    output outputs_21__11 ;
    output outputs_21__10 ;
    output outputs_21__9 ;
    output outputs_21__8 ;
    output outputs_21__7 ;
    output outputs_21__6 ;
    output outputs_21__5 ;
    output outputs_21__4 ;
    output outputs_21__3 ;
    output outputs_21__2 ;
    output outputs_21__1 ;
    output outputs_21__0 ;
    output outputs_20__15 ;
    output outputs_20__14 ;
    output outputs_20__13 ;
    output outputs_20__12 ;
    output outputs_20__11 ;
    output outputs_20__10 ;
    output outputs_20__9 ;
    output outputs_20__8 ;
    output outputs_20__7 ;
    output outputs_20__6 ;
    output outputs_20__5 ;
    output outputs_20__4 ;
    output outputs_20__3 ;
    output outputs_20__2 ;
    output outputs_20__1 ;
    output outputs_20__0 ;
    output outputs_19__15 ;
    output outputs_19__14 ;
    output outputs_19__13 ;
    output outputs_19__12 ;
    output outputs_19__11 ;
    output outputs_19__10 ;
    output outputs_19__9 ;
    output outputs_19__8 ;
    output outputs_19__7 ;
    output outputs_19__6 ;
    output outputs_19__5 ;
    output outputs_19__4 ;
    output outputs_19__3 ;
    output outputs_19__2 ;
    output outputs_19__1 ;
    output outputs_19__0 ;
    output outputs_18__15 ;
    output outputs_18__14 ;
    output outputs_18__13 ;
    output outputs_18__12 ;
    output outputs_18__11 ;
    output outputs_18__10 ;
    output outputs_18__9 ;
    output outputs_18__8 ;
    output outputs_18__7 ;
    output outputs_18__6 ;
    output outputs_18__5 ;
    output outputs_18__4 ;
    output outputs_18__3 ;
    output outputs_18__2 ;
    output outputs_18__1 ;
    output outputs_18__0 ;
    output outputs_17__15 ;
    output outputs_17__14 ;
    output outputs_17__13 ;
    output outputs_17__12 ;
    output outputs_17__11 ;
    output outputs_17__10 ;
    output outputs_17__9 ;
    output outputs_17__8 ;
    output outputs_17__7 ;
    output outputs_17__6 ;
    output outputs_17__5 ;
    output outputs_17__4 ;
    output outputs_17__3 ;
    output outputs_17__2 ;
    output outputs_17__1 ;
    output outputs_17__0 ;
    output outputs_16__15 ;
    output outputs_16__14 ;
    output outputs_16__13 ;
    output outputs_16__12 ;
    output outputs_16__11 ;
    output outputs_16__10 ;
    output outputs_16__9 ;
    output outputs_16__8 ;
    output outputs_16__7 ;
    output outputs_16__6 ;
    output outputs_16__5 ;
    output outputs_16__4 ;
    output outputs_16__3 ;
    output outputs_16__2 ;
    output outputs_16__1 ;
    output outputs_16__0 ;
    output outputs_15__15 ;
    output outputs_15__14 ;
    output outputs_15__13 ;
    output outputs_15__12 ;
    output outputs_15__11 ;
    output outputs_15__10 ;
    output outputs_15__9 ;
    output outputs_15__8 ;
    output outputs_15__7 ;
    output outputs_15__6 ;
    output outputs_15__5 ;
    output outputs_15__4 ;
    output outputs_15__3 ;
    output outputs_15__2 ;
    output outputs_15__1 ;
    output outputs_15__0 ;
    output outputs_14__15 ;
    output outputs_14__14 ;
    output outputs_14__13 ;
    output outputs_14__12 ;
    output outputs_14__11 ;
    output outputs_14__10 ;
    output outputs_14__9 ;
    output outputs_14__8 ;
    output outputs_14__7 ;
    output outputs_14__6 ;
    output outputs_14__5 ;
    output outputs_14__4 ;
    output outputs_14__3 ;
    output outputs_14__2 ;
    output outputs_14__1 ;
    output outputs_14__0 ;
    output outputs_13__15 ;
    output outputs_13__14 ;
    output outputs_13__13 ;
    output outputs_13__12 ;
    output outputs_13__11 ;
    output outputs_13__10 ;
    output outputs_13__9 ;
    output outputs_13__8 ;
    output outputs_13__7 ;
    output outputs_13__6 ;
    output outputs_13__5 ;
    output outputs_13__4 ;
    output outputs_13__3 ;
    output outputs_13__2 ;
    output outputs_13__1 ;
    output outputs_13__0 ;
    output outputs_12__15 ;
    output outputs_12__14 ;
    output outputs_12__13 ;
    output outputs_12__12 ;
    output outputs_12__11 ;
    output outputs_12__10 ;
    output outputs_12__9 ;
    output outputs_12__8 ;
    output outputs_12__7 ;
    output outputs_12__6 ;
    output outputs_12__5 ;
    output outputs_12__4 ;
    output outputs_12__3 ;
    output outputs_12__2 ;
    output outputs_12__1 ;
    output outputs_12__0 ;
    output outputs_11__15 ;
    output outputs_11__14 ;
    output outputs_11__13 ;
    output outputs_11__12 ;
    output outputs_11__11 ;
    output outputs_11__10 ;
    output outputs_11__9 ;
    output outputs_11__8 ;
    output outputs_11__7 ;
    output outputs_11__6 ;
    output outputs_11__5 ;
    output outputs_11__4 ;
    output outputs_11__3 ;
    output outputs_11__2 ;
    output outputs_11__1 ;
    output outputs_11__0 ;
    output outputs_10__15 ;
    output outputs_10__14 ;
    output outputs_10__13 ;
    output outputs_10__12 ;
    output outputs_10__11 ;
    output outputs_10__10 ;
    output outputs_10__9 ;
    output outputs_10__8 ;
    output outputs_10__7 ;
    output outputs_10__6 ;
    output outputs_10__5 ;
    output outputs_10__4 ;
    output outputs_10__3 ;
    output outputs_10__2 ;
    output outputs_10__1 ;
    output outputs_10__0 ;
    output outputs_9__15 ;
    output outputs_9__14 ;
    output outputs_9__13 ;
    output outputs_9__12 ;
    output outputs_9__11 ;
    output outputs_9__10 ;
    output outputs_9__9 ;
    output outputs_9__8 ;
    output outputs_9__7 ;
    output outputs_9__6 ;
    output outputs_9__5 ;
    output outputs_9__4 ;
    output outputs_9__3 ;
    output outputs_9__2 ;
    output outputs_9__1 ;
    output outputs_9__0 ;
    output outputs_8__15 ;
    output outputs_8__14 ;
    output outputs_8__13 ;
    output outputs_8__12 ;
    output outputs_8__11 ;
    output outputs_8__10 ;
    output outputs_8__9 ;
    output outputs_8__8 ;
    output outputs_8__7 ;
    output outputs_8__6 ;
    output outputs_8__5 ;
    output outputs_8__4 ;
    output outputs_8__3 ;
    output outputs_8__2 ;
    output outputs_8__1 ;
    output outputs_8__0 ;
    output outputs_7__15 ;
    output outputs_7__14 ;
    output outputs_7__13 ;
    output outputs_7__12 ;
    output outputs_7__11 ;
    output outputs_7__10 ;
    output outputs_7__9 ;
    output outputs_7__8 ;
    output outputs_7__7 ;
    output outputs_7__6 ;
    output outputs_7__5 ;
    output outputs_7__4 ;
    output outputs_7__3 ;
    output outputs_7__2 ;
    output outputs_7__1 ;
    output outputs_7__0 ;
    output outputs_6__15 ;
    output outputs_6__14 ;
    output outputs_6__13 ;
    output outputs_6__12 ;
    output outputs_6__11 ;
    output outputs_6__10 ;
    output outputs_6__9 ;
    output outputs_6__8 ;
    output outputs_6__7 ;
    output outputs_6__6 ;
    output outputs_6__5 ;
    output outputs_6__4 ;
    output outputs_6__3 ;
    output outputs_6__2 ;
    output outputs_6__1 ;
    output outputs_6__0 ;
    output outputs_5__15 ;
    output outputs_5__14 ;
    output outputs_5__13 ;
    output outputs_5__12 ;
    output outputs_5__11 ;
    output outputs_5__10 ;
    output outputs_5__9 ;
    output outputs_5__8 ;
    output outputs_5__7 ;
    output outputs_5__6 ;
    output outputs_5__5 ;
    output outputs_5__4 ;
    output outputs_5__3 ;
    output outputs_5__2 ;
    output outputs_5__1 ;
    output outputs_5__0 ;
    output outputs_4__15 ;
    output outputs_4__14 ;
    output outputs_4__13 ;
    output outputs_4__12 ;
    output outputs_4__11 ;
    output outputs_4__10 ;
    output outputs_4__9 ;
    output outputs_4__8 ;
    output outputs_4__7 ;
    output outputs_4__6 ;
    output outputs_4__5 ;
    output outputs_4__4 ;
    output outputs_4__3 ;
    output outputs_4__2 ;
    output outputs_4__1 ;
    output outputs_4__0 ;
    output outputs_3__15 ;
    output outputs_3__14 ;
    output outputs_3__13 ;
    output outputs_3__12 ;
    output outputs_3__11 ;
    output outputs_3__10 ;
    output outputs_3__9 ;
    output outputs_3__8 ;
    output outputs_3__7 ;
    output outputs_3__6 ;
    output outputs_3__5 ;
    output outputs_3__4 ;
    output outputs_3__3 ;
    output outputs_3__2 ;
    output outputs_3__1 ;
    output outputs_3__0 ;
    output outputs_2__15 ;
    output outputs_2__14 ;
    output outputs_2__13 ;
    output outputs_2__12 ;
    output outputs_2__11 ;
    output outputs_2__10 ;
    output outputs_2__9 ;
    output outputs_2__8 ;
    output outputs_2__7 ;
    output outputs_2__6 ;
    output outputs_2__5 ;
    output outputs_2__4 ;
    output outputs_2__3 ;
    output outputs_2__2 ;
    output outputs_2__1 ;
    output outputs_2__0 ;
    output outputs_1__15 ;
    output outputs_1__14 ;
    output outputs_1__13 ;
    output outputs_1__12 ;
    output outputs_1__11 ;
    output outputs_1__10 ;
    output outputs_1__9 ;
    output outputs_1__8 ;
    output outputs_1__7 ;
    output outputs_1__6 ;
    output outputs_1__5 ;
    output outputs_1__4 ;
    output outputs_1__3 ;
    output outputs_1__2 ;
    output outputs_1__1 ;
    output outputs_1__0 ;
    output outputs_0__15 ;
    output outputs_0__14 ;
    output outputs_0__13 ;
    output outputs_0__12 ;
    output outputs_0__11 ;
    output outputs_0__10 ;
    output outputs_0__9 ;
    output outputs_0__8 ;
    output outputs_0__7 ;
    output outputs_0__6 ;
    output outputs_0__5 ;
    output outputs_0__4 ;
    output outputs_0__3 ;
    output outputs_0__2 ;
    output outputs_0__1 ;
    output outputs_0__0 ;
    input clk ;
    input start ;
    input rst ;
    output doneOut ;
    output workingOut ;

    wire counter_0, counterRst, restartDetection, firstStart, PWR, nx843, nx845, 
         nx847, nx849, nx851, nx853, nx855, nx857, nx859, nx861, nx863, nx865, 
         nx867, nx869, nx871, nx877, nx879, nx881, nx883, nx885;
    wire [1:0] \$dummy ;




    Mul8x16 gen_24_cmp (.q ({filter_24__7,filter_24__6,filter_24__5,filter_24__4
            ,filter_24__3,filter_24__2,filter_24__1,filter_24__0}), .m ({
            window_24__15,window_24__14,window_24__13,window_24__12,
            window_24__11,window_24__10,window_24__9,window_24__8,window_24__7,
            window_24__6,window_24__5,window_24__4,window_24__3,window_24__2,
            window_24__1,window_24__0}), .f ({outputs_24__15,outputs_24__14,
            outputs_24__13,outputs_24__12,outputs_24__11,outputs_24__10,
            outputs_24__9,outputs_24__8,outputs_24__7,outputs_24__6,
            outputs_24__5,outputs_24__4,outputs_24__3,outputs_24__2,
            outputs_24__1,outputs_24__0}), .clk (nx865), .start (nx879), .rst (
            rst), .sel (nx857), .startAndPause (nx845)) ;
    Mul8x16 gen_23_cmp (.q ({filter_23__7,filter_23__6,filter_23__5,filter_23__4
            ,filter_23__3,filter_23__2,filter_23__1,filter_23__0}), .m ({
            window_23__15,window_23__14,window_23__13,window_23__12,
            window_23__11,window_23__10,window_23__9,window_23__8,window_23__7,
            window_23__6,window_23__5,window_23__4,window_23__3,window_23__2,
            window_23__1,window_23__0}), .f ({outputs_23__15,outputs_23__14,
            outputs_23__13,outputs_23__12,outputs_23__11,outputs_23__10,
            outputs_23__9,outputs_23__8,outputs_23__7,outputs_23__6,
            outputs_23__5,outputs_23__4,outputs_23__3,outputs_23__2,
            outputs_23__1,outputs_23__0}), .clk (nx865), .start (nx879), .rst (
            rst), .sel (nx857), .startAndPause (nx845)) ;
    Mul8x16 gen_22_cmp (.q ({filter_22__7,filter_22__6,filter_22__5,filter_22__4
            ,filter_22__3,filter_22__2,filter_22__1,filter_22__0}), .m ({
            window_22__15,window_22__14,window_22__13,window_22__12,
            window_22__11,window_22__10,window_22__9,window_22__8,window_22__7,
            window_22__6,window_22__5,window_22__4,window_22__3,window_22__2,
            window_22__1,window_22__0}), .f ({outputs_22__15,outputs_22__14,
            outputs_22__13,outputs_22__12,outputs_22__11,outputs_22__10,
            outputs_22__9,outputs_22__8,outputs_22__7,outputs_22__6,
            outputs_22__5,outputs_22__4,outputs_22__3,outputs_22__2,
            outputs_22__1,outputs_22__0}), .clk (nx865), .start (nx879), .rst (
            rst), .sel (nx857), .startAndPause (nx845)) ;
    Mul8x16 gen_21_cmp (.q ({filter_21__7,filter_21__6,filter_21__5,filter_21__4
            ,filter_21__3,filter_21__2,filter_21__1,filter_21__0}), .m ({
            window_21__15,window_21__14,window_21__13,window_21__12,
            window_21__11,window_21__10,window_21__9,window_21__8,window_21__7,
            window_21__6,window_21__5,window_21__4,window_21__3,window_21__2,
            window_21__1,window_21__0}), .f ({outputs_21__15,outputs_21__14,
            outputs_21__13,outputs_21__12,outputs_21__11,outputs_21__10,
            outputs_21__9,outputs_21__8,outputs_21__7,outputs_21__6,
            outputs_21__5,outputs_21__4,outputs_21__3,outputs_21__2,
            outputs_21__1,outputs_21__0}), .clk (nx865), .start (nx879), .rst (
            rst), .sel (nx857), .startAndPause (nx845)) ;
    Mul8x16 gen_20_cmp (.q ({filter_20__7,filter_20__6,filter_20__5,filter_20__4
            ,filter_20__3,filter_20__2,filter_20__1,filter_20__0}), .m ({
            window_20__15,window_20__14,window_20__13,window_20__12,
            window_20__11,window_20__10,window_20__9,window_20__8,window_20__7,
            window_20__6,window_20__5,window_20__4,window_20__3,window_20__2,
            window_20__1,window_20__0}), .f ({outputs_20__15,outputs_20__14,
            outputs_20__13,outputs_20__12,outputs_20__11,outputs_20__10,
            outputs_20__9,outputs_20__8,outputs_20__7,outputs_20__6,
            outputs_20__5,outputs_20__4,outputs_20__3,outputs_20__2,
            outputs_20__1,outputs_20__0}), .clk (nx865), .start (nx879), .rst (
            rst), .sel (nx857), .startAndPause (nx845)) ;
    Mul8x16 gen_19_cmp (.q ({filter_19__7,filter_19__6,filter_19__5,filter_19__4
            ,filter_19__3,filter_19__2,filter_19__1,filter_19__0}), .m ({
            window_19__15,window_19__14,window_19__13,window_19__12,
            window_19__11,window_19__10,window_19__9,window_19__8,window_19__7,
            window_19__6,window_19__5,window_19__4,window_19__3,window_19__2,
            window_19__1,window_19__0}), .f ({outputs_19__15,outputs_19__14,
            outputs_19__13,outputs_19__12,outputs_19__11,outputs_19__10,
            outputs_19__9,outputs_19__8,outputs_19__7,outputs_19__6,
            outputs_19__5,outputs_19__4,outputs_19__3,outputs_19__2,
            outputs_19__1,outputs_19__0}), .clk (nx865), .start (nx879), .rst (
            rst), .sel (nx857), .startAndPause (nx845)) ;
    Mul8x16 gen_18_cmp (.q ({filter_18__7,filter_18__6,filter_18__5,filter_18__4
            ,filter_18__3,filter_18__2,filter_18__1,filter_18__0}), .m ({
            window_18__15,window_18__14,window_18__13,window_18__12,
            window_18__11,window_18__10,window_18__9,window_18__8,window_18__7,
            window_18__6,window_18__5,window_18__4,window_18__3,window_18__2,
            window_18__1,window_18__0}), .f ({outputs_18__15,outputs_18__14,
            outputs_18__13,outputs_18__12,outputs_18__11,outputs_18__10,
            outputs_18__9,outputs_18__8,outputs_18__7,outputs_18__6,
            outputs_18__5,outputs_18__4,outputs_18__3,outputs_18__2,
            outputs_18__1,outputs_18__0}), .clk (nx865), .start (nx879), .rst (
            rst), .sel (nx857), .startAndPause (nx845)) ;
    Mul8x16 gen_17_cmp (.q ({filter_17__7,filter_17__6,filter_17__5,filter_17__4
            ,filter_17__3,filter_17__2,filter_17__1,filter_17__0}), .m ({
            window_17__15,window_17__14,window_17__13,window_17__12,
            window_17__11,window_17__10,window_17__9,window_17__8,window_17__7,
            window_17__6,window_17__5,window_17__4,window_17__3,window_17__2,
            window_17__1,window_17__0}), .f ({outputs_17__15,outputs_17__14,
            outputs_17__13,outputs_17__12,outputs_17__11,outputs_17__10,
            outputs_17__9,outputs_17__8,outputs_17__7,outputs_17__6,
            outputs_17__5,outputs_17__4,outputs_17__3,outputs_17__2,
            outputs_17__1,outputs_17__0}), .clk (nx867), .start (nx881), .rst (
            rst), .sel (nx859), .startAndPause (nx847)) ;
    Mul8x16 gen_16_cmp (.q ({filter_16__7,filter_16__6,filter_16__5,filter_16__4
            ,filter_16__3,filter_16__2,filter_16__1,filter_16__0}), .m ({
            window_16__15,window_16__14,window_16__13,window_16__12,
            window_16__11,window_16__10,window_16__9,window_16__8,window_16__7,
            window_16__6,window_16__5,window_16__4,window_16__3,window_16__2,
            window_16__1,window_16__0}), .f ({outputs_16__15,outputs_16__14,
            outputs_16__13,outputs_16__12,outputs_16__11,outputs_16__10,
            outputs_16__9,outputs_16__8,outputs_16__7,outputs_16__6,
            outputs_16__5,outputs_16__4,outputs_16__3,outputs_16__2,
            outputs_16__1,outputs_16__0}), .clk (nx867), .start (nx881), .rst (
            rst), .sel (nx859), .startAndPause (nx847)) ;
    Mul8x16 gen_15_cmp (.q ({filter_15__7,filter_15__6,filter_15__5,filter_15__4
            ,filter_15__3,filter_15__2,filter_15__1,filter_15__0}), .m ({
            window_15__15,window_15__14,window_15__13,window_15__12,
            window_15__11,window_15__10,window_15__9,window_15__8,window_15__7,
            window_15__6,window_15__5,window_15__4,window_15__3,window_15__2,
            window_15__1,window_15__0}), .f ({outputs_15__15,outputs_15__14,
            outputs_15__13,outputs_15__12,outputs_15__11,outputs_15__10,
            outputs_15__9,outputs_15__8,outputs_15__7,outputs_15__6,
            outputs_15__5,outputs_15__4,outputs_15__3,outputs_15__2,
            outputs_15__1,outputs_15__0}), .clk (nx867), .start (nx881), .rst (
            rst), .sel (nx859), .startAndPause (nx847)) ;
    Mul8x16 gen_14_cmp (.q ({filter_14__7,filter_14__6,filter_14__5,filter_14__4
            ,filter_14__3,filter_14__2,filter_14__1,filter_14__0}), .m ({
            window_14__15,window_14__14,window_14__13,window_14__12,
            window_14__11,window_14__10,window_14__9,window_14__8,window_14__7,
            window_14__6,window_14__5,window_14__4,window_14__3,window_14__2,
            window_14__1,window_14__0}), .f ({outputs_14__15,outputs_14__14,
            outputs_14__13,outputs_14__12,outputs_14__11,outputs_14__10,
            outputs_14__9,outputs_14__8,outputs_14__7,outputs_14__6,
            outputs_14__5,outputs_14__4,outputs_14__3,outputs_14__2,
            outputs_14__1,outputs_14__0}), .clk (nx867), .start (nx881), .rst (
            rst), .sel (nx859), .startAndPause (nx847)) ;
    Mul8x16 gen_13_cmp (.q ({filter_13__7,filter_13__6,filter_13__5,filter_13__4
            ,filter_13__3,filter_13__2,filter_13__1,filter_13__0}), .m ({
            window_13__15,window_13__14,window_13__13,window_13__12,
            window_13__11,window_13__10,window_13__9,window_13__8,window_13__7,
            window_13__6,window_13__5,window_13__4,window_13__3,window_13__2,
            window_13__1,window_13__0}), .f ({outputs_13__15,outputs_13__14,
            outputs_13__13,outputs_13__12,outputs_13__11,outputs_13__10,
            outputs_13__9,outputs_13__8,outputs_13__7,outputs_13__6,
            outputs_13__5,outputs_13__4,outputs_13__3,outputs_13__2,
            outputs_13__1,outputs_13__0}), .clk (nx867), .start (nx881), .rst (
            rst), .sel (nx859), .startAndPause (nx847)) ;
    Mul8x16 gen_12_cmp (.q ({filter_12__7,filter_12__6,filter_12__5,filter_12__4
            ,filter_12__3,filter_12__2,filter_12__1,filter_12__0}), .m ({
            window_12__15,window_12__14,window_12__13,window_12__12,
            window_12__11,window_12__10,window_12__9,window_12__8,window_12__7,
            window_12__6,window_12__5,window_12__4,window_12__3,window_12__2,
            window_12__1,window_12__0}), .f ({outputs_12__15,outputs_12__14,
            outputs_12__13,outputs_12__12,outputs_12__11,outputs_12__10,
            outputs_12__9,outputs_12__8,outputs_12__7,outputs_12__6,
            outputs_12__5,outputs_12__4,outputs_12__3,outputs_12__2,
            outputs_12__1,outputs_12__0}), .clk (nx867), .start (nx881), .rst (
            rst), .sel (nx859), .startAndPause (nx847)) ;
    Mul8x16 gen_11_cmp (.q ({filter_11__7,filter_11__6,filter_11__5,filter_11__4
            ,filter_11__3,filter_11__2,filter_11__1,filter_11__0}), .m ({
            window_11__15,window_11__14,window_11__13,window_11__12,
            window_11__11,window_11__10,window_11__9,window_11__8,window_11__7,
            window_11__6,window_11__5,window_11__4,window_11__3,window_11__2,
            window_11__1,window_11__0}), .f ({outputs_11__15,outputs_11__14,
            outputs_11__13,outputs_11__12,outputs_11__11,outputs_11__10,
            outputs_11__9,outputs_11__8,outputs_11__7,outputs_11__6,
            outputs_11__5,outputs_11__4,outputs_11__3,outputs_11__2,
            outputs_11__1,outputs_11__0}), .clk (nx867), .start (nx881), .rst (
            rst), .sel (nx859), .startAndPause (nx847)) ;
    Mul8x16 gen_10_cmp (.q ({filter_10__7,filter_10__6,filter_10__5,filter_10__4
            ,filter_10__3,filter_10__2,filter_10__1,filter_10__0}), .m ({
            window_10__15,window_10__14,window_10__13,window_10__12,
            window_10__11,window_10__10,window_10__9,window_10__8,window_10__7,
            window_10__6,window_10__5,window_10__4,window_10__3,window_10__2,
            window_10__1,window_10__0}), .f ({outputs_10__15,outputs_10__14,
            outputs_10__13,outputs_10__12,outputs_10__11,outputs_10__10,
            outputs_10__9,outputs_10__8,outputs_10__7,outputs_10__6,
            outputs_10__5,outputs_10__4,outputs_10__3,outputs_10__2,
            outputs_10__1,outputs_10__0}), .clk (nx869), .start (nx883), .rst (
            rst), .sel (nx861), .startAndPause (nx849)) ;
    Mul8x16 gen_9_cmp (.q ({filter_9__7,filter_9__6,filter_9__5,filter_9__4,
            filter_9__3,filter_9__2,filter_9__1,filter_9__0}), .m ({window_9__15
            ,window_9__14,window_9__13,window_9__12,window_9__11,window_9__10,
            window_9__9,window_9__8,window_9__7,window_9__6,window_9__5,
            window_9__4,window_9__3,window_9__2,window_9__1,window_9__0}), .f ({
            outputs_9__15,outputs_9__14,outputs_9__13,outputs_9__12,
            outputs_9__11,outputs_9__10,outputs_9__9,outputs_9__8,outputs_9__7,
            outputs_9__6,outputs_9__5,outputs_9__4,outputs_9__3,outputs_9__2,
            outputs_9__1,outputs_9__0}), .clk (nx869), .start (nx883), .rst (rst
            ), .sel (nx861), .startAndPause (nx849)) ;
    Mul8x16 gen_8_cmp (.q ({filter_8__7,filter_8__6,filter_8__5,filter_8__4,
            filter_8__3,filter_8__2,filter_8__1,filter_8__0}), .m ({window_8__15
            ,window_8__14,window_8__13,window_8__12,window_8__11,window_8__10,
            window_8__9,window_8__8,window_8__7,window_8__6,window_8__5,
            window_8__4,window_8__3,window_8__2,window_8__1,window_8__0}), .f ({
            outputs_8__15,outputs_8__14,outputs_8__13,outputs_8__12,
            outputs_8__11,outputs_8__10,outputs_8__9,outputs_8__8,outputs_8__7,
            outputs_8__6,outputs_8__5,outputs_8__4,outputs_8__3,outputs_8__2,
            outputs_8__1,outputs_8__0}), .clk (nx869), .start (nx883), .rst (rst
            ), .sel (nx861), .startAndPause (nx849)) ;
    Mul8x16 gen_7_cmp (.q ({filter_7__7,filter_7__6,filter_7__5,filter_7__4,
            filter_7__3,filter_7__2,filter_7__1,filter_7__0}), .m ({window_7__15
            ,window_7__14,window_7__13,window_7__12,window_7__11,window_7__10,
            window_7__9,window_7__8,window_7__7,window_7__6,window_7__5,
            window_7__4,window_7__3,window_7__2,window_7__1,window_7__0}), .f ({
            outputs_7__15,outputs_7__14,outputs_7__13,outputs_7__12,
            outputs_7__11,outputs_7__10,outputs_7__9,outputs_7__8,outputs_7__7,
            outputs_7__6,outputs_7__5,outputs_7__4,outputs_7__3,outputs_7__2,
            outputs_7__1,outputs_7__0}), .clk (nx869), .start (nx883), .rst (rst
            ), .sel (nx861), .startAndPause (nx849)) ;
    Mul8x16 gen_6_cmp (.q ({filter_6__7,filter_6__6,filter_6__5,filter_6__4,
            filter_6__3,filter_6__2,filter_6__1,filter_6__0}), .m ({window_6__15
            ,window_6__14,window_6__13,window_6__12,window_6__11,window_6__10,
            window_6__9,window_6__8,window_6__7,window_6__6,window_6__5,
            window_6__4,window_6__3,window_6__2,window_6__1,window_6__0}), .f ({
            outputs_6__15,outputs_6__14,outputs_6__13,outputs_6__12,
            outputs_6__11,outputs_6__10,outputs_6__9,outputs_6__8,outputs_6__7,
            outputs_6__6,outputs_6__5,outputs_6__4,outputs_6__3,outputs_6__2,
            outputs_6__1,outputs_6__0}), .clk (nx869), .start (nx883), .rst (rst
            ), .sel (nx861), .startAndPause (nx849)) ;
    Mul8x16 gen_5_cmp (.q ({filter_5__7,filter_5__6,filter_5__5,filter_5__4,
            filter_5__3,filter_5__2,filter_5__1,filter_5__0}), .m ({window_5__15
            ,window_5__14,window_5__13,window_5__12,window_5__11,window_5__10,
            window_5__9,window_5__8,window_5__7,window_5__6,window_5__5,
            window_5__4,window_5__3,window_5__2,window_5__1,window_5__0}), .f ({
            outputs_5__15,outputs_5__14,outputs_5__13,outputs_5__12,
            outputs_5__11,outputs_5__10,outputs_5__9,outputs_5__8,outputs_5__7,
            outputs_5__6,outputs_5__5,outputs_5__4,outputs_5__3,outputs_5__2,
            outputs_5__1,outputs_5__0}), .clk (nx869), .start (nx883), .rst (rst
            ), .sel (nx861), .startAndPause (nx849)) ;
    Mul8x16 gen_4_cmp (.q ({filter_4__7,filter_4__6,filter_4__5,filter_4__4,
            filter_4__3,filter_4__2,filter_4__1,filter_4__0}), .m ({window_4__15
            ,window_4__14,window_4__13,window_4__12,window_4__11,window_4__10,
            window_4__9,window_4__8,window_4__7,window_4__6,window_4__5,
            window_4__4,window_4__3,window_4__2,window_4__1,window_4__0}), .f ({
            outputs_4__15,outputs_4__14,outputs_4__13,outputs_4__12,
            outputs_4__11,outputs_4__10,outputs_4__9,outputs_4__8,outputs_4__7,
            outputs_4__6,outputs_4__5,outputs_4__4,outputs_4__3,outputs_4__2,
            outputs_4__1,outputs_4__0}), .clk (nx869), .start (nx883), .rst (rst
            ), .sel (nx861), .startAndPause (nx849)) ;
    Mul8x16 gen_3_cmp (.q ({filter_3__7,filter_3__6,filter_3__5,filter_3__4,
            filter_3__3,filter_3__2,filter_3__1,filter_3__0}), .m ({window_3__15
            ,window_3__14,window_3__13,window_3__12,window_3__11,window_3__10,
            window_3__9,window_3__8,window_3__7,window_3__6,window_3__5,
            window_3__4,window_3__3,window_3__2,window_3__1,window_3__0}), .f ({
            outputs_3__15,outputs_3__14,outputs_3__13,outputs_3__12,
            outputs_3__11,outputs_3__10,outputs_3__9,outputs_3__8,outputs_3__7,
            outputs_3__6,outputs_3__5,outputs_3__4,outputs_3__3,outputs_3__2,
            outputs_3__1,outputs_3__0}), .clk (nx871), .start (nx885), .rst (rst
            ), .sel (nx863), .startAndPause (nx851)) ;
    Mul8x16 gen_2_cmp (.q ({filter_2__7,filter_2__6,filter_2__5,filter_2__4,
            filter_2__3,filter_2__2,filter_2__1,filter_2__0}), .m ({window_2__15
            ,window_2__14,window_2__13,window_2__12,window_2__11,window_2__10,
            window_2__9,window_2__8,window_2__7,window_2__6,window_2__5,
            window_2__4,window_2__3,window_2__2,window_2__1,window_2__0}), .f ({
            outputs_2__15,outputs_2__14,outputs_2__13,outputs_2__12,
            outputs_2__11,outputs_2__10,outputs_2__9,outputs_2__8,outputs_2__7,
            outputs_2__6,outputs_2__5,outputs_2__4,outputs_2__3,outputs_2__2,
            outputs_2__1,outputs_2__0}), .clk (nx871), .start (nx885), .rst (rst
            ), .sel (nx863), .startAndPause (nx851)) ;
    Mul8x16 gen_1_cmp (.q ({filter_1__7,filter_1__6,filter_1__5,filter_1__4,
            filter_1__3,filter_1__2,filter_1__1,filter_1__0}), .m ({window_1__15
            ,window_1__14,window_1__13,window_1__12,window_1__11,window_1__10,
            window_1__9,window_1__8,window_1__7,window_1__6,window_1__5,
            window_1__4,window_1__3,window_1__2,window_1__1,window_1__0}), .f ({
            outputs_1__15,outputs_1__14,outputs_1__13,outputs_1__12,
            outputs_1__11,outputs_1__10,outputs_1__9,outputs_1__8,outputs_1__7,
            outputs_1__6,outputs_1__5,outputs_1__4,outputs_1__3,outputs_1__2,
            outputs_1__1,outputs_1__0}), .clk (nx871), .start (nx885), .rst (rst
            ), .sel (nx863), .startAndPause (nx851)) ;
    Mul8x16 gen_0_cmp (.q ({filter_0__7,filter_0__6,filter_0__5,filter_0__4,
            filter_0__3,filter_0__2,filter_0__1,filter_0__0}), .m ({window_0__15
            ,window_0__14,window_0__13,window_0__12,window_0__11,window_0__10,
            window_0__9,window_0__8,window_0__7,window_0__6,window_0__5,
            window_0__4,window_0__3,window_0__2,window_0__1,window_0__0}), .f ({
            outputs_0__15,outputs_0__14,outputs_0__13,outputs_0__12,
            outputs_0__11,outputs_0__10,outputs_0__9,outputs_0__8,outputs_0__7,
            outputs_0__6,outputs_0__5,outputs_0__4,outputs_0__3,outputs_0__2,
            outputs_0__1,outputs_0__0}), .clk (nx871), .start (nx885), .rst (rst
            ), .sel (nx863), .startAndPause (nx851)) ;
    TransitionDetector StartCaptuerCmp (.edge (nx885), .clk (clk), .rst (rst), .f (
                       restartDetection)) ;
    ShiftReg_3 CounterCmp (.outp ({doneOut,\$dummy [0],\$dummy [1],counter_0}), 
               .clk (clk), .en (nx853), .rst (counterRst)) ;
    Reg_1 firtStartLachCmp (.D ({PWR}), .en (PWR), .clk (nx885), .rst (rst), .Q (
          {firstStart})) ;
    fake_vcc ix822 (.Y (PWR)) ;
    or02 ix3 (.Y (counterRst), .A0 (rst), .A1 (restartDetection)) ;
    nor02ii ix7 (.Y (workingOut), .A0 (doneOut), .A1 (firstStart)) ;
    inv01 ix842 (.Y (nx843), .A (workingOut)) ;
    inv01 ix844 (.Y (nx845), .A (nx843)) ;
    inv01 ix846 (.Y (nx847), .A (nx843)) ;
    inv01 ix848 (.Y (nx849), .A (nx843)) ;
    inv01 ix850 (.Y (nx851), .A (nx843)) ;
    inv01 ix852 (.Y (nx853), .A (nx843)) ;
    inv01 ix854 (.Y (nx855), .A (counter_0)) ;
    inv01 ix856 (.Y (nx857), .A (nx855)) ;
    inv01 ix858 (.Y (nx859), .A (nx855)) ;
    inv01 ix860 (.Y (nx861), .A (nx855)) ;
    inv01 ix862 (.Y (nx863), .A (nx855)) ;
    inv01 ix864 (.Y (nx865), .A (clk)) ;
    inv01 ix866 (.Y (nx867), .A (clk)) ;
    inv01 ix868 (.Y (nx869), .A (clk)) ;
    inv01 ix870 (.Y (nx871), .A (clk)) ;
    inv01 ix876 (.Y (nx877), .A (start)) ;
    inv01 ix878 (.Y (nx879), .A (nx877)) ;
    inv01 ix880 (.Y (nx881), .A (nx877)) ;
    inv01 ix882 (.Y (nx883), .A (nx877)) ;
    inv01 ix884 (.Y (nx885), .A (nx877)) ;
endmodule


module Reg_1 ( D, en, clk, rst, Q ) ;

    input [0:0]D ;
    input en ;
    input clk ;
    input rst ;
    output [0:0]Q ;

    wire nx48;
    wire [0:0] \$dummy ;




    dffr reg_Q_0 (.Q (Q[0]), .QB (\$dummy [0]), .D (nx48), .CLK (clk), .R (rst)
         ) ;
    mux21_ni ix49 (.Y (nx48), .A0 (Q[0]), .A1 (D[0]), .S0 (en)) ;
endmodule


module ShiftReg_3 ( outp, clk, en, rst ) ;

    inout [3:0]outp ;
    input clk ;
    input en ;
    input rst ;

    wire nx80, nx94, nx104, nx114;
    wire [3:0] \$dummy ;




    dffs_ni reg_outp_0 (.Q (outp[0]), .QB (\$dummy [0]), .D (nx80), .CLK (clk), 
            .S (rst)) ;
    nor02ii ix81 (.Y (nx80), .A0 (en), .A1 (outp[0])) ;
    dffr reg_outp_1 (.Q (outp[1]), .QB (\$dummy [1]), .D (nx94), .CLK (clk), .R (
         rst)) ;
    mux21_ni ix95 (.Y (nx94), .A0 (outp[1]), .A1 (outp[0]), .S0 (en)) ;
    dffr reg_outp_2 (.Q (outp[2]), .QB (\$dummy [2]), .D (nx104), .CLK (clk), .R (
         rst)) ;
    mux21_ni ix105 (.Y (nx104), .A0 (outp[2]), .A1 (outp[1]), .S0 (en)) ;
    dffr reg_outp_3 (.Q (outp[3]), .QB (\$dummy [3]), .D (nx114), .CLK (clk), .R (
         rst)) ;
    mux21_ni ix115 (.Y (nx114), .A0 (outp[3]), .A1 (outp[2]), .S0 (en)) ;
endmodule


module TransitionDetector ( edge, clk, rst, f ) ;

    input edge ;
    input clk ;
    input rst ;
    inout f ;

    wire nx0, d, NOT_clk, nx10;
    wire [1:0] \$dummy ;




    fake_vcc ix1 (.Y (nx0)) ;
    dffr reg_f (.Q (f), .QB (\$dummy [0]), .D (nx0), .CLK (edge), .R (nx10)) ;
    or02 ix11 (.Y (nx10), .A0 (d), .A1 (rst)) ;
    dff reg_d (.Q (d), .QB (\$dummy [1]), .D (f), .CLK (NOT_clk)) ;
    inv01 ix31 (.Y (NOT_clk), .A (clk)) ;
endmodule


module Mul8x16 ( q, m, f, clk, start, rst, sel, startAndPause ) ;

    input [7:0]q ;
    input [15:0]m ;
    output [15:0]f ;
    input clk ;
    input start ;
    input rst ;
    input sel ;
    input startAndPause ;

    wire pBs_32, pBs_30, pBs_29, pBs_28, pBs_27, pBs_26, pBs_25, pBs_24, pBs_23, 
         pMux_32, pMux_31, pMux_30, pMux_29, pMux_28, pMux_27, pMux_26, pMux_25, 
         pMux_24, pMux_23, pMux_22, pMux_21, pMux_20, pMux_19, pMux_18, pMux_17, 
         pMux_16, pMux_15, pMux_14, pMux_13, pMux_12, pMux_11, pMux_10, pMux_9, 
         pMux_8, pMux_7, pMux_6, pMux_5, pMux_4, pMux_3, pMux_2, pMux_1, pMux_0, 
         pReg_32, pReg_31, pReg_30, pReg_29, pReg_28, pReg_27, pReg_26, pReg_25, 
         pReg_24, pReg_23, pReg_22, pReg_21, pReg_20, pReg_19, pReg_18, pReg_17, 
         pReg_16, pReg_15, pReg_14, pReg_13, pReg_12, pReg_11, pReg_10, pReg_9, 
         pReg_8, pReg_7, pReg_6, pReg_5, pReg_4, pReg_3, pReg_2, pReg_1, pReg_0, 
         mReg_15, mReg_14, mReg_13, mReg_12, mReg_11, mReg_10, mReg_9, mReg_8, 
         mReg_7, mReg_6, mReg_5, mReg_4, mReg_3, mReg_2, mReg_1, mReg_0, PWR, 
         pInit_32, nx196, nx198, nx200, nx202, nx204, nx206, nx208, nx210, nx212
         ;
    wire [7:0] \$dummy ;




    Reg_33 pRegCmp (.D ({pBs_32,pBs_32,pBs_30,pBs_29,pBs_28,pBs_27,pBs_26,pBs_25
           ,pBs_24,pBs_23,f[15],f[14],f[13],f[12],f[11],f[10],f[9],f[8],f[7],
           f[6],f[5],f[4],f[3],f[2],f[1],f[0],pMux_8,pMux_7,pMux_6,pMux_5,pMux_4
           ,pMux_3,pMux_2}), .en (startAndPause), .clk (clk), .rst (rst), .Q ({
           pReg_32,pReg_31,pReg_30,pReg_29,pReg_28,pReg_27,pReg_26,pReg_25,
           pReg_24,pReg_23,pReg_22,pReg_21,pReg_20,pReg_19,pReg_18,pReg_17,
           pReg_16,pReg_15,pReg_14,pReg_13,pReg_12,pReg_11,pReg_10,pReg_9,pReg_8
           ,pReg_7,pReg_6,pReg_5,pReg_4,pReg_3,pReg_2,pReg_1,pReg_0})) ;
    Reg_16 mRegCmp (.D ({m[15],m[14],m[13],m[12],m[11],m[10],m[9],m[8],m[7],m[6]
           ,m[5],m[4],m[3],m[2],m[1],m[0]}), .en (PWR), .clk (start), .rst (rst)
           , .Q ({mReg_15,mReg_14,mReg_13,mReg_12,mReg_11,mReg_10,mReg_9,mReg_8,
           mReg_7,mReg_6,mReg_5,mReg_4,mReg_3,mReg_2,mReg_1,mReg_0})) ;
    BinaryMux_33 MuxCmp (.a ({pReg_32,pReg_31,pReg_30,pReg_29,pReg_28,pReg_27,
                 pReg_26,pReg_25,pReg_24,pReg_23,pReg_22,pReg_21,pReg_20,pReg_19
                 ,pReg_18,pReg_17,pReg_16,pReg_15,pReg_14,pReg_13,pReg_12,
                 pReg_11,pReg_10,pReg_9,pReg_8,pReg_7,pReg_6,pReg_5,pReg_4,
                 pReg_3,pReg_2,pReg_1,pReg_0}), .b ({pInit_32,pInit_32,pInit_32,
                 pInit_32,pInit_32,pInit_32,pInit_32,pInit_32,pInit_32,pInit_32,
                 pInit_32,pInit_32,pInit_32,pInit_32,pInit_32,pInit_32,pInit_32,
                 pInit_32,pInit_32,pInit_32,pInit_32,pInit_32,pInit_32,pInit_32,
                 q[7],q[6],q[5],q[4],q[3],q[2],q[1],q[0],pInit_32}), .sel (sel)
                 , .f ({pMux_32,pMux_31,pMux_30,pMux_29,pMux_28,pMux_27,pMux_26,
                 pMux_25,pMux_24,pMux_23,pMux_22,pMux_21,pMux_20,pMux_19,pMux_18
                 ,pMux_17,pMux_16,pMux_15,pMux_14,pMux_13,pMux_12,pMux_11,
                 pMux_10,pMux_9,pMux_8,pMux_7,pMux_6,pMux_5,pMux_4,pMux_3,pMux_2
                 ,pMux_1,pMux_0})) ;
    BoothStep BSCmp (.p ({pMux_32,pMux_31,pMux_30,pMux_29,pMux_28,pMux_27,
              pMux_26,pMux_25,pMux_24,pMux_23,pMux_22,pMux_21,pMux_20,pMux_19,
              pMux_18,pMux_17,pMux_16,pMux_15,pMux_14,pMux_13,pMux_12,pMux_11,
              pMux_10,pMux_9,pMux_8,pMux_7,pMux_6,pMux_5,pMux_4,pMux_3,pMux_2,
              pMux_1,pMux_0}), .x ({nx198,nx198,nx200,nx202,nx204,nx206,nx208,
              nx210,nx212,mReg_14,mReg_13,mReg_12,mReg_11,mReg_10,mReg_9,mReg_8,
              mReg_7,mReg_6,mReg_5,mReg_4,mReg_3,mReg_2,mReg_1,mReg_0}), .f ({
              pBs_32,\$dummy [0],pBs_30,pBs_29,pBs_28,pBs_27,pBs_26,pBs_25,
              pBs_24,pBs_23,f[15],f[14],f[13],f[12],f[11],f[10],f[9],f[8],f[7],
              f[6],f[5],f[4],f[3],f[2],f[1],f[0],\$dummy [1],\$dummy [2],
              \$dummy [3],\$dummy [4],\$dummy [5],\$dummy [6],\$dummy [7]})) ;
    fake_gnd ix188 (.Y (pInit_32)) ;
    fake_vcc ix186 (.Y (PWR)) ;
    inv01 ix195 (.Y (nx196), .A (mReg_15)) ;
    inv01 ix197 (.Y (nx198), .A (nx196)) ;
    inv01 ix199 (.Y (nx200), .A (nx196)) ;
    inv01 ix201 (.Y (nx202), .A (nx196)) ;
    inv01 ix203 (.Y (nx204), .A (nx196)) ;
    inv01 ix205 (.Y (nx206), .A (nx196)) ;
    inv01 ix207 (.Y (nx208), .A (nx196)) ;
    inv01 ix209 (.Y (nx210), .A (nx196)) ;
    inv01 ix211 (.Y (nx212), .A (nx196)) ;
endmodule


module BoothStep ( p, x, f ) ;

    input [32:0]p ;
    input [23:0]x ;
    output [32:0]f ;

    wire op2_0, carryIn, op2_23, op2_22, op2_21, op2_20, op2_19, op2_18, op2_17, 
         op2_16, op2_15, op2_14, op2_13, op2_12, op2_11, op2_10, op2_9, op2_8, 
         op2_7, op2_6, op2_5, op2_4, op2_3, op2_2, op2_1, nx28, nx305, nx307, 
         nx311, nx317, nx321, nx325, nx329, nx333, nx337, nx341, nx345, nx349, 
         nx353, nx357, nx361, nx365, nx369, nx373, nx377, nx381, nx385, nx389, 
         nx393, nx397, nx401, nx405, nx407, nx414, nx416, nx418, nx421, nx423, 
         nx425, nx427, nx429, nx431, nx433, nx435, nx437, nx439, nx441, nx443, 
         nx445, nx447, nx449, nx451, nx458;
    wire [0:0] \$dummy ;




    assign f[31] = f[32] ;
    assign f[6] = p[8] ;
    assign f[5] = p[7] ;
    assign f[4] = p[6] ;
    assign f[3] = p[5] ;
    assign f[2] = p[4] ;
    assign f[1] = p[3] ;
    assign f[0] = p[2] ;
    NBitAdder_24 AdderCmp (.a ({p[32],p[31],p[30],p[29],p[28],p[27],p[26],p[25],
                 p[24],p[23],p[22],p[21],p[20],p[19],p[18],p[17],p[16],p[15],
                 p[14],p[13],p[12],p[11],p[10],p[9]}), .b ({op2_23,op2_22,op2_21
                 ,op2_20,op2_19,op2_18,op2_17,op2_16,op2_15,op2_14,op2_13,op2_12
                 ,op2_11,op2_10,op2_9,op2_8,op2_7,op2_6,op2_5,op2_4,op2_3,op2_2,
                 op2_1,op2_0}), .carryIn (carryIn), .sum ({f[30],f[29],f[28],
                 f[27],f[26],f[25],f[24],f[23],f[22],f[21],f[20],f[19],f[18],
                 f[17],f[16],f[15],f[14],f[13],f[12],f[11],f[10],f[9],f[8],f[7]}
                 ), .carryOut (\$dummy [0])) ;
    fake_gnd ix256 (.Y (f[32])) ;
    oai221 ix59 (.Y (op2_1), .A0 (x[0]), .A1 (nx435), .B0 (x[1]), .B1 (nx445), .C0 (
           nx307)) ;
    aoi21 ix15 (.Y (carryIn), .A0 (p[1]), .A1 (p[0]), .B0 (nx305)) ;
    inv01 ix306 (.Y (nx305), .A (p[2])) ;
    aoi22 ix308 (.Y (nx307), .A0 (x[1]), .A1 (nx414), .B0 (x[0]), .B1 (nx425)) ;
    nor02_2x ix29 (.Y (nx28), .A0 (p[2]), .A1 (nx311)) ;
    xnor2 ix312 (.Y (nx311), .A0 (p[0]), .A1 (p[1])) ;
    oai221 ix77 (.Y (op2_2), .A0 (x[1]), .A1 (nx435), .B0 (x[2]), .B1 (nx445), .C0 (
           nx317)) ;
    aoi22 ix318 (.Y (nx317), .A0 (x[2]), .A1 (nx414), .B0 (x[1]), .B1 (nx425)) ;
    oai221 ix95 (.Y (op2_3), .A0 (x[2]), .A1 (nx435), .B0 (x[3]), .B1 (nx445), .C0 (
           nx321)) ;
    aoi22 ix322 (.Y (nx321), .A0 (x[3]), .A1 (nx414), .B0 (x[2]), .B1 (nx425)) ;
    oai221 ix113 (.Y (op2_4), .A0 (x[3]), .A1 (nx435), .B0 (x[4]), .B1 (nx445), 
           .C0 (nx325)) ;
    aoi22 ix326 (.Y (nx325), .A0 (x[4]), .A1 (nx414), .B0 (x[3]), .B1 (nx425)) ;
    oai221 ix131 (.Y (op2_5), .A0 (x[4]), .A1 (nx435), .B0 (x[5]), .B1 (nx445), 
           .C0 (nx329)) ;
    aoi22 ix330 (.Y (nx329), .A0 (x[5]), .A1 (nx414), .B0 (x[4]), .B1 (nx425)) ;
    oai221 ix149 (.Y (op2_6), .A0 (x[5]), .A1 (nx435), .B0 (x[6]), .B1 (nx445), 
           .C0 (nx333)) ;
    aoi22 ix334 (.Y (nx333), .A0 (x[6]), .A1 (nx414), .B0 (x[5]), .B1 (nx425)) ;
    oai221 ix167 (.Y (op2_7), .A0 (x[6]), .A1 (nx437), .B0 (x[7]), .B1 (nx445), 
           .C0 (nx337)) ;
    aoi22 ix338 (.Y (nx337), .A0 (x[7]), .A1 (nx414), .B0 (x[6]), .B1 (nx425)) ;
    oai221 ix185 (.Y (op2_8), .A0 (x[7]), .A1 (nx437), .B0 (x[8]), .B1 (nx447), 
           .C0 (nx341)) ;
    aoi22 ix342 (.Y (nx341), .A0 (x[8]), .A1 (nx416), .B0 (x[7]), .B1 (nx427)) ;
    oai221 ix203 (.Y (op2_9), .A0 (x[8]), .A1 (nx437), .B0 (x[9]), .B1 (nx447), 
           .C0 (nx345)) ;
    aoi22 ix346 (.Y (nx345), .A0 (x[9]), .A1 (nx416), .B0 (x[8]), .B1 (nx427)) ;
    oai221 ix221 (.Y (op2_10), .A0 (x[9]), .A1 (nx437), .B0 (x[10]), .B1 (nx447)
           , .C0 (nx349)) ;
    aoi22 ix350 (.Y (nx349), .A0 (x[10]), .A1 (nx416), .B0 (x[9]), .B1 (nx427)
          ) ;
    oai221 ix239 (.Y (op2_11), .A0 (x[10]), .A1 (nx437), .B0 (x[11]), .B1 (nx447
           ), .C0 (nx353)) ;
    aoi22 ix354 (.Y (nx353), .A0 (x[11]), .A1 (nx416), .B0 (x[10]), .B1 (nx427)
          ) ;
    oai221 ix257 (.Y (op2_12), .A0 (x[11]), .A1 (nx437), .B0 (x[12]), .B1 (nx447
           ), .C0 (nx357)) ;
    aoi22 ix358 (.Y (nx357), .A0 (x[12]), .A1 (nx416), .B0 (x[11]), .B1 (nx427)
          ) ;
    oai221 ix275 (.Y (op2_13), .A0 (x[12]), .A1 (nx437), .B0 (x[13]), .B1 (nx447
           ), .C0 (nx361)) ;
    aoi22 ix362 (.Y (nx361), .A0 (x[13]), .A1 (nx416), .B0 (x[12]), .B1 (nx427)
          ) ;
    oai221 ix293 (.Y (op2_14), .A0 (x[13]), .A1 (nx439), .B0 (x[14]), .B1 (nx447
           ), .C0 (nx365)) ;
    aoi22 ix366 (.Y (nx365), .A0 (x[14]), .A1 (nx416), .B0 (x[13]), .B1 (nx427)
          ) ;
    oai221 ix311 (.Y (op2_15), .A0 (x[14]), .A1 (nx439), .B0 (x[15]), .B1 (nx449
           ), .C0 (nx369)) ;
    aoi22 ix370 (.Y (nx369), .A0 (x[15]), .A1 (nx418), .B0 (x[14]), .B1 (nx429)
          ) ;
    oai221 ix329 (.Y (op2_16), .A0 (x[15]), .A1 (nx439), .B0 (x[16]), .B1 (nx449
           ), .C0 (nx373)) ;
    aoi22 ix374 (.Y (nx373), .A0 (x[16]), .A1 (nx418), .B0 (x[15]), .B1 (nx429)
          ) ;
    oai221 ix347 (.Y (op2_17), .A0 (x[16]), .A1 (nx439), .B0 (x[17]), .B1 (nx449
           ), .C0 (nx377)) ;
    aoi22 ix378 (.Y (nx377), .A0 (x[17]), .A1 (nx418), .B0 (x[16]), .B1 (nx429)
          ) ;
    oai221 ix365 (.Y (op2_18), .A0 (x[17]), .A1 (nx439), .B0 (x[18]), .B1 (nx449
           ), .C0 (nx381)) ;
    aoi22 ix382 (.Y (nx381), .A0 (x[18]), .A1 (nx418), .B0 (x[17]), .B1 (nx429)
          ) ;
    oai221 ix383 (.Y (op2_19), .A0 (x[18]), .A1 (nx439), .B0 (x[19]), .B1 (nx449
           ), .C0 (nx385)) ;
    aoi22 ix386 (.Y (nx385), .A0 (x[19]), .A1 (nx418), .B0 (x[18]), .B1 (nx429)
          ) ;
    oai221 ix401 (.Y (op2_20), .A0 (x[19]), .A1 (nx439), .B0 (x[20]), .B1 (nx449
           ), .C0 (nx389)) ;
    aoi22 ix390 (.Y (nx389), .A0 (x[20]), .A1 (nx418), .B0 (x[19]), .B1 (nx429)
          ) ;
    oai221 ix419 (.Y (op2_21), .A0 (x[20]), .A1 (nx441), .B0 (x[21]), .B1 (nx449
           ), .C0 (nx393)) ;
    aoi22 ix394 (.Y (nx393), .A0 (x[21]), .A1 (nx418), .B0 (x[20]), .B1 (nx429)
          ) ;
    oai221 ix437 (.Y (op2_22), .A0 (x[21]), .A1 (nx441), .B0 (x[22]), .B1 (nx451
           ), .C0 (nx397)) ;
    aoi22 ix398 (.Y (nx397), .A0 (x[22]), .A1 (nx421), .B0 (x[21]), .B1 (nx431)
          ) ;
    oai221 ix455 (.Y (op2_23), .A0 (x[22]), .A1 (nx441), .B0 (x[23]), .B1 (nx451
           ), .C0 (nx401)) ;
    aoi22 ix402 (.Y (nx401), .A0 (x[23]), .A1 (nx421), .B0 (x[22]), .B1 (nx431)
          ) ;
    nand02 ix35 (.Y (op2_0), .A0 (nx405), .A1 (nx441)) ;
    inv01 ix408 (.Y (nx407), .A (nx28)) ;
    inv02 ix413 (.Y (nx414), .A (nx407)) ;
    inv02 ix415 (.Y (nx416), .A (nx407)) ;
    inv02 ix417 (.Y (nx418), .A (nx407)) ;
    inv02 ix420 (.Y (nx421), .A (nx407)) ;
    inv02 ix424 (.Y (nx425), .A (nx423)) ;
    inv02 ix426 (.Y (nx427), .A (nx423)) ;
    inv02 ix428 (.Y (nx429), .A (nx423)) ;
    inv02 ix430 (.Y (nx431), .A (nx423)) ;
    inv02 ix434 (.Y (nx435), .A (nx433)) ;
    inv02 ix436 (.Y (nx437), .A (nx433)) ;
    inv02 ix438 (.Y (nx439), .A (nx433)) ;
    inv02 ix440 (.Y (nx441), .A (nx433)) ;
    inv02 ix444 (.Y (nx445), .A (nx443)) ;
    inv02 ix446 (.Y (nx447), .A (nx458)) ;
    inv02 ix448 (.Y (nx449), .A (nx458)) ;
    inv02 ix450 (.Y (nx451), .A (nx458)) ;
    nor03_2x ix296 (.Y (nx433), .A0 (p[1]), .A1 (nx305), .A2 (p[0])) ;
    nor02ii ix302 (.Y (nx443), .A0 (nx433), .A1 (carryIn)) ;
    nand03 ix51 (.Y (nx423), .A0 (p[1]), .A1 (nx305), .A2 (p[0])) ;
    mux21 ix406 (.Y (nx405), .A0 (nx458), .A1 (nx28), .S0 (x[0])) ;
    inv01 ix457 (.Y (nx458), .A (nx445)) ;
endmodule


module NBitAdder_24 ( a, b, carryIn, sum, carryOut ) ;

    input [23:0]a ;
    input [23:0]b ;
    input carryIn ;
    output [23:0]sum ;
    output carryOut ;

    wire temp_22, temp_21, temp_20, temp_19, temp_18, temp_17, temp_16, temp_15, 
         temp_14, temp_13, temp_12, temp_11, temp_10, temp_9, temp_8, temp_7, 
         temp_6, temp_5, temp_4, temp_3, temp_2, temp_1, temp_0;



    FullAdder f0 (.a (a[0]), .b (b[0]), .cin (carryIn), .s (sum[0]), .cout (
              temp_0)) ;
    FullAdder loop1_1_fx (.a (a[1]), .b (b[1]), .cin (temp_0), .s (sum[1]), .cout (
              temp_1)) ;
    FullAdder loop1_2_fx (.a (a[2]), .b (b[2]), .cin (temp_1), .s (sum[2]), .cout (
              temp_2)) ;
    FullAdder loop1_3_fx (.a (a[3]), .b (b[3]), .cin (temp_2), .s (sum[3]), .cout (
              temp_3)) ;
    FullAdder loop1_4_fx (.a (a[4]), .b (b[4]), .cin (temp_3), .s (sum[4]), .cout (
              temp_4)) ;
    FullAdder loop1_5_fx (.a (a[5]), .b (b[5]), .cin (temp_4), .s (sum[5]), .cout (
              temp_5)) ;
    FullAdder loop1_6_fx (.a (a[6]), .b (b[6]), .cin (temp_5), .s (sum[6]), .cout (
              temp_6)) ;
    FullAdder loop1_7_fx (.a (a[7]), .b (b[7]), .cin (temp_6), .s (sum[7]), .cout (
              temp_7)) ;
    FullAdder loop1_8_fx (.a (a[8]), .b (b[8]), .cin (temp_7), .s (sum[8]), .cout (
              temp_8)) ;
    FullAdder loop1_9_fx (.a (a[9]), .b (b[9]), .cin (temp_8), .s (sum[9]), .cout (
              temp_9)) ;
    FullAdder loop1_10_fx (.a (a[10]), .b (b[10]), .cin (temp_9), .s (sum[10]), 
              .cout (temp_10)) ;
    FullAdder loop1_11_fx (.a (a[11]), .b (b[11]), .cin (temp_10), .s (sum[11])
              , .cout (temp_11)) ;
    FullAdder loop1_12_fx (.a (a[12]), .b (b[12]), .cin (temp_11), .s (sum[12])
              , .cout (temp_12)) ;
    FullAdder loop1_13_fx (.a (a[13]), .b (b[13]), .cin (temp_12), .s (sum[13])
              , .cout (temp_13)) ;
    FullAdder loop1_14_fx (.a (a[14]), .b (b[14]), .cin (temp_13), .s (sum[14])
              , .cout (temp_14)) ;
    FullAdder loop1_15_fx (.a (a[15]), .b (b[15]), .cin (temp_14), .s (sum[15])
              , .cout (temp_15)) ;
    FullAdder loop1_16_fx (.a (a[16]), .b (b[16]), .cin (temp_15), .s (sum[16])
              , .cout (temp_16)) ;
    FullAdder loop1_17_fx (.a (a[17]), .b (b[17]), .cin (temp_16), .s (sum[17])
              , .cout (temp_17)) ;
    FullAdder loop1_18_fx (.a (a[18]), .b (b[18]), .cin (temp_17), .s (sum[18])
              , .cout (temp_18)) ;
    FullAdder loop1_19_fx (.a (a[19]), .b (b[19]), .cin (temp_18), .s (sum[19])
              , .cout (temp_19)) ;
    FullAdder loop1_20_fx (.a (a[20]), .b (b[20]), .cin (temp_19), .s (sum[20])
              , .cout (temp_20)) ;
    FullAdder loop1_21_fx (.a (a[21]), .b (b[21]), .cin (temp_20), .s (sum[21])
              , .cout (temp_21)) ;
    FullAdder loop1_22_fx (.a (a[22]), .b (b[22]), .cin (temp_21), .s (sum[22])
              , .cout (temp_22)) ;
    FullAdder loop1_23_fx (.a (a[23]), .b (b[23]), .cin (temp_22), .s (sum[23])
              , .cout (carryOut)) ;
endmodule


module FullAdder ( a, b, cin, s, cout ) ;

    input a ;
    input b ;
    input cin ;
    output s ;
    output cout ;

    wire nx0, nx69;



    ao22 ix7 (.Y (cout), .A0 (b), .A1 (a), .B0 (cin), .B1 (nx0)) ;
    xnor2 ix9 (.Y (s), .A0 (nx69), .A1 (cin)) ;
    xnor2 ix70 (.Y (nx69), .A0 (a), .A1 (b)) ;
    inv01 ix1 (.Y (nx0), .A (nx69)) ;
endmodule


module BinaryMux_33 ( a, b, sel, f ) ;

    input [32:0]a ;
    input [32:0]b ;
    input sel ;
    output [32:0]f ;

    wire nx298, nx300, nx302, nx304, nx306, nx308;



    mux21_ni ix7 (.Y (f[0]), .A0 (a[0]), .A1 (b[0]), .S0 (nx300)) ;
    mux21_ni ix15 (.Y (f[1]), .A0 (a[1]), .A1 (b[1]), .S0 (nx300)) ;
    mux21_ni ix23 (.Y (f[2]), .A0 (a[2]), .A1 (b[2]), .S0 (nx300)) ;
    mux21_ni ix31 (.Y (f[3]), .A0 (a[3]), .A1 (b[3]), .S0 (nx300)) ;
    mux21_ni ix39 (.Y (f[4]), .A0 (a[4]), .A1 (b[4]), .S0 (nx300)) ;
    mux21_ni ix47 (.Y (f[5]), .A0 (a[5]), .A1 (b[5]), .S0 (nx300)) ;
    mux21_ni ix55 (.Y (f[6]), .A0 (a[6]), .A1 (b[6]), .S0 (nx300)) ;
    mux21_ni ix63 (.Y (f[7]), .A0 (a[7]), .A1 (b[7]), .S0 (nx302)) ;
    mux21_ni ix71 (.Y (f[8]), .A0 (a[8]), .A1 (b[8]), .S0 (nx302)) ;
    mux21_ni ix79 (.Y (f[9]), .A0 (a[9]), .A1 (b[9]), .S0 (nx302)) ;
    mux21_ni ix87 (.Y (f[10]), .A0 (a[10]), .A1 (b[10]), .S0 (nx302)) ;
    mux21_ni ix95 (.Y (f[11]), .A0 (a[11]), .A1 (b[11]), .S0 (nx302)) ;
    mux21_ni ix103 (.Y (f[12]), .A0 (a[12]), .A1 (b[12]), .S0 (nx302)) ;
    mux21_ni ix111 (.Y (f[13]), .A0 (a[13]), .A1 (b[13]), .S0 (nx302)) ;
    mux21_ni ix119 (.Y (f[14]), .A0 (a[14]), .A1 (b[14]), .S0 (nx304)) ;
    mux21_ni ix127 (.Y (f[15]), .A0 (a[15]), .A1 (b[15]), .S0 (nx304)) ;
    mux21_ni ix135 (.Y (f[16]), .A0 (a[16]), .A1 (b[16]), .S0 (nx304)) ;
    mux21_ni ix143 (.Y (f[17]), .A0 (a[17]), .A1 (b[17]), .S0 (nx304)) ;
    mux21_ni ix151 (.Y (f[18]), .A0 (a[18]), .A1 (b[18]), .S0 (nx304)) ;
    mux21_ni ix159 (.Y (f[19]), .A0 (a[19]), .A1 (b[19]), .S0 (nx304)) ;
    mux21_ni ix167 (.Y (f[20]), .A0 (a[20]), .A1 (b[20]), .S0 (nx304)) ;
    mux21_ni ix175 (.Y (f[21]), .A0 (a[21]), .A1 (b[21]), .S0 (nx306)) ;
    mux21_ni ix183 (.Y (f[22]), .A0 (a[22]), .A1 (b[22]), .S0 (nx306)) ;
    mux21_ni ix191 (.Y (f[23]), .A0 (a[23]), .A1 (b[23]), .S0 (nx306)) ;
    mux21_ni ix199 (.Y (f[24]), .A0 (a[24]), .A1 (b[24]), .S0 (nx306)) ;
    mux21_ni ix207 (.Y (f[25]), .A0 (a[25]), .A1 (b[25]), .S0 (nx306)) ;
    mux21_ni ix215 (.Y (f[26]), .A0 (a[26]), .A1 (b[26]), .S0 (nx306)) ;
    mux21_ni ix223 (.Y (f[27]), .A0 (a[27]), .A1 (b[27]), .S0 (nx306)) ;
    mux21_ni ix231 (.Y (f[28]), .A0 (a[28]), .A1 (b[28]), .S0 (nx308)) ;
    mux21_ni ix239 (.Y (f[29]), .A0 (a[29]), .A1 (b[29]), .S0 (nx308)) ;
    mux21_ni ix247 (.Y (f[30]), .A0 (a[30]), .A1 (b[30]), .S0 (nx308)) ;
    mux21_ni ix255 (.Y (f[31]), .A0 (a[31]), .A1 (b[31]), .S0 (nx308)) ;
    mux21_ni ix263 (.Y (f[32]), .A0 (a[32]), .A1 (b[32]), .S0 (nx308)) ;
    inv01 ix297 (.Y (nx298), .A (sel)) ;
    inv02 ix299 (.Y (nx300), .A (nx298)) ;
    inv02 ix301 (.Y (nx302), .A (nx298)) ;
    inv02 ix303 (.Y (nx304), .A (nx298)) ;
    inv02 ix305 (.Y (nx306), .A (nx298)) ;
    inv02 ix307 (.Y (nx308), .A (nx298)) ;
endmodule


module Reg_33 ( D, en, clk, rst, Q ) ;

    input [32:0]D ;
    input en ;
    input clk ;
    input rst ;
    output [32:0]Q ;

    wire nx432, nx442, nx452, nx462, nx472, nx482, nx492, nx502, nx512, nx522, 
         nx532, nx542, nx552, nx562, nx572, nx582, nx592, nx602, nx612, nx622, 
         nx632, nx642, nx652, nx662, nx672, nx682, nx692, nx702, nx712, nx722, 
         nx732, nx742, nx752, nx866, nx868, nx870, nx872, nx874, nx876, nx878, 
         nx880, nx882, nx884, nx886, nx888;
    wire [32:0] \$dummy ;




    dffr reg_Q_0 (.Q (Q[0]), .QB (\$dummy [0]), .D (nx432), .CLK (nx880), .R (
         rst)) ;
    mux21_ni ix433 (.Y (nx432), .A0 (Q[0]), .A1 (D[0]), .S0 (nx868)) ;
    dffr reg_Q_1 (.Q (Q[1]), .QB (\$dummy [1]), .D (nx442), .CLK (nx880), .R (
         rst)) ;
    mux21_ni ix443 (.Y (nx442), .A0 (Q[1]), .A1 (D[1]), .S0 (nx868)) ;
    dffr reg_Q_2 (.Q (Q[2]), .QB (\$dummy [2]), .D (nx452), .CLK (nx880), .R (
         rst)) ;
    mux21_ni ix453 (.Y (nx452), .A0 (Q[2]), .A1 (D[2]), .S0 (nx868)) ;
    dffr reg_Q_3 (.Q (Q[3]), .QB (\$dummy [3]), .D (nx462), .CLK (nx880), .R (
         rst)) ;
    mux21_ni ix463 (.Y (nx462), .A0 (Q[3]), .A1 (D[3]), .S0 (nx868)) ;
    dffr reg_Q_4 (.Q (Q[4]), .QB (\$dummy [4]), .D (nx472), .CLK (nx880), .R (
         rst)) ;
    mux21_ni ix473 (.Y (nx472), .A0 (Q[4]), .A1 (D[4]), .S0 (nx868)) ;
    dffr reg_Q_5 (.Q (Q[5]), .QB (\$dummy [5]), .D (nx482), .CLK (nx880), .R (
         rst)) ;
    mux21_ni ix483 (.Y (nx482), .A0 (Q[5]), .A1 (D[5]), .S0 (nx868)) ;
    dffr reg_Q_6 (.Q (Q[6]), .QB (\$dummy [6]), .D (nx492), .CLK (nx880), .R (
         rst)) ;
    mux21_ni ix493 (.Y (nx492), .A0 (Q[6]), .A1 (D[6]), .S0 (nx868)) ;
    dffr reg_Q_7 (.Q (Q[7]), .QB (\$dummy [7]), .D (nx502), .CLK (nx882), .R (
         rst)) ;
    mux21_ni ix503 (.Y (nx502), .A0 (Q[7]), .A1 (D[7]), .S0 (nx870)) ;
    dffr reg_Q_8 (.Q (Q[8]), .QB (\$dummy [8]), .D (nx512), .CLK (nx882), .R (
         rst)) ;
    mux21_ni ix513 (.Y (nx512), .A0 (Q[8]), .A1 (D[8]), .S0 (nx870)) ;
    dffr reg_Q_9 (.Q (Q[9]), .QB (\$dummy [9]), .D (nx522), .CLK (nx882), .R (
         rst)) ;
    mux21_ni ix523 (.Y (nx522), .A0 (Q[9]), .A1 (D[9]), .S0 (nx870)) ;
    dffr reg_Q_10 (.Q (Q[10]), .QB (\$dummy [10]), .D (nx532), .CLK (nx882), .R (
         rst)) ;
    mux21_ni ix533 (.Y (nx532), .A0 (Q[10]), .A1 (D[10]), .S0 (nx870)) ;
    dffr reg_Q_11 (.Q (Q[11]), .QB (\$dummy [11]), .D (nx542), .CLK (nx882), .R (
         rst)) ;
    mux21_ni ix543 (.Y (nx542), .A0 (Q[11]), .A1 (D[11]), .S0 (nx870)) ;
    dffr reg_Q_12 (.Q (Q[12]), .QB (\$dummy [12]), .D (nx552), .CLK (nx882), .R (
         rst)) ;
    mux21_ni ix553 (.Y (nx552), .A0 (Q[12]), .A1 (D[12]), .S0 (nx870)) ;
    dffr reg_Q_13 (.Q (Q[13]), .QB (\$dummy [13]), .D (nx562), .CLK (nx882), .R (
         rst)) ;
    mux21_ni ix563 (.Y (nx562), .A0 (Q[13]), .A1 (D[13]), .S0 (nx870)) ;
    dffr reg_Q_14 (.Q (Q[14]), .QB (\$dummy [14]), .D (nx572), .CLK (nx884), .R (
         rst)) ;
    mux21_ni ix573 (.Y (nx572), .A0 (Q[14]), .A1 (D[14]), .S0 (nx872)) ;
    dffr reg_Q_15 (.Q (Q[15]), .QB (\$dummy [15]), .D (nx582), .CLK (nx884), .R (
         rst)) ;
    mux21_ni ix583 (.Y (nx582), .A0 (Q[15]), .A1 (D[15]), .S0 (nx872)) ;
    dffr reg_Q_16 (.Q (Q[16]), .QB (\$dummy [16]), .D (nx592), .CLK (nx884), .R (
         rst)) ;
    mux21_ni ix593 (.Y (nx592), .A0 (Q[16]), .A1 (D[16]), .S0 (nx872)) ;
    dffr reg_Q_17 (.Q (Q[17]), .QB (\$dummy [17]), .D (nx602), .CLK (nx884), .R (
         rst)) ;
    mux21_ni ix603 (.Y (nx602), .A0 (Q[17]), .A1 (D[17]), .S0 (nx872)) ;
    dffr reg_Q_18 (.Q (Q[18]), .QB (\$dummy [18]), .D (nx612), .CLK (nx884), .R (
         rst)) ;
    mux21_ni ix613 (.Y (nx612), .A0 (Q[18]), .A1 (D[18]), .S0 (nx872)) ;
    dffr reg_Q_19 (.Q (Q[19]), .QB (\$dummy [19]), .D (nx622), .CLK (nx884), .R (
         rst)) ;
    mux21_ni ix623 (.Y (nx622), .A0 (Q[19]), .A1 (D[19]), .S0 (nx872)) ;
    dffr reg_Q_20 (.Q (Q[20]), .QB (\$dummy [20]), .D (nx632), .CLK (nx884), .R (
         rst)) ;
    mux21_ni ix633 (.Y (nx632), .A0 (Q[20]), .A1 (D[20]), .S0 (nx872)) ;
    dffr reg_Q_21 (.Q (Q[21]), .QB (\$dummy [21]), .D (nx642), .CLK (nx886), .R (
         rst)) ;
    mux21_ni ix643 (.Y (nx642), .A0 (Q[21]), .A1 (D[21]), .S0 (nx874)) ;
    dffr reg_Q_22 (.Q (Q[22]), .QB (\$dummy [22]), .D (nx652), .CLK (nx886), .R (
         rst)) ;
    mux21_ni ix653 (.Y (nx652), .A0 (Q[22]), .A1 (D[22]), .S0 (nx874)) ;
    dffr reg_Q_23 (.Q (Q[23]), .QB (\$dummy [23]), .D (nx662), .CLK (nx886), .R (
         rst)) ;
    mux21_ni ix663 (.Y (nx662), .A0 (Q[23]), .A1 (D[23]), .S0 (nx874)) ;
    dffr reg_Q_24 (.Q (Q[24]), .QB (\$dummy [24]), .D (nx672), .CLK (nx886), .R (
         rst)) ;
    mux21_ni ix673 (.Y (nx672), .A0 (Q[24]), .A1 (D[24]), .S0 (nx874)) ;
    dffr reg_Q_25 (.Q (Q[25]), .QB (\$dummy [25]), .D (nx682), .CLK (nx886), .R (
         rst)) ;
    mux21_ni ix683 (.Y (nx682), .A0 (Q[25]), .A1 (D[25]), .S0 (nx874)) ;
    dffr reg_Q_26 (.Q (Q[26]), .QB (\$dummy [26]), .D (nx692), .CLK (nx886), .R (
         rst)) ;
    mux21_ni ix693 (.Y (nx692), .A0 (Q[26]), .A1 (D[26]), .S0 (nx874)) ;
    dffr reg_Q_27 (.Q (Q[27]), .QB (\$dummy [27]), .D (nx702), .CLK (nx886), .R (
         rst)) ;
    mux21_ni ix703 (.Y (nx702), .A0 (Q[27]), .A1 (D[27]), .S0 (nx874)) ;
    dffr reg_Q_28 (.Q (Q[28]), .QB (\$dummy [28]), .D (nx712), .CLK (nx888), .R (
         rst)) ;
    mux21_ni ix713 (.Y (nx712), .A0 (Q[28]), .A1 (D[28]), .S0 (nx876)) ;
    dffr reg_Q_29 (.Q (Q[29]), .QB (\$dummy [29]), .D (nx722), .CLK (nx888), .R (
         rst)) ;
    mux21_ni ix723 (.Y (nx722), .A0 (Q[29]), .A1 (D[29]), .S0 (nx876)) ;
    dffr reg_Q_30 (.Q (Q[30]), .QB (\$dummy [30]), .D (nx732), .CLK (nx888), .R (
         rst)) ;
    mux21_ni ix733 (.Y (nx732), .A0 (Q[30]), .A1 (D[30]), .S0 (nx876)) ;
    dffr reg_Q_31 (.Q (Q[31]), .QB (\$dummy [31]), .D (nx742), .CLK (nx888), .R (
         rst)) ;
    mux21_ni ix743 (.Y (nx742), .A0 (Q[31]), .A1 (D[31]), .S0 (nx876)) ;
    dffr reg_Q_32 (.Q (Q[32]), .QB (\$dummy [32]), .D (nx752), .CLK (nx888), .R (
         rst)) ;
    mux21_ni ix753 (.Y (nx752), .A0 (Q[32]), .A1 (D[32]), .S0 (nx876)) ;
    inv01 ix865 (.Y (nx866), .A (en)) ;
    inv02 ix867 (.Y (nx868), .A (nx866)) ;
    inv02 ix869 (.Y (nx870), .A (nx866)) ;
    inv02 ix871 (.Y (nx872), .A (nx866)) ;
    inv02 ix873 (.Y (nx874), .A (nx866)) ;
    inv02 ix875 (.Y (nx876), .A (nx866)) ;
    inv01 ix877 (.Y (nx878), .A (clk)) ;
    inv02 ix879 (.Y (nx880), .A (nx878)) ;
    inv02 ix881 (.Y (nx882), .A (nx878)) ;
    inv02 ix883 (.Y (nx884), .A (nx878)) ;
    inv02 ix885 (.Y (nx886), .A (nx878)) ;
    inv02 ix887 (.Y (nx888), .A (nx878)) ;
endmodule


module RegFile_8_16_5_5_3_3 ( filterBus, windowBus, decoderRow, clk, rst, 
                              enablePage1Read, enablePage2Read, enableFilterRead, 
                              shift2To1, shift1To2, pageTurn, pagesOuts_0__15, 
                              pagesOuts_0__14, pagesOuts_0__13, pagesOuts_0__12, 
                              pagesOuts_0__11, pagesOuts_0__10, pagesOuts_0__9, 
                              pagesOuts_0__8, pagesOuts_0__7, pagesOuts_0__6, 
                              pagesOuts_0__5, pagesOuts_0__4, pagesOuts_0__3, 
                              pagesOuts_0__2, pagesOuts_0__1, pagesOuts_0__0, 
                              pagesOuts_1__15, pagesOuts_1__14, pagesOuts_1__13, 
                              pagesOuts_1__12, pagesOuts_1__11, pagesOuts_1__10, 
                              pagesOuts_1__9, pagesOuts_1__8, pagesOuts_1__7, 
                              pagesOuts_1__6, pagesOuts_1__5, pagesOuts_1__4, 
                              pagesOuts_1__3, pagesOuts_1__2, pagesOuts_1__1, 
                              pagesOuts_1__0, pagesOuts_2__15, pagesOuts_2__14, 
                              pagesOuts_2__13, pagesOuts_2__12, pagesOuts_2__11, 
                              pagesOuts_2__10, pagesOuts_2__9, pagesOuts_2__8, 
                              pagesOuts_2__7, pagesOuts_2__6, pagesOuts_2__5, 
                              pagesOuts_2__4, pagesOuts_2__3, pagesOuts_2__2, 
                              pagesOuts_2__1, pagesOuts_2__0, pagesOuts_3__15, 
                              pagesOuts_3__14, pagesOuts_3__13, pagesOuts_3__12, 
                              pagesOuts_3__11, pagesOuts_3__10, pagesOuts_3__9, 
                              pagesOuts_3__8, pagesOuts_3__7, pagesOuts_3__6, 
                              pagesOuts_3__5, pagesOuts_3__4, pagesOuts_3__3, 
                              pagesOuts_3__2, pagesOuts_3__1, pagesOuts_3__0, 
                              pagesOuts_4__15, pagesOuts_4__14, pagesOuts_4__13, 
                              pagesOuts_4__12, pagesOuts_4__11, pagesOuts_4__10, 
                              pagesOuts_4__9, pagesOuts_4__8, pagesOuts_4__7, 
                              pagesOuts_4__6, pagesOuts_4__5, pagesOuts_4__4, 
                              pagesOuts_4__3, pagesOuts_4__2, pagesOuts_4__1, 
                              pagesOuts_4__0, pagesOuts_5__15, pagesOuts_5__14, 
                              pagesOuts_5__13, pagesOuts_5__12, pagesOuts_5__11, 
                              pagesOuts_5__10, pagesOuts_5__9, pagesOuts_5__8, 
                              pagesOuts_5__7, pagesOuts_5__6, pagesOuts_5__5, 
                              pagesOuts_5__4, pagesOuts_5__3, pagesOuts_5__2, 
                              pagesOuts_5__1, pagesOuts_5__0, pagesOuts_6__15, 
                              pagesOuts_6__14, pagesOuts_6__13, pagesOuts_6__12, 
                              pagesOuts_6__11, pagesOuts_6__10, pagesOuts_6__9, 
                              pagesOuts_6__8, pagesOuts_6__7, pagesOuts_6__6, 
                              pagesOuts_6__5, pagesOuts_6__4, pagesOuts_6__3, 
                              pagesOuts_6__2, pagesOuts_6__1, pagesOuts_6__0, 
                              pagesOuts_7__15, pagesOuts_7__14, pagesOuts_7__13, 
                              pagesOuts_7__12, pagesOuts_7__11, pagesOuts_7__10, 
                              pagesOuts_7__9, pagesOuts_7__8, pagesOuts_7__7, 
                              pagesOuts_7__6, pagesOuts_7__5, pagesOuts_7__4, 
                              pagesOuts_7__3, pagesOuts_7__2, pagesOuts_7__1, 
                              pagesOuts_7__0, pagesOuts_8__15, pagesOuts_8__14, 
                              pagesOuts_8__13, pagesOuts_8__12, pagesOuts_8__11, 
                              pagesOuts_8__10, pagesOuts_8__9, pagesOuts_8__8, 
                              pagesOuts_8__7, pagesOuts_8__6, pagesOuts_8__5, 
                              pagesOuts_8__4, pagesOuts_8__3, pagesOuts_8__2, 
                              pagesOuts_8__1, pagesOuts_8__0, pagesOuts_9__15, 
                              pagesOuts_9__14, pagesOuts_9__13, pagesOuts_9__12, 
                              pagesOuts_9__11, pagesOuts_9__10, pagesOuts_9__9, 
                              pagesOuts_9__8, pagesOuts_9__7, pagesOuts_9__6, 
                              pagesOuts_9__5, pagesOuts_9__4, pagesOuts_9__3, 
                              pagesOuts_9__2, pagesOuts_9__1, pagesOuts_9__0, 
                              pagesOuts_10__15, pagesOuts_10__14, 
                              pagesOuts_10__13, pagesOuts_10__12, 
                              pagesOuts_10__11, pagesOuts_10__10, 
                              pagesOuts_10__9, pagesOuts_10__8, pagesOuts_10__7, 
                              pagesOuts_10__6, pagesOuts_10__5, pagesOuts_10__4, 
                              pagesOuts_10__3, pagesOuts_10__2, pagesOuts_10__1, 
                              pagesOuts_10__0, pagesOuts_11__15, 
                              pagesOuts_11__14, pagesOuts_11__13, 
                              pagesOuts_11__12, pagesOuts_11__11, 
                              pagesOuts_11__10, pagesOuts_11__9, pagesOuts_11__8, 
                              pagesOuts_11__7, pagesOuts_11__6, pagesOuts_11__5, 
                              pagesOuts_11__4, pagesOuts_11__3, pagesOuts_11__2, 
                              pagesOuts_11__1, pagesOuts_11__0, pagesOuts_12__15, 
                              pagesOuts_12__14, pagesOuts_12__13, 
                              pagesOuts_12__12, pagesOuts_12__11, 
                              pagesOuts_12__10, pagesOuts_12__9, pagesOuts_12__8, 
                              pagesOuts_12__7, pagesOuts_12__6, pagesOuts_12__5, 
                              pagesOuts_12__4, pagesOuts_12__3, pagesOuts_12__2, 
                              pagesOuts_12__1, pagesOuts_12__0, pagesOuts_13__15, 
                              pagesOuts_13__14, pagesOuts_13__13, 
                              pagesOuts_13__12, pagesOuts_13__11, 
                              pagesOuts_13__10, pagesOuts_13__9, pagesOuts_13__8, 
                              pagesOuts_13__7, pagesOuts_13__6, pagesOuts_13__5, 
                              pagesOuts_13__4, pagesOuts_13__3, pagesOuts_13__2, 
                              pagesOuts_13__1, pagesOuts_13__0, pagesOuts_14__15, 
                              pagesOuts_14__14, pagesOuts_14__13, 
                              pagesOuts_14__12, pagesOuts_14__11, 
                              pagesOuts_14__10, pagesOuts_14__9, pagesOuts_14__8, 
                              pagesOuts_14__7, pagesOuts_14__6, pagesOuts_14__5, 
                              pagesOuts_14__4, pagesOuts_14__3, pagesOuts_14__2, 
                              pagesOuts_14__1, pagesOuts_14__0, pagesOuts_15__15, 
                              pagesOuts_15__14, pagesOuts_15__13, 
                              pagesOuts_15__12, pagesOuts_15__11, 
                              pagesOuts_15__10, pagesOuts_15__9, pagesOuts_15__8, 
                              pagesOuts_15__7, pagesOuts_15__6, pagesOuts_15__5, 
                              pagesOuts_15__4, pagesOuts_15__3, pagesOuts_15__2, 
                              pagesOuts_15__1, pagesOuts_15__0, pagesOuts_16__15, 
                              pagesOuts_16__14, pagesOuts_16__13, 
                              pagesOuts_16__12, pagesOuts_16__11, 
                              pagesOuts_16__10, pagesOuts_16__9, pagesOuts_16__8, 
                              pagesOuts_16__7, pagesOuts_16__6, pagesOuts_16__5, 
                              pagesOuts_16__4, pagesOuts_16__3, pagesOuts_16__2, 
                              pagesOuts_16__1, pagesOuts_16__0, pagesOuts_17__15, 
                              pagesOuts_17__14, pagesOuts_17__13, 
                              pagesOuts_17__12, pagesOuts_17__11, 
                              pagesOuts_17__10, pagesOuts_17__9, pagesOuts_17__8, 
                              pagesOuts_17__7, pagesOuts_17__6, pagesOuts_17__5, 
                              pagesOuts_17__4, pagesOuts_17__3, pagesOuts_17__2, 
                              pagesOuts_17__1, pagesOuts_17__0, pagesOuts_18__15, 
                              pagesOuts_18__14, pagesOuts_18__13, 
                              pagesOuts_18__12, pagesOuts_18__11, 
                              pagesOuts_18__10, pagesOuts_18__9, pagesOuts_18__8, 
                              pagesOuts_18__7, pagesOuts_18__6, pagesOuts_18__5, 
                              pagesOuts_18__4, pagesOuts_18__3, pagesOuts_18__2, 
                              pagesOuts_18__1, pagesOuts_18__0, pagesOuts_19__15, 
                              pagesOuts_19__14, pagesOuts_19__13, 
                              pagesOuts_19__12, pagesOuts_19__11, 
                              pagesOuts_19__10, pagesOuts_19__9, pagesOuts_19__8, 
                              pagesOuts_19__7, pagesOuts_19__6, pagesOuts_19__5, 
                              pagesOuts_19__4, pagesOuts_19__3, pagesOuts_19__2, 
                              pagesOuts_19__1, pagesOuts_19__0, pagesOuts_20__15, 
                              pagesOuts_20__14, pagesOuts_20__13, 
                              pagesOuts_20__12, pagesOuts_20__11, 
                              pagesOuts_20__10, pagesOuts_20__9, pagesOuts_20__8, 
                              pagesOuts_20__7, pagesOuts_20__6, pagesOuts_20__5, 
                              pagesOuts_20__4, pagesOuts_20__3, pagesOuts_20__2, 
                              pagesOuts_20__1, pagesOuts_20__0, pagesOuts_21__15, 
                              pagesOuts_21__14, pagesOuts_21__13, 
                              pagesOuts_21__12, pagesOuts_21__11, 
                              pagesOuts_21__10, pagesOuts_21__9, pagesOuts_21__8, 
                              pagesOuts_21__7, pagesOuts_21__6, pagesOuts_21__5, 
                              pagesOuts_21__4, pagesOuts_21__3, pagesOuts_21__2, 
                              pagesOuts_21__1, pagesOuts_21__0, pagesOuts_22__15, 
                              pagesOuts_22__14, pagesOuts_22__13, 
                              pagesOuts_22__12, pagesOuts_22__11, 
                              pagesOuts_22__10, pagesOuts_22__9, pagesOuts_22__8, 
                              pagesOuts_22__7, pagesOuts_22__6, pagesOuts_22__5, 
                              pagesOuts_22__4, pagesOuts_22__3, pagesOuts_22__2, 
                              pagesOuts_22__1, pagesOuts_22__0, pagesOuts_23__15, 
                              pagesOuts_23__14, pagesOuts_23__13, 
                              pagesOuts_23__12, pagesOuts_23__11, 
                              pagesOuts_23__10, pagesOuts_23__9, pagesOuts_23__8, 
                              pagesOuts_23__7, pagesOuts_23__6, pagesOuts_23__5, 
                              pagesOuts_23__4, pagesOuts_23__3, pagesOuts_23__2, 
                              pagesOuts_23__1, pagesOuts_23__0, pagesOuts_24__15, 
                              pagesOuts_24__14, pagesOuts_24__13, 
                              pagesOuts_24__12, pagesOuts_24__11, 
                              pagesOuts_24__10, pagesOuts_24__9, pagesOuts_24__8, 
                              pagesOuts_24__7, pagesOuts_24__6, pagesOuts_24__5, 
                              pagesOuts_24__4, pagesOuts_24__3, pagesOuts_24__2, 
                              pagesOuts_24__1, pagesOuts_24__0, filtersOuts_0__7, 
                              filtersOuts_0__6, filtersOuts_0__5, 
                              filtersOuts_0__4, filtersOuts_0__3, 
                              filtersOuts_0__2, filtersOuts_0__1, 
                              filtersOuts_0__0, filtersOuts_1__7, 
                              filtersOuts_1__6, filtersOuts_1__5, 
                              filtersOuts_1__4, filtersOuts_1__3, 
                              filtersOuts_1__2, filtersOuts_1__1, 
                              filtersOuts_1__0, filtersOuts_2__7, 
                              filtersOuts_2__6, filtersOuts_2__5, 
                              filtersOuts_2__4, filtersOuts_2__3, 
                              filtersOuts_2__2, filtersOuts_2__1, 
                              filtersOuts_2__0, filtersOuts_3__7, 
                              filtersOuts_3__6, filtersOuts_3__5, 
                              filtersOuts_3__4, filtersOuts_3__3, 
                              filtersOuts_3__2, filtersOuts_3__1, 
                              filtersOuts_3__0, filtersOuts_4__7, 
                              filtersOuts_4__6, filtersOuts_4__5, 
                              filtersOuts_4__4, filtersOuts_4__3, 
                              filtersOuts_4__2, filtersOuts_4__1, 
                              filtersOuts_4__0, filtersOuts_5__7, 
                              filtersOuts_5__6, filtersOuts_5__5, 
                              filtersOuts_5__4, filtersOuts_5__3, 
                              filtersOuts_5__2, filtersOuts_5__1, 
                              filtersOuts_5__0, filtersOuts_6__7, 
                              filtersOuts_6__6, filtersOuts_6__5, 
                              filtersOuts_6__4, filtersOuts_6__3, 
                              filtersOuts_6__2, filtersOuts_6__1, 
                              filtersOuts_6__0, filtersOuts_7__7, 
                              filtersOuts_7__6, filtersOuts_7__5, 
                              filtersOuts_7__4, filtersOuts_7__3, 
                              filtersOuts_7__2, filtersOuts_7__1, 
                              filtersOuts_7__0, filtersOuts_8__7, 
                              filtersOuts_8__6, filtersOuts_8__5, 
                              filtersOuts_8__4, filtersOuts_8__3, 
                              filtersOuts_8__2, filtersOuts_8__1, 
                              filtersOuts_8__0, filtersOuts_9__7, 
                              filtersOuts_9__6, filtersOuts_9__5, 
                              filtersOuts_9__4, filtersOuts_9__3, 
                              filtersOuts_9__2, filtersOuts_9__1, 
                              filtersOuts_9__0, filtersOuts_10__7, 
                              filtersOuts_10__6, filtersOuts_10__5, 
                              filtersOuts_10__4, filtersOuts_10__3, 
                              filtersOuts_10__2, filtersOuts_10__1, 
                              filtersOuts_10__0, filtersOuts_11__7, 
                              filtersOuts_11__6, filtersOuts_11__5, 
                              filtersOuts_11__4, filtersOuts_11__3, 
                              filtersOuts_11__2, filtersOuts_11__1, 
                              filtersOuts_11__0, filtersOuts_12__7, 
                              filtersOuts_12__6, filtersOuts_12__5, 
                              filtersOuts_12__4, filtersOuts_12__3, 
                              filtersOuts_12__2, filtersOuts_12__1, 
                              filtersOuts_12__0, filtersOuts_13__7, 
                              filtersOuts_13__6, filtersOuts_13__5, 
                              filtersOuts_13__4, filtersOuts_13__3, 
                              filtersOuts_13__2, filtersOuts_13__1, 
                              filtersOuts_13__0, filtersOuts_14__7, 
                              filtersOuts_14__6, filtersOuts_14__5, 
                              filtersOuts_14__4, filtersOuts_14__3, 
                              filtersOuts_14__2, filtersOuts_14__1, 
                              filtersOuts_14__0, filtersOuts_15__7, 
                              filtersOuts_15__6, filtersOuts_15__5, 
                              filtersOuts_15__4, filtersOuts_15__3, 
                              filtersOuts_15__2, filtersOuts_15__1, 
                              filtersOuts_15__0, filtersOuts_16__7, 
                              filtersOuts_16__6, filtersOuts_16__5, 
                              filtersOuts_16__4, filtersOuts_16__3, 
                              filtersOuts_16__2, filtersOuts_16__1, 
                              filtersOuts_16__0, filtersOuts_17__7, 
                              filtersOuts_17__6, filtersOuts_17__5, 
                              filtersOuts_17__4, filtersOuts_17__3, 
                              filtersOuts_17__2, filtersOuts_17__1, 
                              filtersOuts_17__0, filtersOuts_18__7, 
                              filtersOuts_18__6, filtersOuts_18__5, 
                              filtersOuts_18__4, filtersOuts_18__3, 
                              filtersOuts_18__2, filtersOuts_18__1, 
                              filtersOuts_18__0, filtersOuts_19__7, 
                              filtersOuts_19__6, filtersOuts_19__5, 
                              filtersOuts_19__4, filtersOuts_19__3, 
                              filtersOuts_19__2, filtersOuts_19__1, 
                              filtersOuts_19__0, filtersOuts_20__7, 
                              filtersOuts_20__6, filtersOuts_20__5, 
                              filtersOuts_20__4, filtersOuts_20__3, 
                              filtersOuts_20__2, filtersOuts_20__1, 
                              filtersOuts_20__0, filtersOuts_21__7, 
                              filtersOuts_21__6, filtersOuts_21__5, 
                              filtersOuts_21__4, filtersOuts_21__3, 
                              filtersOuts_21__2, filtersOuts_21__1, 
                              filtersOuts_21__0, filtersOuts_22__7, 
                              filtersOuts_22__6, filtersOuts_22__5, 
                              filtersOuts_22__4, filtersOuts_22__3, 
                              filtersOuts_22__2, filtersOuts_22__1, 
                              filtersOuts_22__0, filtersOuts_23__7, 
                              filtersOuts_23__6, filtersOuts_23__5, 
                              filtersOuts_23__4, filtersOuts_23__3, 
                              filtersOuts_23__2, filtersOuts_23__1, 
                              filtersOuts_23__0, filtersOuts_24__7, 
                              filtersOuts_24__6, filtersOuts_24__5, 
                              filtersOuts_24__4, filtersOuts_24__3, 
                              filtersOuts_24__2, filtersOuts_24__1, 
                              filtersOuts_24__0 ) ;

    input [39:0]filterBus ;
    input [79:0]windowBus ;
    input [2:0]decoderRow ;
    input clk ;
    input rst ;
    input enablePage1Read ;
    input enablePage2Read ;
    input enableFilterRead ;
    input shift2To1 ;
    input shift1To2 ;
    input pageTurn ;
    output pagesOuts_0__15 ;
    output pagesOuts_0__14 ;
    output pagesOuts_0__13 ;
    output pagesOuts_0__12 ;
    output pagesOuts_0__11 ;
    output pagesOuts_0__10 ;
    output pagesOuts_0__9 ;
    output pagesOuts_0__8 ;
    output pagesOuts_0__7 ;
    output pagesOuts_0__6 ;
    output pagesOuts_0__5 ;
    output pagesOuts_0__4 ;
    output pagesOuts_0__3 ;
    output pagesOuts_0__2 ;
    output pagesOuts_0__1 ;
    output pagesOuts_0__0 ;
    output pagesOuts_1__15 ;
    output pagesOuts_1__14 ;
    output pagesOuts_1__13 ;
    output pagesOuts_1__12 ;
    output pagesOuts_1__11 ;
    output pagesOuts_1__10 ;
    output pagesOuts_1__9 ;
    output pagesOuts_1__8 ;
    output pagesOuts_1__7 ;
    output pagesOuts_1__6 ;
    output pagesOuts_1__5 ;
    output pagesOuts_1__4 ;
    output pagesOuts_1__3 ;
    output pagesOuts_1__2 ;
    output pagesOuts_1__1 ;
    output pagesOuts_1__0 ;
    output pagesOuts_2__15 ;
    output pagesOuts_2__14 ;
    output pagesOuts_2__13 ;
    output pagesOuts_2__12 ;
    output pagesOuts_2__11 ;
    output pagesOuts_2__10 ;
    output pagesOuts_2__9 ;
    output pagesOuts_2__8 ;
    output pagesOuts_2__7 ;
    output pagesOuts_2__6 ;
    output pagesOuts_2__5 ;
    output pagesOuts_2__4 ;
    output pagesOuts_2__3 ;
    output pagesOuts_2__2 ;
    output pagesOuts_2__1 ;
    output pagesOuts_2__0 ;
    output pagesOuts_3__15 ;
    output pagesOuts_3__14 ;
    output pagesOuts_3__13 ;
    output pagesOuts_3__12 ;
    output pagesOuts_3__11 ;
    output pagesOuts_3__10 ;
    output pagesOuts_3__9 ;
    output pagesOuts_3__8 ;
    output pagesOuts_3__7 ;
    output pagesOuts_3__6 ;
    output pagesOuts_3__5 ;
    output pagesOuts_3__4 ;
    output pagesOuts_3__3 ;
    output pagesOuts_3__2 ;
    output pagesOuts_3__1 ;
    output pagesOuts_3__0 ;
    output pagesOuts_4__15 ;
    output pagesOuts_4__14 ;
    output pagesOuts_4__13 ;
    output pagesOuts_4__12 ;
    output pagesOuts_4__11 ;
    output pagesOuts_4__10 ;
    output pagesOuts_4__9 ;
    output pagesOuts_4__8 ;
    output pagesOuts_4__7 ;
    output pagesOuts_4__6 ;
    output pagesOuts_4__5 ;
    output pagesOuts_4__4 ;
    output pagesOuts_4__3 ;
    output pagesOuts_4__2 ;
    output pagesOuts_4__1 ;
    output pagesOuts_4__0 ;
    output pagesOuts_5__15 ;
    output pagesOuts_5__14 ;
    output pagesOuts_5__13 ;
    output pagesOuts_5__12 ;
    output pagesOuts_5__11 ;
    output pagesOuts_5__10 ;
    output pagesOuts_5__9 ;
    output pagesOuts_5__8 ;
    output pagesOuts_5__7 ;
    output pagesOuts_5__6 ;
    output pagesOuts_5__5 ;
    output pagesOuts_5__4 ;
    output pagesOuts_5__3 ;
    output pagesOuts_5__2 ;
    output pagesOuts_5__1 ;
    output pagesOuts_5__0 ;
    output pagesOuts_6__15 ;
    output pagesOuts_6__14 ;
    output pagesOuts_6__13 ;
    output pagesOuts_6__12 ;
    output pagesOuts_6__11 ;
    output pagesOuts_6__10 ;
    output pagesOuts_6__9 ;
    output pagesOuts_6__8 ;
    output pagesOuts_6__7 ;
    output pagesOuts_6__6 ;
    output pagesOuts_6__5 ;
    output pagesOuts_6__4 ;
    output pagesOuts_6__3 ;
    output pagesOuts_6__2 ;
    output pagesOuts_6__1 ;
    output pagesOuts_6__0 ;
    output pagesOuts_7__15 ;
    output pagesOuts_7__14 ;
    output pagesOuts_7__13 ;
    output pagesOuts_7__12 ;
    output pagesOuts_7__11 ;
    output pagesOuts_7__10 ;
    output pagesOuts_7__9 ;
    output pagesOuts_7__8 ;
    output pagesOuts_7__7 ;
    output pagesOuts_7__6 ;
    output pagesOuts_7__5 ;
    output pagesOuts_7__4 ;
    output pagesOuts_7__3 ;
    output pagesOuts_7__2 ;
    output pagesOuts_7__1 ;
    output pagesOuts_7__0 ;
    output pagesOuts_8__15 ;
    output pagesOuts_8__14 ;
    output pagesOuts_8__13 ;
    output pagesOuts_8__12 ;
    output pagesOuts_8__11 ;
    output pagesOuts_8__10 ;
    output pagesOuts_8__9 ;
    output pagesOuts_8__8 ;
    output pagesOuts_8__7 ;
    output pagesOuts_8__6 ;
    output pagesOuts_8__5 ;
    output pagesOuts_8__4 ;
    output pagesOuts_8__3 ;
    output pagesOuts_8__2 ;
    output pagesOuts_8__1 ;
    output pagesOuts_8__0 ;
    output pagesOuts_9__15 ;
    output pagesOuts_9__14 ;
    output pagesOuts_9__13 ;
    output pagesOuts_9__12 ;
    output pagesOuts_9__11 ;
    output pagesOuts_9__10 ;
    output pagesOuts_9__9 ;
    output pagesOuts_9__8 ;
    output pagesOuts_9__7 ;
    output pagesOuts_9__6 ;
    output pagesOuts_9__5 ;
    output pagesOuts_9__4 ;
    output pagesOuts_9__3 ;
    output pagesOuts_9__2 ;
    output pagesOuts_9__1 ;
    output pagesOuts_9__0 ;
    output pagesOuts_10__15 ;
    output pagesOuts_10__14 ;
    output pagesOuts_10__13 ;
    output pagesOuts_10__12 ;
    output pagesOuts_10__11 ;
    output pagesOuts_10__10 ;
    output pagesOuts_10__9 ;
    output pagesOuts_10__8 ;
    output pagesOuts_10__7 ;
    output pagesOuts_10__6 ;
    output pagesOuts_10__5 ;
    output pagesOuts_10__4 ;
    output pagesOuts_10__3 ;
    output pagesOuts_10__2 ;
    output pagesOuts_10__1 ;
    output pagesOuts_10__0 ;
    output pagesOuts_11__15 ;
    output pagesOuts_11__14 ;
    output pagesOuts_11__13 ;
    output pagesOuts_11__12 ;
    output pagesOuts_11__11 ;
    output pagesOuts_11__10 ;
    output pagesOuts_11__9 ;
    output pagesOuts_11__8 ;
    output pagesOuts_11__7 ;
    output pagesOuts_11__6 ;
    output pagesOuts_11__5 ;
    output pagesOuts_11__4 ;
    output pagesOuts_11__3 ;
    output pagesOuts_11__2 ;
    output pagesOuts_11__1 ;
    output pagesOuts_11__0 ;
    output pagesOuts_12__15 ;
    output pagesOuts_12__14 ;
    output pagesOuts_12__13 ;
    output pagesOuts_12__12 ;
    output pagesOuts_12__11 ;
    output pagesOuts_12__10 ;
    output pagesOuts_12__9 ;
    output pagesOuts_12__8 ;
    output pagesOuts_12__7 ;
    output pagesOuts_12__6 ;
    output pagesOuts_12__5 ;
    output pagesOuts_12__4 ;
    output pagesOuts_12__3 ;
    output pagesOuts_12__2 ;
    output pagesOuts_12__1 ;
    output pagesOuts_12__0 ;
    output pagesOuts_13__15 ;
    output pagesOuts_13__14 ;
    output pagesOuts_13__13 ;
    output pagesOuts_13__12 ;
    output pagesOuts_13__11 ;
    output pagesOuts_13__10 ;
    output pagesOuts_13__9 ;
    output pagesOuts_13__8 ;
    output pagesOuts_13__7 ;
    output pagesOuts_13__6 ;
    output pagesOuts_13__5 ;
    output pagesOuts_13__4 ;
    output pagesOuts_13__3 ;
    output pagesOuts_13__2 ;
    output pagesOuts_13__1 ;
    output pagesOuts_13__0 ;
    output pagesOuts_14__15 ;
    output pagesOuts_14__14 ;
    output pagesOuts_14__13 ;
    output pagesOuts_14__12 ;
    output pagesOuts_14__11 ;
    output pagesOuts_14__10 ;
    output pagesOuts_14__9 ;
    output pagesOuts_14__8 ;
    output pagesOuts_14__7 ;
    output pagesOuts_14__6 ;
    output pagesOuts_14__5 ;
    output pagesOuts_14__4 ;
    output pagesOuts_14__3 ;
    output pagesOuts_14__2 ;
    output pagesOuts_14__1 ;
    output pagesOuts_14__0 ;
    output pagesOuts_15__15 ;
    output pagesOuts_15__14 ;
    output pagesOuts_15__13 ;
    output pagesOuts_15__12 ;
    output pagesOuts_15__11 ;
    output pagesOuts_15__10 ;
    output pagesOuts_15__9 ;
    output pagesOuts_15__8 ;
    output pagesOuts_15__7 ;
    output pagesOuts_15__6 ;
    output pagesOuts_15__5 ;
    output pagesOuts_15__4 ;
    output pagesOuts_15__3 ;
    output pagesOuts_15__2 ;
    output pagesOuts_15__1 ;
    output pagesOuts_15__0 ;
    output pagesOuts_16__15 ;
    output pagesOuts_16__14 ;
    output pagesOuts_16__13 ;
    output pagesOuts_16__12 ;
    output pagesOuts_16__11 ;
    output pagesOuts_16__10 ;
    output pagesOuts_16__9 ;
    output pagesOuts_16__8 ;
    output pagesOuts_16__7 ;
    output pagesOuts_16__6 ;
    output pagesOuts_16__5 ;
    output pagesOuts_16__4 ;
    output pagesOuts_16__3 ;
    output pagesOuts_16__2 ;
    output pagesOuts_16__1 ;
    output pagesOuts_16__0 ;
    output pagesOuts_17__15 ;
    output pagesOuts_17__14 ;
    output pagesOuts_17__13 ;
    output pagesOuts_17__12 ;
    output pagesOuts_17__11 ;
    output pagesOuts_17__10 ;
    output pagesOuts_17__9 ;
    output pagesOuts_17__8 ;
    output pagesOuts_17__7 ;
    output pagesOuts_17__6 ;
    output pagesOuts_17__5 ;
    output pagesOuts_17__4 ;
    output pagesOuts_17__3 ;
    output pagesOuts_17__2 ;
    output pagesOuts_17__1 ;
    output pagesOuts_17__0 ;
    output pagesOuts_18__15 ;
    output pagesOuts_18__14 ;
    output pagesOuts_18__13 ;
    output pagesOuts_18__12 ;
    output pagesOuts_18__11 ;
    output pagesOuts_18__10 ;
    output pagesOuts_18__9 ;
    output pagesOuts_18__8 ;
    output pagesOuts_18__7 ;
    output pagesOuts_18__6 ;
    output pagesOuts_18__5 ;
    output pagesOuts_18__4 ;
    output pagesOuts_18__3 ;
    output pagesOuts_18__2 ;
    output pagesOuts_18__1 ;
    output pagesOuts_18__0 ;
    output pagesOuts_19__15 ;
    output pagesOuts_19__14 ;
    output pagesOuts_19__13 ;
    output pagesOuts_19__12 ;
    output pagesOuts_19__11 ;
    output pagesOuts_19__10 ;
    output pagesOuts_19__9 ;
    output pagesOuts_19__8 ;
    output pagesOuts_19__7 ;
    output pagesOuts_19__6 ;
    output pagesOuts_19__5 ;
    output pagesOuts_19__4 ;
    output pagesOuts_19__3 ;
    output pagesOuts_19__2 ;
    output pagesOuts_19__1 ;
    output pagesOuts_19__0 ;
    output pagesOuts_20__15 ;
    output pagesOuts_20__14 ;
    output pagesOuts_20__13 ;
    output pagesOuts_20__12 ;
    output pagesOuts_20__11 ;
    output pagesOuts_20__10 ;
    output pagesOuts_20__9 ;
    output pagesOuts_20__8 ;
    output pagesOuts_20__7 ;
    output pagesOuts_20__6 ;
    output pagesOuts_20__5 ;
    output pagesOuts_20__4 ;
    output pagesOuts_20__3 ;
    output pagesOuts_20__2 ;
    output pagesOuts_20__1 ;
    output pagesOuts_20__0 ;
    output pagesOuts_21__15 ;
    output pagesOuts_21__14 ;
    output pagesOuts_21__13 ;
    output pagesOuts_21__12 ;
    output pagesOuts_21__11 ;
    output pagesOuts_21__10 ;
    output pagesOuts_21__9 ;
    output pagesOuts_21__8 ;
    output pagesOuts_21__7 ;
    output pagesOuts_21__6 ;
    output pagesOuts_21__5 ;
    output pagesOuts_21__4 ;
    output pagesOuts_21__3 ;
    output pagesOuts_21__2 ;
    output pagesOuts_21__1 ;
    output pagesOuts_21__0 ;
    output pagesOuts_22__15 ;
    output pagesOuts_22__14 ;
    output pagesOuts_22__13 ;
    output pagesOuts_22__12 ;
    output pagesOuts_22__11 ;
    output pagesOuts_22__10 ;
    output pagesOuts_22__9 ;
    output pagesOuts_22__8 ;
    output pagesOuts_22__7 ;
    output pagesOuts_22__6 ;
    output pagesOuts_22__5 ;
    output pagesOuts_22__4 ;
    output pagesOuts_22__3 ;
    output pagesOuts_22__2 ;
    output pagesOuts_22__1 ;
    output pagesOuts_22__0 ;
    output pagesOuts_23__15 ;
    output pagesOuts_23__14 ;
    output pagesOuts_23__13 ;
    output pagesOuts_23__12 ;
    output pagesOuts_23__11 ;
    output pagesOuts_23__10 ;
    output pagesOuts_23__9 ;
    output pagesOuts_23__8 ;
    output pagesOuts_23__7 ;
    output pagesOuts_23__6 ;
    output pagesOuts_23__5 ;
    output pagesOuts_23__4 ;
    output pagesOuts_23__3 ;
    output pagesOuts_23__2 ;
    output pagesOuts_23__1 ;
    output pagesOuts_23__0 ;
    output pagesOuts_24__15 ;
    output pagesOuts_24__14 ;
    output pagesOuts_24__13 ;
    output pagesOuts_24__12 ;
    output pagesOuts_24__11 ;
    output pagesOuts_24__10 ;
    output pagesOuts_24__9 ;
    output pagesOuts_24__8 ;
    output pagesOuts_24__7 ;
    output pagesOuts_24__6 ;
    output pagesOuts_24__5 ;
    output pagesOuts_24__4 ;
    output pagesOuts_24__3 ;
    output pagesOuts_24__2 ;
    output pagesOuts_24__1 ;
    output pagesOuts_24__0 ;
    output filtersOuts_0__7 ;
    output filtersOuts_0__6 ;
    output filtersOuts_0__5 ;
    output filtersOuts_0__4 ;
    output filtersOuts_0__3 ;
    output filtersOuts_0__2 ;
    output filtersOuts_0__1 ;
    output filtersOuts_0__0 ;
    output filtersOuts_1__7 ;
    output filtersOuts_1__6 ;
    output filtersOuts_1__5 ;
    output filtersOuts_1__4 ;
    output filtersOuts_1__3 ;
    output filtersOuts_1__2 ;
    output filtersOuts_1__1 ;
    output filtersOuts_1__0 ;
    output filtersOuts_2__7 ;
    output filtersOuts_2__6 ;
    output filtersOuts_2__5 ;
    output filtersOuts_2__4 ;
    output filtersOuts_2__3 ;
    output filtersOuts_2__2 ;
    output filtersOuts_2__1 ;
    output filtersOuts_2__0 ;
    output filtersOuts_3__7 ;
    output filtersOuts_3__6 ;
    output filtersOuts_3__5 ;
    output filtersOuts_3__4 ;
    output filtersOuts_3__3 ;
    output filtersOuts_3__2 ;
    output filtersOuts_3__1 ;
    output filtersOuts_3__0 ;
    output filtersOuts_4__7 ;
    output filtersOuts_4__6 ;
    output filtersOuts_4__5 ;
    output filtersOuts_4__4 ;
    output filtersOuts_4__3 ;
    output filtersOuts_4__2 ;
    output filtersOuts_4__1 ;
    output filtersOuts_4__0 ;
    output filtersOuts_5__7 ;
    output filtersOuts_5__6 ;
    output filtersOuts_5__5 ;
    output filtersOuts_5__4 ;
    output filtersOuts_5__3 ;
    output filtersOuts_5__2 ;
    output filtersOuts_5__1 ;
    output filtersOuts_5__0 ;
    output filtersOuts_6__7 ;
    output filtersOuts_6__6 ;
    output filtersOuts_6__5 ;
    output filtersOuts_6__4 ;
    output filtersOuts_6__3 ;
    output filtersOuts_6__2 ;
    output filtersOuts_6__1 ;
    output filtersOuts_6__0 ;
    output filtersOuts_7__7 ;
    output filtersOuts_7__6 ;
    output filtersOuts_7__5 ;
    output filtersOuts_7__4 ;
    output filtersOuts_7__3 ;
    output filtersOuts_7__2 ;
    output filtersOuts_7__1 ;
    output filtersOuts_7__0 ;
    output filtersOuts_8__7 ;
    output filtersOuts_8__6 ;
    output filtersOuts_8__5 ;
    output filtersOuts_8__4 ;
    output filtersOuts_8__3 ;
    output filtersOuts_8__2 ;
    output filtersOuts_8__1 ;
    output filtersOuts_8__0 ;
    output filtersOuts_9__7 ;
    output filtersOuts_9__6 ;
    output filtersOuts_9__5 ;
    output filtersOuts_9__4 ;
    output filtersOuts_9__3 ;
    output filtersOuts_9__2 ;
    output filtersOuts_9__1 ;
    output filtersOuts_9__0 ;
    output filtersOuts_10__7 ;
    output filtersOuts_10__6 ;
    output filtersOuts_10__5 ;
    output filtersOuts_10__4 ;
    output filtersOuts_10__3 ;
    output filtersOuts_10__2 ;
    output filtersOuts_10__1 ;
    output filtersOuts_10__0 ;
    output filtersOuts_11__7 ;
    output filtersOuts_11__6 ;
    output filtersOuts_11__5 ;
    output filtersOuts_11__4 ;
    output filtersOuts_11__3 ;
    output filtersOuts_11__2 ;
    output filtersOuts_11__1 ;
    output filtersOuts_11__0 ;
    output filtersOuts_12__7 ;
    output filtersOuts_12__6 ;
    output filtersOuts_12__5 ;
    output filtersOuts_12__4 ;
    output filtersOuts_12__3 ;
    output filtersOuts_12__2 ;
    output filtersOuts_12__1 ;
    output filtersOuts_12__0 ;
    output filtersOuts_13__7 ;
    output filtersOuts_13__6 ;
    output filtersOuts_13__5 ;
    output filtersOuts_13__4 ;
    output filtersOuts_13__3 ;
    output filtersOuts_13__2 ;
    output filtersOuts_13__1 ;
    output filtersOuts_13__0 ;
    output filtersOuts_14__7 ;
    output filtersOuts_14__6 ;
    output filtersOuts_14__5 ;
    output filtersOuts_14__4 ;
    output filtersOuts_14__3 ;
    output filtersOuts_14__2 ;
    output filtersOuts_14__1 ;
    output filtersOuts_14__0 ;
    output filtersOuts_15__7 ;
    output filtersOuts_15__6 ;
    output filtersOuts_15__5 ;
    output filtersOuts_15__4 ;
    output filtersOuts_15__3 ;
    output filtersOuts_15__2 ;
    output filtersOuts_15__1 ;
    output filtersOuts_15__0 ;
    output filtersOuts_16__7 ;
    output filtersOuts_16__6 ;
    output filtersOuts_16__5 ;
    output filtersOuts_16__4 ;
    output filtersOuts_16__3 ;
    output filtersOuts_16__2 ;
    output filtersOuts_16__1 ;
    output filtersOuts_16__0 ;
    output filtersOuts_17__7 ;
    output filtersOuts_17__6 ;
    output filtersOuts_17__5 ;
    output filtersOuts_17__4 ;
    output filtersOuts_17__3 ;
    output filtersOuts_17__2 ;
    output filtersOuts_17__1 ;
    output filtersOuts_17__0 ;
    output filtersOuts_18__7 ;
    output filtersOuts_18__6 ;
    output filtersOuts_18__5 ;
    output filtersOuts_18__4 ;
    output filtersOuts_18__3 ;
    output filtersOuts_18__2 ;
    output filtersOuts_18__1 ;
    output filtersOuts_18__0 ;
    output filtersOuts_19__7 ;
    output filtersOuts_19__6 ;
    output filtersOuts_19__5 ;
    output filtersOuts_19__4 ;
    output filtersOuts_19__3 ;
    output filtersOuts_19__2 ;
    output filtersOuts_19__1 ;
    output filtersOuts_19__0 ;
    output filtersOuts_20__7 ;
    output filtersOuts_20__6 ;
    output filtersOuts_20__5 ;
    output filtersOuts_20__4 ;
    output filtersOuts_20__3 ;
    output filtersOuts_20__2 ;
    output filtersOuts_20__1 ;
    output filtersOuts_20__0 ;
    output filtersOuts_21__7 ;
    output filtersOuts_21__6 ;
    output filtersOuts_21__5 ;
    output filtersOuts_21__4 ;
    output filtersOuts_21__3 ;
    output filtersOuts_21__2 ;
    output filtersOuts_21__1 ;
    output filtersOuts_21__0 ;
    output filtersOuts_22__7 ;
    output filtersOuts_22__6 ;
    output filtersOuts_22__5 ;
    output filtersOuts_22__4 ;
    output filtersOuts_22__3 ;
    output filtersOuts_22__2 ;
    output filtersOuts_22__1 ;
    output filtersOuts_22__0 ;
    output filtersOuts_23__7 ;
    output filtersOuts_23__6 ;
    output filtersOuts_23__5 ;
    output filtersOuts_23__4 ;
    output filtersOuts_23__3 ;
    output filtersOuts_23__2 ;
    output filtersOuts_23__1 ;
    output filtersOuts_23__0 ;
    output filtersOuts_24__7 ;
    output filtersOuts_24__6 ;
    output filtersOuts_24__5 ;
    output filtersOuts_24__4 ;
    output filtersOuts_24__3 ;
    output filtersOuts_24__2 ;
    output filtersOuts_24__1 ;
    output filtersOuts_24__0 ;

    wire page1Out_5__15, page1Out_5__14, page1Out_5__13, page1Out_5__12, 
         page1Out_5__11, page1Out_5__10, page1Out_5__9, page1Out_5__8, 
         page1Out_5__7, page1Out_5__6, page1Out_5__5, page1Out_5__4, 
         page1Out_5__3, page1Out_5__2, page1Out_5__1, page1Out_5__0, 
         page1Out_6__15, page1Out_6__14, page1Out_6__13, page1Out_6__12, 
         page1Out_6__11, page1Out_6__10, page1Out_6__9, page1Out_6__8, 
         page1Out_6__7, page1Out_6__6, page1Out_6__5, page1Out_6__4, 
         page1Out_6__3, page1Out_6__2, page1Out_6__1, page1Out_6__0, 
         page1Out_7__15, page1Out_7__14, page1Out_7__13, page1Out_7__12, 
         page1Out_7__11, page1Out_7__10, page1Out_7__9, page1Out_7__8, 
         page1Out_7__7, page1Out_7__6, page1Out_7__5, page1Out_7__4, 
         page1Out_7__3, page1Out_7__2, page1Out_7__1, page1Out_7__0, 
         page1Out_8__15, page1Out_8__14, page1Out_8__13, page1Out_8__12, 
         page1Out_8__11, page1Out_8__10, page1Out_8__9, page1Out_8__8, 
         page1Out_8__7, page1Out_8__6, page1Out_8__5, page1Out_8__4, 
         page1Out_8__3, page1Out_8__2, page1Out_8__1, page1Out_8__0, 
         page1Out_9__15, page1Out_9__14, page1Out_9__13, page1Out_9__12, 
         page1Out_9__11, page1Out_9__10, page1Out_9__9, page1Out_9__8, 
         page1Out_9__7, page1Out_9__6, page1Out_9__5, page1Out_9__4, 
         page1Out_9__3, page1Out_9__2, page1Out_9__1, page1Out_9__0, 
         page1Out_10__15, page1Out_10__14, page1Out_10__13, page1Out_10__12, 
         page1Out_10__11, page1Out_10__10, page1Out_10__9, page1Out_10__8, 
         page1Out_10__7, page1Out_10__6, page1Out_10__5, page1Out_10__4, 
         page1Out_10__3, page1Out_10__2, page1Out_10__1, page1Out_10__0, 
         page1Out_11__15, page1Out_11__14, page1Out_11__13, page1Out_11__12, 
         page1Out_11__11, page1Out_11__10, page1Out_11__9, page1Out_11__8, 
         page1Out_11__7, page1Out_11__6, page1Out_11__5, page1Out_11__4, 
         page1Out_11__3, page1Out_11__2, page1Out_11__1, page1Out_11__0, 
         page1Out_12__15, page1Out_12__14, page1Out_12__13, page1Out_12__12, 
         page1Out_12__11, page1Out_12__10, page1Out_12__9, page1Out_12__8, 
         page1Out_12__7, page1Out_12__6, page1Out_12__5, page1Out_12__4, 
         page1Out_12__3, page1Out_12__2, page1Out_12__1, page1Out_12__0, 
         page1Out_13__15, page1Out_13__14, page1Out_13__13, page1Out_13__12, 
         page1Out_13__11, page1Out_13__10, page1Out_13__9, page1Out_13__8, 
         page1Out_13__7, page1Out_13__6, page1Out_13__5, page1Out_13__4, 
         page1Out_13__3, page1Out_13__2, page1Out_13__1, page1Out_13__0, 
         page1Out_14__15, page1Out_14__14, page1Out_14__13, page1Out_14__12, 
         page1Out_14__11, page1Out_14__10, page1Out_14__9, page1Out_14__8, 
         page1Out_14__7, page1Out_14__6, page1Out_14__5, page1Out_14__4, 
         page1Out_14__3, page1Out_14__2, page1Out_14__1, page1Out_14__0, 
         page1Out_15__15, page1Out_15__14, page1Out_15__13, page1Out_15__12, 
         page1Out_15__11, page1Out_15__10, page1Out_15__9, page1Out_15__8, 
         page1Out_15__7, page1Out_15__6, page1Out_15__5, page1Out_15__4, 
         page1Out_15__3, page1Out_15__2, page1Out_15__1, page1Out_15__0, 
         page1Out_16__15, page1Out_16__14, page1Out_16__13, page1Out_16__12, 
         page1Out_16__11, page1Out_16__10, page1Out_16__9, page1Out_16__8, 
         page1Out_16__7, page1Out_16__6, page1Out_16__5, page1Out_16__4, 
         page1Out_16__3, page1Out_16__2, page1Out_16__1, page1Out_16__0, 
         page1Out_17__15, page1Out_17__14, page1Out_17__13, page1Out_17__12, 
         page1Out_17__11, page1Out_17__10, page1Out_17__9, page1Out_17__8, 
         page1Out_17__7, page1Out_17__6, page1Out_17__5, page1Out_17__4, 
         page1Out_17__3, page1Out_17__2, page1Out_17__1, page1Out_17__0, 
         page1Out_18__15, page1Out_18__14, page1Out_18__13, page1Out_18__12, 
         page1Out_18__11, page1Out_18__10, page1Out_18__9, page1Out_18__8, 
         page1Out_18__7, page1Out_18__6, page1Out_18__5, page1Out_18__4, 
         page1Out_18__3, page1Out_18__2, page1Out_18__1, page1Out_18__0, 
         page1Out_19__15, page1Out_19__14, page1Out_19__13, page1Out_19__12, 
         page1Out_19__11, page1Out_19__10, page1Out_19__9, page1Out_19__8, 
         page1Out_19__7, page1Out_19__6, page1Out_19__5, page1Out_19__4, 
         page1Out_19__3, page1Out_19__2, page1Out_19__1, page1Out_19__0, 
         page1Out_20__15, page1Out_20__14, page1Out_20__13, page1Out_20__12, 
         page1Out_20__11, page1Out_20__10, page1Out_20__9, page1Out_20__8, 
         page1Out_20__7, page1Out_20__6, page1Out_20__5, page1Out_20__4, 
         page1Out_20__3, page1Out_20__2, page1Out_20__1, page1Out_20__0, 
         page1Out_21__15, page1Out_21__14, page1Out_21__13, page1Out_21__12, 
         page1Out_21__11, page1Out_21__10, page1Out_21__9, page1Out_21__8, 
         page1Out_21__7, page1Out_21__6, page1Out_21__5, page1Out_21__4, 
         page1Out_21__3, page1Out_21__2, page1Out_21__1, page1Out_21__0, 
         page1Out_22__15, page1Out_22__14, page1Out_22__13, page1Out_22__12, 
         page1Out_22__11, page1Out_22__10, page1Out_22__9, page1Out_22__8, 
         page1Out_22__7, page1Out_22__6, page1Out_22__5, page1Out_22__4, 
         page1Out_22__3, page1Out_22__2, page1Out_22__1, page1Out_22__0, 
         page1Out_23__15, page1Out_23__14, page1Out_23__13, page1Out_23__12, 
         page1Out_23__11, page1Out_23__10, page1Out_23__9, page1Out_23__8, 
         page1Out_23__7, page1Out_23__6, page1Out_23__5, page1Out_23__4, 
         page1Out_23__3, page1Out_23__2, page1Out_23__1, page1Out_23__0, 
         page1Out_24__15, page1Out_24__14, page1Out_24__13, page1Out_24__12, 
         page1Out_24__11, page1Out_24__10, page1Out_24__9, page1Out_24__8, 
         page1Out_24__7, page1Out_24__6, page1Out_24__5, page1Out_24__4, 
         page1Out_24__3, page1Out_24__2, page1Out_24__1, page1Out_24__0, 
         page2Out_5__15, page2Out_5__14, page2Out_5__13, page2Out_5__12, 
         page2Out_5__11, page2Out_5__10, page2Out_5__9, page2Out_5__8, 
         page2Out_5__7, page2Out_5__6, page2Out_5__5, page2Out_5__4, 
         page2Out_5__3, page2Out_5__2, page2Out_5__1, page2Out_5__0, 
         page2Out_6__15, page2Out_6__14, page2Out_6__13, page2Out_6__12, 
         page2Out_6__11, page2Out_6__10, page2Out_6__9, page2Out_6__8, 
         page2Out_6__7, page2Out_6__6, page2Out_6__5, page2Out_6__4, 
         page2Out_6__3, page2Out_6__2, page2Out_6__1, page2Out_6__0, 
         page2Out_7__15, page2Out_7__14, page2Out_7__13, page2Out_7__12, 
         page2Out_7__11, page2Out_7__10, page2Out_7__9, page2Out_7__8, 
         page2Out_7__7, page2Out_7__6, page2Out_7__5, page2Out_7__4, 
         page2Out_7__3, page2Out_7__2, page2Out_7__1, page2Out_7__0, 
         page2Out_8__15, page2Out_8__14, page2Out_8__13, page2Out_8__12, 
         page2Out_8__11, page2Out_8__10, page2Out_8__9, page2Out_8__8, 
         page2Out_8__7, page2Out_8__6, page2Out_8__5, page2Out_8__4, 
         page2Out_8__3, page2Out_8__2, page2Out_8__1, page2Out_8__0, 
         page2Out_9__15, page2Out_9__14, page2Out_9__13, page2Out_9__12, 
         page2Out_9__11, page2Out_9__10, page2Out_9__9, page2Out_9__8, 
         page2Out_9__7, page2Out_9__6, page2Out_9__5, page2Out_9__4, 
         page2Out_9__3, page2Out_9__2, page2Out_9__1, page2Out_9__0, 
         page2Out_10__15, page2Out_10__14, page2Out_10__13, page2Out_10__12, 
         page2Out_10__11, page2Out_10__10, page2Out_10__9, page2Out_10__8, 
         page2Out_10__7, page2Out_10__6, page2Out_10__5, page2Out_10__4, 
         page2Out_10__3, page2Out_10__2, page2Out_10__1, page2Out_10__0, 
         page2Out_11__15, page2Out_11__14, page2Out_11__13, page2Out_11__12, 
         page2Out_11__11, page2Out_11__10, page2Out_11__9, page2Out_11__8, 
         page2Out_11__7, page2Out_11__6, page2Out_11__5, page2Out_11__4, 
         page2Out_11__3, page2Out_11__2, page2Out_11__1, page2Out_11__0, 
         page2Out_12__15, page2Out_12__14, page2Out_12__13, page2Out_12__12, 
         page2Out_12__11, page2Out_12__10, page2Out_12__9, page2Out_12__8, 
         page2Out_12__7, page2Out_12__6, page2Out_12__5, page2Out_12__4, 
         page2Out_12__3, page2Out_12__2, page2Out_12__1, page2Out_12__0, 
         page2Out_13__15, page2Out_13__14, page2Out_13__13, page2Out_13__12, 
         page2Out_13__11, page2Out_13__10, page2Out_13__9, page2Out_13__8, 
         page2Out_13__7, page2Out_13__6, page2Out_13__5, page2Out_13__4, 
         page2Out_13__3, page2Out_13__2, page2Out_13__1, page2Out_13__0, 
         page2Out_14__15, page2Out_14__14, page2Out_14__13, page2Out_14__12, 
         page2Out_14__11, page2Out_14__10, page2Out_14__9, page2Out_14__8, 
         page2Out_14__7, page2Out_14__6, page2Out_14__5, page2Out_14__4, 
         page2Out_14__3, page2Out_14__2, page2Out_14__1, page2Out_14__0, 
         page2Out_15__15, page2Out_15__14, page2Out_15__13, page2Out_15__12, 
         page2Out_15__11, page2Out_15__10, page2Out_15__9, page2Out_15__8, 
         page2Out_15__7, page2Out_15__6, page2Out_15__5, page2Out_15__4, 
         page2Out_15__3, page2Out_15__2, page2Out_15__1, page2Out_15__0, 
         page2Out_16__15, page2Out_16__14, page2Out_16__13, page2Out_16__12, 
         page2Out_16__11, page2Out_16__10, page2Out_16__9, page2Out_16__8, 
         page2Out_16__7, page2Out_16__6, page2Out_16__5, page2Out_16__4, 
         page2Out_16__3, page2Out_16__2, page2Out_16__1, page2Out_16__0, 
         page2Out_17__15, page2Out_17__14, page2Out_17__13, page2Out_17__12, 
         page2Out_17__11, page2Out_17__10, page2Out_17__9, page2Out_17__8, 
         page2Out_17__7, page2Out_17__6, page2Out_17__5, page2Out_17__4, 
         page2Out_17__3, page2Out_17__2, page2Out_17__1, page2Out_17__0, 
         page2Out_18__15, page2Out_18__14, page2Out_18__13, page2Out_18__12, 
         page2Out_18__11, page2Out_18__10, page2Out_18__9, page2Out_18__8, 
         page2Out_18__7, page2Out_18__6, page2Out_18__5, page2Out_18__4, 
         page2Out_18__3, page2Out_18__2, page2Out_18__1, page2Out_18__0, 
         page2Out_19__15, page2Out_19__14, page2Out_19__13, page2Out_19__12, 
         page2Out_19__11, page2Out_19__10, page2Out_19__9, page2Out_19__8, 
         page2Out_19__7, page2Out_19__6, page2Out_19__5, page2Out_19__4, 
         page2Out_19__3, page2Out_19__2, page2Out_19__1, page2Out_19__0, 
         page2Out_20__15, page2Out_20__14, page2Out_20__13, page2Out_20__12, 
         page2Out_20__11, page2Out_20__10, page2Out_20__9, page2Out_20__8, 
         page2Out_20__7, page2Out_20__6, page2Out_20__5, page2Out_20__4, 
         page2Out_20__3, page2Out_20__2, page2Out_20__1, page2Out_20__0, 
         page2Out_21__15, page2Out_21__14, page2Out_21__13, page2Out_21__12, 
         page2Out_21__11, page2Out_21__10, page2Out_21__9, page2Out_21__8, 
         page2Out_21__7, page2Out_21__6, page2Out_21__5, page2Out_21__4, 
         page2Out_21__3, page2Out_21__2, page2Out_21__1, page2Out_21__0, 
         page2Out_22__15, page2Out_22__14, page2Out_22__13, page2Out_22__12, 
         page2Out_22__11, page2Out_22__10, page2Out_22__9, page2Out_22__8, 
         page2Out_22__7, page2Out_22__6, page2Out_22__5, page2Out_22__4, 
         page2Out_22__3, page2Out_22__2, page2Out_22__1, page2Out_22__0, 
         page2Out_23__15, page2Out_23__14, page2Out_23__13, page2Out_23__12, 
         page2Out_23__11, page2Out_23__10, page2Out_23__9, page2Out_23__8, 
         page2Out_23__7, page2Out_23__6, page2Out_23__5, page2Out_23__4, 
         page2Out_23__3, page2Out_23__2, page2Out_23__1, page2Out_23__0, 
         page2Out_24__15, page2Out_24__14, page2Out_24__13, page2Out_24__12, 
         page2Out_24__11, page2Out_24__10, page2Out_24__9, page2Out_24__8, 
         page2Out_24__7, page2Out_24__6, page2Out_24__5, page2Out_24__4, 
         page2Out_24__3, page2Out_24__2, page2Out_24__1, page2Out_24__0, 
         page1Enables_0, page1Enables_1, page1Enables_2, page1Enables_3, 
         page1Enables_4, page2Enables_0, page2Enables_1, page2Enables_2, 
         page2Enables_3, page2Enables_4, filterEnables_0, filterEnables_1, 
         filterEnables_2, filterEnables_3, filterEnables_4, decodedRow_4, 
         decodedRow_3, decodedRow_2, decodedRow_1, decodedRow_0, 
         decoderRowEnable, page1Out_25__15, nx2788, nx2790, nx2792, nx2794, 
         nx2796, nx2798, nx2800, nx2802, nx2804, nx2806, nx2808, nx2810, nx2812, 
         nx2814, nx2816, nx2818, nx2820, nx2822, nx2824, nx2826, nx2828, nx2830, 
         nx2832, nx2834, nx2836, nx2838, nx2840, nx2842, nx2844, nx2846, nx2848, 
         nx2850, nx2852, nx2854, nx2856, nx2858, nx2860, nx2862, nx2864, nx2866, 
         nx2868, nx2870, nx2872, nx2874, nx2876, nx2878, nx2880, nx2882, nx2884, 
         nx2886, nx2888, nx2890, nx2892, nx2894, nx2896, nx2898, nx2900, nx2902, 
         nx2904, nx2906, nx2908, nx2910, nx2912, nx2914, nx2916, nx2918, nx2920, 
         nx2922, nx2924, nx2926, nx2928, nx2930, nx2932, nx2934, nx2936, nx2938, 
         nx2940, nx2942, nx2944, nx2946, nx2948, nx2950, nx2952, nx2954, nx2956, 
         nx2958, nx2960, nx2962, nx2964, nx2966, nx2968, nx2970, nx2972, nx2974, 
         nx2976, nx2978, nx2980, nx2982, nx2984, nx2986, nx2988, nx2990, nx2992, 
         nx2994, nx2996, nx2998, nx3000, nx3002, nx3004, nx3006, nx3008, nx3010, 
         nx3012, nx3014, nx3016, nx3018, nx3020, nx3022, nx3024, nx3026, nx3028, 
         nx3030, nx3032, nx3034, nx3036, nx3038, nx3040, nx3042, nx3044, nx3046, 
         nx3048, nx3050, nx3052, nx3054, nx3056, nx3058, nx3060, nx3062, nx3064, 
         nx3066, nx3068, nx3070, nx3072, nx3074, nx3076, nx3078, nx3080, nx3082, 
         nx3084, nx3086, nx3088, nx3090, nx3092, nx3094, nx3096, nx3098, nx3100, 
         nx3102, nx3104, nx3106, nx3108, nx3110, nx3112, nx3114, nx3116, nx3118, 
         nx3120, nx3122, nx3124, nx3126;
    wire [162:0] \$dummy ;




    Decoder_3 decoderRowMap (.T ({decoderRow[2],decoderRow[1],decoderRow[0]}), .en (
              decoderRowEnable), .decoded ({\$dummy [0],\$dummy [1],\$dummy [2],
              decodedRow_4,decodedRow_3,decodedRow_2,decodedRow_1,decodedRow_0})
              ) ;
    RegRow_8_16_5_3 loop1_0_regRowMap (.filterBus ({filterBus[39],filterBus[38],
                    filterBus[37],filterBus[36],filterBus[35],filterBus[34],
                    filterBus[33],filterBus[32],filterBus[31],filterBus[30],
                    filterBus[29],filterBus[28],filterBus[27],filterBus[26],
                    filterBus[25],filterBus[24],filterBus[23],filterBus[22],
                    filterBus[21],filterBus[20],filterBus[19],filterBus[18],
                    filterBus[17],filterBus[16],filterBus[15],filterBus[14],
                    filterBus[13],filterBus[12],filterBus[11],filterBus[10],
                    filterBus[9],filterBus[8],filterBus[7],filterBus[6],
                    filterBus[5],filterBus[4],filterBus[3],filterBus[2],
                    filterBus[1],filterBus[0]}), .windowBus ({nx2800,nx2804,
                    nx2808,nx2812,nx2816,nx2820,nx2824,nx2828,nx2832,nx2836,
                    nx2840,nx2844,nx2848,nx2852,nx2856,nx2860,nx2864,nx2868,
                    nx2872,nx2876,nx2880,nx2884,nx2888,nx2892,nx2896,nx2900,
                    nx2904,nx2908,nx2912,nx2916,nx2920,nx2924,nx2928,nx2932,
                    nx2936,nx2940,nx2944,nx2948,nx2952,nx2956,nx2960,nx2964,
                    nx2968,nx2972,nx2976,nx2980,nx2984,nx2988,nx2992,nx2996,
                    nx3000,nx3004,nx3008,nx3012,nx3016,nx3020,nx3024,nx3028,
                    nx3032,nx3036,nx3040,nx3044,nx3048,nx3052,nx3056,nx3060,
                    nx3064,nx3068,nx3072,nx3076,nx3080,nx3084,nx3088,nx3092,
                    nx3096,nx3100,nx3104,nx3108,nx3112,nx3116}), .page1NextRow_0__15 (
                    page1Out_5__15), .page1NextRow_0__14 (page1Out_5__14), .page1NextRow_0__13 (
                    page1Out_5__13), .page1NextRow_0__12 (page1Out_5__12), .page1NextRow_0__11 (
                    page1Out_5__11), .page1NextRow_0__10 (page1Out_5__10), .page1NextRow_0__9 (
                    page1Out_5__9), .page1NextRow_0__8 (page1Out_5__8), .page1NextRow_0__7 (
                    page1Out_5__7), .page1NextRow_0__6 (page1Out_5__6), .page1NextRow_0__5 (
                    page1Out_5__5), .page1NextRow_0__4 (page1Out_5__4), .page1NextRow_0__3 (
                    page1Out_5__3), .page1NextRow_0__2 (page1Out_5__2), .page1NextRow_0__1 (
                    page1Out_5__1), .page1NextRow_0__0 (page1Out_5__0), .page1NextRow_1__15 (
                    page1Out_6__15), .page1NextRow_1__14 (page1Out_6__14), .page1NextRow_1__13 (
                    page1Out_6__13), .page1NextRow_1__12 (page1Out_6__12), .page1NextRow_1__11 (
                    page1Out_6__11), .page1NextRow_1__10 (page1Out_6__10), .page1NextRow_1__9 (
                    page1Out_6__9), .page1NextRow_1__8 (page1Out_6__8), .page1NextRow_1__7 (
                    page1Out_6__7), .page1NextRow_1__6 (page1Out_6__6), .page1NextRow_1__5 (
                    page1Out_6__5), .page1NextRow_1__4 (page1Out_6__4), .page1NextRow_1__3 (
                    page1Out_6__3), .page1NextRow_1__2 (page1Out_6__2), .page1NextRow_1__1 (
                    page1Out_6__1), .page1NextRow_1__0 (page1Out_6__0), .page1NextRow_2__15 (
                    page1Out_7__15), .page1NextRow_2__14 (page1Out_7__14), .page1NextRow_2__13 (
                    page1Out_7__13), .page1NextRow_2__12 (page1Out_7__12), .page1NextRow_2__11 (
                    page1Out_7__11), .page1NextRow_2__10 (page1Out_7__10), .page1NextRow_2__9 (
                    page1Out_7__9), .page1NextRow_2__8 (page1Out_7__8), .page1NextRow_2__7 (
                    page1Out_7__7), .page1NextRow_2__6 (page1Out_7__6), .page1NextRow_2__5 (
                    page1Out_7__5), .page1NextRow_2__4 (page1Out_7__4), .page1NextRow_2__3 (
                    page1Out_7__3), .page1NextRow_2__2 (page1Out_7__2), .page1NextRow_2__1 (
                    page1Out_7__1), .page1NextRow_2__0 (page1Out_7__0), .page1NextRow_3__15 (
                    page1Out_8__15), .page1NextRow_3__14 (page1Out_8__14), .page1NextRow_3__13 (
                    page1Out_8__13), .page1NextRow_3__12 (page1Out_8__12), .page1NextRow_3__11 (
                    page1Out_8__11), .page1NextRow_3__10 (page1Out_8__10), .page1NextRow_3__9 (
                    page1Out_8__9), .page1NextRow_3__8 (page1Out_8__8), .page1NextRow_3__7 (
                    page1Out_8__7), .page1NextRow_3__6 (page1Out_8__6), .page1NextRow_3__5 (
                    page1Out_8__5), .page1NextRow_3__4 (page1Out_8__4), .page1NextRow_3__3 (
                    page1Out_8__3), .page1NextRow_3__2 (page1Out_8__2), .page1NextRow_3__1 (
                    page1Out_8__1), .page1NextRow_3__0 (page1Out_8__0), .page1NextRow_4__15 (
                    page1Out_9__15), .page1NextRow_4__14 (page1Out_9__14), .page1NextRow_4__13 (
                    page1Out_9__13), .page1NextRow_4__12 (page1Out_9__12), .page1NextRow_4__11 (
                    page1Out_9__11), .page1NextRow_4__10 (page1Out_9__10), .page1NextRow_4__9 (
                    page1Out_9__9), .page1NextRow_4__8 (page1Out_9__8), .page1NextRow_4__7 (
                    page1Out_9__7), .page1NextRow_4__6 (page1Out_9__6), .page1NextRow_4__5 (
                    page1Out_9__5), .page1NextRow_4__4 (page1Out_9__4), .page1NextRow_4__3 (
                    page1Out_9__3), .page1NextRow_4__2 (page1Out_9__2), .page1NextRow_4__1 (
                    page1Out_9__1), .page1NextRow_4__0 (page1Out_9__0), .page2NextRow_0__15 (
                    page2Out_5__15), .page2NextRow_0__14 (page2Out_5__14), .page2NextRow_0__13 (
                    page2Out_5__13), .page2NextRow_0__12 (page2Out_5__12), .page2NextRow_0__11 (
                    page2Out_5__11), .page2NextRow_0__10 (page2Out_5__10), .page2NextRow_0__9 (
                    page2Out_5__9), .page2NextRow_0__8 (page2Out_5__8), .page2NextRow_0__7 (
                    page2Out_5__7), .page2NextRow_0__6 (page2Out_5__6), .page2NextRow_0__5 (
                    page2Out_5__5), .page2NextRow_0__4 (page2Out_5__4), .page2NextRow_0__3 (
                    page2Out_5__3), .page2NextRow_0__2 (page2Out_5__2), .page2NextRow_0__1 (
                    page2Out_5__1), .page2NextRow_0__0 (page2Out_5__0), .page2NextRow_1__15 (
                    page2Out_6__15), .page2NextRow_1__14 (page2Out_6__14), .page2NextRow_1__13 (
                    page2Out_6__13), .page2NextRow_1__12 (page2Out_6__12), .page2NextRow_1__11 (
                    page2Out_6__11), .page2NextRow_1__10 (page2Out_6__10), .page2NextRow_1__9 (
                    page2Out_6__9), .page2NextRow_1__8 (page2Out_6__8), .page2NextRow_1__7 (
                    page2Out_6__7), .page2NextRow_1__6 (page2Out_6__6), .page2NextRow_1__5 (
                    page2Out_6__5), .page2NextRow_1__4 (page2Out_6__4), .page2NextRow_1__3 (
                    page2Out_6__3), .page2NextRow_1__2 (page2Out_6__2), .page2NextRow_1__1 (
                    page2Out_6__1), .page2NextRow_1__0 (page2Out_6__0), .page2NextRow_2__15 (
                    page2Out_7__15), .page2NextRow_2__14 (page2Out_7__14), .page2NextRow_2__13 (
                    page2Out_7__13), .page2NextRow_2__12 (page2Out_7__12), .page2NextRow_2__11 (
                    page2Out_7__11), .page2NextRow_2__10 (page2Out_7__10), .page2NextRow_2__9 (
                    page2Out_7__9), .page2NextRow_2__8 (page2Out_7__8), .page2NextRow_2__7 (
                    page2Out_7__7), .page2NextRow_2__6 (page2Out_7__6), .page2NextRow_2__5 (
                    page2Out_7__5), .page2NextRow_2__4 (page2Out_7__4), .page2NextRow_2__3 (
                    page2Out_7__3), .page2NextRow_2__2 (page2Out_7__2), .page2NextRow_2__1 (
                    page2Out_7__1), .page2NextRow_2__0 (page2Out_7__0), .page2NextRow_3__15 (
                    page2Out_8__15), .page2NextRow_3__14 (page2Out_8__14), .page2NextRow_3__13 (
                    page2Out_8__13), .page2NextRow_3__12 (page2Out_8__12), .page2NextRow_3__11 (
                    page2Out_8__11), .page2NextRow_3__10 (page2Out_8__10), .page2NextRow_3__9 (
                    page2Out_8__9), .page2NextRow_3__8 (page2Out_8__8), .page2NextRow_3__7 (
                    page2Out_8__7), .page2NextRow_3__6 (page2Out_8__6), .page2NextRow_3__5 (
                    page2Out_8__5), .page2NextRow_3__4 (page2Out_8__4), .page2NextRow_3__3 (
                    page2Out_8__3), .page2NextRow_3__2 (page2Out_8__2), .page2NextRow_3__1 (
                    page2Out_8__1), .page2NextRow_3__0 (page2Out_8__0), .page2NextRow_4__15 (
                    page2Out_9__15), .page2NextRow_4__14 (page2Out_9__14), .page2NextRow_4__13 (
                    page2Out_9__13), .page2NextRow_4__12 (page2Out_9__12), .page2NextRow_4__11 (
                    page2Out_9__11), .page2NextRow_4__10 (page2Out_9__10), .page2NextRow_4__9 (
                    page2Out_9__9), .page2NextRow_4__8 (page2Out_9__8), .page2NextRow_4__7 (
                    page2Out_9__7), .page2NextRow_4__6 (page2Out_9__6), .page2NextRow_4__5 (
                    page2Out_9__5), .page2NextRow_4__4 (page2Out_9__4), .page2NextRow_4__3 (
                    page2Out_9__3), .page2NextRow_4__2 (page2Out_9__2), .page2NextRow_4__1 (
                    page2Out_9__1), .page2NextRow_4__0 (page2Out_9__0), .clk (
                    clk), .rst (rst), .enablePage1Read (page1Enables_0), .enablePage2Read (
                    page2Enables_0), .enableFilterRead (filterEnables_0), .shift2To1 (
                    nx3120), .shift1To2 (nx3124), .pageTurn (nx2790), .page1Out_0__15 (
                    \$dummy [3]), .page1Out_0__14 (\$dummy [4]), .page1Out_0__13 (
                    \$dummy [5]), .page1Out_0__12 (\$dummy [6]), .page1Out_0__11 (
                    \$dummy [7]), .page1Out_0__10 (\$dummy [8]), .page1Out_0__9 (
                    \$dummy [9]), .page1Out_0__8 (\$dummy [10]), .page1Out_0__7 (
                    \$dummy [11]), .page1Out_0__6 (\$dummy [12]), .page1Out_0__5 (
                    \$dummy [13]), .page1Out_0__4 (\$dummy [14]), .page1Out_0__3 (
                    \$dummy [15]), .page1Out_0__2 (\$dummy [16]), .page1Out_0__1 (
                    \$dummy [17]), .page1Out_0__0 (\$dummy [18]), .page1Out_1__15 (
                    \$dummy [19]), .page1Out_1__14 (\$dummy [20]), .page1Out_1__13 (
                    \$dummy [21]), .page1Out_1__12 (\$dummy [22]), .page1Out_1__11 (
                    \$dummy [23]), .page1Out_1__10 (\$dummy [24]), .page1Out_1__9 (
                    \$dummy [25]), .page1Out_1__8 (\$dummy [26]), .page1Out_1__7 (
                    \$dummy [27]), .page1Out_1__6 (\$dummy [28]), .page1Out_1__5 (
                    \$dummy [29]), .page1Out_1__4 (\$dummy [30]), .page1Out_1__3 (
                    \$dummy [31]), .page1Out_1__2 (\$dummy [32]), .page1Out_1__1 (
                    \$dummy [33]), .page1Out_1__0 (\$dummy [34]), .page1Out_2__15 (
                    \$dummy [35]), .page1Out_2__14 (\$dummy [36]), .page1Out_2__13 (
                    \$dummy [37]), .page1Out_2__12 (\$dummy [38]), .page1Out_2__11 (
                    \$dummy [39]), .page1Out_2__10 (\$dummy [40]), .page1Out_2__9 (
                    \$dummy [41]), .page1Out_2__8 (\$dummy [42]), .page1Out_2__7 (
                    \$dummy [43]), .page1Out_2__6 (\$dummy [44]), .page1Out_2__5 (
                    \$dummy [45]), .page1Out_2__4 (\$dummy [46]), .page1Out_2__3 (
                    \$dummy [47]), .page1Out_2__2 (\$dummy [48]), .page1Out_2__1 (
                    \$dummy [49]), .page1Out_2__0 (\$dummy [50]), .page1Out_3__15 (
                    \$dummy [51]), .page1Out_3__14 (\$dummy [52]), .page1Out_3__13 (
                    \$dummy [53]), .page1Out_3__12 (\$dummy [54]), .page1Out_3__11 (
                    \$dummy [55]), .page1Out_3__10 (\$dummy [56]), .page1Out_3__9 (
                    \$dummy [57]), .page1Out_3__8 (\$dummy [58]), .page1Out_3__7 (
                    \$dummy [59]), .page1Out_3__6 (\$dummy [60]), .page1Out_3__5 (
                    \$dummy [61]), .page1Out_3__4 (\$dummy [62]), .page1Out_3__3 (
                    \$dummy [63]), .page1Out_3__2 (\$dummy [64]), .page1Out_3__1 (
                    \$dummy [65]), .page1Out_3__0 (\$dummy [66]), .page1Out_4__15 (
                    \$dummy [67]), .page1Out_4__14 (\$dummy [68]), .page1Out_4__13 (
                    \$dummy [69]), .page1Out_4__12 (\$dummy [70]), .page1Out_4__11 (
                    \$dummy [71]), .page1Out_4__10 (\$dummy [72]), .page1Out_4__9 (
                    \$dummy [73]), .page1Out_4__8 (\$dummy [74]), .page1Out_4__7 (
                    \$dummy [75]), .page1Out_4__6 (\$dummy [76]), .page1Out_4__5 (
                    \$dummy [77]), .page1Out_4__4 (\$dummy [78]), .page1Out_4__3 (
                    \$dummy [79]), .page1Out_4__2 (\$dummy [80]), .page1Out_4__1 (
                    \$dummy [81]), .page1Out_4__0 (\$dummy [82]), .page2Out_0__15 (
                    \$dummy [83]), .page2Out_0__14 (\$dummy [84]), .page2Out_0__13 (
                    \$dummy [85]), .page2Out_0__12 (\$dummy [86]), .page2Out_0__11 (
                    \$dummy [87]), .page2Out_0__10 (\$dummy [88]), .page2Out_0__9 (
                    \$dummy [89]), .page2Out_0__8 (\$dummy [90]), .page2Out_0__7 (
                    \$dummy [91]), .page2Out_0__6 (\$dummy [92]), .page2Out_0__5 (
                    \$dummy [93]), .page2Out_0__4 (\$dummy [94]), .page2Out_0__3 (
                    \$dummy [95]), .page2Out_0__2 (\$dummy [96]), .page2Out_0__1 (
                    \$dummy [97]), .page2Out_0__0 (\$dummy [98]), .page2Out_1__15 (
                    \$dummy [99]), .page2Out_1__14 (\$dummy [100]), .page2Out_1__13 (
                    \$dummy [101]), .page2Out_1__12 (\$dummy [102]), .page2Out_1__11 (
                    \$dummy [103]), .page2Out_1__10 (\$dummy [104]), .page2Out_1__9 (
                    \$dummy [105]), .page2Out_1__8 (\$dummy [106]), .page2Out_1__7 (
                    \$dummy [107]), .page2Out_1__6 (\$dummy [108]), .page2Out_1__5 (
                    \$dummy [109]), .page2Out_1__4 (\$dummy [110]), .page2Out_1__3 (
                    \$dummy [111]), .page2Out_1__2 (\$dummy [112]), .page2Out_1__1 (
                    \$dummy [113]), .page2Out_1__0 (\$dummy [114]), .page2Out_2__15 (
                    \$dummy [115]), .page2Out_2__14 (\$dummy [116]), .page2Out_2__13 (
                    \$dummy [117]), .page2Out_2__12 (\$dummy [118]), .page2Out_2__11 (
                    \$dummy [119]), .page2Out_2__10 (\$dummy [120]), .page2Out_2__9 (
                    \$dummy [121]), .page2Out_2__8 (\$dummy [122]), .page2Out_2__7 (
                    \$dummy [123]), .page2Out_2__6 (\$dummy [124]), .page2Out_2__5 (
                    \$dummy [125]), .page2Out_2__4 (\$dummy [126]), .page2Out_2__3 (
                    \$dummy [127]), .page2Out_2__2 (\$dummy [128]), .page2Out_2__1 (
                    \$dummy [129]), .page2Out_2__0 (\$dummy [130]), .page2Out_3__15 (
                    \$dummy [131]), .page2Out_3__14 (\$dummy [132]), .page2Out_3__13 (
                    \$dummy [133]), .page2Out_3__12 (\$dummy [134]), .page2Out_3__11 (
                    \$dummy [135]), .page2Out_3__10 (\$dummy [136]), .page2Out_3__9 (
                    \$dummy [137]), .page2Out_3__8 (\$dummy [138]), .page2Out_3__7 (
                    \$dummy [139]), .page2Out_3__6 (\$dummy [140]), .page2Out_3__5 (
                    \$dummy [141]), .page2Out_3__4 (\$dummy [142]), .page2Out_3__3 (
                    \$dummy [143]), .page2Out_3__2 (\$dummy [144]), .page2Out_3__1 (
                    \$dummy [145]), .page2Out_3__0 (\$dummy [146]), .page2Out_4__15 (
                    \$dummy [147]), .page2Out_4__14 (\$dummy [148]), .page2Out_4__13 (
                    \$dummy [149]), .page2Out_4__12 (\$dummy [150]), .page2Out_4__11 (
                    \$dummy [151]), .page2Out_4__10 (\$dummy [152]), .page2Out_4__9 (
                    \$dummy [153]), .page2Out_4__8 (\$dummy [154]), .page2Out_4__7 (
                    \$dummy [155]), .page2Out_4__6 (\$dummy [156]), .page2Out_4__5 (
                    \$dummy [157]), .page2Out_4__4 (\$dummy [158]), .page2Out_4__3 (
                    \$dummy [159]), .page2Out_4__2 (\$dummy [160]), .page2Out_4__1 (
                    \$dummy [161]), .page2Out_4__0 (\$dummy [162]), .pagesOutsPrimary_0__15 (
                    pagesOuts_0__15), .pagesOutsPrimary_0__14 (pagesOuts_0__14)
                    , .pagesOutsPrimary_0__13 (pagesOuts_0__13), .pagesOutsPrimary_0__12 (
                    pagesOuts_0__12), .pagesOutsPrimary_0__11 (pagesOuts_0__11)
                    , .pagesOutsPrimary_0__10 (pagesOuts_0__10), .pagesOutsPrimary_0__9 (
                    pagesOuts_0__9), .pagesOutsPrimary_0__8 (pagesOuts_0__8), .pagesOutsPrimary_0__7 (
                    pagesOuts_0__7), .pagesOutsPrimary_0__6 (pagesOuts_0__6), .pagesOutsPrimary_0__5 (
                    pagesOuts_0__5), .pagesOutsPrimary_0__4 (pagesOuts_0__4), .pagesOutsPrimary_0__3 (
                    pagesOuts_0__3), .pagesOutsPrimary_0__2 (pagesOuts_0__2), .pagesOutsPrimary_0__1 (
                    pagesOuts_0__1), .pagesOutsPrimary_0__0 (pagesOuts_0__0), .pagesOutsPrimary_1__15 (
                    pagesOuts_1__15), .pagesOutsPrimary_1__14 (pagesOuts_1__14)
                    , .pagesOutsPrimary_1__13 (pagesOuts_1__13), .pagesOutsPrimary_1__12 (
                    pagesOuts_1__12), .pagesOutsPrimary_1__11 (pagesOuts_1__11)
                    , .pagesOutsPrimary_1__10 (pagesOuts_1__10), .pagesOutsPrimary_1__9 (
                    pagesOuts_1__9), .pagesOutsPrimary_1__8 (pagesOuts_1__8), .pagesOutsPrimary_1__7 (
                    pagesOuts_1__7), .pagesOutsPrimary_1__6 (pagesOuts_1__6), .pagesOutsPrimary_1__5 (
                    pagesOuts_1__5), .pagesOutsPrimary_1__4 (pagesOuts_1__4), .pagesOutsPrimary_1__3 (
                    pagesOuts_1__3), .pagesOutsPrimary_1__2 (pagesOuts_1__2), .pagesOutsPrimary_1__1 (
                    pagesOuts_1__1), .pagesOutsPrimary_1__0 (pagesOuts_1__0), .pagesOutsPrimary_2__15 (
                    pagesOuts_2__15), .pagesOutsPrimary_2__14 (pagesOuts_2__14)
                    , .pagesOutsPrimary_2__13 (pagesOuts_2__13), .pagesOutsPrimary_2__12 (
                    pagesOuts_2__12), .pagesOutsPrimary_2__11 (pagesOuts_2__11)
                    , .pagesOutsPrimary_2__10 (pagesOuts_2__10), .pagesOutsPrimary_2__9 (
                    pagesOuts_2__9), .pagesOutsPrimary_2__8 (pagesOuts_2__8), .pagesOutsPrimary_2__7 (
                    pagesOuts_2__7), .pagesOutsPrimary_2__6 (pagesOuts_2__6), .pagesOutsPrimary_2__5 (
                    pagesOuts_2__5), .pagesOutsPrimary_2__4 (pagesOuts_2__4), .pagesOutsPrimary_2__3 (
                    pagesOuts_2__3), .pagesOutsPrimary_2__2 (pagesOuts_2__2), .pagesOutsPrimary_2__1 (
                    pagesOuts_2__1), .pagesOutsPrimary_2__0 (pagesOuts_2__0), .pagesOutsSecondary_0__15 (
                    pagesOuts_15__15), .pagesOutsSecondary_0__14 (
                    pagesOuts_15__14), .pagesOutsSecondary_0__13 (
                    pagesOuts_15__13), .pagesOutsSecondary_0__12 (
                    pagesOuts_15__12), .pagesOutsSecondary_0__11 (
                    pagesOuts_15__11), .pagesOutsSecondary_0__10 (
                    pagesOuts_15__10), .pagesOutsSecondary_0__9 (pagesOuts_15__9
                    ), .pagesOutsSecondary_0__8 (pagesOuts_15__8), .pagesOutsSecondary_0__7 (
                    pagesOuts_15__7), .pagesOutsSecondary_0__6 (pagesOuts_15__6)
                    , .pagesOutsSecondary_0__5 (pagesOuts_15__5), .pagesOutsSecondary_0__4 (
                    pagesOuts_15__4), .pagesOutsSecondary_0__3 (pagesOuts_15__3)
                    , .pagesOutsSecondary_0__2 (pagesOuts_15__2), .pagesOutsSecondary_0__1 (
                    pagesOuts_15__1), .pagesOutsSecondary_0__0 (pagesOuts_15__0)
                    , .pagesOutsSecondary_1__15 (pagesOuts_16__15), .pagesOutsSecondary_1__14 (
                    pagesOuts_16__14), .pagesOutsSecondary_1__13 (
                    pagesOuts_16__13), .pagesOutsSecondary_1__12 (
                    pagesOuts_16__12), .pagesOutsSecondary_1__11 (
                    pagesOuts_16__11), .pagesOutsSecondary_1__10 (
                    pagesOuts_16__10), .pagesOutsSecondary_1__9 (pagesOuts_16__9
                    ), .pagesOutsSecondary_1__8 (pagesOuts_16__8), .pagesOutsSecondary_1__7 (
                    pagesOuts_16__7), .pagesOutsSecondary_1__6 (pagesOuts_16__6)
                    , .pagesOutsSecondary_1__5 (pagesOuts_16__5), .pagesOutsSecondary_1__4 (
                    pagesOuts_16__4), .pagesOutsSecondary_1__3 (pagesOuts_16__3)
                    , .pagesOutsSecondary_1__2 (pagesOuts_16__2), .pagesOutsSecondary_1__1 (
                    pagesOuts_16__1), .pagesOutsSecondary_1__0 (pagesOuts_16__0)
                    , .filtersOutsPrimary_0__7 (filtersOuts_0__7), .filtersOutsPrimary_0__6 (
                    filtersOuts_0__6), .filtersOutsPrimary_0__5 (
                    filtersOuts_0__5), .filtersOutsPrimary_0__4 (
                    filtersOuts_0__4), .filtersOutsPrimary_0__3 (
                    filtersOuts_0__3), .filtersOutsPrimary_0__2 (
                    filtersOuts_0__2), .filtersOutsPrimary_0__1 (
                    filtersOuts_0__1), .filtersOutsPrimary_0__0 (
                    filtersOuts_0__0), .filtersOutsPrimary_1__7 (
                    filtersOuts_1__7), .filtersOutsPrimary_1__6 (
                    filtersOuts_1__6), .filtersOutsPrimary_1__5 (
                    filtersOuts_1__5), .filtersOutsPrimary_1__4 (
                    filtersOuts_1__4), .filtersOutsPrimary_1__3 (
                    filtersOuts_1__3), .filtersOutsPrimary_1__2 (
                    filtersOuts_1__2), .filtersOutsPrimary_1__1 (
                    filtersOuts_1__1), .filtersOutsPrimary_1__0 (
                    filtersOuts_1__0), .filtersOutsPrimary_2__7 (
                    filtersOuts_2__7), .filtersOutsPrimary_2__6 (
                    filtersOuts_2__6), .filtersOutsPrimary_2__5 (
                    filtersOuts_2__5), .filtersOutsPrimary_2__4 (
                    filtersOuts_2__4), .filtersOutsPrimary_2__3 (
                    filtersOuts_2__3), .filtersOutsPrimary_2__2 (
                    filtersOuts_2__2), .filtersOutsPrimary_2__1 (
                    filtersOuts_2__1), .filtersOutsPrimary_2__0 (
                    filtersOuts_2__0), .filtersOutsSecondary_0__7 (
                    filtersOuts_15__7), .filtersOutsSecondary_0__6 (
                    filtersOuts_15__6), .filtersOutsSecondary_0__5 (
                    filtersOuts_15__5), .filtersOutsSecondary_0__4 (
                    filtersOuts_15__4), .filtersOutsSecondary_0__3 (
                    filtersOuts_15__3), .filtersOutsSecondary_0__2 (
                    filtersOuts_15__2), .filtersOutsSecondary_0__1 (
                    filtersOuts_15__1), .filtersOutsSecondary_0__0 (
                    filtersOuts_15__0), .filtersOutsSecondary_1__7 (
                    filtersOuts_16__7), .filtersOutsSecondary_1__6 (
                    filtersOuts_16__6), .filtersOutsSecondary_1__5 (
                    filtersOuts_16__5), .filtersOutsSecondary_1__4 (
                    filtersOuts_16__4), .filtersOutsSecondary_1__3 (
                    filtersOuts_16__3), .filtersOutsSecondary_1__2 (
                    filtersOuts_16__2), .filtersOutsSecondary_1__1 (
                    filtersOuts_16__1), .filtersOutsSecondary_1__0 (
                    filtersOuts_16__0)) ;
    RegRow_8_16_5_3 loop1_1_regRowMap (.filterBus ({filterBus[39],filterBus[38],
                    filterBus[37],filterBus[36],filterBus[35],filterBus[34],
                    filterBus[33],filterBus[32],filterBus[31],filterBus[30],
                    filterBus[29],filterBus[28],filterBus[27],filterBus[26],
                    filterBus[25],filterBus[24],filterBus[23],filterBus[22],
                    filterBus[21],filterBus[20],filterBus[19],filterBus[18],
                    filterBus[17],filterBus[16],filterBus[15],filterBus[14],
                    filterBus[13],filterBus[12],filterBus[11],filterBus[10],
                    filterBus[9],filterBus[8],filterBus[7],filterBus[6],
                    filterBus[5],filterBus[4],filterBus[3],filterBus[2],
                    filterBus[1],filterBus[0]}), .windowBus ({nx2800,nx2804,
                    nx2808,nx2812,nx2816,nx2820,nx2824,nx2828,nx2832,nx2836,
                    nx2840,nx2844,nx2848,nx2852,nx2856,nx2860,nx2864,nx2868,
                    nx2872,nx2876,nx2880,nx2884,nx2888,nx2892,nx2896,nx2900,
                    nx2904,nx2908,nx2912,nx2916,nx2920,nx2924,nx2928,nx2932,
                    nx2936,nx2940,nx2944,nx2948,nx2952,nx2956,nx2960,nx2964,
                    nx2968,nx2972,nx2976,nx2980,nx2984,nx2988,nx2992,nx2996,
                    nx3000,nx3004,nx3008,nx3012,nx3016,nx3020,nx3024,nx3028,
                    nx3032,nx3036,nx3040,nx3044,nx3048,nx3052,nx3056,nx3060,
                    nx3064,nx3068,nx3072,nx3076,nx3080,nx3084,nx3088,nx3092,
                    nx3096,nx3100,nx3104,nx3108,nx3112,nx3116}), .page1NextRow_0__15 (
                    page1Out_10__15), .page1NextRow_0__14 (page1Out_10__14), .page1NextRow_0__13 (
                    page1Out_10__13), .page1NextRow_0__12 (page1Out_10__12), .page1NextRow_0__11 (
                    page1Out_10__11), .page1NextRow_0__10 (page1Out_10__10), .page1NextRow_0__9 (
                    page1Out_10__9), .page1NextRow_0__8 (page1Out_10__8), .page1NextRow_0__7 (
                    page1Out_10__7), .page1NextRow_0__6 (page1Out_10__6), .page1NextRow_0__5 (
                    page1Out_10__5), .page1NextRow_0__4 (page1Out_10__4), .page1NextRow_0__3 (
                    page1Out_10__3), .page1NextRow_0__2 (page1Out_10__2), .page1NextRow_0__1 (
                    page1Out_10__1), .page1NextRow_0__0 (page1Out_10__0), .page1NextRow_1__15 (
                    page1Out_11__15), .page1NextRow_1__14 (page1Out_11__14), .page1NextRow_1__13 (
                    page1Out_11__13), .page1NextRow_1__12 (page1Out_11__12), .page1NextRow_1__11 (
                    page1Out_11__11), .page1NextRow_1__10 (page1Out_11__10), .page1NextRow_1__9 (
                    page1Out_11__9), .page1NextRow_1__8 (page1Out_11__8), .page1NextRow_1__7 (
                    page1Out_11__7), .page1NextRow_1__6 (page1Out_11__6), .page1NextRow_1__5 (
                    page1Out_11__5), .page1NextRow_1__4 (page1Out_11__4), .page1NextRow_1__3 (
                    page1Out_11__3), .page1NextRow_1__2 (page1Out_11__2), .page1NextRow_1__1 (
                    page1Out_11__1), .page1NextRow_1__0 (page1Out_11__0), .page1NextRow_2__15 (
                    page1Out_12__15), .page1NextRow_2__14 (page1Out_12__14), .page1NextRow_2__13 (
                    page1Out_12__13), .page1NextRow_2__12 (page1Out_12__12), .page1NextRow_2__11 (
                    page1Out_12__11), .page1NextRow_2__10 (page1Out_12__10), .page1NextRow_2__9 (
                    page1Out_12__9), .page1NextRow_2__8 (page1Out_12__8), .page1NextRow_2__7 (
                    page1Out_12__7), .page1NextRow_2__6 (page1Out_12__6), .page1NextRow_2__5 (
                    page1Out_12__5), .page1NextRow_2__4 (page1Out_12__4), .page1NextRow_2__3 (
                    page1Out_12__3), .page1NextRow_2__2 (page1Out_12__2), .page1NextRow_2__1 (
                    page1Out_12__1), .page1NextRow_2__0 (page1Out_12__0), .page1NextRow_3__15 (
                    page1Out_13__15), .page1NextRow_3__14 (page1Out_13__14), .page1NextRow_3__13 (
                    page1Out_13__13), .page1NextRow_3__12 (page1Out_13__12), .page1NextRow_3__11 (
                    page1Out_13__11), .page1NextRow_3__10 (page1Out_13__10), .page1NextRow_3__9 (
                    page1Out_13__9), .page1NextRow_3__8 (page1Out_13__8), .page1NextRow_3__7 (
                    page1Out_13__7), .page1NextRow_3__6 (page1Out_13__6), .page1NextRow_3__5 (
                    page1Out_13__5), .page1NextRow_3__4 (page1Out_13__4), .page1NextRow_3__3 (
                    page1Out_13__3), .page1NextRow_3__2 (page1Out_13__2), .page1NextRow_3__1 (
                    page1Out_13__1), .page1NextRow_3__0 (page1Out_13__0), .page1NextRow_4__15 (
                    page1Out_14__15), .page1NextRow_4__14 (page1Out_14__14), .page1NextRow_4__13 (
                    page1Out_14__13), .page1NextRow_4__12 (page1Out_14__12), .page1NextRow_4__11 (
                    page1Out_14__11), .page1NextRow_4__10 (page1Out_14__10), .page1NextRow_4__9 (
                    page1Out_14__9), .page1NextRow_4__8 (page1Out_14__8), .page1NextRow_4__7 (
                    page1Out_14__7), .page1NextRow_4__6 (page1Out_14__6), .page1NextRow_4__5 (
                    page1Out_14__5), .page1NextRow_4__4 (page1Out_14__4), .page1NextRow_4__3 (
                    page1Out_14__3), .page1NextRow_4__2 (page1Out_14__2), .page1NextRow_4__1 (
                    page1Out_14__1), .page1NextRow_4__0 (page1Out_14__0), .page2NextRow_0__15 (
                    page2Out_10__15), .page2NextRow_0__14 (page2Out_10__14), .page2NextRow_0__13 (
                    page2Out_10__13), .page2NextRow_0__12 (page2Out_10__12), .page2NextRow_0__11 (
                    page2Out_10__11), .page2NextRow_0__10 (page2Out_10__10), .page2NextRow_0__9 (
                    page2Out_10__9), .page2NextRow_0__8 (page2Out_10__8), .page2NextRow_0__7 (
                    page2Out_10__7), .page2NextRow_0__6 (page2Out_10__6), .page2NextRow_0__5 (
                    page2Out_10__5), .page2NextRow_0__4 (page2Out_10__4), .page2NextRow_0__3 (
                    page2Out_10__3), .page2NextRow_0__2 (page2Out_10__2), .page2NextRow_0__1 (
                    page2Out_10__1), .page2NextRow_0__0 (page2Out_10__0), .page2NextRow_1__15 (
                    page2Out_11__15), .page2NextRow_1__14 (page2Out_11__14), .page2NextRow_1__13 (
                    page2Out_11__13), .page2NextRow_1__12 (page2Out_11__12), .page2NextRow_1__11 (
                    page2Out_11__11), .page2NextRow_1__10 (page2Out_11__10), .page2NextRow_1__9 (
                    page2Out_11__9), .page2NextRow_1__8 (page2Out_11__8), .page2NextRow_1__7 (
                    page2Out_11__7), .page2NextRow_1__6 (page2Out_11__6), .page2NextRow_1__5 (
                    page2Out_11__5), .page2NextRow_1__4 (page2Out_11__4), .page2NextRow_1__3 (
                    page2Out_11__3), .page2NextRow_1__2 (page2Out_11__2), .page2NextRow_1__1 (
                    page2Out_11__1), .page2NextRow_1__0 (page2Out_11__0), .page2NextRow_2__15 (
                    page2Out_12__15), .page2NextRow_2__14 (page2Out_12__14), .page2NextRow_2__13 (
                    page2Out_12__13), .page2NextRow_2__12 (page2Out_12__12), .page2NextRow_2__11 (
                    page2Out_12__11), .page2NextRow_2__10 (page2Out_12__10), .page2NextRow_2__9 (
                    page2Out_12__9), .page2NextRow_2__8 (page2Out_12__8), .page2NextRow_2__7 (
                    page2Out_12__7), .page2NextRow_2__6 (page2Out_12__6), .page2NextRow_2__5 (
                    page2Out_12__5), .page2NextRow_2__4 (page2Out_12__4), .page2NextRow_2__3 (
                    page2Out_12__3), .page2NextRow_2__2 (page2Out_12__2), .page2NextRow_2__1 (
                    page2Out_12__1), .page2NextRow_2__0 (page2Out_12__0), .page2NextRow_3__15 (
                    page2Out_13__15), .page2NextRow_3__14 (page2Out_13__14), .page2NextRow_3__13 (
                    page2Out_13__13), .page2NextRow_3__12 (page2Out_13__12), .page2NextRow_3__11 (
                    page2Out_13__11), .page2NextRow_3__10 (page2Out_13__10), .page2NextRow_3__9 (
                    page2Out_13__9), .page2NextRow_3__8 (page2Out_13__8), .page2NextRow_3__7 (
                    page2Out_13__7), .page2NextRow_3__6 (page2Out_13__6), .page2NextRow_3__5 (
                    page2Out_13__5), .page2NextRow_3__4 (page2Out_13__4), .page2NextRow_3__3 (
                    page2Out_13__3), .page2NextRow_3__2 (page2Out_13__2), .page2NextRow_3__1 (
                    page2Out_13__1), .page2NextRow_3__0 (page2Out_13__0), .page2NextRow_4__15 (
                    page2Out_14__15), .page2NextRow_4__14 (page2Out_14__14), .page2NextRow_4__13 (
                    page2Out_14__13), .page2NextRow_4__12 (page2Out_14__12), .page2NextRow_4__11 (
                    page2Out_14__11), .page2NextRow_4__10 (page2Out_14__10), .page2NextRow_4__9 (
                    page2Out_14__9), .page2NextRow_4__8 (page2Out_14__8), .page2NextRow_4__7 (
                    page2Out_14__7), .page2NextRow_4__6 (page2Out_14__6), .page2NextRow_4__5 (
                    page2Out_14__5), .page2NextRow_4__4 (page2Out_14__4), .page2NextRow_4__3 (
                    page2Out_14__3), .page2NextRow_4__2 (page2Out_14__2), .page2NextRow_4__1 (
                    page2Out_14__1), .page2NextRow_4__0 (page2Out_14__0), .clk (
                    clk), .rst (rst), .enablePage1Read (page1Enables_1), .enablePage2Read (
                    page2Enables_1), .enableFilterRead (filterEnables_1), .shift2To1 (
                    nx3120), .shift1To2 (nx3124), .pageTurn (nx2792), .page1Out_0__15 (
                    page1Out_5__15), .page1Out_0__14 (page1Out_5__14), .page1Out_0__13 (
                    page1Out_5__13), .page1Out_0__12 (page1Out_5__12), .page1Out_0__11 (
                    page1Out_5__11), .page1Out_0__10 (page1Out_5__10), .page1Out_0__9 (
                    page1Out_5__9), .page1Out_0__8 (page1Out_5__8), .page1Out_0__7 (
                    page1Out_5__7), .page1Out_0__6 (page1Out_5__6), .page1Out_0__5 (
                    page1Out_5__5), .page1Out_0__4 (page1Out_5__4), .page1Out_0__3 (
                    page1Out_5__3), .page1Out_0__2 (page1Out_5__2), .page1Out_0__1 (
                    page1Out_5__1), .page1Out_0__0 (page1Out_5__0), .page1Out_1__15 (
                    page1Out_6__15), .page1Out_1__14 (page1Out_6__14), .page1Out_1__13 (
                    page1Out_6__13), .page1Out_1__12 (page1Out_6__12), .page1Out_1__11 (
                    page1Out_6__11), .page1Out_1__10 (page1Out_6__10), .page1Out_1__9 (
                    page1Out_6__9), .page1Out_1__8 (page1Out_6__8), .page1Out_1__7 (
                    page1Out_6__7), .page1Out_1__6 (page1Out_6__6), .page1Out_1__5 (
                    page1Out_6__5), .page1Out_1__4 (page1Out_6__4), .page1Out_1__3 (
                    page1Out_6__3), .page1Out_1__2 (page1Out_6__2), .page1Out_1__1 (
                    page1Out_6__1), .page1Out_1__0 (page1Out_6__0), .page1Out_2__15 (
                    page1Out_7__15), .page1Out_2__14 (page1Out_7__14), .page1Out_2__13 (
                    page1Out_7__13), .page1Out_2__12 (page1Out_7__12), .page1Out_2__11 (
                    page1Out_7__11), .page1Out_2__10 (page1Out_7__10), .page1Out_2__9 (
                    page1Out_7__9), .page1Out_2__8 (page1Out_7__8), .page1Out_2__7 (
                    page1Out_7__7), .page1Out_2__6 (page1Out_7__6), .page1Out_2__5 (
                    page1Out_7__5), .page1Out_2__4 (page1Out_7__4), .page1Out_2__3 (
                    page1Out_7__3), .page1Out_2__2 (page1Out_7__2), .page1Out_2__1 (
                    page1Out_7__1), .page1Out_2__0 (page1Out_7__0), .page1Out_3__15 (
                    page1Out_8__15), .page1Out_3__14 (page1Out_8__14), .page1Out_3__13 (
                    page1Out_8__13), .page1Out_3__12 (page1Out_8__12), .page1Out_3__11 (
                    page1Out_8__11), .page1Out_3__10 (page1Out_8__10), .page1Out_3__9 (
                    page1Out_8__9), .page1Out_3__8 (page1Out_8__8), .page1Out_3__7 (
                    page1Out_8__7), .page1Out_3__6 (page1Out_8__6), .page1Out_3__5 (
                    page1Out_8__5), .page1Out_3__4 (page1Out_8__4), .page1Out_3__3 (
                    page1Out_8__3), .page1Out_3__2 (page1Out_8__2), .page1Out_3__1 (
                    page1Out_8__1), .page1Out_3__0 (page1Out_8__0), .page1Out_4__15 (
                    page1Out_9__15), .page1Out_4__14 (page1Out_9__14), .page1Out_4__13 (
                    page1Out_9__13), .page1Out_4__12 (page1Out_9__12), .page1Out_4__11 (
                    page1Out_9__11), .page1Out_4__10 (page1Out_9__10), .page1Out_4__9 (
                    page1Out_9__9), .page1Out_4__8 (page1Out_9__8), .page1Out_4__7 (
                    page1Out_9__7), .page1Out_4__6 (page1Out_9__6), .page1Out_4__5 (
                    page1Out_9__5), .page1Out_4__4 (page1Out_9__4), .page1Out_4__3 (
                    page1Out_9__3), .page1Out_4__2 (page1Out_9__2), .page1Out_4__1 (
                    page1Out_9__1), .page1Out_4__0 (page1Out_9__0), .page2Out_0__15 (
                    page2Out_5__15), .page2Out_0__14 (page2Out_5__14), .page2Out_0__13 (
                    page2Out_5__13), .page2Out_0__12 (page2Out_5__12), .page2Out_0__11 (
                    page2Out_5__11), .page2Out_0__10 (page2Out_5__10), .page2Out_0__9 (
                    page2Out_5__9), .page2Out_0__8 (page2Out_5__8), .page2Out_0__7 (
                    page2Out_5__7), .page2Out_0__6 (page2Out_5__6), .page2Out_0__5 (
                    page2Out_5__5), .page2Out_0__4 (page2Out_5__4), .page2Out_0__3 (
                    page2Out_5__3), .page2Out_0__2 (page2Out_5__2), .page2Out_0__1 (
                    page2Out_5__1), .page2Out_0__0 (page2Out_5__0), .page2Out_1__15 (
                    page2Out_6__15), .page2Out_1__14 (page2Out_6__14), .page2Out_1__13 (
                    page2Out_6__13), .page2Out_1__12 (page2Out_6__12), .page2Out_1__11 (
                    page2Out_6__11), .page2Out_1__10 (page2Out_6__10), .page2Out_1__9 (
                    page2Out_6__9), .page2Out_1__8 (page2Out_6__8), .page2Out_1__7 (
                    page2Out_6__7), .page2Out_1__6 (page2Out_6__6), .page2Out_1__5 (
                    page2Out_6__5), .page2Out_1__4 (page2Out_6__4), .page2Out_1__3 (
                    page2Out_6__3), .page2Out_1__2 (page2Out_6__2), .page2Out_1__1 (
                    page2Out_6__1), .page2Out_1__0 (page2Out_6__0), .page2Out_2__15 (
                    page2Out_7__15), .page2Out_2__14 (page2Out_7__14), .page2Out_2__13 (
                    page2Out_7__13), .page2Out_2__12 (page2Out_7__12), .page2Out_2__11 (
                    page2Out_7__11), .page2Out_2__10 (page2Out_7__10), .page2Out_2__9 (
                    page2Out_7__9), .page2Out_2__8 (page2Out_7__8), .page2Out_2__7 (
                    page2Out_7__7), .page2Out_2__6 (page2Out_7__6), .page2Out_2__5 (
                    page2Out_7__5), .page2Out_2__4 (page2Out_7__4), .page2Out_2__3 (
                    page2Out_7__3), .page2Out_2__2 (page2Out_7__2), .page2Out_2__1 (
                    page2Out_7__1), .page2Out_2__0 (page2Out_7__0), .page2Out_3__15 (
                    page2Out_8__15), .page2Out_3__14 (page2Out_8__14), .page2Out_3__13 (
                    page2Out_8__13), .page2Out_3__12 (page2Out_8__12), .page2Out_3__11 (
                    page2Out_8__11), .page2Out_3__10 (page2Out_8__10), .page2Out_3__9 (
                    page2Out_8__9), .page2Out_3__8 (page2Out_8__8), .page2Out_3__7 (
                    page2Out_8__7), .page2Out_3__6 (page2Out_8__6), .page2Out_3__5 (
                    page2Out_8__5), .page2Out_3__4 (page2Out_8__4), .page2Out_3__3 (
                    page2Out_8__3), .page2Out_3__2 (page2Out_8__2), .page2Out_3__1 (
                    page2Out_8__1), .page2Out_3__0 (page2Out_8__0), .page2Out_4__15 (
                    page2Out_9__15), .page2Out_4__14 (page2Out_9__14), .page2Out_4__13 (
                    page2Out_9__13), .page2Out_4__12 (page2Out_9__12), .page2Out_4__11 (
                    page2Out_9__11), .page2Out_4__10 (page2Out_9__10), .page2Out_4__9 (
                    page2Out_9__9), .page2Out_4__8 (page2Out_9__8), .page2Out_4__7 (
                    page2Out_9__7), .page2Out_4__6 (page2Out_9__6), .page2Out_4__5 (
                    page2Out_9__5), .page2Out_4__4 (page2Out_9__4), .page2Out_4__3 (
                    page2Out_9__3), .page2Out_4__2 (page2Out_9__2), .page2Out_4__1 (
                    page2Out_9__1), .page2Out_4__0 (page2Out_9__0), .pagesOutsPrimary_0__15 (
                    pagesOuts_3__15), .pagesOutsPrimary_0__14 (pagesOuts_3__14)
                    , .pagesOutsPrimary_0__13 (pagesOuts_3__13), .pagesOutsPrimary_0__12 (
                    pagesOuts_3__12), .pagesOutsPrimary_0__11 (pagesOuts_3__11)
                    , .pagesOutsPrimary_0__10 (pagesOuts_3__10), .pagesOutsPrimary_0__9 (
                    pagesOuts_3__9), .pagesOutsPrimary_0__8 (pagesOuts_3__8), .pagesOutsPrimary_0__7 (
                    pagesOuts_3__7), .pagesOutsPrimary_0__6 (pagesOuts_3__6), .pagesOutsPrimary_0__5 (
                    pagesOuts_3__5), .pagesOutsPrimary_0__4 (pagesOuts_3__4), .pagesOutsPrimary_0__3 (
                    pagesOuts_3__3), .pagesOutsPrimary_0__2 (pagesOuts_3__2), .pagesOutsPrimary_0__1 (
                    pagesOuts_3__1), .pagesOutsPrimary_0__0 (pagesOuts_3__0), .pagesOutsPrimary_1__15 (
                    pagesOuts_4__15), .pagesOutsPrimary_1__14 (pagesOuts_4__14)
                    , .pagesOutsPrimary_1__13 (pagesOuts_4__13), .pagesOutsPrimary_1__12 (
                    pagesOuts_4__12), .pagesOutsPrimary_1__11 (pagesOuts_4__11)
                    , .pagesOutsPrimary_1__10 (pagesOuts_4__10), .pagesOutsPrimary_1__9 (
                    pagesOuts_4__9), .pagesOutsPrimary_1__8 (pagesOuts_4__8), .pagesOutsPrimary_1__7 (
                    pagesOuts_4__7), .pagesOutsPrimary_1__6 (pagesOuts_4__6), .pagesOutsPrimary_1__5 (
                    pagesOuts_4__5), .pagesOutsPrimary_1__4 (pagesOuts_4__4), .pagesOutsPrimary_1__3 (
                    pagesOuts_4__3), .pagesOutsPrimary_1__2 (pagesOuts_4__2), .pagesOutsPrimary_1__1 (
                    pagesOuts_4__1), .pagesOutsPrimary_1__0 (pagesOuts_4__0), .pagesOutsPrimary_2__15 (
                    pagesOuts_5__15), .pagesOutsPrimary_2__14 (pagesOuts_5__14)
                    , .pagesOutsPrimary_2__13 (pagesOuts_5__13), .pagesOutsPrimary_2__12 (
                    pagesOuts_5__12), .pagesOutsPrimary_2__11 (pagesOuts_5__11)
                    , .pagesOutsPrimary_2__10 (pagesOuts_5__10), .pagesOutsPrimary_2__9 (
                    pagesOuts_5__9), .pagesOutsPrimary_2__8 (pagesOuts_5__8), .pagesOutsPrimary_2__7 (
                    pagesOuts_5__7), .pagesOutsPrimary_2__6 (pagesOuts_5__6), .pagesOutsPrimary_2__5 (
                    pagesOuts_5__5), .pagesOutsPrimary_2__4 (pagesOuts_5__4), .pagesOutsPrimary_2__3 (
                    pagesOuts_5__3), .pagesOutsPrimary_2__2 (pagesOuts_5__2), .pagesOutsPrimary_2__1 (
                    pagesOuts_5__1), .pagesOutsPrimary_2__0 (pagesOuts_5__0), .pagesOutsSecondary_0__15 (
                    pagesOuts_17__15), .pagesOutsSecondary_0__14 (
                    pagesOuts_17__14), .pagesOutsSecondary_0__13 (
                    pagesOuts_17__13), .pagesOutsSecondary_0__12 (
                    pagesOuts_17__12), .pagesOutsSecondary_0__11 (
                    pagesOuts_17__11), .pagesOutsSecondary_0__10 (
                    pagesOuts_17__10), .pagesOutsSecondary_0__9 (pagesOuts_17__9
                    ), .pagesOutsSecondary_0__8 (pagesOuts_17__8), .pagesOutsSecondary_0__7 (
                    pagesOuts_17__7), .pagesOutsSecondary_0__6 (pagesOuts_17__6)
                    , .pagesOutsSecondary_0__5 (pagesOuts_17__5), .pagesOutsSecondary_0__4 (
                    pagesOuts_17__4), .pagesOutsSecondary_0__3 (pagesOuts_17__3)
                    , .pagesOutsSecondary_0__2 (pagesOuts_17__2), .pagesOutsSecondary_0__1 (
                    pagesOuts_17__1), .pagesOutsSecondary_0__0 (pagesOuts_17__0)
                    , .pagesOutsSecondary_1__15 (pagesOuts_18__15), .pagesOutsSecondary_1__14 (
                    pagesOuts_18__14), .pagesOutsSecondary_1__13 (
                    pagesOuts_18__13), .pagesOutsSecondary_1__12 (
                    pagesOuts_18__12), .pagesOutsSecondary_1__11 (
                    pagesOuts_18__11), .pagesOutsSecondary_1__10 (
                    pagesOuts_18__10), .pagesOutsSecondary_1__9 (pagesOuts_18__9
                    ), .pagesOutsSecondary_1__8 (pagesOuts_18__8), .pagesOutsSecondary_1__7 (
                    pagesOuts_18__7), .pagesOutsSecondary_1__6 (pagesOuts_18__6)
                    , .pagesOutsSecondary_1__5 (pagesOuts_18__5), .pagesOutsSecondary_1__4 (
                    pagesOuts_18__4), .pagesOutsSecondary_1__3 (pagesOuts_18__3)
                    , .pagesOutsSecondary_1__2 (pagesOuts_18__2), .pagesOutsSecondary_1__1 (
                    pagesOuts_18__1), .pagesOutsSecondary_1__0 (pagesOuts_18__0)
                    , .filtersOutsPrimary_0__7 (filtersOuts_3__7), .filtersOutsPrimary_0__6 (
                    filtersOuts_3__6), .filtersOutsPrimary_0__5 (
                    filtersOuts_3__5), .filtersOutsPrimary_0__4 (
                    filtersOuts_3__4), .filtersOutsPrimary_0__3 (
                    filtersOuts_3__3), .filtersOutsPrimary_0__2 (
                    filtersOuts_3__2), .filtersOutsPrimary_0__1 (
                    filtersOuts_3__1), .filtersOutsPrimary_0__0 (
                    filtersOuts_3__0), .filtersOutsPrimary_1__7 (
                    filtersOuts_4__7), .filtersOutsPrimary_1__6 (
                    filtersOuts_4__6), .filtersOutsPrimary_1__5 (
                    filtersOuts_4__5), .filtersOutsPrimary_1__4 (
                    filtersOuts_4__4), .filtersOutsPrimary_1__3 (
                    filtersOuts_4__3), .filtersOutsPrimary_1__2 (
                    filtersOuts_4__2), .filtersOutsPrimary_1__1 (
                    filtersOuts_4__1), .filtersOutsPrimary_1__0 (
                    filtersOuts_4__0), .filtersOutsPrimary_2__7 (
                    filtersOuts_5__7), .filtersOutsPrimary_2__6 (
                    filtersOuts_5__6), .filtersOutsPrimary_2__5 (
                    filtersOuts_5__5), .filtersOutsPrimary_2__4 (
                    filtersOuts_5__4), .filtersOutsPrimary_2__3 (
                    filtersOuts_5__3), .filtersOutsPrimary_2__2 (
                    filtersOuts_5__2), .filtersOutsPrimary_2__1 (
                    filtersOuts_5__1), .filtersOutsPrimary_2__0 (
                    filtersOuts_5__0), .filtersOutsSecondary_0__7 (
                    filtersOuts_17__7), .filtersOutsSecondary_0__6 (
                    filtersOuts_17__6), .filtersOutsSecondary_0__5 (
                    filtersOuts_17__5), .filtersOutsSecondary_0__4 (
                    filtersOuts_17__4), .filtersOutsSecondary_0__3 (
                    filtersOuts_17__3), .filtersOutsSecondary_0__2 (
                    filtersOuts_17__2), .filtersOutsSecondary_0__1 (
                    filtersOuts_17__1), .filtersOutsSecondary_0__0 (
                    filtersOuts_17__0), .filtersOutsSecondary_1__7 (
                    filtersOuts_18__7), .filtersOutsSecondary_1__6 (
                    filtersOuts_18__6), .filtersOutsSecondary_1__5 (
                    filtersOuts_18__5), .filtersOutsSecondary_1__4 (
                    filtersOuts_18__4), .filtersOutsSecondary_1__3 (
                    filtersOuts_18__3), .filtersOutsSecondary_1__2 (
                    filtersOuts_18__2), .filtersOutsSecondary_1__1 (
                    filtersOuts_18__1), .filtersOutsSecondary_1__0 (
                    filtersOuts_18__0)) ;
    RegRow_8_16_5_3 loop1_2_regRowMap (.filterBus ({filterBus[39],filterBus[38],
                    filterBus[37],filterBus[36],filterBus[35],filterBus[34],
                    filterBus[33],filterBus[32],filterBus[31],filterBus[30],
                    filterBus[29],filterBus[28],filterBus[27],filterBus[26],
                    filterBus[25],filterBus[24],filterBus[23],filterBus[22],
                    filterBus[21],filterBus[20],filterBus[19],filterBus[18],
                    filterBus[17],filterBus[16],filterBus[15],filterBus[14],
                    filterBus[13],filterBus[12],filterBus[11],filterBus[10],
                    filterBus[9],filterBus[8],filterBus[7],filterBus[6],
                    filterBus[5],filterBus[4],filterBus[3],filterBus[2],
                    filterBus[1],filterBus[0]}), .windowBus ({nx2800,nx2804,
                    nx2808,nx2812,nx2816,nx2820,nx2824,nx2828,nx2832,nx2836,
                    nx2840,nx2844,nx2848,nx2852,nx2856,nx2860,nx2864,nx2868,
                    nx2872,nx2876,nx2880,nx2884,nx2888,nx2892,nx2896,nx2900,
                    nx2904,nx2908,nx2912,nx2916,nx2920,nx2924,nx2928,nx2932,
                    nx2936,nx2940,nx2944,nx2948,nx2952,nx2956,nx2960,nx2964,
                    nx2968,nx2972,nx2976,nx2980,nx2984,nx2988,nx2992,nx2996,
                    nx3000,nx3004,nx3008,nx3012,nx3016,nx3020,nx3024,nx3028,
                    nx3032,nx3036,nx3040,nx3044,nx3048,nx3052,nx3056,nx3060,
                    nx3064,nx3068,nx3072,nx3076,nx3080,nx3084,nx3088,nx3092,
                    nx3096,nx3100,nx3104,nx3108,nx3112,nx3116}), .page1NextRow_0__15 (
                    page1Out_15__15), .page1NextRow_0__14 (page1Out_15__14), .page1NextRow_0__13 (
                    page1Out_15__13), .page1NextRow_0__12 (page1Out_15__12), .page1NextRow_0__11 (
                    page1Out_15__11), .page1NextRow_0__10 (page1Out_15__10), .page1NextRow_0__9 (
                    page1Out_15__9), .page1NextRow_0__8 (page1Out_15__8), .page1NextRow_0__7 (
                    page1Out_15__7), .page1NextRow_0__6 (page1Out_15__6), .page1NextRow_0__5 (
                    page1Out_15__5), .page1NextRow_0__4 (page1Out_15__4), .page1NextRow_0__3 (
                    page1Out_15__3), .page1NextRow_0__2 (page1Out_15__2), .page1NextRow_0__1 (
                    page1Out_15__1), .page1NextRow_0__0 (page1Out_15__0), .page1NextRow_1__15 (
                    page1Out_16__15), .page1NextRow_1__14 (page1Out_16__14), .page1NextRow_1__13 (
                    page1Out_16__13), .page1NextRow_1__12 (page1Out_16__12), .page1NextRow_1__11 (
                    page1Out_16__11), .page1NextRow_1__10 (page1Out_16__10), .page1NextRow_1__9 (
                    page1Out_16__9), .page1NextRow_1__8 (page1Out_16__8), .page1NextRow_1__7 (
                    page1Out_16__7), .page1NextRow_1__6 (page1Out_16__6), .page1NextRow_1__5 (
                    page1Out_16__5), .page1NextRow_1__4 (page1Out_16__4), .page1NextRow_1__3 (
                    page1Out_16__3), .page1NextRow_1__2 (page1Out_16__2), .page1NextRow_1__1 (
                    page1Out_16__1), .page1NextRow_1__0 (page1Out_16__0), .page1NextRow_2__15 (
                    page1Out_17__15), .page1NextRow_2__14 (page1Out_17__14), .page1NextRow_2__13 (
                    page1Out_17__13), .page1NextRow_2__12 (page1Out_17__12), .page1NextRow_2__11 (
                    page1Out_17__11), .page1NextRow_2__10 (page1Out_17__10), .page1NextRow_2__9 (
                    page1Out_17__9), .page1NextRow_2__8 (page1Out_17__8), .page1NextRow_2__7 (
                    page1Out_17__7), .page1NextRow_2__6 (page1Out_17__6), .page1NextRow_2__5 (
                    page1Out_17__5), .page1NextRow_2__4 (page1Out_17__4), .page1NextRow_2__3 (
                    page1Out_17__3), .page1NextRow_2__2 (page1Out_17__2), .page1NextRow_2__1 (
                    page1Out_17__1), .page1NextRow_2__0 (page1Out_17__0), .page1NextRow_3__15 (
                    page1Out_18__15), .page1NextRow_3__14 (page1Out_18__14), .page1NextRow_3__13 (
                    page1Out_18__13), .page1NextRow_3__12 (page1Out_18__12), .page1NextRow_3__11 (
                    page1Out_18__11), .page1NextRow_3__10 (page1Out_18__10), .page1NextRow_3__9 (
                    page1Out_18__9), .page1NextRow_3__8 (page1Out_18__8), .page1NextRow_3__7 (
                    page1Out_18__7), .page1NextRow_3__6 (page1Out_18__6), .page1NextRow_3__5 (
                    page1Out_18__5), .page1NextRow_3__4 (page1Out_18__4), .page1NextRow_3__3 (
                    page1Out_18__3), .page1NextRow_3__2 (page1Out_18__2), .page1NextRow_3__1 (
                    page1Out_18__1), .page1NextRow_3__0 (page1Out_18__0), .page1NextRow_4__15 (
                    page1Out_19__15), .page1NextRow_4__14 (page1Out_19__14), .page1NextRow_4__13 (
                    page1Out_19__13), .page1NextRow_4__12 (page1Out_19__12), .page1NextRow_4__11 (
                    page1Out_19__11), .page1NextRow_4__10 (page1Out_19__10), .page1NextRow_4__9 (
                    page1Out_19__9), .page1NextRow_4__8 (page1Out_19__8), .page1NextRow_4__7 (
                    page1Out_19__7), .page1NextRow_4__6 (page1Out_19__6), .page1NextRow_4__5 (
                    page1Out_19__5), .page1NextRow_4__4 (page1Out_19__4), .page1NextRow_4__3 (
                    page1Out_19__3), .page1NextRow_4__2 (page1Out_19__2), .page1NextRow_4__1 (
                    page1Out_19__1), .page1NextRow_4__0 (page1Out_19__0), .page2NextRow_0__15 (
                    page2Out_15__15), .page2NextRow_0__14 (page2Out_15__14), .page2NextRow_0__13 (
                    page2Out_15__13), .page2NextRow_0__12 (page2Out_15__12), .page2NextRow_0__11 (
                    page2Out_15__11), .page2NextRow_0__10 (page2Out_15__10), .page2NextRow_0__9 (
                    page2Out_15__9), .page2NextRow_0__8 (page2Out_15__8), .page2NextRow_0__7 (
                    page2Out_15__7), .page2NextRow_0__6 (page2Out_15__6), .page2NextRow_0__5 (
                    page2Out_15__5), .page2NextRow_0__4 (page2Out_15__4), .page2NextRow_0__3 (
                    page2Out_15__3), .page2NextRow_0__2 (page2Out_15__2), .page2NextRow_0__1 (
                    page2Out_15__1), .page2NextRow_0__0 (page2Out_15__0), .page2NextRow_1__15 (
                    page2Out_16__15), .page2NextRow_1__14 (page2Out_16__14), .page2NextRow_1__13 (
                    page2Out_16__13), .page2NextRow_1__12 (page2Out_16__12), .page2NextRow_1__11 (
                    page2Out_16__11), .page2NextRow_1__10 (page2Out_16__10), .page2NextRow_1__9 (
                    page2Out_16__9), .page2NextRow_1__8 (page2Out_16__8), .page2NextRow_1__7 (
                    page2Out_16__7), .page2NextRow_1__6 (page2Out_16__6), .page2NextRow_1__5 (
                    page2Out_16__5), .page2NextRow_1__4 (page2Out_16__4), .page2NextRow_1__3 (
                    page2Out_16__3), .page2NextRow_1__2 (page2Out_16__2), .page2NextRow_1__1 (
                    page2Out_16__1), .page2NextRow_1__0 (page2Out_16__0), .page2NextRow_2__15 (
                    page2Out_17__15), .page2NextRow_2__14 (page2Out_17__14), .page2NextRow_2__13 (
                    page2Out_17__13), .page2NextRow_2__12 (page2Out_17__12), .page2NextRow_2__11 (
                    page2Out_17__11), .page2NextRow_2__10 (page2Out_17__10), .page2NextRow_2__9 (
                    page2Out_17__9), .page2NextRow_2__8 (page2Out_17__8), .page2NextRow_2__7 (
                    page2Out_17__7), .page2NextRow_2__6 (page2Out_17__6), .page2NextRow_2__5 (
                    page2Out_17__5), .page2NextRow_2__4 (page2Out_17__4), .page2NextRow_2__3 (
                    page2Out_17__3), .page2NextRow_2__2 (page2Out_17__2), .page2NextRow_2__1 (
                    page2Out_17__1), .page2NextRow_2__0 (page2Out_17__0), .page2NextRow_3__15 (
                    page2Out_18__15), .page2NextRow_3__14 (page2Out_18__14), .page2NextRow_3__13 (
                    page2Out_18__13), .page2NextRow_3__12 (page2Out_18__12), .page2NextRow_3__11 (
                    page2Out_18__11), .page2NextRow_3__10 (page2Out_18__10), .page2NextRow_3__9 (
                    page2Out_18__9), .page2NextRow_3__8 (page2Out_18__8), .page2NextRow_3__7 (
                    page2Out_18__7), .page2NextRow_3__6 (page2Out_18__6), .page2NextRow_3__5 (
                    page2Out_18__5), .page2NextRow_3__4 (page2Out_18__4), .page2NextRow_3__3 (
                    page2Out_18__3), .page2NextRow_3__2 (page2Out_18__2), .page2NextRow_3__1 (
                    page2Out_18__1), .page2NextRow_3__0 (page2Out_18__0), .page2NextRow_4__15 (
                    page2Out_19__15), .page2NextRow_4__14 (page2Out_19__14), .page2NextRow_4__13 (
                    page2Out_19__13), .page2NextRow_4__12 (page2Out_19__12), .page2NextRow_4__11 (
                    page2Out_19__11), .page2NextRow_4__10 (page2Out_19__10), .page2NextRow_4__9 (
                    page2Out_19__9), .page2NextRow_4__8 (page2Out_19__8), .page2NextRow_4__7 (
                    page2Out_19__7), .page2NextRow_4__6 (page2Out_19__6), .page2NextRow_4__5 (
                    page2Out_19__5), .page2NextRow_4__4 (page2Out_19__4), .page2NextRow_4__3 (
                    page2Out_19__3), .page2NextRow_4__2 (page2Out_19__2), .page2NextRow_4__1 (
                    page2Out_19__1), .page2NextRow_4__0 (page2Out_19__0), .clk (
                    clk), .rst (rst), .enablePage1Read (page1Enables_2), .enablePage2Read (
                    page2Enables_2), .enableFilterRead (filterEnables_2), .shift2To1 (
                    nx3120), .shift1To2 (nx3124), .pageTurn (nx2794), .page1Out_0__15 (
                    page1Out_10__15), .page1Out_0__14 (page1Out_10__14), .page1Out_0__13 (
                    page1Out_10__13), .page1Out_0__12 (page1Out_10__12), .page1Out_0__11 (
                    page1Out_10__11), .page1Out_0__10 (page1Out_10__10), .page1Out_0__9 (
                    page1Out_10__9), .page1Out_0__8 (page1Out_10__8), .page1Out_0__7 (
                    page1Out_10__7), .page1Out_0__6 (page1Out_10__6), .page1Out_0__5 (
                    page1Out_10__5), .page1Out_0__4 (page1Out_10__4), .page1Out_0__3 (
                    page1Out_10__3), .page1Out_0__2 (page1Out_10__2), .page1Out_0__1 (
                    page1Out_10__1), .page1Out_0__0 (page1Out_10__0), .page1Out_1__15 (
                    page1Out_11__15), .page1Out_1__14 (page1Out_11__14), .page1Out_1__13 (
                    page1Out_11__13), .page1Out_1__12 (page1Out_11__12), .page1Out_1__11 (
                    page1Out_11__11), .page1Out_1__10 (page1Out_11__10), .page1Out_1__9 (
                    page1Out_11__9), .page1Out_1__8 (page1Out_11__8), .page1Out_1__7 (
                    page1Out_11__7), .page1Out_1__6 (page1Out_11__6), .page1Out_1__5 (
                    page1Out_11__5), .page1Out_1__4 (page1Out_11__4), .page1Out_1__3 (
                    page1Out_11__3), .page1Out_1__2 (page1Out_11__2), .page1Out_1__1 (
                    page1Out_11__1), .page1Out_1__0 (page1Out_11__0), .page1Out_2__15 (
                    page1Out_12__15), .page1Out_2__14 (page1Out_12__14), .page1Out_2__13 (
                    page1Out_12__13), .page1Out_2__12 (page1Out_12__12), .page1Out_2__11 (
                    page1Out_12__11), .page1Out_2__10 (page1Out_12__10), .page1Out_2__9 (
                    page1Out_12__9), .page1Out_2__8 (page1Out_12__8), .page1Out_2__7 (
                    page1Out_12__7), .page1Out_2__6 (page1Out_12__6), .page1Out_2__5 (
                    page1Out_12__5), .page1Out_2__4 (page1Out_12__4), .page1Out_2__3 (
                    page1Out_12__3), .page1Out_2__2 (page1Out_12__2), .page1Out_2__1 (
                    page1Out_12__1), .page1Out_2__0 (page1Out_12__0), .page1Out_3__15 (
                    page1Out_13__15), .page1Out_3__14 (page1Out_13__14), .page1Out_3__13 (
                    page1Out_13__13), .page1Out_3__12 (page1Out_13__12), .page1Out_3__11 (
                    page1Out_13__11), .page1Out_3__10 (page1Out_13__10), .page1Out_3__9 (
                    page1Out_13__9), .page1Out_3__8 (page1Out_13__8), .page1Out_3__7 (
                    page1Out_13__7), .page1Out_3__6 (page1Out_13__6), .page1Out_3__5 (
                    page1Out_13__5), .page1Out_3__4 (page1Out_13__4), .page1Out_3__3 (
                    page1Out_13__3), .page1Out_3__2 (page1Out_13__2), .page1Out_3__1 (
                    page1Out_13__1), .page1Out_3__0 (page1Out_13__0), .page1Out_4__15 (
                    page1Out_14__15), .page1Out_4__14 (page1Out_14__14), .page1Out_4__13 (
                    page1Out_14__13), .page1Out_4__12 (page1Out_14__12), .page1Out_4__11 (
                    page1Out_14__11), .page1Out_4__10 (page1Out_14__10), .page1Out_4__9 (
                    page1Out_14__9), .page1Out_4__8 (page1Out_14__8), .page1Out_4__7 (
                    page1Out_14__7), .page1Out_4__6 (page1Out_14__6), .page1Out_4__5 (
                    page1Out_14__5), .page1Out_4__4 (page1Out_14__4), .page1Out_4__3 (
                    page1Out_14__3), .page1Out_4__2 (page1Out_14__2), .page1Out_4__1 (
                    page1Out_14__1), .page1Out_4__0 (page1Out_14__0), .page2Out_0__15 (
                    page2Out_10__15), .page2Out_0__14 (page2Out_10__14), .page2Out_0__13 (
                    page2Out_10__13), .page2Out_0__12 (page2Out_10__12), .page2Out_0__11 (
                    page2Out_10__11), .page2Out_0__10 (page2Out_10__10), .page2Out_0__9 (
                    page2Out_10__9), .page2Out_0__8 (page2Out_10__8), .page2Out_0__7 (
                    page2Out_10__7), .page2Out_0__6 (page2Out_10__6), .page2Out_0__5 (
                    page2Out_10__5), .page2Out_0__4 (page2Out_10__4), .page2Out_0__3 (
                    page2Out_10__3), .page2Out_0__2 (page2Out_10__2), .page2Out_0__1 (
                    page2Out_10__1), .page2Out_0__0 (page2Out_10__0), .page2Out_1__15 (
                    page2Out_11__15), .page2Out_1__14 (page2Out_11__14), .page2Out_1__13 (
                    page2Out_11__13), .page2Out_1__12 (page2Out_11__12), .page2Out_1__11 (
                    page2Out_11__11), .page2Out_1__10 (page2Out_11__10), .page2Out_1__9 (
                    page2Out_11__9), .page2Out_1__8 (page2Out_11__8), .page2Out_1__7 (
                    page2Out_11__7), .page2Out_1__6 (page2Out_11__6), .page2Out_1__5 (
                    page2Out_11__5), .page2Out_1__4 (page2Out_11__4), .page2Out_1__3 (
                    page2Out_11__3), .page2Out_1__2 (page2Out_11__2), .page2Out_1__1 (
                    page2Out_11__1), .page2Out_1__0 (page2Out_11__0), .page2Out_2__15 (
                    page2Out_12__15), .page2Out_2__14 (page2Out_12__14), .page2Out_2__13 (
                    page2Out_12__13), .page2Out_2__12 (page2Out_12__12), .page2Out_2__11 (
                    page2Out_12__11), .page2Out_2__10 (page2Out_12__10), .page2Out_2__9 (
                    page2Out_12__9), .page2Out_2__8 (page2Out_12__8), .page2Out_2__7 (
                    page2Out_12__7), .page2Out_2__6 (page2Out_12__6), .page2Out_2__5 (
                    page2Out_12__5), .page2Out_2__4 (page2Out_12__4), .page2Out_2__3 (
                    page2Out_12__3), .page2Out_2__2 (page2Out_12__2), .page2Out_2__1 (
                    page2Out_12__1), .page2Out_2__0 (page2Out_12__0), .page2Out_3__15 (
                    page2Out_13__15), .page2Out_3__14 (page2Out_13__14), .page2Out_3__13 (
                    page2Out_13__13), .page2Out_3__12 (page2Out_13__12), .page2Out_3__11 (
                    page2Out_13__11), .page2Out_3__10 (page2Out_13__10), .page2Out_3__9 (
                    page2Out_13__9), .page2Out_3__8 (page2Out_13__8), .page2Out_3__7 (
                    page2Out_13__7), .page2Out_3__6 (page2Out_13__6), .page2Out_3__5 (
                    page2Out_13__5), .page2Out_3__4 (page2Out_13__4), .page2Out_3__3 (
                    page2Out_13__3), .page2Out_3__2 (page2Out_13__2), .page2Out_3__1 (
                    page2Out_13__1), .page2Out_3__0 (page2Out_13__0), .page2Out_4__15 (
                    page2Out_14__15), .page2Out_4__14 (page2Out_14__14), .page2Out_4__13 (
                    page2Out_14__13), .page2Out_4__12 (page2Out_14__12), .page2Out_4__11 (
                    page2Out_14__11), .page2Out_4__10 (page2Out_14__10), .page2Out_4__9 (
                    page2Out_14__9), .page2Out_4__8 (page2Out_14__8), .page2Out_4__7 (
                    page2Out_14__7), .page2Out_4__6 (page2Out_14__6), .page2Out_4__5 (
                    page2Out_14__5), .page2Out_4__4 (page2Out_14__4), .page2Out_4__3 (
                    page2Out_14__3), .page2Out_4__2 (page2Out_14__2), .page2Out_4__1 (
                    page2Out_14__1), .page2Out_4__0 (page2Out_14__0), .pagesOutsPrimary_0__15 (
                    pagesOuts_6__15), .pagesOutsPrimary_0__14 (pagesOuts_6__14)
                    , .pagesOutsPrimary_0__13 (pagesOuts_6__13), .pagesOutsPrimary_0__12 (
                    pagesOuts_6__12), .pagesOutsPrimary_0__11 (pagesOuts_6__11)
                    , .pagesOutsPrimary_0__10 (pagesOuts_6__10), .pagesOutsPrimary_0__9 (
                    pagesOuts_6__9), .pagesOutsPrimary_0__8 (pagesOuts_6__8), .pagesOutsPrimary_0__7 (
                    pagesOuts_6__7), .pagesOutsPrimary_0__6 (pagesOuts_6__6), .pagesOutsPrimary_0__5 (
                    pagesOuts_6__5), .pagesOutsPrimary_0__4 (pagesOuts_6__4), .pagesOutsPrimary_0__3 (
                    pagesOuts_6__3), .pagesOutsPrimary_0__2 (pagesOuts_6__2), .pagesOutsPrimary_0__1 (
                    pagesOuts_6__1), .pagesOutsPrimary_0__0 (pagesOuts_6__0), .pagesOutsPrimary_1__15 (
                    pagesOuts_7__15), .pagesOutsPrimary_1__14 (pagesOuts_7__14)
                    , .pagesOutsPrimary_1__13 (pagesOuts_7__13), .pagesOutsPrimary_1__12 (
                    pagesOuts_7__12), .pagesOutsPrimary_1__11 (pagesOuts_7__11)
                    , .pagesOutsPrimary_1__10 (pagesOuts_7__10), .pagesOutsPrimary_1__9 (
                    pagesOuts_7__9), .pagesOutsPrimary_1__8 (pagesOuts_7__8), .pagesOutsPrimary_1__7 (
                    pagesOuts_7__7), .pagesOutsPrimary_1__6 (pagesOuts_7__6), .pagesOutsPrimary_1__5 (
                    pagesOuts_7__5), .pagesOutsPrimary_1__4 (pagesOuts_7__4), .pagesOutsPrimary_1__3 (
                    pagesOuts_7__3), .pagesOutsPrimary_1__2 (pagesOuts_7__2), .pagesOutsPrimary_1__1 (
                    pagesOuts_7__1), .pagesOutsPrimary_1__0 (pagesOuts_7__0), .pagesOutsPrimary_2__15 (
                    pagesOuts_8__15), .pagesOutsPrimary_2__14 (pagesOuts_8__14)
                    , .pagesOutsPrimary_2__13 (pagesOuts_8__13), .pagesOutsPrimary_2__12 (
                    pagesOuts_8__12), .pagesOutsPrimary_2__11 (pagesOuts_8__11)
                    , .pagesOutsPrimary_2__10 (pagesOuts_8__10), .pagesOutsPrimary_2__9 (
                    pagesOuts_8__9), .pagesOutsPrimary_2__8 (pagesOuts_8__8), .pagesOutsPrimary_2__7 (
                    pagesOuts_8__7), .pagesOutsPrimary_2__6 (pagesOuts_8__6), .pagesOutsPrimary_2__5 (
                    pagesOuts_8__5), .pagesOutsPrimary_2__4 (pagesOuts_8__4), .pagesOutsPrimary_2__3 (
                    pagesOuts_8__3), .pagesOutsPrimary_2__2 (pagesOuts_8__2), .pagesOutsPrimary_2__1 (
                    pagesOuts_8__1), .pagesOutsPrimary_2__0 (pagesOuts_8__0), .pagesOutsSecondary_0__15 (
                    pagesOuts_19__15), .pagesOutsSecondary_0__14 (
                    pagesOuts_19__14), .pagesOutsSecondary_0__13 (
                    pagesOuts_19__13), .pagesOutsSecondary_0__12 (
                    pagesOuts_19__12), .pagesOutsSecondary_0__11 (
                    pagesOuts_19__11), .pagesOutsSecondary_0__10 (
                    pagesOuts_19__10), .pagesOutsSecondary_0__9 (pagesOuts_19__9
                    ), .pagesOutsSecondary_0__8 (pagesOuts_19__8), .pagesOutsSecondary_0__7 (
                    pagesOuts_19__7), .pagesOutsSecondary_0__6 (pagesOuts_19__6)
                    , .pagesOutsSecondary_0__5 (pagesOuts_19__5), .pagesOutsSecondary_0__4 (
                    pagesOuts_19__4), .pagesOutsSecondary_0__3 (pagesOuts_19__3)
                    , .pagesOutsSecondary_0__2 (pagesOuts_19__2), .pagesOutsSecondary_0__1 (
                    pagesOuts_19__1), .pagesOutsSecondary_0__0 (pagesOuts_19__0)
                    , .pagesOutsSecondary_1__15 (pagesOuts_20__15), .pagesOutsSecondary_1__14 (
                    pagesOuts_20__14), .pagesOutsSecondary_1__13 (
                    pagesOuts_20__13), .pagesOutsSecondary_1__12 (
                    pagesOuts_20__12), .pagesOutsSecondary_1__11 (
                    pagesOuts_20__11), .pagesOutsSecondary_1__10 (
                    pagesOuts_20__10), .pagesOutsSecondary_1__9 (pagesOuts_20__9
                    ), .pagesOutsSecondary_1__8 (pagesOuts_20__8), .pagesOutsSecondary_1__7 (
                    pagesOuts_20__7), .pagesOutsSecondary_1__6 (pagesOuts_20__6)
                    , .pagesOutsSecondary_1__5 (pagesOuts_20__5), .pagesOutsSecondary_1__4 (
                    pagesOuts_20__4), .pagesOutsSecondary_1__3 (pagesOuts_20__3)
                    , .pagesOutsSecondary_1__2 (pagesOuts_20__2), .pagesOutsSecondary_1__1 (
                    pagesOuts_20__1), .pagesOutsSecondary_1__0 (pagesOuts_20__0)
                    , .filtersOutsPrimary_0__7 (filtersOuts_6__7), .filtersOutsPrimary_0__6 (
                    filtersOuts_6__6), .filtersOutsPrimary_0__5 (
                    filtersOuts_6__5), .filtersOutsPrimary_0__4 (
                    filtersOuts_6__4), .filtersOutsPrimary_0__3 (
                    filtersOuts_6__3), .filtersOutsPrimary_0__2 (
                    filtersOuts_6__2), .filtersOutsPrimary_0__1 (
                    filtersOuts_6__1), .filtersOutsPrimary_0__0 (
                    filtersOuts_6__0), .filtersOutsPrimary_1__7 (
                    filtersOuts_7__7), .filtersOutsPrimary_1__6 (
                    filtersOuts_7__6), .filtersOutsPrimary_1__5 (
                    filtersOuts_7__5), .filtersOutsPrimary_1__4 (
                    filtersOuts_7__4), .filtersOutsPrimary_1__3 (
                    filtersOuts_7__3), .filtersOutsPrimary_1__2 (
                    filtersOuts_7__2), .filtersOutsPrimary_1__1 (
                    filtersOuts_7__1), .filtersOutsPrimary_1__0 (
                    filtersOuts_7__0), .filtersOutsPrimary_2__7 (
                    filtersOuts_8__7), .filtersOutsPrimary_2__6 (
                    filtersOuts_8__6), .filtersOutsPrimary_2__5 (
                    filtersOuts_8__5), .filtersOutsPrimary_2__4 (
                    filtersOuts_8__4), .filtersOutsPrimary_2__3 (
                    filtersOuts_8__3), .filtersOutsPrimary_2__2 (
                    filtersOuts_8__2), .filtersOutsPrimary_2__1 (
                    filtersOuts_8__1), .filtersOutsPrimary_2__0 (
                    filtersOuts_8__0), .filtersOutsSecondary_0__7 (
                    filtersOuts_19__7), .filtersOutsSecondary_0__6 (
                    filtersOuts_19__6), .filtersOutsSecondary_0__5 (
                    filtersOuts_19__5), .filtersOutsSecondary_0__4 (
                    filtersOuts_19__4), .filtersOutsSecondary_0__3 (
                    filtersOuts_19__3), .filtersOutsSecondary_0__2 (
                    filtersOuts_19__2), .filtersOutsSecondary_0__1 (
                    filtersOuts_19__1), .filtersOutsSecondary_0__0 (
                    filtersOuts_19__0), .filtersOutsSecondary_1__7 (
                    filtersOuts_20__7), .filtersOutsSecondary_1__6 (
                    filtersOuts_20__6), .filtersOutsSecondary_1__5 (
                    filtersOuts_20__5), .filtersOutsSecondary_1__4 (
                    filtersOuts_20__4), .filtersOutsSecondary_1__3 (
                    filtersOuts_20__3), .filtersOutsSecondary_1__2 (
                    filtersOuts_20__2), .filtersOutsSecondary_1__1 (
                    filtersOuts_20__1), .filtersOutsSecondary_1__0 (
                    filtersOuts_20__0)) ;
    RegRow_8_16_5_3 loop1_3_regRowMap (.filterBus ({filterBus[39],filterBus[38],
                    filterBus[37],filterBus[36],filterBus[35],filterBus[34],
                    filterBus[33],filterBus[32],filterBus[31],filterBus[30],
                    filterBus[29],filterBus[28],filterBus[27],filterBus[26],
                    filterBus[25],filterBus[24],filterBus[23],filterBus[22],
                    filterBus[21],filterBus[20],filterBus[19],filterBus[18],
                    filterBus[17],filterBus[16],filterBus[15],filterBus[14],
                    filterBus[13],filterBus[12],filterBus[11],filterBus[10],
                    filterBus[9],filterBus[8],filterBus[7],filterBus[6],
                    filterBus[5],filterBus[4],filterBus[3],filterBus[2],
                    filterBus[1],filterBus[0]}), .windowBus ({nx2802,nx2806,
                    nx2810,nx2814,nx2818,nx2822,nx2826,nx2830,nx2834,nx2838,
                    nx2842,nx2846,nx2850,nx2854,nx2858,nx2862,nx2866,nx2870,
                    nx2874,nx2878,nx2882,nx2886,nx2890,nx2894,nx2898,nx2902,
                    nx2906,nx2910,nx2914,nx2918,nx2922,nx2926,nx2930,nx2934,
                    nx2938,nx2942,nx2946,nx2950,nx2954,nx2958,nx2962,nx2966,
                    nx2970,nx2974,nx2978,nx2982,nx2986,nx2990,nx2994,nx2998,
                    nx3002,nx3006,nx3010,nx3014,nx3018,nx3022,nx3026,nx3030,
                    nx3034,nx3038,nx3042,nx3046,nx3050,nx3054,nx3058,nx3062,
                    nx3066,nx3070,nx3074,nx3078,nx3082,nx3086,nx3090,nx3094,
                    nx3098,nx3102,nx3106,nx3110,nx3114,nx3118}), .page1NextRow_0__15 (
                    page1Out_20__15), .page1NextRow_0__14 (page1Out_20__14), .page1NextRow_0__13 (
                    page1Out_20__13), .page1NextRow_0__12 (page1Out_20__12), .page1NextRow_0__11 (
                    page1Out_20__11), .page1NextRow_0__10 (page1Out_20__10), .page1NextRow_0__9 (
                    page1Out_20__9), .page1NextRow_0__8 (page1Out_20__8), .page1NextRow_0__7 (
                    page1Out_20__7), .page1NextRow_0__6 (page1Out_20__6), .page1NextRow_0__5 (
                    page1Out_20__5), .page1NextRow_0__4 (page1Out_20__4), .page1NextRow_0__3 (
                    page1Out_20__3), .page1NextRow_0__2 (page1Out_20__2), .page1NextRow_0__1 (
                    page1Out_20__1), .page1NextRow_0__0 (page1Out_20__0), .page1NextRow_1__15 (
                    page1Out_21__15), .page1NextRow_1__14 (page1Out_21__14), .page1NextRow_1__13 (
                    page1Out_21__13), .page1NextRow_1__12 (page1Out_21__12), .page1NextRow_1__11 (
                    page1Out_21__11), .page1NextRow_1__10 (page1Out_21__10), .page1NextRow_1__9 (
                    page1Out_21__9), .page1NextRow_1__8 (page1Out_21__8), .page1NextRow_1__7 (
                    page1Out_21__7), .page1NextRow_1__6 (page1Out_21__6), .page1NextRow_1__5 (
                    page1Out_21__5), .page1NextRow_1__4 (page1Out_21__4), .page1NextRow_1__3 (
                    page1Out_21__3), .page1NextRow_1__2 (page1Out_21__2), .page1NextRow_1__1 (
                    page1Out_21__1), .page1NextRow_1__0 (page1Out_21__0), .page1NextRow_2__15 (
                    page1Out_22__15), .page1NextRow_2__14 (page1Out_22__14), .page1NextRow_2__13 (
                    page1Out_22__13), .page1NextRow_2__12 (page1Out_22__12), .page1NextRow_2__11 (
                    page1Out_22__11), .page1NextRow_2__10 (page1Out_22__10), .page1NextRow_2__9 (
                    page1Out_22__9), .page1NextRow_2__8 (page1Out_22__8), .page1NextRow_2__7 (
                    page1Out_22__7), .page1NextRow_2__6 (page1Out_22__6), .page1NextRow_2__5 (
                    page1Out_22__5), .page1NextRow_2__4 (page1Out_22__4), .page1NextRow_2__3 (
                    page1Out_22__3), .page1NextRow_2__2 (page1Out_22__2), .page1NextRow_2__1 (
                    page1Out_22__1), .page1NextRow_2__0 (page1Out_22__0), .page1NextRow_3__15 (
                    page1Out_23__15), .page1NextRow_3__14 (page1Out_23__14), .page1NextRow_3__13 (
                    page1Out_23__13), .page1NextRow_3__12 (page1Out_23__12), .page1NextRow_3__11 (
                    page1Out_23__11), .page1NextRow_3__10 (page1Out_23__10), .page1NextRow_3__9 (
                    page1Out_23__9), .page1NextRow_3__8 (page1Out_23__8), .page1NextRow_3__7 (
                    page1Out_23__7), .page1NextRow_3__6 (page1Out_23__6), .page1NextRow_3__5 (
                    page1Out_23__5), .page1NextRow_3__4 (page1Out_23__4), .page1NextRow_3__3 (
                    page1Out_23__3), .page1NextRow_3__2 (page1Out_23__2), .page1NextRow_3__1 (
                    page1Out_23__1), .page1NextRow_3__0 (page1Out_23__0), .page1NextRow_4__15 (
                    page1Out_24__15), .page1NextRow_4__14 (page1Out_24__14), .page1NextRow_4__13 (
                    page1Out_24__13), .page1NextRow_4__12 (page1Out_24__12), .page1NextRow_4__11 (
                    page1Out_24__11), .page1NextRow_4__10 (page1Out_24__10), .page1NextRow_4__9 (
                    page1Out_24__9), .page1NextRow_4__8 (page1Out_24__8), .page1NextRow_4__7 (
                    page1Out_24__7), .page1NextRow_4__6 (page1Out_24__6), .page1NextRow_4__5 (
                    page1Out_24__5), .page1NextRow_4__4 (page1Out_24__4), .page1NextRow_4__3 (
                    page1Out_24__3), .page1NextRow_4__2 (page1Out_24__2), .page1NextRow_4__1 (
                    page1Out_24__1), .page1NextRow_4__0 (page1Out_24__0), .page2NextRow_0__15 (
                    page2Out_20__15), .page2NextRow_0__14 (page2Out_20__14), .page2NextRow_0__13 (
                    page2Out_20__13), .page2NextRow_0__12 (page2Out_20__12), .page2NextRow_0__11 (
                    page2Out_20__11), .page2NextRow_0__10 (page2Out_20__10), .page2NextRow_0__9 (
                    page2Out_20__9), .page2NextRow_0__8 (page2Out_20__8), .page2NextRow_0__7 (
                    page2Out_20__7), .page2NextRow_0__6 (page2Out_20__6), .page2NextRow_0__5 (
                    page2Out_20__5), .page2NextRow_0__4 (page2Out_20__4), .page2NextRow_0__3 (
                    page2Out_20__3), .page2NextRow_0__2 (page2Out_20__2), .page2NextRow_0__1 (
                    page2Out_20__1), .page2NextRow_0__0 (page2Out_20__0), .page2NextRow_1__15 (
                    page2Out_21__15), .page2NextRow_1__14 (page2Out_21__14), .page2NextRow_1__13 (
                    page2Out_21__13), .page2NextRow_1__12 (page2Out_21__12), .page2NextRow_1__11 (
                    page2Out_21__11), .page2NextRow_1__10 (page2Out_21__10), .page2NextRow_1__9 (
                    page2Out_21__9), .page2NextRow_1__8 (page2Out_21__8), .page2NextRow_1__7 (
                    page2Out_21__7), .page2NextRow_1__6 (page2Out_21__6), .page2NextRow_1__5 (
                    page2Out_21__5), .page2NextRow_1__4 (page2Out_21__4), .page2NextRow_1__3 (
                    page2Out_21__3), .page2NextRow_1__2 (page2Out_21__2), .page2NextRow_1__1 (
                    page2Out_21__1), .page2NextRow_1__0 (page2Out_21__0), .page2NextRow_2__15 (
                    page2Out_22__15), .page2NextRow_2__14 (page2Out_22__14), .page2NextRow_2__13 (
                    page2Out_22__13), .page2NextRow_2__12 (page2Out_22__12), .page2NextRow_2__11 (
                    page2Out_22__11), .page2NextRow_2__10 (page2Out_22__10), .page2NextRow_2__9 (
                    page2Out_22__9), .page2NextRow_2__8 (page2Out_22__8), .page2NextRow_2__7 (
                    page2Out_22__7), .page2NextRow_2__6 (page2Out_22__6), .page2NextRow_2__5 (
                    page2Out_22__5), .page2NextRow_2__4 (page2Out_22__4), .page2NextRow_2__3 (
                    page2Out_22__3), .page2NextRow_2__2 (page2Out_22__2), .page2NextRow_2__1 (
                    page2Out_22__1), .page2NextRow_2__0 (page2Out_22__0), .page2NextRow_3__15 (
                    page2Out_23__15), .page2NextRow_3__14 (page2Out_23__14), .page2NextRow_3__13 (
                    page2Out_23__13), .page2NextRow_3__12 (page2Out_23__12), .page2NextRow_3__11 (
                    page2Out_23__11), .page2NextRow_3__10 (page2Out_23__10), .page2NextRow_3__9 (
                    page2Out_23__9), .page2NextRow_3__8 (page2Out_23__8), .page2NextRow_3__7 (
                    page2Out_23__7), .page2NextRow_3__6 (page2Out_23__6), .page2NextRow_3__5 (
                    page2Out_23__5), .page2NextRow_3__4 (page2Out_23__4), .page2NextRow_3__3 (
                    page2Out_23__3), .page2NextRow_3__2 (page2Out_23__2), .page2NextRow_3__1 (
                    page2Out_23__1), .page2NextRow_3__0 (page2Out_23__0), .page2NextRow_4__15 (
                    page2Out_24__15), .page2NextRow_4__14 (page2Out_24__14), .page2NextRow_4__13 (
                    page2Out_24__13), .page2NextRow_4__12 (page2Out_24__12), .page2NextRow_4__11 (
                    page2Out_24__11), .page2NextRow_4__10 (page2Out_24__10), .page2NextRow_4__9 (
                    page2Out_24__9), .page2NextRow_4__8 (page2Out_24__8), .page2NextRow_4__7 (
                    page2Out_24__7), .page2NextRow_4__6 (page2Out_24__6), .page2NextRow_4__5 (
                    page2Out_24__5), .page2NextRow_4__4 (page2Out_24__4), .page2NextRow_4__3 (
                    page2Out_24__3), .page2NextRow_4__2 (page2Out_24__2), .page2NextRow_4__1 (
                    page2Out_24__1), .page2NextRow_4__0 (page2Out_24__0), .clk (
                    clk), .rst (rst), .enablePage1Read (page1Enables_3), .enablePage2Read (
                    page2Enables_3), .enableFilterRead (filterEnables_3), .shift2To1 (
                    nx3122), .shift1To2 (nx3126), .pageTurn (nx2796), .page1Out_0__15 (
                    page1Out_15__15), .page1Out_0__14 (page1Out_15__14), .page1Out_0__13 (
                    page1Out_15__13), .page1Out_0__12 (page1Out_15__12), .page1Out_0__11 (
                    page1Out_15__11), .page1Out_0__10 (page1Out_15__10), .page1Out_0__9 (
                    page1Out_15__9), .page1Out_0__8 (page1Out_15__8), .page1Out_0__7 (
                    page1Out_15__7), .page1Out_0__6 (page1Out_15__6), .page1Out_0__5 (
                    page1Out_15__5), .page1Out_0__4 (page1Out_15__4), .page1Out_0__3 (
                    page1Out_15__3), .page1Out_0__2 (page1Out_15__2), .page1Out_0__1 (
                    page1Out_15__1), .page1Out_0__0 (page1Out_15__0), .page1Out_1__15 (
                    page1Out_16__15), .page1Out_1__14 (page1Out_16__14), .page1Out_1__13 (
                    page1Out_16__13), .page1Out_1__12 (page1Out_16__12), .page1Out_1__11 (
                    page1Out_16__11), .page1Out_1__10 (page1Out_16__10), .page1Out_1__9 (
                    page1Out_16__9), .page1Out_1__8 (page1Out_16__8), .page1Out_1__7 (
                    page1Out_16__7), .page1Out_1__6 (page1Out_16__6), .page1Out_1__5 (
                    page1Out_16__5), .page1Out_1__4 (page1Out_16__4), .page1Out_1__3 (
                    page1Out_16__3), .page1Out_1__2 (page1Out_16__2), .page1Out_1__1 (
                    page1Out_16__1), .page1Out_1__0 (page1Out_16__0), .page1Out_2__15 (
                    page1Out_17__15), .page1Out_2__14 (page1Out_17__14), .page1Out_2__13 (
                    page1Out_17__13), .page1Out_2__12 (page1Out_17__12), .page1Out_2__11 (
                    page1Out_17__11), .page1Out_2__10 (page1Out_17__10), .page1Out_2__9 (
                    page1Out_17__9), .page1Out_2__8 (page1Out_17__8), .page1Out_2__7 (
                    page1Out_17__7), .page1Out_2__6 (page1Out_17__6), .page1Out_2__5 (
                    page1Out_17__5), .page1Out_2__4 (page1Out_17__4), .page1Out_2__3 (
                    page1Out_17__3), .page1Out_2__2 (page1Out_17__2), .page1Out_2__1 (
                    page1Out_17__1), .page1Out_2__0 (page1Out_17__0), .page1Out_3__15 (
                    page1Out_18__15), .page1Out_3__14 (page1Out_18__14), .page1Out_3__13 (
                    page1Out_18__13), .page1Out_3__12 (page1Out_18__12), .page1Out_3__11 (
                    page1Out_18__11), .page1Out_3__10 (page1Out_18__10), .page1Out_3__9 (
                    page1Out_18__9), .page1Out_3__8 (page1Out_18__8), .page1Out_3__7 (
                    page1Out_18__7), .page1Out_3__6 (page1Out_18__6), .page1Out_3__5 (
                    page1Out_18__5), .page1Out_3__4 (page1Out_18__4), .page1Out_3__3 (
                    page1Out_18__3), .page1Out_3__2 (page1Out_18__2), .page1Out_3__1 (
                    page1Out_18__1), .page1Out_3__0 (page1Out_18__0), .page1Out_4__15 (
                    page1Out_19__15), .page1Out_4__14 (page1Out_19__14), .page1Out_4__13 (
                    page1Out_19__13), .page1Out_4__12 (page1Out_19__12), .page1Out_4__11 (
                    page1Out_19__11), .page1Out_4__10 (page1Out_19__10), .page1Out_4__9 (
                    page1Out_19__9), .page1Out_4__8 (page1Out_19__8), .page1Out_4__7 (
                    page1Out_19__7), .page1Out_4__6 (page1Out_19__6), .page1Out_4__5 (
                    page1Out_19__5), .page1Out_4__4 (page1Out_19__4), .page1Out_4__3 (
                    page1Out_19__3), .page1Out_4__2 (page1Out_19__2), .page1Out_4__1 (
                    page1Out_19__1), .page1Out_4__0 (page1Out_19__0), .page2Out_0__15 (
                    page2Out_15__15), .page2Out_0__14 (page2Out_15__14), .page2Out_0__13 (
                    page2Out_15__13), .page2Out_0__12 (page2Out_15__12), .page2Out_0__11 (
                    page2Out_15__11), .page2Out_0__10 (page2Out_15__10), .page2Out_0__9 (
                    page2Out_15__9), .page2Out_0__8 (page2Out_15__8), .page2Out_0__7 (
                    page2Out_15__7), .page2Out_0__6 (page2Out_15__6), .page2Out_0__5 (
                    page2Out_15__5), .page2Out_0__4 (page2Out_15__4), .page2Out_0__3 (
                    page2Out_15__3), .page2Out_0__2 (page2Out_15__2), .page2Out_0__1 (
                    page2Out_15__1), .page2Out_0__0 (page2Out_15__0), .page2Out_1__15 (
                    page2Out_16__15), .page2Out_1__14 (page2Out_16__14), .page2Out_1__13 (
                    page2Out_16__13), .page2Out_1__12 (page2Out_16__12), .page2Out_1__11 (
                    page2Out_16__11), .page2Out_1__10 (page2Out_16__10), .page2Out_1__9 (
                    page2Out_16__9), .page2Out_1__8 (page2Out_16__8), .page2Out_1__7 (
                    page2Out_16__7), .page2Out_1__6 (page2Out_16__6), .page2Out_1__5 (
                    page2Out_16__5), .page2Out_1__4 (page2Out_16__4), .page2Out_1__3 (
                    page2Out_16__3), .page2Out_1__2 (page2Out_16__2), .page2Out_1__1 (
                    page2Out_16__1), .page2Out_1__0 (page2Out_16__0), .page2Out_2__15 (
                    page2Out_17__15), .page2Out_2__14 (page2Out_17__14), .page2Out_2__13 (
                    page2Out_17__13), .page2Out_2__12 (page2Out_17__12), .page2Out_2__11 (
                    page2Out_17__11), .page2Out_2__10 (page2Out_17__10), .page2Out_2__9 (
                    page2Out_17__9), .page2Out_2__8 (page2Out_17__8), .page2Out_2__7 (
                    page2Out_17__7), .page2Out_2__6 (page2Out_17__6), .page2Out_2__5 (
                    page2Out_17__5), .page2Out_2__4 (page2Out_17__4), .page2Out_2__3 (
                    page2Out_17__3), .page2Out_2__2 (page2Out_17__2), .page2Out_2__1 (
                    page2Out_17__1), .page2Out_2__0 (page2Out_17__0), .page2Out_3__15 (
                    page2Out_18__15), .page2Out_3__14 (page2Out_18__14), .page2Out_3__13 (
                    page2Out_18__13), .page2Out_3__12 (page2Out_18__12), .page2Out_3__11 (
                    page2Out_18__11), .page2Out_3__10 (page2Out_18__10), .page2Out_3__9 (
                    page2Out_18__9), .page2Out_3__8 (page2Out_18__8), .page2Out_3__7 (
                    page2Out_18__7), .page2Out_3__6 (page2Out_18__6), .page2Out_3__5 (
                    page2Out_18__5), .page2Out_3__4 (page2Out_18__4), .page2Out_3__3 (
                    page2Out_18__3), .page2Out_3__2 (page2Out_18__2), .page2Out_3__1 (
                    page2Out_18__1), .page2Out_3__0 (page2Out_18__0), .page2Out_4__15 (
                    page2Out_19__15), .page2Out_4__14 (page2Out_19__14), .page2Out_4__13 (
                    page2Out_19__13), .page2Out_4__12 (page2Out_19__12), .page2Out_4__11 (
                    page2Out_19__11), .page2Out_4__10 (page2Out_19__10), .page2Out_4__9 (
                    page2Out_19__9), .page2Out_4__8 (page2Out_19__8), .page2Out_4__7 (
                    page2Out_19__7), .page2Out_4__6 (page2Out_19__6), .page2Out_4__5 (
                    page2Out_19__5), .page2Out_4__4 (page2Out_19__4), .page2Out_4__3 (
                    page2Out_19__3), .page2Out_4__2 (page2Out_19__2), .page2Out_4__1 (
                    page2Out_19__1), .page2Out_4__0 (page2Out_19__0), .pagesOutsPrimary_0__15 (
                    pagesOuts_9__15), .pagesOutsPrimary_0__14 (pagesOuts_9__14)
                    , .pagesOutsPrimary_0__13 (pagesOuts_9__13), .pagesOutsPrimary_0__12 (
                    pagesOuts_9__12), .pagesOutsPrimary_0__11 (pagesOuts_9__11)
                    , .pagesOutsPrimary_0__10 (pagesOuts_9__10), .pagesOutsPrimary_0__9 (
                    pagesOuts_9__9), .pagesOutsPrimary_0__8 (pagesOuts_9__8), .pagesOutsPrimary_0__7 (
                    pagesOuts_9__7), .pagesOutsPrimary_0__6 (pagesOuts_9__6), .pagesOutsPrimary_0__5 (
                    pagesOuts_9__5), .pagesOutsPrimary_0__4 (pagesOuts_9__4), .pagesOutsPrimary_0__3 (
                    pagesOuts_9__3), .pagesOutsPrimary_0__2 (pagesOuts_9__2), .pagesOutsPrimary_0__1 (
                    pagesOuts_9__1), .pagesOutsPrimary_0__0 (pagesOuts_9__0), .pagesOutsPrimary_1__15 (
                    pagesOuts_10__15), .pagesOutsPrimary_1__14 (pagesOuts_10__14
                    ), .pagesOutsPrimary_1__13 (pagesOuts_10__13), .pagesOutsPrimary_1__12 (
                    pagesOuts_10__12), .pagesOutsPrimary_1__11 (pagesOuts_10__11
                    ), .pagesOutsPrimary_1__10 (pagesOuts_10__10), .pagesOutsPrimary_1__9 (
                    pagesOuts_10__9), .pagesOutsPrimary_1__8 (pagesOuts_10__8), 
                    .pagesOutsPrimary_1__7 (pagesOuts_10__7), .pagesOutsPrimary_1__6 (
                    pagesOuts_10__6), .pagesOutsPrimary_1__5 (pagesOuts_10__5), 
                    .pagesOutsPrimary_1__4 (pagesOuts_10__4), .pagesOutsPrimary_1__3 (
                    pagesOuts_10__3), .pagesOutsPrimary_1__2 (pagesOuts_10__2), 
                    .pagesOutsPrimary_1__1 (pagesOuts_10__1), .pagesOutsPrimary_1__0 (
                    pagesOuts_10__0), .pagesOutsPrimary_2__15 (pagesOuts_11__15)
                    , .pagesOutsPrimary_2__14 (pagesOuts_11__14), .pagesOutsPrimary_2__13 (
                    pagesOuts_11__13), .pagesOutsPrimary_2__12 (pagesOuts_11__12
                    ), .pagesOutsPrimary_2__11 (pagesOuts_11__11), .pagesOutsPrimary_2__10 (
                    pagesOuts_11__10), .pagesOutsPrimary_2__9 (pagesOuts_11__9)
                    , .pagesOutsPrimary_2__8 (pagesOuts_11__8), .pagesOutsPrimary_2__7 (
                    pagesOuts_11__7), .pagesOutsPrimary_2__6 (pagesOuts_11__6), 
                    .pagesOutsPrimary_2__5 (pagesOuts_11__5), .pagesOutsPrimary_2__4 (
                    pagesOuts_11__4), .pagesOutsPrimary_2__3 (pagesOuts_11__3), 
                    .pagesOutsPrimary_2__2 (pagesOuts_11__2), .pagesOutsPrimary_2__1 (
                    pagesOuts_11__1), .pagesOutsPrimary_2__0 (pagesOuts_11__0), 
                    .pagesOutsSecondary_0__15 (pagesOuts_21__15), .pagesOutsSecondary_0__14 (
                    pagesOuts_21__14), .pagesOutsSecondary_0__13 (
                    pagesOuts_21__13), .pagesOutsSecondary_0__12 (
                    pagesOuts_21__12), .pagesOutsSecondary_0__11 (
                    pagesOuts_21__11), .pagesOutsSecondary_0__10 (
                    pagesOuts_21__10), .pagesOutsSecondary_0__9 (pagesOuts_21__9
                    ), .pagesOutsSecondary_0__8 (pagesOuts_21__8), .pagesOutsSecondary_0__7 (
                    pagesOuts_21__7), .pagesOutsSecondary_0__6 (pagesOuts_21__6)
                    , .pagesOutsSecondary_0__5 (pagesOuts_21__5), .pagesOutsSecondary_0__4 (
                    pagesOuts_21__4), .pagesOutsSecondary_0__3 (pagesOuts_21__3)
                    , .pagesOutsSecondary_0__2 (pagesOuts_21__2), .pagesOutsSecondary_0__1 (
                    pagesOuts_21__1), .pagesOutsSecondary_0__0 (pagesOuts_21__0)
                    , .pagesOutsSecondary_1__15 (pagesOuts_22__15), .pagesOutsSecondary_1__14 (
                    pagesOuts_22__14), .pagesOutsSecondary_1__13 (
                    pagesOuts_22__13), .pagesOutsSecondary_1__12 (
                    pagesOuts_22__12), .pagesOutsSecondary_1__11 (
                    pagesOuts_22__11), .pagesOutsSecondary_1__10 (
                    pagesOuts_22__10), .pagesOutsSecondary_1__9 (pagesOuts_22__9
                    ), .pagesOutsSecondary_1__8 (pagesOuts_22__8), .pagesOutsSecondary_1__7 (
                    pagesOuts_22__7), .pagesOutsSecondary_1__6 (pagesOuts_22__6)
                    , .pagesOutsSecondary_1__5 (pagesOuts_22__5), .pagesOutsSecondary_1__4 (
                    pagesOuts_22__4), .pagesOutsSecondary_1__3 (pagesOuts_22__3)
                    , .pagesOutsSecondary_1__2 (pagesOuts_22__2), .pagesOutsSecondary_1__1 (
                    pagesOuts_22__1), .pagesOutsSecondary_1__0 (pagesOuts_22__0)
                    , .filtersOutsPrimary_0__7 (filtersOuts_9__7), .filtersOutsPrimary_0__6 (
                    filtersOuts_9__6), .filtersOutsPrimary_0__5 (
                    filtersOuts_9__5), .filtersOutsPrimary_0__4 (
                    filtersOuts_9__4), .filtersOutsPrimary_0__3 (
                    filtersOuts_9__3), .filtersOutsPrimary_0__2 (
                    filtersOuts_9__2), .filtersOutsPrimary_0__1 (
                    filtersOuts_9__1), .filtersOutsPrimary_0__0 (
                    filtersOuts_9__0), .filtersOutsPrimary_1__7 (
                    filtersOuts_10__7), .filtersOutsPrimary_1__6 (
                    filtersOuts_10__6), .filtersOutsPrimary_1__5 (
                    filtersOuts_10__5), .filtersOutsPrimary_1__4 (
                    filtersOuts_10__4), .filtersOutsPrimary_1__3 (
                    filtersOuts_10__3), .filtersOutsPrimary_1__2 (
                    filtersOuts_10__2), .filtersOutsPrimary_1__1 (
                    filtersOuts_10__1), .filtersOutsPrimary_1__0 (
                    filtersOuts_10__0), .filtersOutsPrimary_2__7 (
                    filtersOuts_11__7), .filtersOutsPrimary_2__6 (
                    filtersOuts_11__6), .filtersOutsPrimary_2__5 (
                    filtersOuts_11__5), .filtersOutsPrimary_2__4 (
                    filtersOuts_11__4), .filtersOutsPrimary_2__3 (
                    filtersOuts_11__3), .filtersOutsPrimary_2__2 (
                    filtersOuts_11__2), .filtersOutsPrimary_2__1 (
                    filtersOuts_11__1), .filtersOutsPrimary_2__0 (
                    filtersOuts_11__0), .filtersOutsSecondary_0__7 (
                    filtersOuts_21__7), .filtersOutsSecondary_0__6 (
                    filtersOuts_21__6), .filtersOutsSecondary_0__5 (
                    filtersOuts_21__5), .filtersOutsSecondary_0__4 (
                    filtersOuts_21__4), .filtersOutsSecondary_0__3 (
                    filtersOuts_21__3), .filtersOutsSecondary_0__2 (
                    filtersOuts_21__2), .filtersOutsSecondary_0__1 (
                    filtersOuts_21__1), .filtersOutsSecondary_0__0 (
                    filtersOuts_21__0), .filtersOutsSecondary_1__7 (
                    filtersOuts_22__7), .filtersOutsSecondary_1__6 (
                    filtersOuts_22__6), .filtersOutsSecondary_1__5 (
                    filtersOuts_22__5), .filtersOutsSecondary_1__4 (
                    filtersOuts_22__4), .filtersOutsSecondary_1__3 (
                    filtersOuts_22__3), .filtersOutsSecondary_1__2 (
                    filtersOuts_22__2), .filtersOutsSecondary_1__1 (
                    filtersOuts_22__1), .filtersOutsSecondary_1__0 (
                    filtersOuts_22__0)) ;
    RegRow_8_16_5_3 loop1_4_regRowMap (.filterBus ({filterBus[39],filterBus[38],
                    filterBus[37],filterBus[36],filterBus[35],filterBus[34],
                    filterBus[33],filterBus[32],filterBus[31],filterBus[30],
                    filterBus[29],filterBus[28],filterBus[27],filterBus[26],
                    filterBus[25],filterBus[24],filterBus[23],filterBus[22],
                    filterBus[21],filterBus[20],filterBus[19],filterBus[18],
                    filterBus[17],filterBus[16],filterBus[15],filterBus[14],
                    filterBus[13],filterBus[12],filterBus[11],filterBus[10],
                    filterBus[9],filterBus[8],filterBus[7],filterBus[6],
                    filterBus[5],filterBus[4],filterBus[3],filterBus[2],
                    filterBus[1],filterBus[0]}), .windowBus ({nx2802,nx2806,
                    nx2810,nx2814,nx2818,nx2822,nx2826,nx2830,nx2834,nx2838,
                    nx2842,nx2846,nx2850,nx2854,nx2858,nx2862,nx2866,nx2870,
                    nx2874,nx2878,nx2882,nx2886,nx2890,nx2894,nx2898,nx2902,
                    nx2906,nx2910,nx2914,nx2918,nx2922,nx2926,nx2930,nx2934,
                    nx2938,nx2942,nx2946,nx2950,nx2954,nx2958,nx2962,nx2966,
                    nx2970,nx2974,nx2978,nx2982,nx2986,nx2990,nx2994,nx2998,
                    nx3002,nx3006,nx3010,nx3014,nx3018,nx3022,nx3026,nx3030,
                    nx3034,nx3038,nx3042,nx3046,nx3050,nx3054,nx3058,nx3062,
                    nx3066,nx3070,nx3074,nx3078,nx3082,nx3086,nx3090,nx3094,
                    nx3098,nx3102,nx3106,nx3110,nx3114,nx3118}), .page1NextRow_0__15 (
                    page1Out_25__15), .page1NextRow_0__14 (page1Out_25__15), .page1NextRow_0__13 (
                    page1Out_25__15), .page1NextRow_0__12 (page1Out_25__15), .page1NextRow_0__11 (
                    page1Out_25__15), .page1NextRow_0__10 (page1Out_25__15), .page1NextRow_0__9 (
                    page1Out_25__15), .page1NextRow_0__8 (page1Out_25__15), .page1NextRow_0__7 (
                    page1Out_25__15), .page1NextRow_0__6 (page1Out_25__15), .page1NextRow_0__5 (
                    page1Out_25__15), .page1NextRow_0__4 (page1Out_25__15), .page1NextRow_0__3 (
                    page1Out_25__15), .page1NextRow_0__2 (page1Out_25__15), .page1NextRow_0__1 (
                    page1Out_25__15), .page1NextRow_0__0 (page1Out_25__15), .page1NextRow_1__15 (
                    page1Out_25__15), .page1NextRow_1__14 (page1Out_25__15), .page1NextRow_1__13 (
                    page1Out_25__15), .page1NextRow_1__12 (page1Out_25__15), .page1NextRow_1__11 (
                    page1Out_25__15), .page1NextRow_1__10 (page1Out_25__15), .page1NextRow_1__9 (
                    page1Out_25__15), .page1NextRow_1__8 (page1Out_25__15), .page1NextRow_1__7 (
                    page1Out_25__15), .page1NextRow_1__6 (page1Out_25__15), .page1NextRow_1__5 (
                    page1Out_25__15), .page1NextRow_1__4 (page1Out_25__15), .page1NextRow_1__3 (
                    page1Out_25__15), .page1NextRow_1__2 (page1Out_25__15), .page1NextRow_1__1 (
                    page1Out_25__15), .page1NextRow_1__0 (page1Out_25__15), .page1NextRow_2__15 (
                    page1Out_25__15), .page1NextRow_2__14 (page1Out_25__15), .page1NextRow_2__13 (
                    page1Out_25__15), .page1NextRow_2__12 (page1Out_25__15), .page1NextRow_2__11 (
                    page1Out_25__15), .page1NextRow_2__10 (page1Out_25__15), .page1NextRow_2__9 (
                    page1Out_25__15), .page1NextRow_2__8 (page1Out_25__15), .page1NextRow_2__7 (
                    page1Out_25__15), .page1NextRow_2__6 (page1Out_25__15), .page1NextRow_2__5 (
                    page1Out_25__15), .page1NextRow_2__4 (page1Out_25__15), .page1NextRow_2__3 (
                    page1Out_25__15), .page1NextRow_2__2 (page1Out_25__15), .page1NextRow_2__1 (
                    page1Out_25__15), .page1NextRow_2__0 (page1Out_25__15), .page1NextRow_3__15 (
                    page1Out_25__15), .page1NextRow_3__14 (page1Out_25__15), .page1NextRow_3__13 (
                    page1Out_25__15), .page1NextRow_3__12 (page1Out_25__15), .page1NextRow_3__11 (
                    page1Out_25__15), .page1NextRow_3__10 (page1Out_25__15), .page1NextRow_3__9 (
                    page1Out_25__15), .page1NextRow_3__8 (page1Out_25__15), .page1NextRow_3__7 (
                    page1Out_25__15), .page1NextRow_3__6 (page1Out_25__15), .page1NextRow_3__5 (
                    page1Out_25__15), .page1NextRow_3__4 (page1Out_25__15), .page1NextRow_3__3 (
                    page1Out_25__15), .page1NextRow_3__2 (page1Out_25__15), .page1NextRow_3__1 (
                    page1Out_25__15), .page1NextRow_3__0 (page1Out_25__15), .page1NextRow_4__15 (
                    page1Out_25__15), .page1NextRow_4__14 (page1Out_25__15), .page1NextRow_4__13 (
                    page1Out_25__15), .page1NextRow_4__12 (page1Out_25__15), .page1NextRow_4__11 (
                    page1Out_25__15), .page1NextRow_4__10 (page1Out_25__15), .page1NextRow_4__9 (
                    page1Out_25__15), .page1NextRow_4__8 (page1Out_25__15), .page1NextRow_4__7 (
                    page1Out_25__15), .page1NextRow_4__6 (page1Out_25__15), .page1NextRow_4__5 (
                    page1Out_25__15), .page1NextRow_4__4 (page1Out_25__15), .page1NextRow_4__3 (
                    page1Out_25__15), .page1NextRow_4__2 (page1Out_25__15), .page1NextRow_4__1 (
                    page1Out_25__15), .page1NextRow_4__0 (page1Out_25__15), .page2NextRow_0__15 (
                    page1Out_25__15), .page2NextRow_0__14 (page1Out_25__15), .page2NextRow_0__13 (
                    page1Out_25__15), .page2NextRow_0__12 (page1Out_25__15), .page2NextRow_0__11 (
                    page1Out_25__15), .page2NextRow_0__10 (page1Out_25__15), .page2NextRow_0__9 (
                    page1Out_25__15), .page2NextRow_0__8 (page1Out_25__15), .page2NextRow_0__7 (
                    page1Out_25__15), .page2NextRow_0__6 (page1Out_25__15), .page2NextRow_0__5 (
                    page1Out_25__15), .page2NextRow_0__4 (page1Out_25__15), .page2NextRow_0__3 (
                    page1Out_25__15), .page2NextRow_0__2 (page1Out_25__15), .page2NextRow_0__1 (
                    page1Out_25__15), .page2NextRow_0__0 (page1Out_25__15), .page2NextRow_1__15 (
                    page1Out_25__15), .page2NextRow_1__14 (page1Out_25__15), .page2NextRow_1__13 (
                    page1Out_25__15), .page2NextRow_1__12 (page1Out_25__15), .page2NextRow_1__11 (
                    page1Out_25__15), .page2NextRow_1__10 (page1Out_25__15), .page2NextRow_1__9 (
                    page1Out_25__15), .page2NextRow_1__8 (page1Out_25__15), .page2NextRow_1__7 (
                    page1Out_25__15), .page2NextRow_1__6 (page1Out_25__15), .page2NextRow_1__5 (
                    page1Out_25__15), .page2NextRow_1__4 (page1Out_25__15), .page2NextRow_1__3 (
                    page1Out_25__15), .page2NextRow_1__2 (page1Out_25__15), .page2NextRow_1__1 (
                    page1Out_25__15), .page2NextRow_1__0 (page1Out_25__15), .page2NextRow_2__15 (
                    page1Out_25__15), .page2NextRow_2__14 (page1Out_25__15), .page2NextRow_2__13 (
                    page1Out_25__15), .page2NextRow_2__12 (page1Out_25__15), .page2NextRow_2__11 (
                    page1Out_25__15), .page2NextRow_2__10 (page1Out_25__15), .page2NextRow_2__9 (
                    page1Out_25__15), .page2NextRow_2__8 (page1Out_25__15), .page2NextRow_2__7 (
                    page1Out_25__15), .page2NextRow_2__6 (page1Out_25__15), .page2NextRow_2__5 (
                    page1Out_25__15), .page2NextRow_2__4 (page1Out_25__15), .page2NextRow_2__3 (
                    page1Out_25__15), .page2NextRow_2__2 (page1Out_25__15), .page2NextRow_2__1 (
                    page1Out_25__15), .page2NextRow_2__0 (page1Out_25__15), .page2NextRow_3__15 (
                    page1Out_25__15), .page2NextRow_3__14 (page1Out_25__15), .page2NextRow_3__13 (
                    page1Out_25__15), .page2NextRow_3__12 (page1Out_25__15), .page2NextRow_3__11 (
                    page1Out_25__15), .page2NextRow_3__10 (page1Out_25__15), .page2NextRow_3__9 (
                    page1Out_25__15), .page2NextRow_3__8 (page1Out_25__15), .page2NextRow_3__7 (
                    page1Out_25__15), .page2NextRow_3__6 (page1Out_25__15), .page2NextRow_3__5 (
                    page1Out_25__15), .page2NextRow_3__4 (page1Out_25__15), .page2NextRow_3__3 (
                    page1Out_25__15), .page2NextRow_3__2 (page1Out_25__15), .page2NextRow_3__1 (
                    page1Out_25__15), .page2NextRow_3__0 (page1Out_25__15), .page2NextRow_4__15 (
                    page1Out_25__15), .page2NextRow_4__14 (page1Out_25__15), .page2NextRow_4__13 (
                    page1Out_25__15), .page2NextRow_4__12 (page1Out_25__15), .page2NextRow_4__11 (
                    page1Out_25__15), .page2NextRow_4__10 (page1Out_25__15), .page2NextRow_4__9 (
                    page1Out_25__15), .page2NextRow_4__8 (page1Out_25__15), .page2NextRow_4__7 (
                    page1Out_25__15), .page2NextRow_4__6 (page1Out_25__15), .page2NextRow_4__5 (
                    page1Out_25__15), .page2NextRow_4__4 (page1Out_25__15), .page2NextRow_4__3 (
                    page1Out_25__15), .page2NextRow_4__2 (page1Out_25__15), .page2NextRow_4__1 (
                    page1Out_25__15), .page2NextRow_4__0 (page1Out_25__15), .clk (
                    clk), .rst (rst), .enablePage1Read (page1Enables_4), .enablePage2Read (
                    page2Enables_4), .enableFilterRead (filterEnables_4), .shift2To1 (
                    nx3122), .shift1To2 (nx3126), .pageTurn (nx2798), .page1Out_0__15 (
                    page1Out_20__15), .page1Out_0__14 (page1Out_20__14), .page1Out_0__13 (
                    page1Out_20__13), .page1Out_0__12 (page1Out_20__12), .page1Out_0__11 (
                    page1Out_20__11), .page1Out_0__10 (page1Out_20__10), .page1Out_0__9 (
                    page1Out_20__9), .page1Out_0__8 (page1Out_20__8), .page1Out_0__7 (
                    page1Out_20__7), .page1Out_0__6 (page1Out_20__6), .page1Out_0__5 (
                    page1Out_20__5), .page1Out_0__4 (page1Out_20__4), .page1Out_0__3 (
                    page1Out_20__3), .page1Out_0__2 (page1Out_20__2), .page1Out_0__1 (
                    page1Out_20__1), .page1Out_0__0 (page1Out_20__0), .page1Out_1__15 (
                    page1Out_21__15), .page1Out_1__14 (page1Out_21__14), .page1Out_1__13 (
                    page1Out_21__13), .page1Out_1__12 (page1Out_21__12), .page1Out_1__11 (
                    page1Out_21__11), .page1Out_1__10 (page1Out_21__10), .page1Out_1__9 (
                    page1Out_21__9), .page1Out_1__8 (page1Out_21__8), .page1Out_1__7 (
                    page1Out_21__7), .page1Out_1__6 (page1Out_21__6), .page1Out_1__5 (
                    page1Out_21__5), .page1Out_1__4 (page1Out_21__4), .page1Out_1__3 (
                    page1Out_21__3), .page1Out_1__2 (page1Out_21__2), .page1Out_1__1 (
                    page1Out_21__1), .page1Out_1__0 (page1Out_21__0), .page1Out_2__15 (
                    page1Out_22__15), .page1Out_2__14 (page1Out_22__14), .page1Out_2__13 (
                    page1Out_22__13), .page1Out_2__12 (page1Out_22__12), .page1Out_2__11 (
                    page1Out_22__11), .page1Out_2__10 (page1Out_22__10), .page1Out_2__9 (
                    page1Out_22__9), .page1Out_2__8 (page1Out_22__8), .page1Out_2__7 (
                    page1Out_22__7), .page1Out_2__6 (page1Out_22__6), .page1Out_2__5 (
                    page1Out_22__5), .page1Out_2__4 (page1Out_22__4), .page1Out_2__3 (
                    page1Out_22__3), .page1Out_2__2 (page1Out_22__2), .page1Out_2__1 (
                    page1Out_22__1), .page1Out_2__0 (page1Out_22__0), .page1Out_3__15 (
                    page1Out_23__15), .page1Out_3__14 (page1Out_23__14), .page1Out_3__13 (
                    page1Out_23__13), .page1Out_3__12 (page1Out_23__12), .page1Out_3__11 (
                    page1Out_23__11), .page1Out_3__10 (page1Out_23__10), .page1Out_3__9 (
                    page1Out_23__9), .page1Out_3__8 (page1Out_23__8), .page1Out_3__7 (
                    page1Out_23__7), .page1Out_3__6 (page1Out_23__6), .page1Out_3__5 (
                    page1Out_23__5), .page1Out_3__4 (page1Out_23__4), .page1Out_3__3 (
                    page1Out_23__3), .page1Out_3__2 (page1Out_23__2), .page1Out_3__1 (
                    page1Out_23__1), .page1Out_3__0 (page1Out_23__0), .page1Out_4__15 (
                    page1Out_24__15), .page1Out_4__14 (page1Out_24__14), .page1Out_4__13 (
                    page1Out_24__13), .page1Out_4__12 (page1Out_24__12), .page1Out_4__11 (
                    page1Out_24__11), .page1Out_4__10 (page1Out_24__10), .page1Out_4__9 (
                    page1Out_24__9), .page1Out_4__8 (page1Out_24__8), .page1Out_4__7 (
                    page1Out_24__7), .page1Out_4__6 (page1Out_24__6), .page1Out_4__5 (
                    page1Out_24__5), .page1Out_4__4 (page1Out_24__4), .page1Out_4__3 (
                    page1Out_24__3), .page1Out_4__2 (page1Out_24__2), .page1Out_4__1 (
                    page1Out_24__1), .page1Out_4__0 (page1Out_24__0), .page2Out_0__15 (
                    page2Out_20__15), .page2Out_0__14 (page2Out_20__14), .page2Out_0__13 (
                    page2Out_20__13), .page2Out_0__12 (page2Out_20__12), .page2Out_0__11 (
                    page2Out_20__11), .page2Out_0__10 (page2Out_20__10), .page2Out_0__9 (
                    page2Out_20__9), .page2Out_0__8 (page2Out_20__8), .page2Out_0__7 (
                    page2Out_20__7), .page2Out_0__6 (page2Out_20__6), .page2Out_0__5 (
                    page2Out_20__5), .page2Out_0__4 (page2Out_20__4), .page2Out_0__3 (
                    page2Out_20__3), .page2Out_0__2 (page2Out_20__2), .page2Out_0__1 (
                    page2Out_20__1), .page2Out_0__0 (page2Out_20__0), .page2Out_1__15 (
                    page2Out_21__15), .page2Out_1__14 (page2Out_21__14), .page2Out_1__13 (
                    page2Out_21__13), .page2Out_1__12 (page2Out_21__12), .page2Out_1__11 (
                    page2Out_21__11), .page2Out_1__10 (page2Out_21__10), .page2Out_1__9 (
                    page2Out_21__9), .page2Out_1__8 (page2Out_21__8), .page2Out_1__7 (
                    page2Out_21__7), .page2Out_1__6 (page2Out_21__6), .page2Out_1__5 (
                    page2Out_21__5), .page2Out_1__4 (page2Out_21__4), .page2Out_1__3 (
                    page2Out_21__3), .page2Out_1__2 (page2Out_21__2), .page2Out_1__1 (
                    page2Out_21__1), .page2Out_1__0 (page2Out_21__0), .page2Out_2__15 (
                    page2Out_22__15), .page2Out_2__14 (page2Out_22__14), .page2Out_2__13 (
                    page2Out_22__13), .page2Out_2__12 (page2Out_22__12), .page2Out_2__11 (
                    page2Out_22__11), .page2Out_2__10 (page2Out_22__10), .page2Out_2__9 (
                    page2Out_22__9), .page2Out_2__8 (page2Out_22__8), .page2Out_2__7 (
                    page2Out_22__7), .page2Out_2__6 (page2Out_22__6), .page2Out_2__5 (
                    page2Out_22__5), .page2Out_2__4 (page2Out_22__4), .page2Out_2__3 (
                    page2Out_22__3), .page2Out_2__2 (page2Out_22__2), .page2Out_2__1 (
                    page2Out_22__1), .page2Out_2__0 (page2Out_22__0), .page2Out_3__15 (
                    page2Out_23__15), .page2Out_3__14 (page2Out_23__14), .page2Out_3__13 (
                    page2Out_23__13), .page2Out_3__12 (page2Out_23__12), .page2Out_3__11 (
                    page2Out_23__11), .page2Out_3__10 (page2Out_23__10), .page2Out_3__9 (
                    page2Out_23__9), .page2Out_3__8 (page2Out_23__8), .page2Out_3__7 (
                    page2Out_23__7), .page2Out_3__6 (page2Out_23__6), .page2Out_3__5 (
                    page2Out_23__5), .page2Out_3__4 (page2Out_23__4), .page2Out_3__3 (
                    page2Out_23__3), .page2Out_3__2 (page2Out_23__2), .page2Out_3__1 (
                    page2Out_23__1), .page2Out_3__0 (page2Out_23__0), .page2Out_4__15 (
                    page2Out_24__15), .page2Out_4__14 (page2Out_24__14), .page2Out_4__13 (
                    page2Out_24__13), .page2Out_4__12 (page2Out_24__12), .page2Out_4__11 (
                    page2Out_24__11), .page2Out_4__10 (page2Out_24__10), .page2Out_4__9 (
                    page2Out_24__9), .page2Out_4__8 (page2Out_24__8), .page2Out_4__7 (
                    page2Out_24__7), .page2Out_4__6 (page2Out_24__6), .page2Out_4__5 (
                    page2Out_24__5), .page2Out_4__4 (page2Out_24__4), .page2Out_4__3 (
                    page2Out_24__3), .page2Out_4__2 (page2Out_24__2), .page2Out_4__1 (
                    page2Out_24__1), .page2Out_4__0 (page2Out_24__0), .pagesOutsPrimary_0__15 (
                    pagesOuts_12__15), .pagesOutsPrimary_0__14 (pagesOuts_12__14
                    ), .pagesOutsPrimary_0__13 (pagesOuts_12__13), .pagesOutsPrimary_0__12 (
                    pagesOuts_12__12), .pagesOutsPrimary_0__11 (pagesOuts_12__11
                    ), .pagesOutsPrimary_0__10 (pagesOuts_12__10), .pagesOutsPrimary_0__9 (
                    pagesOuts_12__9), .pagesOutsPrimary_0__8 (pagesOuts_12__8), 
                    .pagesOutsPrimary_0__7 (pagesOuts_12__7), .pagesOutsPrimary_0__6 (
                    pagesOuts_12__6), .pagesOutsPrimary_0__5 (pagesOuts_12__5), 
                    .pagesOutsPrimary_0__4 (pagesOuts_12__4), .pagesOutsPrimary_0__3 (
                    pagesOuts_12__3), .pagesOutsPrimary_0__2 (pagesOuts_12__2), 
                    .pagesOutsPrimary_0__1 (pagesOuts_12__1), .pagesOutsPrimary_0__0 (
                    pagesOuts_12__0), .pagesOutsPrimary_1__15 (pagesOuts_13__15)
                    , .pagesOutsPrimary_1__14 (pagesOuts_13__14), .pagesOutsPrimary_1__13 (
                    pagesOuts_13__13), .pagesOutsPrimary_1__12 (pagesOuts_13__12
                    ), .pagesOutsPrimary_1__11 (pagesOuts_13__11), .pagesOutsPrimary_1__10 (
                    pagesOuts_13__10), .pagesOutsPrimary_1__9 (pagesOuts_13__9)
                    , .pagesOutsPrimary_1__8 (pagesOuts_13__8), .pagesOutsPrimary_1__7 (
                    pagesOuts_13__7), .pagesOutsPrimary_1__6 (pagesOuts_13__6), 
                    .pagesOutsPrimary_1__5 (pagesOuts_13__5), .pagesOutsPrimary_1__4 (
                    pagesOuts_13__4), .pagesOutsPrimary_1__3 (pagesOuts_13__3), 
                    .pagesOutsPrimary_1__2 (pagesOuts_13__2), .pagesOutsPrimary_1__1 (
                    pagesOuts_13__1), .pagesOutsPrimary_1__0 (pagesOuts_13__0), 
                    .pagesOutsPrimary_2__15 (pagesOuts_14__15), .pagesOutsPrimary_2__14 (
                    pagesOuts_14__14), .pagesOutsPrimary_2__13 (pagesOuts_14__13
                    ), .pagesOutsPrimary_2__12 (pagesOuts_14__12), .pagesOutsPrimary_2__11 (
                    pagesOuts_14__11), .pagesOutsPrimary_2__10 (pagesOuts_14__10
                    ), .pagesOutsPrimary_2__9 (pagesOuts_14__9), .pagesOutsPrimary_2__8 (
                    pagesOuts_14__8), .pagesOutsPrimary_2__7 (pagesOuts_14__7), 
                    .pagesOutsPrimary_2__6 (pagesOuts_14__6), .pagesOutsPrimary_2__5 (
                    pagesOuts_14__5), .pagesOutsPrimary_2__4 (pagesOuts_14__4), 
                    .pagesOutsPrimary_2__3 (pagesOuts_14__3), .pagesOutsPrimary_2__2 (
                    pagesOuts_14__2), .pagesOutsPrimary_2__1 (pagesOuts_14__1), 
                    .pagesOutsPrimary_2__0 (pagesOuts_14__0), .pagesOutsSecondary_0__15 (
                    pagesOuts_23__15), .pagesOutsSecondary_0__14 (
                    pagesOuts_23__14), .pagesOutsSecondary_0__13 (
                    pagesOuts_23__13), .pagesOutsSecondary_0__12 (
                    pagesOuts_23__12), .pagesOutsSecondary_0__11 (
                    pagesOuts_23__11), .pagesOutsSecondary_0__10 (
                    pagesOuts_23__10), .pagesOutsSecondary_0__9 (pagesOuts_23__9
                    ), .pagesOutsSecondary_0__8 (pagesOuts_23__8), .pagesOutsSecondary_0__7 (
                    pagesOuts_23__7), .pagesOutsSecondary_0__6 (pagesOuts_23__6)
                    , .pagesOutsSecondary_0__5 (pagesOuts_23__5), .pagesOutsSecondary_0__4 (
                    pagesOuts_23__4), .pagesOutsSecondary_0__3 (pagesOuts_23__3)
                    , .pagesOutsSecondary_0__2 (pagesOuts_23__2), .pagesOutsSecondary_0__1 (
                    pagesOuts_23__1), .pagesOutsSecondary_0__0 (pagesOuts_23__0)
                    , .pagesOutsSecondary_1__15 (pagesOuts_24__15), .pagesOutsSecondary_1__14 (
                    pagesOuts_24__14), .pagesOutsSecondary_1__13 (
                    pagesOuts_24__13), .pagesOutsSecondary_1__12 (
                    pagesOuts_24__12), .pagesOutsSecondary_1__11 (
                    pagesOuts_24__11), .pagesOutsSecondary_1__10 (
                    pagesOuts_24__10), .pagesOutsSecondary_1__9 (pagesOuts_24__9
                    ), .pagesOutsSecondary_1__8 (pagesOuts_24__8), .pagesOutsSecondary_1__7 (
                    pagesOuts_24__7), .pagesOutsSecondary_1__6 (pagesOuts_24__6)
                    , .pagesOutsSecondary_1__5 (pagesOuts_24__5), .pagesOutsSecondary_1__4 (
                    pagesOuts_24__4), .pagesOutsSecondary_1__3 (pagesOuts_24__3)
                    , .pagesOutsSecondary_1__2 (pagesOuts_24__2), .pagesOutsSecondary_1__1 (
                    pagesOuts_24__1), .pagesOutsSecondary_1__0 (pagesOuts_24__0)
                    , .filtersOutsPrimary_0__7 (filtersOuts_12__7), .filtersOutsPrimary_0__6 (
                    filtersOuts_12__6), .filtersOutsPrimary_0__5 (
                    filtersOuts_12__5), .filtersOutsPrimary_0__4 (
                    filtersOuts_12__4), .filtersOutsPrimary_0__3 (
                    filtersOuts_12__3), .filtersOutsPrimary_0__2 (
                    filtersOuts_12__2), .filtersOutsPrimary_0__1 (
                    filtersOuts_12__1), .filtersOutsPrimary_0__0 (
                    filtersOuts_12__0), .filtersOutsPrimary_1__7 (
                    filtersOuts_13__7), .filtersOutsPrimary_1__6 (
                    filtersOuts_13__6), .filtersOutsPrimary_1__5 (
                    filtersOuts_13__5), .filtersOutsPrimary_1__4 (
                    filtersOuts_13__4), .filtersOutsPrimary_1__3 (
                    filtersOuts_13__3), .filtersOutsPrimary_1__2 (
                    filtersOuts_13__2), .filtersOutsPrimary_1__1 (
                    filtersOuts_13__1), .filtersOutsPrimary_1__0 (
                    filtersOuts_13__0), .filtersOutsPrimary_2__7 (
                    filtersOuts_14__7), .filtersOutsPrimary_2__6 (
                    filtersOuts_14__6), .filtersOutsPrimary_2__5 (
                    filtersOuts_14__5), .filtersOutsPrimary_2__4 (
                    filtersOuts_14__4), .filtersOutsPrimary_2__3 (
                    filtersOuts_14__3), .filtersOutsPrimary_2__2 (
                    filtersOuts_14__2), .filtersOutsPrimary_2__1 (
                    filtersOuts_14__1), .filtersOutsPrimary_2__0 (
                    filtersOuts_14__0), .filtersOutsSecondary_0__7 (
                    filtersOuts_23__7), .filtersOutsSecondary_0__6 (
                    filtersOuts_23__6), .filtersOutsSecondary_0__5 (
                    filtersOuts_23__5), .filtersOutsSecondary_0__4 (
                    filtersOuts_23__4), .filtersOutsSecondary_0__3 (
                    filtersOuts_23__3), .filtersOutsSecondary_0__2 (
                    filtersOuts_23__2), .filtersOutsSecondary_0__1 (
                    filtersOuts_23__1), .filtersOutsSecondary_0__0 (
                    filtersOuts_23__0), .filtersOutsSecondary_1__7 (
                    filtersOuts_24__7), .filtersOutsSecondary_1__6 (
                    filtersOuts_24__6), .filtersOutsSecondary_1__5 (
                    filtersOuts_24__5), .filtersOutsSecondary_1__4 (
                    filtersOuts_24__4), .filtersOutsSecondary_1__3 (
                    filtersOuts_24__3), .filtersOutsSecondary_1__2 (
                    filtersOuts_24__2), .filtersOutsSecondary_1__1 (
                    filtersOuts_24__1), .filtersOutsSecondary_1__0 (
                    filtersOuts_24__0)) ;
    fake_gnd ix2748 (.Y (page1Out_25__15)) ;
    or03 ix33 (.Y (decoderRowEnable), .A0 (enablePage2Read), .A1 (
         enableFilterRead), .A2 (enablePage1Read)) ;
    and02 ix1 (.Y (filterEnables_4), .A0 (decodedRow_4), .A1 (enableFilterRead)
          ) ;
    and02 ix7 (.Y (filterEnables_3), .A0 (decodedRow_3), .A1 (enableFilterRead)
          ) ;
    and02 ix13 (.Y (filterEnables_2), .A0 (decodedRow_2), .A1 (enableFilterRead)
          ) ;
    and02 ix19 (.Y (filterEnables_1), .A0 (decodedRow_1), .A1 (enableFilterRead)
          ) ;
    and02 ix25 (.Y (filterEnables_0), .A0 (decodedRow_0), .A1 (enableFilterRead)
          ) ;
    and02 ix3 (.Y (page2Enables_4), .A0 (decodedRow_4), .A1 (enablePage2Read)) ;
    and02 ix9 (.Y (page2Enables_3), .A0 (decodedRow_3), .A1 (enablePage2Read)) ;
    and02 ix15 (.Y (page2Enables_2), .A0 (decodedRow_2), .A1 (enablePage2Read)
          ) ;
    and02 ix21 (.Y (page2Enables_1), .A0 (decodedRow_1), .A1 (enablePage2Read)
          ) ;
    and02 ix27 (.Y (page2Enables_0), .A0 (decodedRow_0), .A1 (enablePage2Read)
          ) ;
    and02 ix5 (.Y (page1Enables_4), .A0 (decodedRow_4), .A1 (enablePage1Read)) ;
    and02 ix11 (.Y (page1Enables_3), .A0 (decodedRow_3), .A1 (enablePage1Read)
          ) ;
    and02 ix17 (.Y (page1Enables_2), .A0 (decodedRow_2), .A1 (enablePage1Read)
          ) ;
    and02 ix23 (.Y (page1Enables_1), .A0 (decodedRow_1), .A1 (enablePage1Read)
          ) ;
    and02 ix29 (.Y (page1Enables_0), .A0 (decodedRow_0), .A1 (enablePage1Read)
          ) ;
    inv01 ix2787 (.Y (nx2788), .A (pageTurn)) ;
    inv01 ix2789 (.Y (nx2790), .A (nx2788)) ;
    inv01 ix2791 (.Y (nx2792), .A (nx2788)) ;
    inv01 ix2793 (.Y (nx2794), .A (nx2788)) ;
    inv01 ix2795 (.Y (nx2796), .A (nx2788)) ;
    inv01 ix2797 (.Y (nx2798), .A (nx2788)) ;
    buf02 ix2799 (.Y (nx2800), .A (windowBus[79])) ;
    buf02 ix2801 (.Y (nx2802), .A (windowBus[79])) ;
    buf02 ix2803 (.Y (nx2804), .A (windowBus[78])) ;
    buf02 ix2805 (.Y (nx2806), .A (windowBus[78])) ;
    buf02 ix2807 (.Y (nx2808), .A (windowBus[77])) ;
    buf02 ix2809 (.Y (nx2810), .A (windowBus[77])) ;
    buf02 ix2811 (.Y (nx2812), .A (windowBus[76])) ;
    buf02 ix2813 (.Y (nx2814), .A (windowBus[76])) ;
    buf02 ix2815 (.Y (nx2816), .A (windowBus[75])) ;
    buf02 ix2817 (.Y (nx2818), .A (windowBus[75])) ;
    buf02 ix2819 (.Y (nx2820), .A (windowBus[74])) ;
    buf02 ix2821 (.Y (nx2822), .A (windowBus[74])) ;
    buf02 ix2823 (.Y (nx2824), .A (windowBus[73])) ;
    buf02 ix2825 (.Y (nx2826), .A (windowBus[73])) ;
    buf02 ix2827 (.Y (nx2828), .A (windowBus[72])) ;
    buf02 ix2829 (.Y (nx2830), .A (windowBus[72])) ;
    buf02 ix2831 (.Y (nx2832), .A (windowBus[71])) ;
    buf02 ix2833 (.Y (nx2834), .A (windowBus[71])) ;
    buf02 ix2835 (.Y (nx2836), .A (windowBus[70])) ;
    buf02 ix2837 (.Y (nx2838), .A (windowBus[70])) ;
    buf02 ix2839 (.Y (nx2840), .A (windowBus[69])) ;
    buf02 ix2841 (.Y (nx2842), .A (windowBus[69])) ;
    buf02 ix2843 (.Y (nx2844), .A (windowBus[68])) ;
    buf02 ix2845 (.Y (nx2846), .A (windowBus[68])) ;
    buf02 ix2847 (.Y (nx2848), .A (windowBus[67])) ;
    buf02 ix2849 (.Y (nx2850), .A (windowBus[67])) ;
    buf02 ix2851 (.Y (nx2852), .A (windowBus[66])) ;
    buf02 ix2853 (.Y (nx2854), .A (windowBus[66])) ;
    buf02 ix2855 (.Y (nx2856), .A (windowBus[65])) ;
    buf02 ix2857 (.Y (nx2858), .A (windowBus[65])) ;
    buf02 ix2859 (.Y (nx2860), .A (windowBus[64])) ;
    buf02 ix2861 (.Y (nx2862), .A (windowBus[64])) ;
    buf02 ix2863 (.Y (nx2864), .A (windowBus[63])) ;
    buf02 ix2865 (.Y (nx2866), .A (windowBus[63])) ;
    buf02 ix2867 (.Y (nx2868), .A (windowBus[62])) ;
    buf02 ix2869 (.Y (nx2870), .A (windowBus[62])) ;
    buf02 ix2871 (.Y (nx2872), .A (windowBus[61])) ;
    buf02 ix2873 (.Y (nx2874), .A (windowBus[61])) ;
    buf02 ix2875 (.Y (nx2876), .A (windowBus[60])) ;
    buf02 ix2877 (.Y (nx2878), .A (windowBus[60])) ;
    buf02 ix2879 (.Y (nx2880), .A (windowBus[59])) ;
    buf02 ix2881 (.Y (nx2882), .A (windowBus[59])) ;
    buf02 ix2883 (.Y (nx2884), .A (windowBus[58])) ;
    buf02 ix2885 (.Y (nx2886), .A (windowBus[58])) ;
    buf02 ix2887 (.Y (nx2888), .A (windowBus[57])) ;
    buf02 ix2889 (.Y (nx2890), .A (windowBus[57])) ;
    buf02 ix2891 (.Y (nx2892), .A (windowBus[56])) ;
    buf02 ix2893 (.Y (nx2894), .A (windowBus[56])) ;
    buf02 ix2895 (.Y (nx2896), .A (windowBus[55])) ;
    buf02 ix2897 (.Y (nx2898), .A (windowBus[55])) ;
    buf02 ix2899 (.Y (nx2900), .A (windowBus[54])) ;
    buf02 ix2901 (.Y (nx2902), .A (windowBus[54])) ;
    buf02 ix2903 (.Y (nx2904), .A (windowBus[53])) ;
    buf02 ix2905 (.Y (nx2906), .A (windowBus[53])) ;
    buf02 ix2907 (.Y (nx2908), .A (windowBus[52])) ;
    buf02 ix2909 (.Y (nx2910), .A (windowBus[52])) ;
    buf02 ix2911 (.Y (nx2912), .A (windowBus[51])) ;
    buf02 ix2913 (.Y (nx2914), .A (windowBus[51])) ;
    buf02 ix2915 (.Y (nx2916), .A (windowBus[50])) ;
    buf02 ix2917 (.Y (nx2918), .A (windowBus[50])) ;
    buf02 ix2919 (.Y (nx2920), .A (windowBus[49])) ;
    buf02 ix2921 (.Y (nx2922), .A (windowBus[49])) ;
    buf02 ix2923 (.Y (nx2924), .A (windowBus[48])) ;
    buf02 ix2925 (.Y (nx2926), .A (windowBus[48])) ;
    buf02 ix2927 (.Y (nx2928), .A (windowBus[47])) ;
    buf02 ix2929 (.Y (nx2930), .A (windowBus[47])) ;
    buf02 ix2931 (.Y (nx2932), .A (windowBus[46])) ;
    buf02 ix2933 (.Y (nx2934), .A (windowBus[46])) ;
    buf02 ix2935 (.Y (nx2936), .A (windowBus[45])) ;
    buf02 ix2937 (.Y (nx2938), .A (windowBus[45])) ;
    buf02 ix2939 (.Y (nx2940), .A (windowBus[44])) ;
    buf02 ix2941 (.Y (nx2942), .A (windowBus[44])) ;
    buf02 ix2943 (.Y (nx2944), .A (windowBus[43])) ;
    buf02 ix2945 (.Y (nx2946), .A (windowBus[43])) ;
    buf02 ix2947 (.Y (nx2948), .A (windowBus[42])) ;
    buf02 ix2949 (.Y (nx2950), .A (windowBus[42])) ;
    buf02 ix2951 (.Y (nx2952), .A (windowBus[41])) ;
    buf02 ix2953 (.Y (nx2954), .A (windowBus[41])) ;
    buf02 ix2955 (.Y (nx2956), .A (windowBus[40])) ;
    buf02 ix2957 (.Y (nx2958), .A (windowBus[40])) ;
    buf02 ix2959 (.Y (nx2960), .A (windowBus[39])) ;
    buf02 ix2961 (.Y (nx2962), .A (windowBus[39])) ;
    buf02 ix2963 (.Y (nx2964), .A (windowBus[38])) ;
    buf02 ix2965 (.Y (nx2966), .A (windowBus[38])) ;
    buf02 ix2967 (.Y (nx2968), .A (windowBus[37])) ;
    buf02 ix2969 (.Y (nx2970), .A (windowBus[37])) ;
    buf02 ix2971 (.Y (nx2972), .A (windowBus[36])) ;
    buf02 ix2973 (.Y (nx2974), .A (windowBus[36])) ;
    buf02 ix2975 (.Y (nx2976), .A (windowBus[35])) ;
    buf02 ix2977 (.Y (nx2978), .A (windowBus[35])) ;
    buf02 ix2979 (.Y (nx2980), .A (windowBus[34])) ;
    buf02 ix2981 (.Y (nx2982), .A (windowBus[34])) ;
    buf02 ix2983 (.Y (nx2984), .A (windowBus[33])) ;
    buf02 ix2985 (.Y (nx2986), .A (windowBus[33])) ;
    buf02 ix2987 (.Y (nx2988), .A (windowBus[32])) ;
    buf02 ix2989 (.Y (nx2990), .A (windowBus[32])) ;
    buf02 ix2991 (.Y (nx2992), .A (windowBus[31])) ;
    buf02 ix2993 (.Y (nx2994), .A (windowBus[31])) ;
    buf02 ix2995 (.Y (nx2996), .A (windowBus[30])) ;
    buf02 ix2997 (.Y (nx2998), .A (windowBus[30])) ;
    buf02 ix2999 (.Y (nx3000), .A (windowBus[29])) ;
    buf02 ix3001 (.Y (nx3002), .A (windowBus[29])) ;
    buf02 ix3003 (.Y (nx3004), .A (windowBus[28])) ;
    buf02 ix3005 (.Y (nx3006), .A (windowBus[28])) ;
    buf02 ix3007 (.Y (nx3008), .A (windowBus[27])) ;
    buf02 ix3009 (.Y (nx3010), .A (windowBus[27])) ;
    buf02 ix3011 (.Y (nx3012), .A (windowBus[26])) ;
    buf02 ix3013 (.Y (nx3014), .A (windowBus[26])) ;
    buf02 ix3015 (.Y (nx3016), .A (windowBus[25])) ;
    buf02 ix3017 (.Y (nx3018), .A (windowBus[25])) ;
    buf02 ix3019 (.Y (nx3020), .A (windowBus[24])) ;
    buf02 ix3021 (.Y (nx3022), .A (windowBus[24])) ;
    buf02 ix3023 (.Y (nx3024), .A (windowBus[23])) ;
    buf02 ix3025 (.Y (nx3026), .A (windowBus[23])) ;
    buf02 ix3027 (.Y (nx3028), .A (windowBus[22])) ;
    buf02 ix3029 (.Y (nx3030), .A (windowBus[22])) ;
    buf02 ix3031 (.Y (nx3032), .A (windowBus[21])) ;
    buf02 ix3033 (.Y (nx3034), .A (windowBus[21])) ;
    buf02 ix3035 (.Y (nx3036), .A (windowBus[20])) ;
    buf02 ix3037 (.Y (nx3038), .A (windowBus[20])) ;
    buf02 ix3039 (.Y (nx3040), .A (windowBus[19])) ;
    buf02 ix3041 (.Y (nx3042), .A (windowBus[19])) ;
    buf02 ix3043 (.Y (nx3044), .A (windowBus[18])) ;
    buf02 ix3045 (.Y (nx3046), .A (windowBus[18])) ;
    buf02 ix3047 (.Y (nx3048), .A (windowBus[17])) ;
    buf02 ix3049 (.Y (nx3050), .A (windowBus[17])) ;
    buf02 ix3051 (.Y (nx3052), .A (windowBus[16])) ;
    buf02 ix3053 (.Y (nx3054), .A (windowBus[16])) ;
    buf02 ix3055 (.Y (nx3056), .A (windowBus[15])) ;
    buf02 ix3057 (.Y (nx3058), .A (windowBus[15])) ;
    buf02 ix3059 (.Y (nx3060), .A (windowBus[14])) ;
    buf02 ix3061 (.Y (nx3062), .A (windowBus[14])) ;
    buf02 ix3063 (.Y (nx3064), .A (windowBus[13])) ;
    buf02 ix3065 (.Y (nx3066), .A (windowBus[13])) ;
    buf02 ix3067 (.Y (nx3068), .A (windowBus[12])) ;
    buf02 ix3069 (.Y (nx3070), .A (windowBus[12])) ;
    buf02 ix3071 (.Y (nx3072), .A (windowBus[11])) ;
    buf02 ix3073 (.Y (nx3074), .A (windowBus[11])) ;
    buf02 ix3075 (.Y (nx3076), .A (windowBus[10])) ;
    buf02 ix3077 (.Y (nx3078), .A (windowBus[10])) ;
    buf02 ix3079 (.Y (nx3080), .A (windowBus[9])) ;
    buf02 ix3081 (.Y (nx3082), .A (windowBus[9])) ;
    buf02 ix3083 (.Y (nx3084), .A (windowBus[8])) ;
    buf02 ix3085 (.Y (nx3086), .A (windowBus[8])) ;
    buf02 ix3087 (.Y (nx3088), .A (windowBus[7])) ;
    buf02 ix3089 (.Y (nx3090), .A (windowBus[7])) ;
    buf02 ix3091 (.Y (nx3092), .A (windowBus[6])) ;
    buf02 ix3093 (.Y (nx3094), .A (windowBus[6])) ;
    buf02 ix3095 (.Y (nx3096), .A (windowBus[5])) ;
    buf02 ix3097 (.Y (nx3098), .A (windowBus[5])) ;
    buf02 ix3099 (.Y (nx3100), .A (windowBus[4])) ;
    buf02 ix3101 (.Y (nx3102), .A (windowBus[4])) ;
    buf02 ix3103 (.Y (nx3104), .A (windowBus[3])) ;
    buf02 ix3105 (.Y (nx3106), .A (windowBus[3])) ;
    buf02 ix3107 (.Y (nx3108), .A (windowBus[2])) ;
    buf02 ix3109 (.Y (nx3110), .A (windowBus[2])) ;
    buf02 ix3111 (.Y (nx3112), .A (windowBus[1])) ;
    buf02 ix3113 (.Y (nx3114), .A (windowBus[1])) ;
    buf02 ix3115 (.Y (nx3116), .A (windowBus[0])) ;
    buf02 ix3117 (.Y (nx3118), .A (windowBus[0])) ;
    buf02 ix3119 (.Y (nx3120), .A (shift2To1)) ;
    buf02 ix3121 (.Y (nx3122), .A (shift2To1)) ;
    buf02 ix3123 (.Y (nx3124), .A (shift1To2)) ;
    buf02 ix3125 (.Y (nx3126), .A (shift1To2)) ;
endmodule


module RegRow_8_16_5_3 ( filterBus, windowBus, page1NextRow_0__15, 
                         page1NextRow_0__14, page1NextRow_0__13, 
                         page1NextRow_0__12, page1NextRow_0__11, 
                         page1NextRow_0__10, page1NextRow_0__9, 
                         page1NextRow_0__8, page1NextRow_0__7, page1NextRow_0__6, 
                         page1NextRow_0__5, page1NextRow_0__4, page1NextRow_0__3, 
                         page1NextRow_0__2, page1NextRow_0__1, page1NextRow_0__0, 
                         page1NextRow_1__15, page1NextRow_1__14, 
                         page1NextRow_1__13, page1NextRow_1__12, 
                         page1NextRow_1__11, page1NextRow_1__10, 
                         page1NextRow_1__9, page1NextRow_1__8, page1NextRow_1__7, 
                         page1NextRow_1__6, page1NextRow_1__5, page1NextRow_1__4, 
                         page1NextRow_1__3, page1NextRow_1__2, page1NextRow_1__1, 
                         page1NextRow_1__0, page1NextRow_2__15, 
                         page1NextRow_2__14, page1NextRow_2__13, 
                         page1NextRow_2__12, page1NextRow_2__11, 
                         page1NextRow_2__10, page1NextRow_2__9, 
                         page1NextRow_2__8, page1NextRow_2__7, page1NextRow_2__6, 
                         page1NextRow_2__5, page1NextRow_2__4, page1NextRow_2__3, 
                         page1NextRow_2__2, page1NextRow_2__1, page1NextRow_2__0, 
                         page1NextRow_3__15, page1NextRow_3__14, 
                         page1NextRow_3__13, page1NextRow_3__12, 
                         page1NextRow_3__11, page1NextRow_3__10, 
                         page1NextRow_3__9, page1NextRow_3__8, page1NextRow_3__7, 
                         page1NextRow_3__6, page1NextRow_3__5, page1NextRow_3__4, 
                         page1NextRow_3__3, page1NextRow_3__2, page1NextRow_3__1, 
                         page1NextRow_3__0, page1NextRow_4__15, 
                         page1NextRow_4__14, page1NextRow_4__13, 
                         page1NextRow_4__12, page1NextRow_4__11, 
                         page1NextRow_4__10, page1NextRow_4__9, 
                         page1NextRow_4__8, page1NextRow_4__7, page1NextRow_4__6, 
                         page1NextRow_4__5, page1NextRow_4__4, page1NextRow_4__3, 
                         page1NextRow_4__2, page1NextRow_4__1, page1NextRow_4__0, 
                         page2NextRow_0__15, page2NextRow_0__14, 
                         page2NextRow_0__13, page2NextRow_0__12, 
                         page2NextRow_0__11, page2NextRow_0__10, 
                         page2NextRow_0__9, page2NextRow_0__8, page2NextRow_0__7, 
                         page2NextRow_0__6, page2NextRow_0__5, page2NextRow_0__4, 
                         page2NextRow_0__3, page2NextRow_0__2, page2NextRow_0__1, 
                         page2NextRow_0__0, page2NextRow_1__15, 
                         page2NextRow_1__14, page2NextRow_1__13, 
                         page2NextRow_1__12, page2NextRow_1__11, 
                         page2NextRow_1__10, page2NextRow_1__9, 
                         page2NextRow_1__8, page2NextRow_1__7, page2NextRow_1__6, 
                         page2NextRow_1__5, page2NextRow_1__4, page2NextRow_1__3, 
                         page2NextRow_1__2, page2NextRow_1__1, page2NextRow_1__0, 
                         page2NextRow_2__15, page2NextRow_2__14, 
                         page2NextRow_2__13, page2NextRow_2__12, 
                         page2NextRow_2__11, page2NextRow_2__10, 
                         page2NextRow_2__9, page2NextRow_2__8, page2NextRow_2__7, 
                         page2NextRow_2__6, page2NextRow_2__5, page2NextRow_2__4, 
                         page2NextRow_2__3, page2NextRow_2__2, page2NextRow_2__1, 
                         page2NextRow_2__0, page2NextRow_3__15, 
                         page2NextRow_3__14, page2NextRow_3__13, 
                         page2NextRow_3__12, page2NextRow_3__11, 
                         page2NextRow_3__10, page2NextRow_3__9, 
                         page2NextRow_3__8, page2NextRow_3__7, page2NextRow_3__6, 
                         page2NextRow_3__5, page2NextRow_3__4, page2NextRow_3__3, 
                         page2NextRow_3__2, page2NextRow_3__1, page2NextRow_3__0, 
                         page2NextRow_4__15, page2NextRow_4__14, 
                         page2NextRow_4__13, page2NextRow_4__12, 
                         page2NextRow_4__11, page2NextRow_4__10, 
                         page2NextRow_4__9, page2NextRow_4__8, page2NextRow_4__7, 
                         page2NextRow_4__6, page2NextRow_4__5, page2NextRow_4__4, 
                         page2NextRow_4__3, page2NextRow_4__2, page2NextRow_4__1, 
                         page2NextRow_4__0, clk, rst, enablePage1Read, 
                         enablePage2Read, enableFilterRead, shift2To1, shift1To2, 
                         pageTurn, page1Out_0__15, page1Out_0__14, 
                         page1Out_0__13, page1Out_0__12, page1Out_0__11, 
                         page1Out_0__10, page1Out_0__9, page1Out_0__8, 
                         page1Out_0__7, page1Out_0__6, page1Out_0__5, 
                         page1Out_0__4, page1Out_0__3, page1Out_0__2, 
                         page1Out_0__1, page1Out_0__0, page1Out_1__15, 
                         page1Out_1__14, page1Out_1__13, page1Out_1__12, 
                         page1Out_1__11, page1Out_1__10, page1Out_1__9, 
                         page1Out_1__8, page1Out_1__7, page1Out_1__6, 
                         page1Out_1__5, page1Out_1__4, page1Out_1__3, 
                         page1Out_1__2, page1Out_1__1, page1Out_1__0, 
                         page1Out_2__15, page1Out_2__14, page1Out_2__13, 
                         page1Out_2__12, page1Out_2__11, page1Out_2__10, 
                         page1Out_2__9, page1Out_2__8, page1Out_2__7, 
                         page1Out_2__6, page1Out_2__5, page1Out_2__4, 
                         page1Out_2__3, page1Out_2__2, page1Out_2__1, 
                         page1Out_2__0, page1Out_3__15, page1Out_3__14, 
                         page1Out_3__13, page1Out_3__12, page1Out_3__11, 
                         page1Out_3__10, page1Out_3__9, page1Out_3__8, 
                         page1Out_3__7, page1Out_3__6, page1Out_3__5, 
                         page1Out_3__4, page1Out_3__3, page1Out_3__2, 
                         page1Out_3__1, page1Out_3__0, page1Out_4__15, 
                         page1Out_4__14, page1Out_4__13, page1Out_4__12, 
                         page1Out_4__11, page1Out_4__10, page1Out_4__9, 
                         page1Out_4__8, page1Out_4__7, page1Out_4__6, 
                         page1Out_4__5, page1Out_4__4, page1Out_4__3, 
                         page1Out_4__2, page1Out_4__1, page1Out_4__0, 
                         page2Out_0__15, page2Out_0__14, page2Out_0__13, 
                         page2Out_0__12, page2Out_0__11, page2Out_0__10, 
                         page2Out_0__9, page2Out_0__8, page2Out_0__7, 
                         page2Out_0__6, page2Out_0__5, page2Out_0__4, 
                         page2Out_0__3, page2Out_0__2, page2Out_0__1, 
                         page2Out_0__0, page2Out_1__15, page2Out_1__14, 
                         page2Out_1__13, page2Out_1__12, page2Out_1__11, 
                         page2Out_1__10, page2Out_1__9, page2Out_1__8, 
                         page2Out_1__7, page2Out_1__6, page2Out_1__5, 
                         page2Out_1__4, page2Out_1__3, page2Out_1__2, 
                         page2Out_1__1, page2Out_1__0, page2Out_2__15, 
                         page2Out_2__14, page2Out_2__13, page2Out_2__12, 
                         page2Out_2__11, page2Out_2__10, page2Out_2__9, 
                         page2Out_2__8, page2Out_2__7, page2Out_2__6, 
                         page2Out_2__5, page2Out_2__4, page2Out_2__3, 
                         page2Out_2__2, page2Out_2__1, page2Out_2__0, 
                         page2Out_3__15, page2Out_3__14, page2Out_3__13, 
                         page2Out_3__12, page2Out_3__11, page2Out_3__10, 
                         page2Out_3__9, page2Out_3__8, page2Out_3__7, 
                         page2Out_3__6, page2Out_3__5, page2Out_3__4, 
                         page2Out_3__3, page2Out_3__2, page2Out_3__1, 
                         page2Out_3__0, page2Out_4__15, page2Out_4__14, 
                         page2Out_4__13, page2Out_4__12, page2Out_4__11, 
                         page2Out_4__10, page2Out_4__9, page2Out_4__8, 
                         page2Out_4__7, page2Out_4__6, page2Out_4__5, 
                         page2Out_4__4, page2Out_4__3, page2Out_4__2, 
                         page2Out_4__1, page2Out_4__0, pagesOutsPrimary_0__15, 
                         pagesOutsPrimary_0__14, pagesOutsPrimary_0__13, 
                         pagesOutsPrimary_0__12, pagesOutsPrimary_0__11, 
                         pagesOutsPrimary_0__10, pagesOutsPrimary_0__9, 
                         pagesOutsPrimary_0__8, pagesOutsPrimary_0__7, 
                         pagesOutsPrimary_0__6, pagesOutsPrimary_0__5, 
                         pagesOutsPrimary_0__4, pagesOutsPrimary_0__3, 
                         pagesOutsPrimary_0__2, pagesOutsPrimary_0__1, 
                         pagesOutsPrimary_0__0, pagesOutsPrimary_1__15, 
                         pagesOutsPrimary_1__14, pagesOutsPrimary_1__13, 
                         pagesOutsPrimary_1__12, pagesOutsPrimary_1__11, 
                         pagesOutsPrimary_1__10, pagesOutsPrimary_1__9, 
                         pagesOutsPrimary_1__8, pagesOutsPrimary_1__7, 
                         pagesOutsPrimary_1__6, pagesOutsPrimary_1__5, 
                         pagesOutsPrimary_1__4, pagesOutsPrimary_1__3, 
                         pagesOutsPrimary_1__2, pagesOutsPrimary_1__1, 
                         pagesOutsPrimary_1__0, pagesOutsPrimary_2__15, 
                         pagesOutsPrimary_2__14, pagesOutsPrimary_2__13, 
                         pagesOutsPrimary_2__12, pagesOutsPrimary_2__11, 
                         pagesOutsPrimary_2__10, pagesOutsPrimary_2__9, 
                         pagesOutsPrimary_2__8, pagesOutsPrimary_2__7, 
                         pagesOutsPrimary_2__6, pagesOutsPrimary_2__5, 
                         pagesOutsPrimary_2__4, pagesOutsPrimary_2__3, 
                         pagesOutsPrimary_2__2, pagesOutsPrimary_2__1, 
                         pagesOutsPrimary_2__0, pagesOutsSecondary_0__15, 
                         pagesOutsSecondary_0__14, pagesOutsSecondary_0__13, 
                         pagesOutsSecondary_0__12, pagesOutsSecondary_0__11, 
                         pagesOutsSecondary_0__10, pagesOutsSecondary_0__9, 
                         pagesOutsSecondary_0__8, pagesOutsSecondary_0__7, 
                         pagesOutsSecondary_0__6, pagesOutsSecondary_0__5, 
                         pagesOutsSecondary_0__4, pagesOutsSecondary_0__3, 
                         pagesOutsSecondary_0__2, pagesOutsSecondary_0__1, 
                         pagesOutsSecondary_0__0, pagesOutsSecondary_1__15, 
                         pagesOutsSecondary_1__14, pagesOutsSecondary_1__13, 
                         pagesOutsSecondary_1__12, pagesOutsSecondary_1__11, 
                         pagesOutsSecondary_1__10, pagesOutsSecondary_1__9, 
                         pagesOutsSecondary_1__8, pagesOutsSecondary_1__7, 
                         pagesOutsSecondary_1__6, pagesOutsSecondary_1__5, 
                         pagesOutsSecondary_1__4, pagesOutsSecondary_1__3, 
                         pagesOutsSecondary_1__2, pagesOutsSecondary_1__1, 
                         pagesOutsSecondary_1__0, filtersOutsPrimary_0__7, 
                         filtersOutsPrimary_0__6, filtersOutsPrimary_0__5, 
                         filtersOutsPrimary_0__4, filtersOutsPrimary_0__3, 
                         filtersOutsPrimary_0__2, filtersOutsPrimary_0__1, 
                         filtersOutsPrimary_0__0, filtersOutsPrimary_1__7, 
                         filtersOutsPrimary_1__6, filtersOutsPrimary_1__5, 
                         filtersOutsPrimary_1__4, filtersOutsPrimary_1__3, 
                         filtersOutsPrimary_1__2, filtersOutsPrimary_1__1, 
                         filtersOutsPrimary_1__0, filtersOutsPrimary_2__7, 
                         filtersOutsPrimary_2__6, filtersOutsPrimary_2__5, 
                         filtersOutsPrimary_2__4, filtersOutsPrimary_2__3, 
                         filtersOutsPrimary_2__2, filtersOutsPrimary_2__1, 
                         filtersOutsPrimary_2__0, filtersOutsSecondary_0__7, 
                         filtersOutsSecondary_0__6, filtersOutsSecondary_0__5, 
                         filtersOutsSecondary_0__4, filtersOutsSecondary_0__3, 
                         filtersOutsSecondary_0__2, filtersOutsSecondary_0__1, 
                         filtersOutsSecondary_0__0, filtersOutsSecondary_1__7, 
                         filtersOutsSecondary_1__6, filtersOutsSecondary_1__5, 
                         filtersOutsSecondary_1__4, filtersOutsSecondary_1__3, 
                         filtersOutsSecondary_1__2, filtersOutsSecondary_1__1, 
                         filtersOutsSecondary_1__0 ) ;

    input [39:0]filterBus ;
    input [79:0]windowBus ;
    input page1NextRow_0__15 ;
    input page1NextRow_0__14 ;
    input page1NextRow_0__13 ;
    input page1NextRow_0__12 ;
    input page1NextRow_0__11 ;
    input page1NextRow_0__10 ;
    input page1NextRow_0__9 ;
    input page1NextRow_0__8 ;
    input page1NextRow_0__7 ;
    input page1NextRow_0__6 ;
    input page1NextRow_0__5 ;
    input page1NextRow_0__4 ;
    input page1NextRow_0__3 ;
    input page1NextRow_0__2 ;
    input page1NextRow_0__1 ;
    input page1NextRow_0__0 ;
    input page1NextRow_1__15 ;
    input page1NextRow_1__14 ;
    input page1NextRow_1__13 ;
    input page1NextRow_1__12 ;
    input page1NextRow_1__11 ;
    input page1NextRow_1__10 ;
    input page1NextRow_1__9 ;
    input page1NextRow_1__8 ;
    input page1NextRow_1__7 ;
    input page1NextRow_1__6 ;
    input page1NextRow_1__5 ;
    input page1NextRow_1__4 ;
    input page1NextRow_1__3 ;
    input page1NextRow_1__2 ;
    input page1NextRow_1__1 ;
    input page1NextRow_1__0 ;
    input page1NextRow_2__15 ;
    input page1NextRow_2__14 ;
    input page1NextRow_2__13 ;
    input page1NextRow_2__12 ;
    input page1NextRow_2__11 ;
    input page1NextRow_2__10 ;
    input page1NextRow_2__9 ;
    input page1NextRow_2__8 ;
    input page1NextRow_2__7 ;
    input page1NextRow_2__6 ;
    input page1NextRow_2__5 ;
    input page1NextRow_2__4 ;
    input page1NextRow_2__3 ;
    input page1NextRow_2__2 ;
    input page1NextRow_2__1 ;
    input page1NextRow_2__0 ;
    input page1NextRow_3__15 ;
    input page1NextRow_3__14 ;
    input page1NextRow_3__13 ;
    input page1NextRow_3__12 ;
    input page1NextRow_3__11 ;
    input page1NextRow_3__10 ;
    input page1NextRow_3__9 ;
    input page1NextRow_3__8 ;
    input page1NextRow_3__7 ;
    input page1NextRow_3__6 ;
    input page1NextRow_3__5 ;
    input page1NextRow_3__4 ;
    input page1NextRow_3__3 ;
    input page1NextRow_3__2 ;
    input page1NextRow_3__1 ;
    input page1NextRow_3__0 ;
    input page1NextRow_4__15 ;
    input page1NextRow_4__14 ;
    input page1NextRow_4__13 ;
    input page1NextRow_4__12 ;
    input page1NextRow_4__11 ;
    input page1NextRow_4__10 ;
    input page1NextRow_4__9 ;
    input page1NextRow_4__8 ;
    input page1NextRow_4__7 ;
    input page1NextRow_4__6 ;
    input page1NextRow_4__5 ;
    input page1NextRow_4__4 ;
    input page1NextRow_4__3 ;
    input page1NextRow_4__2 ;
    input page1NextRow_4__1 ;
    input page1NextRow_4__0 ;
    input page2NextRow_0__15 ;
    input page2NextRow_0__14 ;
    input page2NextRow_0__13 ;
    input page2NextRow_0__12 ;
    input page2NextRow_0__11 ;
    input page2NextRow_0__10 ;
    input page2NextRow_0__9 ;
    input page2NextRow_0__8 ;
    input page2NextRow_0__7 ;
    input page2NextRow_0__6 ;
    input page2NextRow_0__5 ;
    input page2NextRow_0__4 ;
    input page2NextRow_0__3 ;
    input page2NextRow_0__2 ;
    input page2NextRow_0__1 ;
    input page2NextRow_0__0 ;
    input page2NextRow_1__15 ;
    input page2NextRow_1__14 ;
    input page2NextRow_1__13 ;
    input page2NextRow_1__12 ;
    input page2NextRow_1__11 ;
    input page2NextRow_1__10 ;
    input page2NextRow_1__9 ;
    input page2NextRow_1__8 ;
    input page2NextRow_1__7 ;
    input page2NextRow_1__6 ;
    input page2NextRow_1__5 ;
    input page2NextRow_1__4 ;
    input page2NextRow_1__3 ;
    input page2NextRow_1__2 ;
    input page2NextRow_1__1 ;
    input page2NextRow_1__0 ;
    input page2NextRow_2__15 ;
    input page2NextRow_2__14 ;
    input page2NextRow_2__13 ;
    input page2NextRow_2__12 ;
    input page2NextRow_2__11 ;
    input page2NextRow_2__10 ;
    input page2NextRow_2__9 ;
    input page2NextRow_2__8 ;
    input page2NextRow_2__7 ;
    input page2NextRow_2__6 ;
    input page2NextRow_2__5 ;
    input page2NextRow_2__4 ;
    input page2NextRow_2__3 ;
    input page2NextRow_2__2 ;
    input page2NextRow_2__1 ;
    input page2NextRow_2__0 ;
    input page2NextRow_3__15 ;
    input page2NextRow_3__14 ;
    input page2NextRow_3__13 ;
    input page2NextRow_3__12 ;
    input page2NextRow_3__11 ;
    input page2NextRow_3__10 ;
    input page2NextRow_3__9 ;
    input page2NextRow_3__8 ;
    input page2NextRow_3__7 ;
    input page2NextRow_3__6 ;
    input page2NextRow_3__5 ;
    input page2NextRow_3__4 ;
    input page2NextRow_3__3 ;
    input page2NextRow_3__2 ;
    input page2NextRow_3__1 ;
    input page2NextRow_3__0 ;
    input page2NextRow_4__15 ;
    input page2NextRow_4__14 ;
    input page2NextRow_4__13 ;
    input page2NextRow_4__12 ;
    input page2NextRow_4__11 ;
    input page2NextRow_4__10 ;
    input page2NextRow_4__9 ;
    input page2NextRow_4__8 ;
    input page2NextRow_4__7 ;
    input page2NextRow_4__6 ;
    input page2NextRow_4__5 ;
    input page2NextRow_4__4 ;
    input page2NextRow_4__3 ;
    input page2NextRow_4__2 ;
    input page2NextRow_4__1 ;
    input page2NextRow_4__0 ;
    input clk ;
    input rst ;
    input enablePage1Read ;
    input enablePage2Read ;
    input enableFilterRead ;
    input shift2To1 ;
    input shift1To2 ;
    input pageTurn ;
    output page1Out_0__15 ;
    output page1Out_0__14 ;
    output page1Out_0__13 ;
    output page1Out_0__12 ;
    output page1Out_0__11 ;
    output page1Out_0__10 ;
    output page1Out_0__9 ;
    output page1Out_0__8 ;
    output page1Out_0__7 ;
    output page1Out_0__6 ;
    output page1Out_0__5 ;
    output page1Out_0__4 ;
    output page1Out_0__3 ;
    output page1Out_0__2 ;
    output page1Out_0__1 ;
    output page1Out_0__0 ;
    output page1Out_1__15 ;
    output page1Out_1__14 ;
    output page1Out_1__13 ;
    output page1Out_1__12 ;
    output page1Out_1__11 ;
    output page1Out_1__10 ;
    output page1Out_1__9 ;
    output page1Out_1__8 ;
    output page1Out_1__7 ;
    output page1Out_1__6 ;
    output page1Out_1__5 ;
    output page1Out_1__4 ;
    output page1Out_1__3 ;
    output page1Out_1__2 ;
    output page1Out_1__1 ;
    output page1Out_1__0 ;
    output page1Out_2__15 ;
    output page1Out_2__14 ;
    output page1Out_2__13 ;
    output page1Out_2__12 ;
    output page1Out_2__11 ;
    output page1Out_2__10 ;
    output page1Out_2__9 ;
    output page1Out_2__8 ;
    output page1Out_2__7 ;
    output page1Out_2__6 ;
    output page1Out_2__5 ;
    output page1Out_2__4 ;
    output page1Out_2__3 ;
    output page1Out_2__2 ;
    output page1Out_2__1 ;
    output page1Out_2__0 ;
    output page1Out_3__15 ;
    output page1Out_3__14 ;
    output page1Out_3__13 ;
    output page1Out_3__12 ;
    output page1Out_3__11 ;
    output page1Out_3__10 ;
    output page1Out_3__9 ;
    output page1Out_3__8 ;
    output page1Out_3__7 ;
    output page1Out_3__6 ;
    output page1Out_3__5 ;
    output page1Out_3__4 ;
    output page1Out_3__3 ;
    output page1Out_3__2 ;
    output page1Out_3__1 ;
    output page1Out_3__0 ;
    output page1Out_4__15 ;
    output page1Out_4__14 ;
    output page1Out_4__13 ;
    output page1Out_4__12 ;
    output page1Out_4__11 ;
    output page1Out_4__10 ;
    output page1Out_4__9 ;
    output page1Out_4__8 ;
    output page1Out_4__7 ;
    output page1Out_4__6 ;
    output page1Out_4__5 ;
    output page1Out_4__4 ;
    output page1Out_4__3 ;
    output page1Out_4__2 ;
    output page1Out_4__1 ;
    output page1Out_4__0 ;
    output page2Out_0__15 ;
    output page2Out_0__14 ;
    output page2Out_0__13 ;
    output page2Out_0__12 ;
    output page2Out_0__11 ;
    output page2Out_0__10 ;
    output page2Out_0__9 ;
    output page2Out_0__8 ;
    output page2Out_0__7 ;
    output page2Out_0__6 ;
    output page2Out_0__5 ;
    output page2Out_0__4 ;
    output page2Out_0__3 ;
    output page2Out_0__2 ;
    output page2Out_0__1 ;
    output page2Out_0__0 ;
    output page2Out_1__15 ;
    output page2Out_1__14 ;
    output page2Out_1__13 ;
    output page2Out_1__12 ;
    output page2Out_1__11 ;
    output page2Out_1__10 ;
    output page2Out_1__9 ;
    output page2Out_1__8 ;
    output page2Out_1__7 ;
    output page2Out_1__6 ;
    output page2Out_1__5 ;
    output page2Out_1__4 ;
    output page2Out_1__3 ;
    output page2Out_1__2 ;
    output page2Out_1__1 ;
    output page2Out_1__0 ;
    output page2Out_2__15 ;
    output page2Out_2__14 ;
    output page2Out_2__13 ;
    output page2Out_2__12 ;
    output page2Out_2__11 ;
    output page2Out_2__10 ;
    output page2Out_2__9 ;
    output page2Out_2__8 ;
    output page2Out_2__7 ;
    output page2Out_2__6 ;
    output page2Out_2__5 ;
    output page2Out_2__4 ;
    output page2Out_2__3 ;
    output page2Out_2__2 ;
    output page2Out_2__1 ;
    output page2Out_2__0 ;
    output page2Out_3__15 ;
    output page2Out_3__14 ;
    output page2Out_3__13 ;
    output page2Out_3__12 ;
    output page2Out_3__11 ;
    output page2Out_3__10 ;
    output page2Out_3__9 ;
    output page2Out_3__8 ;
    output page2Out_3__7 ;
    output page2Out_3__6 ;
    output page2Out_3__5 ;
    output page2Out_3__4 ;
    output page2Out_3__3 ;
    output page2Out_3__2 ;
    output page2Out_3__1 ;
    output page2Out_3__0 ;
    output page2Out_4__15 ;
    output page2Out_4__14 ;
    output page2Out_4__13 ;
    output page2Out_4__12 ;
    output page2Out_4__11 ;
    output page2Out_4__10 ;
    output page2Out_4__9 ;
    output page2Out_4__8 ;
    output page2Out_4__7 ;
    output page2Out_4__6 ;
    output page2Out_4__5 ;
    output page2Out_4__4 ;
    output page2Out_4__3 ;
    output page2Out_4__2 ;
    output page2Out_4__1 ;
    output page2Out_4__0 ;
    output pagesOutsPrimary_0__15 ;
    output pagesOutsPrimary_0__14 ;
    output pagesOutsPrimary_0__13 ;
    output pagesOutsPrimary_0__12 ;
    output pagesOutsPrimary_0__11 ;
    output pagesOutsPrimary_0__10 ;
    output pagesOutsPrimary_0__9 ;
    output pagesOutsPrimary_0__8 ;
    output pagesOutsPrimary_0__7 ;
    output pagesOutsPrimary_0__6 ;
    output pagesOutsPrimary_0__5 ;
    output pagesOutsPrimary_0__4 ;
    output pagesOutsPrimary_0__3 ;
    output pagesOutsPrimary_0__2 ;
    output pagesOutsPrimary_0__1 ;
    output pagesOutsPrimary_0__0 ;
    output pagesOutsPrimary_1__15 ;
    output pagesOutsPrimary_1__14 ;
    output pagesOutsPrimary_1__13 ;
    output pagesOutsPrimary_1__12 ;
    output pagesOutsPrimary_1__11 ;
    output pagesOutsPrimary_1__10 ;
    output pagesOutsPrimary_1__9 ;
    output pagesOutsPrimary_1__8 ;
    output pagesOutsPrimary_1__7 ;
    output pagesOutsPrimary_1__6 ;
    output pagesOutsPrimary_1__5 ;
    output pagesOutsPrimary_1__4 ;
    output pagesOutsPrimary_1__3 ;
    output pagesOutsPrimary_1__2 ;
    output pagesOutsPrimary_1__1 ;
    output pagesOutsPrimary_1__0 ;
    output pagesOutsPrimary_2__15 ;
    output pagesOutsPrimary_2__14 ;
    output pagesOutsPrimary_2__13 ;
    output pagesOutsPrimary_2__12 ;
    output pagesOutsPrimary_2__11 ;
    output pagesOutsPrimary_2__10 ;
    output pagesOutsPrimary_2__9 ;
    output pagesOutsPrimary_2__8 ;
    output pagesOutsPrimary_2__7 ;
    output pagesOutsPrimary_2__6 ;
    output pagesOutsPrimary_2__5 ;
    output pagesOutsPrimary_2__4 ;
    output pagesOutsPrimary_2__3 ;
    output pagesOutsPrimary_2__2 ;
    output pagesOutsPrimary_2__1 ;
    output pagesOutsPrimary_2__0 ;
    output pagesOutsSecondary_0__15 ;
    output pagesOutsSecondary_0__14 ;
    output pagesOutsSecondary_0__13 ;
    output pagesOutsSecondary_0__12 ;
    output pagesOutsSecondary_0__11 ;
    output pagesOutsSecondary_0__10 ;
    output pagesOutsSecondary_0__9 ;
    output pagesOutsSecondary_0__8 ;
    output pagesOutsSecondary_0__7 ;
    output pagesOutsSecondary_0__6 ;
    output pagesOutsSecondary_0__5 ;
    output pagesOutsSecondary_0__4 ;
    output pagesOutsSecondary_0__3 ;
    output pagesOutsSecondary_0__2 ;
    output pagesOutsSecondary_0__1 ;
    output pagesOutsSecondary_0__0 ;
    output pagesOutsSecondary_1__15 ;
    output pagesOutsSecondary_1__14 ;
    output pagesOutsSecondary_1__13 ;
    output pagesOutsSecondary_1__12 ;
    output pagesOutsSecondary_1__11 ;
    output pagesOutsSecondary_1__10 ;
    output pagesOutsSecondary_1__9 ;
    output pagesOutsSecondary_1__8 ;
    output pagesOutsSecondary_1__7 ;
    output pagesOutsSecondary_1__6 ;
    output pagesOutsSecondary_1__5 ;
    output pagesOutsSecondary_1__4 ;
    output pagesOutsSecondary_1__3 ;
    output pagesOutsSecondary_1__2 ;
    output pagesOutsSecondary_1__1 ;
    output pagesOutsSecondary_1__0 ;
    output filtersOutsPrimary_0__7 ;
    output filtersOutsPrimary_0__6 ;
    output filtersOutsPrimary_0__5 ;
    output filtersOutsPrimary_0__4 ;
    output filtersOutsPrimary_0__3 ;
    output filtersOutsPrimary_0__2 ;
    output filtersOutsPrimary_0__1 ;
    output filtersOutsPrimary_0__0 ;
    output filtersOutsPrimary_1__7 ;
    output filtersOutsPrimary_1__6 ;
    output filtersOutsPrimary_1__5 ;
    output filtersOutsPrimary_1__4 ;
    output filtersOutsPrimary_1__3 ;
    output filtersOutsPrimary_1__2 ;
    output filtersOutsPrimary_1__1 ;
    output filtersOutsPrimary_1__0 ;
    output filtersOutsPrimary_2__7 ;
    output filtersOutsPrimary_2__6 ;
    output filtersOutsPrimary_2__5 ;
    output filtersOutsPrimary_2__4 ;
    output filtersOutsPrimary_2__3 ;
    output filtersOutsPrimary_2__2 ;
    output filtersOutsPrimary_2__1 ;
    output filtersOutsPrimary_2__0 ;
    output filtersOutsSecondary_0__7 ;
    output filtersOutsSecondary_0__6 ;
    output filtersOutsSecondary_0__5 ;
    output filtersOutsSecondary_0__4 ;
    output filtersOutsSecondary_0__3 ;
    output filtersOutsSecondary_0__2 ;
    output filtersOutsSecondary_0__1 ;
    output filtersOutsSecondary_0__0 ;
    output filtersOutsSecondary_1__7 ;
    output filtersOutsSecondary_1__6 ;
    output filtersOutsSecondary_1__5 ;
    output filtersOutsSecondary_1__4 ;
    output filtersOutsSecondary_1__3 ;
    output filtersOutsSecondary_1__2 ;
    output filtersOutsSecondary_1__1 ;
    output filtersOutsSecondary_1__0 ;

    wire nx559, nx561, nx563, nx565, nx567, nx569;



    RegUnit_8_16 loop1_0_regUnitMap (.filterBus ({filterBus[7],filterBus[6],
                 filterBus[5],filterBus[4],filterBus[3],filterBus[2],
                 filterBus[1],filterBus[0]}), .windowBus ({windowBus[15],
                 windowBus[14],windowBus[13],windowBus[12],windowBus[11],
                 windowBus[10],windowBus[9],windowBus[8],windowBus[7],
                 windowBus[6],windowBus[5],windowBus[4],windowBus[3],
                 windowBus[2],windowBus[1],windowBus[0]}), .regPage1NextUnit ({
                 page1NextRow_0__15,page1NextRow_0__14,page1NextRow_0__13,
                 page1NextRow_0__12,page1NextRow_0__11,page1NextRow_0__10,
                 page1NextRow_0__9,page1NextRow_0__8,page1NextRow_0__7,
                 page1NextRow_0__6,page1NextRow_0__5,page1NextRow_0__4,
                 page1NextRow_0__3,page1NextRow_0__2,page1NextRow_0__1,
                 page1NextRow_0__0}), .regPage2NextUnit ({page2NextRow_0__15,
                 page2NextRow_0__14,page2NextRow_0__13,page2NextRow_0__12,
                 page2NextRow_0__11,page2NextRow_0__10,page2NextRow_0__9,
                 page2NextRow_0__8,page2NextRow_0__7,page2NextRow_0__6,
                 page2NextRow_0__5,page2NextRow_0__4,page2NextRow_0__3,
                 page2NextRow_0__2,page2NextRow_0__1,page2NextRow_0__0}), .clk (
                 clk), .rst (rst), .enableRegPage1 (enablePage1Read), .enableRegPage2 (
                 enablePage2Read), .enableRegFilter (nx559), .page1ReadBusOrPage2 (
                 nx563), .page2ReadBusOrPage1 (nx567), .pageTurn (pageTurn), .outRegPage (
                 {pagesOutsPrimary_0__15,pagesOutsPrimary_0__14,
                 pagesOutsPrimary_0__13,pagesOutsPrimary_0__12,
                 pagesOutsPrimary_0__11,pagesOutsPrimary_0__10,
                 pagesOutsPrimary_0__9,pagesOutsPrimary_0__8,
                 pagesOutsPrimary_0__7,pagesOutsPrimary_0__6,
                 pagesOutsPrimary_0__5,pagesOutsPrimary_0__4,
                 pagesOutsPrimary_0__3,pagesOutsPrimary_0__2,
                 pagesOutsPrimary_0__1,pagesOutsPrimary_0__0}), .outputRegPage1 (
                 {page1Out_0__15,page1Out_0__14,page1Out_0__13,page1Out_0__12,
                 page1Out_0__11,page1Out_0__10,page1Out_0__9,page1Out_0__8,
                 page1Out_0__7,page1Out_0__6,page1Out_0__5,page1Out_0__4,
                 page1Out_0__3,page1Out_0__2,page1Out_0__1,page1Out_0__0}), .outputRegPage2 (
                 {page2Out_0__15,page2Out_0__14,page2Out_0__13,page2Out_0__12,
                 page2Out_0__11,page2Out_0__10,page2Out_0__9,page2Out_0__8,
                 page2Out_0__7,page2Out_0__6,page2Out_0__5,page2Out_0__4,
                 page2Out_0__3,page2Out_0__2,page2Out_0__1,page2Out_0__0}), .outFilter (
                 {filtersOutsPrimary_0__7,filtersOutsPrimary_0__6,
                 filtersOutsPrimary_0__5,filtersOutsPrimary_0__4,
                 filtersOutsPrimary_0__3,filtersOutsPrimary_0__2,
                 filtersOutsPrimary_0__1,filtersOutsPrimary_0__0})) ;
    RegUnit_8_16 loop1_1_regUnitMap (.filterBus ({filterBus[15],filterBus[14],
                 filterBus[13],filterBus[12],filterBus[11],filterBus[10],
                 filterBus[9],filterBus[8]}), .windowBus ({windowBus[31],
                 windowBus[30],windowBus[29],windowBus[28],windowBus[27],
                 windowBus[26],windowBus[25],windowBus[24],windowBus[23],
                 windowBus[22],windowBus[21],windowBus[20],windowBus[19],
                 windowBus[18],windowBus[17],windowBus[16]}), .regPage1NextUnit (
                 {page1NextRow_1__15,page1NextRow_1__14,page1NextRow_1__13,
                 page1NextRow_1__12,page1NextRow_1__11,page1NextRow_1__10,
                 page1NextRow_1__9,page1NextRow_1__8,page1NextRow_1__7,
                 page1NextRow_1__6,page1NextRow_1__5,page1NextRow_1__4,
                 page1NextRow_1__3,page1NextRow_1__2,page1NextRow_1__1,
                 page1NextRow_1__0}), .regPage2NextUnit ({page2NextRow_1__15,
                 page2NextRow_1__14,page2NextRow_1__13,page2NextRow_1__12,
                 page2NextRow_1__11,page2NextRow_1__10,page2NextRow_1__9,
                 page2NextRow_1__8,page2NextRow_1__7,page2NextRow_1__6,
                 page2NextRow_1__5,page2NextRow_1__4,page2NextRow_1__3,
                 page2NextRow_1__2,page2NextRow_1__1,page2NextRow_1__0}), .clk (
                 clk), .rst (rst), .enableRegPage1 (enablePage1Read), .enableRegPage2 (
                 enablePage2Read), .enableRegFilter (nx559), .page1ReadBusOrPage2 (
                 nx563), .page2ReadBusOrPage1 (nx567), .pageTurn (pageTurn), .outRegPage (
                 {pagesOutsPrimary_1__15,pagesOutsPrimary_1__14,
                 pagesOutsPrimary_1__13,pagesOutsPrimary_1__12,
                 pagesOutsPrimary_1__11,pagesOutsPrimary_1__10,
                 pagesOutsPrimary_1__9,pagesOutsPrimary_1__8,
                 pagesOutsPrimary_1__7,pagesOutsPrimary_1__6,
                 pagesOutsPrimary_1__5,pagesOutsPrimary_1__4,
                 pagesOutsPrimary_1__3,pagesOutsPrimary_1__2,
                 pagesOutsPrimary_1__1,pagesOutsPrimary_1__0}), .outputRegPage1 (
                 {page1Out_1__15,page1Out_1__14,page1Out_1__13,page1Out_1__12,
                 page1Out_1__11,page1Out_1__10,page1Out_1__9,page1Out_1__8,
                 page1Out_1__7,page1Out_1__6,page1Out_1__5,page1Out_1__4,
                 page1Out_1__3,page1Out_1__2,page1Out_1__1,page1Out_1__0}), .outputRegPage2 (
                 {page2Out_1__15,page2Out_1__14,page2Out_1__13,page2Out_1__12,
                 page2Out_1__11,page2Out_1__10,page2Out_1__9,page2Out_1__8,
                 page2Out_1__7,page2Out_1__6,page2Out_1__5,page2Out_1__4,
                 page2Out_1__3,page2Out_1__2,page2Out_1__1,page2Out_1__0}), .outFilter (
                 {filtersOutsPrimary_1__7,filtersOutsPrimary_1__6,
                 filtersOutsPrimary_1__5,filtersOutsPrimary_1__4,
                 filtersOutsPrimary_1__3,filtersOutsPrimary_1__2,
                 filtersOutsPrimary_1__1,filtersOutsPrimary_1__0})) ;
    RegUnit_8_16 loop1_2_regUnitMap (.filterBus ({filterBus[23],filterBus[22],
                 filterBus[21],filterBus[20],filterBus[19],filterBus[18],
                 filterBus[17],filterBus[16]}), .windowBus ({windowBus[47],
                 windowBus[46],windowBus[45],windowBus[44],windowBus[43],
                 windowBus[42],windowBus[41],windowBus[40],windowBus[39],
                 windowBus[38],windowBus[37],windowBus[36],windowBus[35],
                 windowBus[34],windowBus[33],windowBus[32]}), .regPage1NextUnit (
                 {page1NextRow_2__15,page1NextRow_2__14,page1NextRow_2__13,
                 page1NextRow_2__12,page1NextRow_2__11,page1NextRow_2__10,
                 page1NextRow_2__9,page1NextRow_2__8,page1NextRow_2__7,
                 page1NextRow_2__6,page1NextRow_2__5,page1NextRow_2__4,
                 page1NextRow_2__3,page1NextRow_2__2,page1NextRow_2__1,
                 page1NextRow_2__0}), .regPage2NextUnit ({page2NextRow_2__15,
                 page2NextRow_2__14,page2NextRow_2__13,page2NextRow_2__12,
                 page2NextRow_2__11,page2NextRow_2__10,page2NextRow_2__9,
                 page2NextRow_2__8,page2NextRow_2__7,page2NextRow_2__6,
                 page2NextRow_2__5,page2NextRow_2__4,page2NextRow_2__3,
                 page2NextRow_2__2,page2NextRow_2__1,page2NextRow_2__0}), .clk (
                 clk), .rst (rst), .enableRegPage1 (enablePage1Read), .enableRegPage2 (
                 enablePage2Read), .enableRegFilter (nx559), .page1ReadBusOrPage2 (
                 nx563), .page2ReadBusOrPage1 (nx567), .pageTurn (pageTurn), .outRegPage (
                 {pagesOutsPrimary_2__15,pagesOutsPrimary_2__14,
                 pagesOutsPrimary_2__13,pagesOutsPrimary_2__12,
                 pagesOutsPrimary_2__11,pagesOutsPrimary_2__10,
                 pagesOutsPrimary_2__9,pagesOutsPrimary_2__8,
                 pagesOutsPrimary_2__7,pagesOutsPrimary_2__6,
                 pagesOutsPrimary_2__5,pagesOutsPrimary_2__4,
                 pagesOutsPrimary_2__3,pagesOutsPrimary_2__2,
                 pagesOutsPrimary_2__1,pagesOutsPrimary_2__0}), .outputRegPage1 (
                 {page1Out_2__15,page1Out_2__14,page1Out_2__13,page1Out_2__12,
                 page1Out_2__11,page1Out_2__10,page1Out_2__9,page1Out_2__8,
                 page1Out_2__7,page1Out_2__6,page1Out_2__5,page1Out_2__4,
                 page1Out_2__3,page1Out_2__2,page1Out_2__1,page1Out_2__0}), .outputRegPage2 (
                 {page2Out_2__15,page2Out_2__14,page2Out_2__13,page2Out_2__12,
                 page2Out_2__11,page2Out_2__10,page2Out_2__9,page2Out_2__8,
                 page2Out_2__7,page2Out_2__6,page2Out_2__5,page2Out_2__4,
                 page2Out_2__3,page2Out_2__2,page2Out_2__1,page2Out_2__0}), .outFilter (
                 {filtersOutsPrimary_2__7,filtersOutsPrimary_2__6,
                 filtersOutsPrimary_2__5,filtersOutsPrimary_2__4,
                 filtersOutsPrimary_2__3,filtersOutsPrimary_2__2,
                 filtersOutsPrimary_2__1,filtersOutsPrimary_2__0})) ;
    RegUnit_8_16 loop1_3_regUnitMap (.filterBus ({filterBus[31],filterBus[30],
                 filterBus[29],filterBus[28],filterBus[27],filterBus[26],
                 filterBus[25],filterBus[24]}), .windowBus ({windowBus[63],
                 windowBus[62],windowBus[61],windowBus[60],windowBus[59],
                 windowBus[58],windowBus[57],windowBus[56],windowBus[55],
                 windowBus[54],windowBus[53],windowBus[52],windowBus[51],
                 windowBus[50],windowBus[49],windowBus[48]}), .regPage1NextUnit (
                 {page1NextRow_3__15,page1NextRow_3__14,page1NextRow_3__13,
                 page1NextRow_3__12,page1NextRow_3__11,page1NextRow_3__10,
                 page1NextRow_3__9,page1NextRow_3__8,page1NextRow_3__7,
                 page1NextRow_3__6,page1NextRow_3__5,page1NextRow_3__4,
                 page1NextRow_3__3,page1NextRow_3__2,page1NextRow_3__1,
                 page1NextRow_3__0}), .regPage2NextUnit ({page2NextRow_3__15,
                 page2NextRow_3__14,page2NextRow_3__13,page2NextRow_3__12,
                 page2NextRow_3__11,page2NextRow_3__10,page2NextRow_3__9,
                 page2NextRow_3__8,page2NextRow_3__7,page2NextRow_3__6,
                 page2NextRow_3__5,page2NextRow_3__4,page2NextRow_3__3,
                 page2NextRow_3__2,page2NextRow_3__1,page2NextRow_3__0}), .clk (
                 clk), .rst (rst), .enableRegPage1 (enablePage1Read), .enableRegPage2 (
                 enablePage2Read), .enableRegFilter (nx561), .page1ReadBusOrPage2 (
                 nx565), .page2ReadBusOrPage1 (nx569), .pageTurn (pageTurn), .outRegPage (
                 {pagesOutsSecondary_0__15,pagesOutsSecondary_0__14,
                 pagesOutsSecondary_0__13,pagesOutsSecondary_0__12,
                 pagesOutsSecondary_0__11,pagesOutsSecondary_0__10,
                 pagesOutsSecondary_0__9,pagesOutsSecondary_0__8,
                 pagesOutsSecondary_0__7,pagesOutsSecondary_0__6,
                 pagesOutsSecondary_0__5,pagesOutsSecondary_0__4,
                 pagesOutsSecondary_0__3,pagesOutsSecondary_0__2,
                 pagesOutsSecondary_0__1,pagesOutsSecondary_0__0}), .outputRegPage1 (
                 {page1Out_3__15,page1Out_3__14,page1Out_3__13,page1Out_3__12,
                 page1Out_3__11,page1Out_3__10,page1Out_3__9,page1Out_3__8,
                 page1Out_3__7,page1Out_3__6,page1Out_3__5,page1Out_3__4,
                 page1Out_3__3,page1Out_3__2,page1Out_3__1,page1Out_3__0}), .outputRegPage2 (
                 {page2Out_3__15,page2Out_3__14,page2Out_3__13,page2Out_3__12,
                 page2Out_3__11,page2Out_3__10,page2Out_3__9,page2Out_3__8,
                 page2Out_3__7,page2Out_3__6,page2Out_3__5,page2Out_3__4,
                 page2Out_3__3,page2Out_3__2,page2Out_3__1,page2Out_3__0}), .outFilter (
                 {filtersOutsSecondary_0__7,filtersOutsSecondary_0__6,
                 filtersOutsSecondary_0__5,filtersOutsSecondary_0__4,
                 filtersOutsSecondary_0__3,filtersOutsSecondary_0__2,
                 filtersOutsSecondary_0__1,filtersOutsSecondary_0__0})) ;
    RegUnit_8_16 loop1_4_regUnitMap (.filterBus ({filterBus[39],filterBus[38],
                 filterBus[37],filterBus[36],filterBus[35],filterBus[34],
                 filterBus[33],filterBus[32]}), .windowBus ({windowBus[79],
                 windowBus[78],windowBus[77],windowBus[76],windowBus[75],
                 windowBus[74],windowBus[73],windowBus[72],windowBus[71],
                 windowBus[70],windowBus[69],windowBus[68],windowBus[67],
                 windowBus[66],windowBus[65],windowBus[64]}), .regPage1NextUnit (
                 {page1NextRow_4__15,page1NextRow_4__14,page1NextRow_4__13,
                 page1NextRow_4__12,page1NextRow_4__11,page1NextRow_4__10,
                 page1NextRow_4__9,page1NextRow_4__8,page1NextRow_4__7,
                 page1NextRow_4__6,page1NextRow_4__5,page1NextRow_4__4,
                 page1NextRow_4__3,page1NextRow_4__2,page1NextRow_4__1,
                 page1NextRow_4__0}), .regPage2NextUnit ({page2NextRow_4__15,
                 page2NextRow_4__14,page2NextRow_4__13,page2NextRow_4__12,
                 page2NextRow_4__11,page2NextRow_4__10,page2NextRow_4__9,
                 page2NextRow_4__8,page2NextRow_4__7,page2NextRow_4__6,
                 page2NextRow_4__5,page2NextRow_4__4,page2NextRow_4__3,
                 page2NextRow_4__2,page2NextRow_4__1,page2NextRow_4__0}), .clk (
                 clk), .rst (rst), .enableRegPage1 (enablePage1Read), .enableRegPage2 (
                 enablePage2Read), .enableRegFilter (nx561), .page1ReadBusOrPage2 (
                 nx565), .page2ReadBusOrPage1 (nx569), .pageTurn (pageTurn), .outRegPage (
                 {pagesOutsSecondary_1__15,pagesOutsSecondary_1__14,
                 pagesOutsSecondary_1__13,pagesOutsSecondary_1__12,
                 pagesOutsSecondary_1__11,pagesOutsSecondary_1__10,
                 pagesOutsSecondary_1__9,pagesOutsSecondary_1__8,
                 pagesOutsSecondary_1__7,pagesOutsSecondary_1__6,
                 pagesOutsSecondary_1__5,pagesOutsSecondary_1__4,
                 pagesOutsSecondary_1__3,pagesOutsSecondary_1__2,
                 pagesOutsSecondary_1__1,pagesOutsSecondary_1__0}), .outputRegPage1 (
                 {page1Out_4__15,page1Out_4__14,page1Out_4__13,page1Out_4__12,
                 page1Out_4__11,page1Out_4__10,page1Out_4__9,page1Out_4__8,
                 page1Out_4__7,page1Out_4__6,page1Out_4__5,page1Out_4__4,
                 page1Out_4__3,page1Out_4__2,page1Out_4__1,page1Out_4__0}), .outputRegPage2 (
                 {page2Out_4__15,page2Out_4__14,page2Out_4__13,page2Out_4__12,
                 page2Out_4__11,page2Out_4__10,page2Out_4__9,page2Out_4__8,
                 page2Out_4__7,page2Out_4__6,page2Out_4__5,page2Out_4__4,
                 page2Out_4__3,page2Out_4__2,page2Out_4__1,page2Out_4__0}), .outFilter (
                 {filtersOutsSecondary_1__7,filtersOutsSecondary_1__6,
                 filtersOutsSecondary_1__5,filtersOutsSecondary_1__4,
                 filtersOutsSecondary_1__3,filtersOutsSecondary_1__2,
                 filtersOutsSecondary_1__1,filtersOutsSecondary_1__0})) ;
    buf02 ix558 (.Y (nx559), .A (enableFilterRead)) ;
    buf02 ix560 (.Y (nx561), .A (enableFilterRead)) ;
    buf02 ix562 (.Y (nx563), .A (shift2To1)) ;
    buf02 ix564 (.Y (nx565), .A (shift2To1)) ;
    buf02 ix566 (.Y (nx567), .A (shift1To2)) ;
    buf02 ix568 (.Y (nx569), .A (shift1To2)) ;
endmodule


module RegUnit_8_16 ( filterBus, windowBus, regPage1NextUnit, regPage2NextUnit, 
                      clk, rst, enableRegPage1, enableRegPage2, enableRegFilter, 
                      page1ReadBusOrPage2, page2ReadBusOrPage1, pageTurn, 
                      outRegPage, outputRegPage1, outputRegPage2, outFilter ) ;

    input [7:0]filterBus ;
    input [15:0]windowBus ;
    input [15:0]regPage1NextUnit ;
    input [15:0]regPage2NextUnit ;
    input clk ;
    input rst ;
    input enableRegPage1 ;
    input enableRegPage2 ;
    input enableRegFilter ;
    input page1ReadBusOrPage2 ;
    input page2ReadBusOrPage1 ;
    input pageTurn ;
    output [15:0]outRegPage ;
    output [15:0]outputRegPage1 ;
    output [15:0]outputRegPage2 ;
    output [7:0]outFilter ;

    wire inputRegPage1_15, inputRegPage1_14, inputRegPage1_13, inputRegPage1_12, 
         inputRegPage1_11, inputRegPage1_10, inputRegPage1_9, inputRegPage1_8, 
         inputRegPage1_7, inputRegPage1_6, inputRegPage1_5, inputRegPage1_4, 
         inputRegPage1_3, inputRegPage1_2, inputRegPage1_1, inputRegPage1_0, 
         inputRegPage2_15, inputRegPage2_14, inputRegPage2_13, inputRegPage2_12, 
         inputRegPage2_11, inputRegPage2_10, inputRegPage2_9, inputRegPage2_8, 
         inputRegPage2_7, inputRegPage2_6, inputRegPage2_5, inputRegPage2_4, 
         inputRegPage2_3, inputRegPage2_2, inputRegPage2_1, inputRegPage2_0, 
         reg1TotalEnable, reg2TotalEnable;



    Mux2_16 inputRegPage1Map (.A ({windowBus[15],windowBus[14],windowBus[13],
            windowBus[12],windowBus[11],windowBus[10],windowBus[9],windowBus[8],
            windowBus[7],windowBus[6],windowBus[5],windowBus[4],windowBus[3],
            windowBus[2],windowBus[1],windowBus[0]}), .B ({regPage2NextUnit[15],
            regPage2NextUnit[14],regPage2NextUnit[13],regPage2NextUnit[12],
            regPage2NextUnit[11],regPage2NextUnit[10],regPage2NextUnit[9],
            regPage2NextUnit[8],regPage2NextUnit[7],regPage2NextUnit[6],
            regPage2NextUnit[5],regPage2NextUnit[4],regPage2NextUnit[3],
            regPage2NextUnit[2],regPage2NextUnit[1],regPage2NextUnit[0]}), .S (
            page1ReadBusOrPage2), .C ({inputRegPage1_15,inputRegPage1_14,
            inputRegPage1_13,inputRegPage1_12,inputRegPage1_11,inputRegPage1_10,
            inputRegPage1_9,inputRegPage1_8,inputRegPage1_7,inputRegPage1_6,
            inputRegPage1_5,inputRegPage1_4,inputRegPage1_3,inputRegPage1_2,
            inputRegPage1_1,inputRegPage1_0})) ;
    Mux2_16 inputRegPage2Map (.A ({windowBus[15],windowBus[14],windowBus[13],
            windowBus[12],windowBus[11],windowBus[10],windowBus[9],windowBus[8],
            windowBus[7],windowBus[6],windowBus[5],windowBus[4],windowBus[3],
            windowBus[2],windowBus[1],windowBus[0]}), .B ({regPage1NextUnit[15],
            regPage1NextUnit[14],regPage1NextUnit[13],regPage1NextUnit[12],
            regPage1NextUnit[11],regPage1NextUnit[10],regPage1NextUnit[9],
            regPage1NextUnit[8],regPage1NextUnit[7],regPage1NextUnit[6],
            regPage1NextUnit[5],regPage1NextUnit[4],regPage1NextUnit[3],
            regPage1NextUnit[2],regPage1NextUnit[1],regPage1NextUnit[0]}), .S (
            page2ReadBusOrPage1), .C ({inputRegPage2_15,inputRegPage2_14,
            inputRegPage2_13,inputRegPage2_12,inputRegPage2_11,inputRegPage2_10,
            inputRegPage2_9,inputRegPage2_8,inputRegPage2_7,inputRegPage2_6,
            inputRegPage2_5,inputRegPage2_4,inputRegPage2_3,inputRegPage2_2,
            inputRegPage2_1,inputRegPage2_0})) ;
    Reg_16 regPage1Map (.D ({inputRegPage1_15,inputRegPage1_14,inputRegPage1_13,
           inputRegPage1_12,inputRegPage1_11,inputRegPage1_10,inputRegPage1_9,
           inputRegPage1_8,inputRegPage1_7,inputRegPage1_6,inputRegPage1_5,
           inputRegPage1_4,inputRegPage1_3,inputRegPage1_2,inputRegPage1_1,
           inputRegPage1_0}), .en (reg1TotalEnable), .clk (clk), .rst (rst), .Q (
           {outputRegPage1[15],outputRegPage1[14],outputRegPage1[13],
           outputRegPage1[12],outputRegPage1[11],outputRegPage1[10],
           outputRegPage1[9],outputRegPage1[8],outputRegPage1[7],
           outputRegPage1[6],outputRegPage1[5],outputRegPage1[4],
           outputRegPage1[3],outputRegPage1[2],outputRegPage1[1],
           outputRegPage1[0]})) ;
    Reg_16 regPage2Map (.D ({inputRegPage2_15,inputRegPage2_14,inputRegPage2_13,
           inputRegPage2_12,inputRegPage2_11,inputRegPage2_10,inputRegPage2_9,
           inputRegPage2_8,inputRegPage2_7,inputRegPage2_6,inputRegPage2_5,
           inputRegPage2_4,inputRegPage2_3,inputRegPage2_2,inputRegPage2_1,
           inputRegPage2_0}), .en (reg2TotalEnable), .clk (clk), .rst (rst), .Q (
           {outputRegPage2[15],outputRegPage2[14],outputRegPage2[13],
           outputRegPage2[12],outputRegPage2[11],outputRegPage2[10],
           outputRegPage2[9],outputRegPage2[8],outputRegPage2[7],
           outputRegPage2[6],outputRegPage2[5],outputRegPage2[4],
           outputRegPage2[3],outputRegPage2[2],outputRegPage2[1],
           outputRegPage2[0]})) ;
    Reg_8 regFilterMap (.D ({filterBus[7],filterBus[6],filterBus[5],filterBus[4]
          ,filterBus[3],filterBus[2],filterBus[1],filterBus[0]}), .en (
          enableRegFilter), .clk (clk), .rst (rst), .Q ({outFilter[7],
          outFilter[6],outFilter[5],outFilter[4],outFilter[3],outFilter[2],
          outFilter[1],outFilter[0]})) ;
    Mux2_16 outPageMap (.A ({outputRegPage1[15],outputRegPage1[14],
            outputRegPage1[13],outputRegPage1[12],outputRegPage1[11],
            outputRegPage1[10],outputRegPage1[9],outputRegPage1[8],
            outputRegPage1[7],outputRegPage1[6],outputRegPage1[5],
            outputRegPage1[4],outputRegPage1[3],outputRegPage1[2],
            outputRegPage1[1],outputRegPage1[0]}), .B ({outputRegPage2[15],
            outputRegPage2[14],outputRegPage2[13],outputRegPage2[12],
            outputRegPage2[11],outputRegPage2[10],outputRegPage2[9],
            outputRegPage2[8],outputRegPage2[7],outputRegPage2[6],
            outputRegPage2[5],outputRegPage2[4],outputRegPage2[3],
            outputRegPage2[2],outputRegPage2[1],outputRegPage2[0]}), .S (
            pageTurn), .C ({outRegPage[15],outRegPage[14],outRegPage[13],
            outRegPage[12],outRegPage[11],outRegPage[10],outRegPage[9],
            outRegPage[8],outRegPage[7],outRegPage[6],outRegPage[5],
            outRegPage[4],outRegPage[3],outRegPage[2],outRegPage[1],
            outRegPage[0]})) ;
    or02 ix1 (.Y (reg2TotalEnable), .A0 (enableRegPage2), .A1 (
         page2ReadBusOrPage1)) ;
    or02 ix3 (.Y (reg1TotalEnable), .A0 (enableRegPage1), .A1 (
         page1ReadBusOrPage2)) ;
endmodule


module Reg_8 ( D, en, clk, rst, Q ) ;

    input [7:0]D ;
    input en ;
    input clk ;
    input rst ;
    output [7:0]Q ;

    wire nx132, nx142, nx152, nx162, nx172, nx182, nx192, nx202, nx241, nx243;
    wire [7:0] \$dummy ;




    dffr reg_Q_0 (.Q (Q[0]), .QB (\$dummy [0]), .D (nx132), .CLK (clk), .R (rst)
         ) ;
    mux21_ni ix133 (.Y (nx132), .A0 (Q[0]), .A1 (D[0]), .S0 (nx241)) ;
    dffr reg_Q_1 (.Q (Q[1]), .QB (\$dummy [1]), .D (nx142), .CLK (clk), .R (rst)
         ) ;
    mux21_ni ix143 (.Y (nx142), .A0 (Q[1]), .A1 (D[1]), .S0 (nx241)) ;
    dffr reg_Q_2 (.Q (Q[2]), .QB (\$dummy [2]), .D (nx152), .CLK (clk), .R (rst)
         ) ;
    mux21_ni ix153 (.Y (nx152), .A0 (Q[2]), .A1 (D[2]), .S0 (nx241)) ;
    dffr reg_Q_3 (.Q (Q[3]), .QB (\$dummy [3]), .D (nx162), .CLK (clk), .R (rst)
         ) ;
    mux21_ni ix163 (.Y (nx162), .A0 (Q[3]), .A1 (D[3]), .S0 (nx241)) ;
    dffr reg_Q_4 (.Q (Q[4]), .QB (\$dummy [4]), .D (nx172), .CLK (clk), .R (rst)
         ) ;
    mux21_ni ix173 (.Y (nx172), .A0 (Q[4]), .A1 (D[4]), .S0 (nx241)) ;
    dffr reg_Q_5 (.Q (Q[5]), .QB (\$dummy [5]), .D (nx182), .CLK (clk), .R (rst)
         ) ;
    mux21_ni ix183 (.Y (nx182), .A0 (Q[5]), .A1 (D[5]), .S0 (nx241)) ;
    dffr reg_Q_6 (.Q (Q[6]), .QB (\$dummy [6]), .D (nx192), .CLK (clk), .R (rst)
         ) ;
    mux21_ni ix193 (.Y (nx192), .A0 (Q[6]), .A1 (D[6]), .S0 (nx241)) ;
    dffr reg_Q_7 (.Q (Q[7]), .QB (\$dummy [7]), .D (nx202), .CLK (clk), .R (rst)
         ) ;
    mux21_ni ix203 (.Y (nx202), .A0 (Q[7]), .A1 (D[7]), .S0 (nx243)) ;
    buf02 ix240 (.Y (nx241), .A (en)) ;
    buf02 ix242 (.Y (nx243), .A (en)) ;
endmodule


module Reg_16 ( D, en, clk, rst, Q ) ;

    input [15:0]D ;
    input en ;
    input clk ;
    input rst ;
    output [15:0]Q ;

    wire nx228, nx238, nx248, nx258, nx268, nx278, nx288, nx298, nx308, nx318, 
         nx328, nx338, nx348, nx358, nx368, nx378, nx441, nx443, nx445, nx447, 
         nx449, nx451, nx453, nx455;
    wire [15:0] \$dummy ;




    dffr reg_Q_0 (.Q (Q[0]), .QB (\$dummy [0]), .D (nx228), .CLK (nx451), .R (
         rst)) ;
    mux21_ni ix229 (.Y (nx228), .A0 (Q[0]), .A1 (D[0]), .S0 (nx443)) ;
    dffr reg_Q_1 (.Q (Q[1]), .QB (\$dummy [1]), .D (nx238), .CLK (nx451), .R (
         rst)) ;
    mux21_ni ix239 (.Y (nx238), .A0 (Q[1]), .A1 (D[1]), .S0 (nx443)) ;
    dffr reg_Q_2 (.Q (Q[2]), .QB (\$dummy [2]), .D (nx248), .CLK (nx451), .R (
         rst)) ;
    mux21_ni ix249 (.Y (nx248), .A0 (Q[2]), .A1 (D[2]), .S0 (nx443)) ;
    dffr reg_Q_3 (.Q (Q[3]), .QB (\$dummy [3]), .D (nx258), .CLK (nx451), .R (
         rst)) ;
    mux21_ni ix259 (.Y (nx258), .A0 (Q[3]), .A1 (D[3]), .S0 (nx443)) ;
    dffr reg_Q_4 (.Q (Q[4]), .QB (\$dummy [4]), .D (nx268), .CLK (nx451), .R (
         rst)) ;
    mux21_ni ix269 (.Y (nx268), .A0 (Q[4]), .A1 (D[4]), .S0 (nx443)) ;
    dffr reg_Q_5 (.Q (Q[5]), .QB (\$dummy [5]), .D (nx278), .CLK (nx451), .R (
         rst)) ;
    mux21_ni ix279 (.Y (nx278), .A0 (Q[5]), .A1 (D[5]), .S0 (nx443)) ;
    dffr reg_Q_6 (.Q (Q[6]), .QB (\$dummy [6]), .D (nx288), .CLK (nx451), .R (
         rst)) ;
    mux21_ni ix289 (.Y (nx288), .A0 (Q[6]), .A1 (D[6]), .S0 (nx443)) ;
    dffr reg_Q_7 (.Q (Q[7]), .QB (\$dummy [7]), .D (nx298), .CLK (nx453), .R (
         rst)) ;
    mux21_ni ix299 (.Y (nx298), .A0 (Q[7]), .A1 (D[7]), .S0 (nx445)) ;
    dffr reg_Q_8 (.Q (Q[8]), .QB (\$dummy [8]), .D (nx308), .CLK (nx453), .R (
         rst)) ;
    mux21_ni ix309 (.Y (nx308), .A0 (Q[8]), .A1 (D[8]), .S0 (nx445)) ;
    dffr reg_Q_9 (.Q (Q[9]), .QB (\$dummy [9]), .D (nx318), .CLK (nx453), .R (
         rst)) ;
    mux21_ni ix319 (.Y (nx318), .A0 (Q[9]), .A1 (D[9]), .S0 (nx445)) ;
    dffr reg_Q_10 (.Q (Q[10]), .QB (\$dummy [10]), .D (nx328), .CLK (nx453), .R (
         rst)) ;
    mux21_ni ix329 (.Y (nx328), .A0 (Q[10]), .A1 (D[10]), .S0 (nx445)) ;
    dffr reg_Q_11 (.Q (Q[11]), .QB (\$dummy [11]), .D (nx338), .CLK (nx453), .R (
         rst)) ;
    mux21_ni ix339 (.Y (nx338), .A0 (Q[11]), .A1 (D[11]), .S0 (nx445)) ;
    dffr reg_Q_12 (.Q (Q[12]), .QB (\$dummy [12]), .D (nx348), .CLK (nx453), .R (
         rst)) ;
    mux21_ni ix349 (.Y (nx348), .A0 (Q[12]), .A1 (D[12]), .S0 (nx445)) ;
    dffr reg_Q_13 (.Q (Q[13]), .QB (\$dummy [13]), .D (nx358), .CLK (nx453), .R (
         rst)) ;
    mux21_ni ix359 (.Y (nx358), .A0 (Q[13]), .A1 (D[13]), .S0 (nx445)) ;
    dffr reg_Q_14 (.Q (Q[14]), .QB (\$dummy [14]), .D (nx368), .CLK (nx455), .R (
         rst)) ;
    mux21_ni ix369 (.Y (nx368), .A0 (Q[14]), .A1 (D[14]), .S0 (nx447)) ;
    dffr reg_Q_15 (.Q (Q[15]), .QB (\$dummy [15]), .D (nx378), .CLK (nx455), .R (
         rst)) ;
    mux21_ni ix379 (.Y (nx378), .A0 (Q[15]), .A1 (D[15]), .S0 (nx447)) ;
    inv01 ix440 (.Y (nx441), .A (en)) ;
    inv02 ix442 (.Y (nx443), .A (nx441)) ;
    inv02 ix444 (.Y (nx445), .A (nx441)) ;
    inv02 ix446 (.Y (nx447), .A (nx441)) ;
    inv01 ix448 (.Y (nx449), .A (clk)) ;
    inv02 ix450 (.Y (nx451), .A (nx449)) ;
    inv02 ix452 (.Y (nx453), .A (nx449)) ;
    inv02 ix454 (.Y (nx455), .A (nx449)) ;
endmodule


module Mux2_16 ( A, B, S, C ) ;

    input [15:0]A ;
    input [15:0]B ;
    input S ;
    output [15:0]C ;

    wire nx173, nx175, nx177, nx179;



    mux21_ni ix7 (.Y (C[0]), .A0 (A[0]), .A1 (B[0]), .S0 (nx175)) ;
    mux21_ni ix15 (.Y (C[1]), .A0 (A[1]), .A1 (B[1]), .S0 (nx175)) ;
    mux21_ni ix23 (.Y (C[2]), .A0 (A[2]), .A1 (B[2]), .S0 (nx175)) ;
    mux21_ni ix31 (.Y (C[3]), .A0 (A[3]), .A1 (B[3]), .S0 (nx175)) ;
    mux21_ni ix39 (.Y (C[4]), .A0 (A[4]), .A1 (B[4]), .S0 (nx175)) ;
    mux21_ni ix47 (.Y (C[5]), .A0 (A[5]), .A1 (B[5]), .S0 (nx175)) ;
    mux21_ni ix55 (.Y (C[6]), .A0 (A[6]), .A1 (B[6]), .S0 (nx175)) ;
    mux21_ni ix63 (.Y (C[7]), .A0 (A[7]), .A1 (B[7]), .S0 (nx177)) ;
    mux21_ni ix71 (.Y (C[8]), .A0 (A[8]), .A1 (B[8]), .S0 (nx177)) ;
    mux21_ni ix79 (.Y (C[9]), .A0 (A[9]), .A1 (B[9]), .S0 (nx177)) ;
    mux21_ni ix87 (.Y (C[10]), .A0 (A[10]), .A1 (B[10]), .S0 (nx177)) ;
    mux21_ni ix95 (.Y (C[11]), .A0 (A[11]), .A1 (B[11]), .S0 (nx177)) ;
    mux21_ni ix103 (.Y (C[12]), .A0 (A[12]), .A1 (B[12]), .S0 (nx177)) ;
    mux21_ni ix111 (.Y (C[13]), .A0 (A[13]), .A1 (B[13]), .S0 (nx177)) ;
    mux21_ni ix119 (.Y (C[14]), .A0 (A[14]), .A1 (B[14]), .S0 (nx179)) ;
    mux21_ni ix127 (.Y (C[15]), .A0 (A[15]), .A1 (B[15]), .S0 (nx179)) ;
    inv01 ix172 (.Y (nx173), .A (S)) ;
    inv02 ix174 (.Y (nx175), .A (nx173)) ;
    inv02 ix176 (.Y (nx177), .A (nx173)) ;
    inv02 ix178 (.Y (nx179), .A (nx173)) ;
endmodule


module Decoder_3 ( T, en, decoded ) ;

    input [2:0]T ;
    input en ;
    output [7:0]decoded ;

    wire nx28, nx108, nx110, nx112, nx120, nx131, nx133;



    nor03_2x ix5 (.Y (decoded[7]), .A0 (nx108), .A1 (nx110), .A2 (nx112)) ;
    nand02 ix109 (.Y (nx108), .A0 (T[2]), .A1 (en)) ;
    inv02 ix111 (.Y (nx110), .A (T[1])) ;
    inv02 ix113 (.Y (nx112), .A (T[0])) ;
    nor03_2x ix11 (.Y (decoded[6]), .A0 (nx108), .A1 (nx110), .A2 (nx133)) ;
    nor03_2x ix17 (.Y (decoded[5]), .A0 (nx108), .A1 (nx131), .A2 (nx112)) ;
    nor03_2x ix25 (.Y (decoded[4]), .A0 (nx108), .A1 (nx131), .A2 (nx133)) ;
    and03 ix33 (.Y (decoded[3]), .A0 (nx28), .A1 (nx131), .A2 (nx133)) ;
    nor02ii ix29 (.Y (nx28), .A0 (T[2]), .A1 (en)) ;
    nor03_2x ix39 (.Y (decoded[2]), .A0 (nx120), .A1 (nx110), .A2 (nx133)) ;
    nor03_2x ix45 (.Y (decoded[1]), .A0 (nx120), .A1 (nx131), .A2 (nx112)) ;
    nor03_2x ix53 (.Y (decoded[0]), .A0 (nx120), .A1 (nx131), .A2 (nx133)) ;
    inv01 ix121 (.Y (nx120), .A (nx28)) ;
    inv02 ix130 (.Y (nx131), .A (nx110)) ;
    inv02 ix132 (.Y (nx133), .A (nx112)) ;
endmodule

