//
// Verilog description for cell RegFile, 
// Wed Apr 10 18:03:36 2019
//
// LeonardoSpectrum Level 3, 2018a.2 
//


module RegFile ( filterBus, windowBus, decoderRow, clk, rst, enablePage1Read, 
                 enablePage2Read, enableFilterRead, shift2To1, shift1To2, 
                 pageTurn, pagesOuts_0__15, pagesOuts_0__14, pagesOuts_0__13, 
                 pagesOuts_0__12, pagesOuts_0__11, pagesOuts_0__10, 
                 pagesOuts_0__9, pagesOuts_0__8, pagesOuts_0__7, pagesOuts_0__6, 
                 pagesOuts_0__5, pagesOuts_0__4, pagesOuts_0__3, pagesOuts_0__2, 
                 pagesOuts_0__1, pagesOuts_0__0, pagesOuts_1__15, 
                 pagesOuts_1__14, pagesOuts_1__13, pagesOuts_1__12, 
                 pagesOuts_1__11, pagesOuts_1__10, pagesOuts_1__9, 
                 pagesOuts_1__8, pagesOuts_1__7, pagesOuts_1__6, pagesOuts_1__5, 
                 pagesOuts_1__4, pagesOuts_1__3, pagesOuts_1__2, pagesOuts_1__1, 
                 pagesOuts_1__0, pagesOuts_2__15, pagesOuts_2__14, 
                 pagesOuts_2__13, pagesOuts_2__12, pagesOuts_2__11, 
                 pagesOuts_2__10, pagesOuts_2__9, pagesOuts_2__8, pagesOuts_2__7, 
                 pagesOuts_2__6, pagesOuts_2__5, pagesOuts_2__4, pagesOuts_2__3, 
                 pagesOuts_2__2, pagesOuts_2__1, pagesOuts_2__0, pagesOuts_3__15, 
                 pagesOuts_3__14, pagesOuts_3__13, pagesOuts_3__12, 
                 pagesOuts_3__11, pagesOuts_3__10, pagesOuts_3__9, 
                 pagesOuts_3__8, pagesOuts_3__7, pagesOuts_3__6, pagesOuts_3__5, 
                 pagesOuts_3__4, pagesOuts_3__3, pagesOuts_3__2, pagesOuts_3__1, 
                 pagesOuts_3__0, pagesOuts_4__15, pagesOuts_4__14, 
                 pagesOuts_4__13, pagesOuts_4__12, pagesOuts_4__11, 
                 pagesOuts_4__10, pagesOuts_4__9, pagesOuts_4__8, pagesOuts_4__7, 
                 pagesOuts_4__6, pagesOuts_4__5, pagesOuts_4__4, pagesOuts_4__3, 
                 pagesOuts_4__2, pagesOuts_4__1, pagesOuts_4__0, pagesOuts_5__15, 
                 pagesOuts_5__14, pagesOuts_5__13, pagesOuts_5__12, 
                 pagesOuts_5__11, pagesOuts_5__10, pagesOuts_5__9, 
                 pagesOuts_5__8, pagesOuts_5__7, pagesOuts_5__6, pagesOuts_5__5, 
                 pagesOuts_5__4, pagesOuts_5__3, pagesOuts_5__2, pagesOuts_5__1, 
                 pagesOuts_5__0, pagesOuts_6__15, pagesOuts_6__14, 
                 pagesOuts_6__13, pagesOuts_6__12, pagesOuts_6__11, 
                 pagesOuts_6__10, pagesOuts_6__9, pagesOuts_6__8, pagesOuts_6__7, 
                 pagesOuts_6__6, pagesOuts_6__5, pagesOuts_6__4, pagesOuts_6__3, 
                 pagesOuts_6__2, pagesOuts_6__1, pagesOuts_6__0, pagesOuts_7__15, 
                 pagesOuts_7__14, pagesOuts_7__13, pagesOuts_7__12, 
                 pagesOuts_7__11, pagesOuts_7__10, pagesOuts_7__9, 
                 pagesOuts_7__8, pagesOuts_7__7, pagesOuts_7__6, pagesOuts_7__5, 
                 pagesOuts_7__4, pagesOuts_7__3, pagesOuts_7__2, pagesOuts_7__1, 
                 pagesOuts_7__0, pagesOuts_8__15, pagesOuts_8__14, 
                 pagesOuts_8__13, pagesOuts_8__12, pagesOuts_8__11, 
                 pagesOuts_8__10, pagesOuts_8__9, pagesOuts_8__8, pagesOuts_8__7, 
                 pagesOuts_8__6, pagesOuts_8__5, pagesOuts_8__4, pagesOuts_8__3, 
                 pagesOuts_8__2, pagesOuts_8__1, pagesOuts_8__0, pagesOuts_9__15, 
                 pagesOuts_9__14, pagesOuts_9__13, pagesOuts_9__12, 
                 pagesOuts_9__11, pagesOuts_9__10, pagesOuts_9__9, 
                 pagesOuts_9__8, pagesOuts_9__7, pagesOuts_9__6, pagesOuts_9__5, 
                 pagesOuts_9__4, pagesOuts_9__3, pagesOuts_9__2, pagesOuts_9__1, 
                 pagesOuts_9__0, pagesOuts_10__15, pagesOuts_10__14, 
                 pagesOuts_10__13, pagesOuts_10__12, pagesOuts_10__11, 
                 pagesOuts_10__10, pagesOuts_10__9, pagesOuts_10__8, 
                 pagesOuts_10__7, pagesOuts_10__6, pagesOuts_10__5, 
                 pagesOuts_10__4, pagesOuts_10__3, pagesOuts_10__2, 
                 pagesOuts_10__1, pagesOuts_10__0, pagesOuts_11__15, 
                 pagesOuts_11__14, pagesOuts_11__13, pagesOuts_11__12, 
                 pagesOuts_11__11, pagesOuts_11__10, pagesOuts_11__9, 
                 pagesOuts_11__8, pagesOuts_11__7, pagesOuts_11__6, 
                 pagesOuts_11__5, pagesOuts_11__4, pagesOuts_11__3, 
                 pagesOuts_11__2, pagesOuts_11__1, pagesOuts_11__0, 
                 pagesOuts_12__15, pagesOuts_12__14, pagesOuts_12__13, 
                 pagesOuts_12__12, pagesOuts_12__11, pagesOuts_12__10, 
                 pagesOuts_12__9, pagesOuts_12__8, pagesOuts_12__7, 
                 pagesOuts_12__6, pagesOuts_12__5, pagesOuts_12__4, 
                 pagesOuts_12__3, pagesOuts_12__2, pagesOuts_12__1, 
                 pagesOuts_12__0, pagesOuts_13__15, pagesOuts_13__14, 
                 pagesOuts_13__13, pagesOuts_13__12, pagesOuts_13__11, 
                 pagesOuts_13__10, pagesOuts_13__9, pagesOuts_13__8, 
                 pagesOuts_13__7, pagesOuts_13__6, pagesOuts_13__5, 
                 pagesOuts_13__4, pagesOuts_13__3, pagesOuts_13__2, 
                 pagesOuts_13__1, pagesOuts_13__0, pagesOuts_14__15, 
                 pagesOuts_14__14, pagesOuts_14__13, pagesOuts_14__12, 
                 pagesOuts_14__11, pagesOuts_14__10, pagesOuts_14__9, 
                 pagesOuts_14__8, pagesOuts_14__7, pagesOuts_14__6, 
                 pagesOuts_14__5, pagesOuts_14__4, pagesOuts_14__3, 
                 pagesOuts_14__2, pagesOuts_14__1, pagesOuts_14__0, 
                 pagesOuts_15__15, pagesOuts_15__14, pagesOuts_15__13, 
                 pagesOuts_15__12, pagesOuts_15__11, pagesOuts_15__10, 
                 pagesOuts_15__9, pagesOuts_15__8, pagesOuts_15__7, 
                 pagesOuts_15__6, pagesOuts_15__5, pagesOuts_15__4, 
                 pagesOuts_15__3, pagesOuts_15__2, pagesOuts_15__1, 
                 pagesOuts_15__0, pagesOuts_16__15, pagesOuts_16__14, 
                 pagesOuts_16__13, pagesOuts_16__12, pagesOuts_16__11, 
                 pagesOuts_16__10, pagesOuts_16__9, pagesOuts_16__8, 
                 pagesOuts_16__7, pagesOuts_16__6, pagesOuts_16__5, 
                 pagesOuts_16__4, pagesOuts_16__3, pagesOuts_16__2, 
                 pagesOuts_16__1, pagesOuts_16__0, pagesOuts_17__15, 
                 pagesOuts_17__14, pagesOuts_17__13, pagesOuts_17__12, 
                 pagesOuts_17__11, pagesOuts_17__10, pagesOuts_17__9, 
                 pagesOuts_17__8, pagesOuts_17__7, pagesOuts_17__6, 
                 pagesOuts_17__5, pagesOuts_17__4, pagesOuts_17__3, 
                 pagesOuts_17__2, pagesOuts_17__1, pagesOuts_17__0, 
                 pagesOuts_18__15, pagesOuts_18__14, pagesOuts_18__13, 
                 pagesOuts_18__12, pagesOuts_18__11, pagesOuts_18__10, 
                 pagesOuts_18__9, pagesOuts_18__8, pagesOuts_18__7, 
                 pagesOuts_18__6, pagesOuts_18__5, pagesOuts_18__4, 
                 pagesOuts_18__3, pagesOuts_18__2, pagesOuts_18__1, 
                 pagesOuts_18__0, pagesOuts_19__15, pagesOuts_19__14, 
                 pagesOuts_19__13, pagesOuts_19__12, pagesOuts_19__11, 
                 pagesOuts_19__10, pagesOuts_19__9, pagesOuts_19__8, 
                 pagesOuts_19__7, pagesOuts_19__6, pagesOuts_19__5, 
                 pagesOuts_19__4, pagesOuts_19__3, pagesOuts_19__2, 
                 pagesOuts_19__1, pagesOuts_19__0, pagesOuts_20__15, 
                 pagesOuts_20__14, pagesOuts_20__13, pagesOuts_20__12, 
                 pagesOuts_20__11, pagesOuts_20__10, pagesOuts_20__9, 
                 pagesOuts_20__8, pagesOuts_20__7, pagesOuts_20__6, 
                 pagesOuts_20__5, pagesOuts_20__4, pagesOuts_20__3, 
                 pagesOuts_20__2, pagesOuts_20__1, pagesOuts_20__0, 
                 pagesOuts_21__15, pagesOuts_21__14, pagesOuts_21__13, 
                 pagesOuts_21__12, pagesOuts_21__11, pagesOuts_21__10, 
                 pagesOuts_21__9, pagesOuts_21__8, pagesOuts_21__7, 
                 pagesOuts_21__6, pagesOuts_21__5, pagesOuts_21__4, 
                 pagesOuts_21__3, pagesOuts_21__2, pagesOuts_21__1, 
                 pagesOuts_21__0, pagesOuts_22__15, pagesOuts_22__14, 
                 pagesOuts_22__13, pagesOuts_22__12, pagesOuts_22__11, 
                 pagesOuts_22__10, pagesOuts_22__9, pagesOuts_22__8, 
                 pagesOuts_22__7, pagesOuts_22__6, pagesOuts_22__5, 
                 pagesOuts_22__4, pagesOuts_22__3, pagesOuts_22__2, 
                 pagesOuts_22__1, pagesOuts_22__0, pagesOuts_23__15, 
                 pagesOuts_23__14, pagesOuts_23__13, pagesOuts_23__12, 
                 pagesOuts_23__11, pagesOuts_23__10, pagesOuts_23__9, 
                 pagesOuts_23__8, pagesOuts_23__7, pagesOuts_23__6, 
                 pagesOuts_23__5, pagesOuts_23__4, pagesOuts_23__3, 
                 pagesOuts_23__2, pagesOuts_23__1, pagesOuts_23__0, 
                 pagesOuts_24__15, pagesOuts_24__14, pagesOuts_24__13, 
                 pagesOuts_24__12, pagesOuts_24__11, pagesOuts_24__10, 
                 pagesOuts_24__9, pagesOuts_24__8, pagesOuts_24__7, 
                 pagesOuts_24__6, pagesOuts_24__5, pagesOuts_24__4, 
                 pagesOuts_24__3, pagesOuts_24__2, pagesOuts_24__1, 
                 pagesOuts_24__0, filtersOuts_0__7, filtersOuts_0__6, 
                 filtersOuts_0__5, filtersOuts_0__4, filtersOuts_0__3, 
                 filtersOuts_0__2, filtersOuts_0__1, filtersOuts_0__0, 
                 filtersOuts_1__7, filtersOuts_1__6, filtersOuts_1__5, 
                 filtersOuts_1__4, filtersOuts_1__3, filtersOuts_1__2, 
                 filtersOuts_1__1, filtersOuts_1__0, filtersOuts_2__7, 
                 filtersOuts_2__6, filtersOuts_2__5, filtersOuts_2__4, 
                 filtersOuts_2__3, filtersOuts_2__2, filtersOuts_2__1, 
                 filtersOuts_2__0, filtersOuts_3__7, filtersOuts_3__6, 
                 filtersOuts_3__5, filtersOuts_3__4, filtersOuts_3__3, 
                 filtersOuts_3__2, filtersOuts_3__1, filtersOuts_3__0, 
                 filtersOuts_4__7, filtersOuts_4__6, filtersOuts_4__5, 
                 filtersOuts_4__4, filtersOuts_4__3, filtersOuts_4__2, 
                 filtersOuts_4__1, filtersOuts_4__0, filtersOuts_5__7, 
                 filtersOuts_5__6, filtersOuts_5__5, filtersOuts_5__4, 
                 filtersOuts_5__3, filtersOuts_5__2, filtersOuts_5__1, 
                 filtersOuts_5__0, filtersOuts_6__7, filtersOuts_6__6, 
                 filtersOuts_6__5, filtersOuts_6__4, filtersOuts_6__3, 
                 filtersOuts_6__2, filtersOuts_6__1, filtersOuts_6__0, 
                 filtersOuts_7__7, filtersOuts_7__6, filtersOuts_7__5, 
                 filtersOuts_7__4, filtersOuts_7__3, filtersOuts_7__2, 
                 filtersOuts_7__1, filtersOuts_7__0, filtersOuts_8__7, 
                 filtersOuts_8__6, filtersOuts_8__5, filtersOuts_8__4, 
                 filtersOuts_8__3, filtersOuts_8__2, filtersOuts_8__1, 
                 filtersOuts_8__0, filtersOuts_9__7, filtersOuts_9__6, 
                 filtersOuts_9__5, filtersOuts_9__4, filtersOuts_9__3, 
                 filtersOuts_9__2, filtersOuts_9__1, filtersOuts_9__0, 
                 filtersOuts_10__7, filtersOuts_10__6, filtersOuts_10__5, 
                 filtersOuts_10__4, filtersOuts_10__3, filtersOuts_10__2, 
                 filtersOuts_10__1, filtersOuts_10__0, filtersOuts_11__7, 
                 filtersOuts_11__6, filtersOuts_11__5, filtersOuts_11__4, 
                 filtersOuts_11__3, filtersOuts_11__2, filtersOuts_11__1, 
                 filtersOuts_11__0, filtersOuts_12__7, filtersOuts_12__6, 
                 filtersOuts_12__5, filtersOuts_12__4, filtersOuts_12__3, 
                 filtersOuts_12__2, filtersOuts_12__1, filtersOuts_12__0, 
                 filtersOuts_13__7, filtersOuts_13__6, filtersOuts_13__5, 
                 filtersOuts_13__4, filtersOuts_13__3, filtersOuts_13__2, 
                 filtersOuts_13__1, filtersOuts_13__0, filtersOuts_14__7, 
                 filtersOuts_14__6, filtersOuts_14__5, filtersOuts_14__4, 
                 filtersOuts_14__3, filtersOuts_14__2, filtersOuts_14__1, 
                 filtersOuts_14__0, filtersOuts_15__7, filtersOuts_15__6, 
                 filtersOuts_15__5, filtersOuts_15__4, filtersOuts_15__3, 
                 filtersOuts_15__2, filtersOuts_15__1, filtersOuts_15__0, 
                 filtersOuts_16__7, filtersOuts_16__6, filtersOuts_16__5, 
                 filtersOuts_16__4, filtersOuts_16__3, filtersOuts_16__2, 
                 filtersOuts_16__1, filtersOuts_16__0, filtersOuts_17__7, 
                 filtersOuts_17__6, filtersOuts_17__5, filtersOuts_17__4, 
                 filtersOuts_17__3, filtersOuts_17__2, filtersOuts_17__1, 
                 filtersOuts_17__0, filtersOuts_18__7, filtersOuts_18__6, 
                 filtersOuts_18__5, filtersOuts_18__4, filtersOuts_18__3, 
                 filtersOuts_18__2, filtersOuts_18__1, filtersOuts_18__0, 
                 filtersOuts_19__7, filtersOuts_19__6, filtersOuts_19__5, 
                 filtersOuts_19__4, filtersOuts_19__3, filtersOuts_19__2, 
                 filtersOuts_19__1, filtersOuts_19__0, filtersOuts_20__7, 
                 filtersOuts_20__6, filtersOuts_20__5, filtersOuts_20__4, 
                 filtersOuts_20__3, filtersOuts_20__2, filtersOuts_20__1, 
                 filtersOuts_20__0, filtersOuts_21__7, filtersOuts_21__6, 
                 filtersOuts_21__5, filtersOuts_21__4, filtersOuts_21__3, 
                 filtersOuts_21__2, filtersOuts_21__1, filtersOuts_21__0, 
                 filtersOuts_22__7, filtersOuts_22__6, filtersOuts_22__5, 
                 filtersOuts_22__4, filtersOuts_22__3, filtersOuts_22__2, 
                 filtersOuts_22__1, filtersOuts_22__0, filtersOuts_23__7, 
                 filtersOuts_23__6, filtersOuts_23__5, filtersOuts_23__4, 
                 filtersOuts_23__3, filtersOuts_23__2, filtersOuts_23__1, 
                 filtersOuts_23__0, filtersOuts_24__7, filtersOuts_24__6, 
                 filtersOuts_24__5, filtersOuts_24__4, filtersOuts_24__3, 
                 filtersOuts_24__2, filtersOuts_24__1, filtersOuts_24__0 ) ;

    input [39:0]filterBus ;
    input [79:0]windowBus ;
    input [2:0]decoderRow ;
    input clk ;
    input rst ;
    input enablePage1Read ;
    input enablePage2Read ;
    input enableFilterRead ;
    input shift2To1 ;
    input shift1To2 ;
    input pageTurn ;
    output pagesOuts_0__15 ;
    output pagesOuts_0__14 ;
    output pagesOuts_0__13 ;
    output pagesOuts_0__12 ;
    output pagesOuts_0__11 ;
    output pagesOuts_0__10 ;
    output pagesOuts_0__9 ;
    output pagesOuts_0__8 ;
    output pagesOuts_0__7 ;
    output pagesOuts_0__6 ;
    output pagesOuts_0__5 ;
    output pagesOuts_0__4 ;
    output pagesOuts_0__3 ;
    output pagesOuts_0__2 ;
    output pagesOuts_0__1 ;
    output pagesOuts_0__0 ;
    output pagesOuts_1__15 ;
    output pagesOuts_1__14 ;
    output pagesOuts_1__13 ;
    output pagesOuts_1__12 ;
    output pagesOuts_1__11 ;
    output pagesOuts_1__10 ;
    output pagesOuts_1__9 ;
    output pagesOuts_1__8 ;
    output pagesOuts_1__7 ;
    output pagesOuts_1__6 ;
    output pagesOuts_1__5 ;
    output pagesOuts_1__4 ;
    output pagesOuts_1__3 ;
    output pagesOuts_1__2 ;
    output pagesOuts_1__1 ;
    output pagesOuts_1__0 ;
    output pagesOuts_2__15 ;
    output pagesOuts_2__14 ;
    output pagesOuts_2__13 ;
    output pagesOuts_2__12 ;
    output pagesOuts_2__11 ;
    output pagesOuts_2__10 ;
    output pagesOuts_2__9 ;
    output pagesOuts_2__8 ;
    output pagesOuts_2__7 ;
    output pagesOuts_2__6 ;
    output pagesOuts_2__5 ;
    output pagesOuts_2__4 ;
    output pagesOuts_2__3 ;
    output pagesOuts_2__2 ;
    output pagesOuts_2__1 ;
    output pagesOuts_2__0 ;
    output pagesOuts_3__15 ;
    output pagesOuts_3__14 ;
    output pagesOuts_3__13 ;
    output pagesOuts_3__12 ;
    output pagesOuts_3__11 ;
    output pagesOuts_3__10 ;
    output pagesOuts_3__9 ;
    output pagesOuts_3__8 ;
    output pagesOuts_3__7 ;
    output pagesOuts_3__6 ;
    output pagesOuts_3__5 ;
    output pagesOuts_3__4 ;
    output pagesOuts_3__3 ;
    output pagesOuts_3__2 ;
    output pagesOuts_3__1 ;
    output pagesOuts_3__0 ;
    output pagesOuts_4__15 ;
    output pagesOuts_4__14 ;
    output pagesOuts_4__13 ;
    output pagesOuts_4__12 ;
    output pagesOuts_4__11 ;
    output pagesOuts_4__10 ;
    output pagesOuts_4__9 ;
    output pagesOuts_4__8 ;
    output pagesOuts_4__7 ;
    output pagesOuts_4__6 ;
    output pagesOuts_4__5 ;
    output pagesOuts_4__4 ;
    output pagesOuts_4__3 ;
    output pagesOuts_4__2 ;
    output pagesOuts_4__1 ;
    output pagesOuts_4__0 ;
    output pagesOuts_5__15 ;
    output pagesOuts_5__14 ;
    output pagesOuts_5__13 ;
    output pagesOuts_5__12 ;
    output pagesOuts_5__11 ;
    output pagesOuts_5__10 ;
    output pagesOuts_5__9 ;
    output pagesOuts_5__8 ;
    output pagesOuts_5__7 ;
    output pagesOuts_5__6 ;
    output pagesOuts_5__5 ;
    output pagesOuts_5__4 ;
    output pagesOuts_5__3 ;
    output pagesOuts_5__2 ;
    output pagesOuts_5__1 ;
    output pagesOuts_5__0 ;
    output pagesOuts_6__15 ;
    output pagesOuts_6__14 ;
    output pagesOuts_6__13 ;
    output pagesOuts_6__12 ;
    output pagesOuts_6__11 ;
    output pagesOuts_6__10 ;
    output pagesOuts_6__9 ;
    output pagesOuts_6__8 ;
    output pagesOuts_6__7 ;
    output pagesOuts_6__6 ;
    output pagesOuts_6__5 ;
    output pagesOuts_6__4 ;
    output pagesOuts_6__3 ;
    output pagesOuts_6__2 ;
    output pagesOuts_6__1 ;
    output pagesOuts_6__0 ;
    output pagesOuts_7__15 ;
    output pagesOuts_7__14 ;
    output pagesOuts_7__13 ;
    output pagesOuts_7__12 ;
    output pagesOuts_7__11 ;
    output pagesOuts_7__10 ;
    output pagesOuts_7__9 ;
    output pagesOuts_7__8 ;
    output pagesOuts_7__7 ;
    output pagesOuts_7__6 ;
    output pagesOuts_7__5 ;
    output pagesOuts_7__4 ;
    output pagesOuts_7__3 ;
    output pagesOuts_7__2 ;
    output pagesOuts_7__1 ;
    output pagesOuts_7__0 ;
    output pagesOuts_8__15 ;
    output pagesOuts_8__14 ;
    output pagesOuts_8__13 ;
    output pagesOuts_8__12 ;
    output pagesOuts_8__11 ;
    output pagesOuts_8__10 ;
    output pagesOuts_8__9 ;
    output pagesOuts_8__8 ;
    output pagesOuts_8__7 ;
    output pagesOuts_8__6 ;
    output pagesOuts_8__5 ;
    output pagesOuts_8__4 ;
    output pagesOuts_8__3 ;
    output pagesOuts_8__2 ;
    output pagesOuts_8__1 ;
    output pagesOuts_8__0 ;
    output pagesOuts_9__15 ;
    output pagesOuts_9__14 ;
    output pagesOuts_9__13 ;
    output pagesOuts_9__12 ;
    output pagesOuts_9__11 ;
    output pagesOuts_9__10 ;
    output pagesOuts_9__9 ;
    output pagesOuts_9__8 ;
    output pagesOuts_9__7 ;
    output pagesOuts_9__6 ;
    output pagesOuts_9__5 ;
    output pagesOuts_9__4 ;
    output pagesOuts_9__3 ;
    output pagesOuts_9__2 ;
    output pagesOuts_9__1 ;
    output pagesOuts_9__0 ;
    output pagesOuts_10__15 ;
    output pagesOuts_10__14 ;
    output pagesOuts_10__13 ;
    output pagesOuts_10__12 ;
    output pagesOuts_10__11 ;
    output pagesOuts_10__10 ;
    output pagesOuts_10__9 ;
    output pagesOuts_10__8 ;
    output pagesOuts_10__7 ;
    output pagesOuts_10__6 ;
    output pagesOuts_10__5 ;
    output pagesOuts_10__4 ;
    output pagesOuts_10__3 ;
    output pagesOuts_10__2 ;
    output pagesOuts_10__1 ;
    output pagesOuts_10__0 ;
    output pagesOuts_11__15 ;
    output pagesOuts_11__14 ;
    output pagesOuts_11__13 ;
    output pagesOuts_11__12 ;
    output pagesOuts_11__11 ;
    output pagesOuts_11__10 ;
    output pagesOuts_11__9 ;
    output pagesOuts_11__8 ;
    output pagesOuts_11__7 ;
    output pagesOuts_11__6 ;
    output pagesOuts_11__5 ;
    output pagesOuts_11__4 ;
    output pagesOuts_11__3 ;
    output pagesOuts_11__2 ;
    output pagesOuts_11__1 ;
    output pagesOuts_11__0 ;
    output pagesOuts_12__15 ;
    output pagesOuts_12__14 ;
    output pagesOuts_12__13 ;
    output pagesOuts_12__12 ;
    output pagesOuts_12__11 ;
    output pagesOuts_12__10 ;
    output pagesOuts_12__9 ;
    output pagesOuts_12__8 ;
    output pagesOuts_12__7 ;
    output pagesOuts_12__6 ;
    output pagesOuts_12__5 ;
    output pagesOuts_12__4 ;
    output pagesOuts_12__3 ;
    output pagesOuts_12__2 ;
    output pagesOuts_12__1 ;
    output pagesOuts_12__0 ;
    output pagesOuts_13__15 ;
    output pagesOuts_13__14 ;
    output pagesOuts_13__13 ;
    output pagesOuts_13__12 ;
    output pagesOuts_13__11 ;
    output pagesOuts_13__10 ;
    output pagesOuts_13__9 ;
    output pagesOuts_13__8 ;
    output pagesOuts_13__7 ;
    output pagesOuts_13__6 ;
    output pagesOuts_13__5 ;
    output pagesOuts_13__4 ;
    output pagesOuts_13__3 ;
    output pagesOuts_13__2 ;
    output pagesOuts_13__1 ;
    output pagesOuts_13__0 ;
    output pagesOuts_14__15 ;
    output pagesOuts_14__14 ;
    output pagesOuts_14__13 ;
    output pagesOuts_14__12 ;
    output pagesOuts_14__11 ;
    output pagesOuts_14__10 ;
    output pagesOuts_14__9 ;
    output pagesOuts_14__8 ;
    output pagesOuts_14__7 ;
    output pagesOuts_14__6 ;
    output pagesOuts_14__5 ;
    output pagesOuts_14__4 ;
    output pagesOuts_14__3 ;
    output pagesOuts_14__2 ;
    output pagesOuts_14__1 ;
    output pagesOuts_14__0 ;
    output pagesOuts_15__15 ;
    output pagesOuts_15__14 ;
    output pagesOuts_15__13 ;
    output pagesOuts_15__12 ;
    output pagesOuts_15__11 ;
    output pagesOuts_15__10 ;
    output pagesOuts_15__9 ;
    output pagesOuts_15__8 ;
    output pagesOuts_15__7 ;
    output pagesOuts_15__6 ;
    output pagesOuts_15__5 ;
    output pagesOuts_15__4 ;
    output pagesOuts_15__3 ;
    output pagesOuts_15__2 ;
    output pagesOuts_15__1 ;
    output pagesOuts_15__0 ;
    output pagesOuts_16__15 ;
    output pagesOuts_16__14 ;
    output pagesOuts_16__13 ;
    output pagesOuts_16__12 ;
    output pagesOuts_16__11 ;
    output pagesOuts_16__10 ;
    output pagesOuts_16__9 ;
    output pagesOuts_16__8 ;
    output pagesOuts_16__7 ;
    output pagesOuts_16__6 ;
    output pagesOuts_16__5 ;
    output pagesOuts_16__4 ;
    output pagesOuts_16__3 ;
    output pagesOuts_16__2 ;
    output pagesOuts_16__1 ;
    output pagesOuts_16__0 ;
    output pagesOuts_17__15 ;
    output pagesOuts_17__14 ;
    output pagesOuts_17__13 ;
    output pagesOuts_17__12 ;
    output pagesOuts_17__11 ;
    output pagesOuts_17__10 ;
    output pagesOuts_17__9 ;
    output pagesOuts_17__8 ;
    output pagesOuts_17__7 ;
    output pagesOuts_17__6 ;
    output pagesOuts_17__5 ;
    output pagesOuts_17__4 ;
    output pagesOuts_17__3 ;
    output pagesOuts_17__2 ;
    output pagesOuts_17__1 ;
    output pagesOuts_17__0 ;
    output pagesOuts_18__15 ;
    output pagesOuts_18__14 ;
    output pagesOuts_18__13 ;
    output pagesOuts_18__12 ;
    output pagesOuts_18__11 ;
    output pagesOuts_18__10 ;
    output pagesOuts_18__9 ;
    output pagesOuts_18__8 ;
    output pagesOuts_18__7 ;
    output pagesOuts_18__6 ;
    output pagesOuts_18__5 ;
    output pagesOuts_18__4 ;
    output pagesOuts_18__3 ;
    output pagesOuts_18__2 ;
    output pagesOuts_18__1 ;
    output pagesOuts_18__0 ;
    output pagesOuts_19__15 ;
    output pagesOuts_19__14 ;
    output pagesOuts_19__13 ;
    output pagesOuts_19__12 ;
    output pagesOuts_19__11 ;
    output pagesOuts_19__10 ;
    output pagesOuts_19__9 ;
    output pagesOuts_19__8 ;
    output pagesOuts_19__7 ;
    output pagesOuts_19__6 ;
    output pagesOuts_19__5 ;
    output pagesOuts_19__4 ;
    output pagesOuts_19__3 ;
    output pagesOuts_19__2 ;
    output pagesOuts_19__1 ;
    output pagesOuts_19__0 ;
    output pagesOuts_20__15 ;
    output pagesOuts_20__14 ;
    output pagesOuts_20__13 ;
    output pagesOuts_20__12 ;
    output pagesOuts_20__11 ;
    output pagesOuts_20__10 ;
    output pagesOuts_20__9 ;
    output pagesOuts_20__8 ;
    output pagesOuts_20__7 ;
    output pagesOuts_20__6 ;
    output pagesOuts_20__5 ;
    output pagesOuts_20__4 ;
    output pagesOuts_20__3 ;
    output pagesOuts_20__2 ;
    output pagesOuts_20__1 ;
    output pagesOuts_20__0 ;
    output pagesOuts_21__15 ;
    output pagesOuts_21__14 ;
    output pagesOuts_21__13 ;
    output pagesOuts_21__12 ;
    output pagesOuts_21__11 ;
    output pagesOuts_21__10 ;
    output pagesOuts_21__9 ;
    output pagesOuts_21__8 ;
    output pagesOuts_21__7 ;
    output pagesOuts_21__6 ;
    output pagesOuts_21__5 ;
    output pagesOuts_21__4 ;
    output pagesOuts_21__3 ;
    output pagesOuts_21__2 ;
    output pagesOuts_21__1 ;
    output pagesOuts_21__0 ;
    output pagesOuts_22__15 ;
    output pagesOuts_22__14 ;
    output pagesOuts_22__13 ;
    output pagesOuts_22__12 ;
    output pagesOuts_22__11 ;
    output pagesOuts_22__10 ;
    output pagesOuts_22__9 ;
    output pagesOuts_22__8 ;
    output pagesOuts_22__7 ;
    output pagesOuts_22__6 ;
    output pagesOuts_22__5 ;
    output pagesOuts_22__4 ;
    output pagesOuts_22__3 ;
    output pagesOuts_22__2 ;
    output pagesOuts_22__1 ;
    output pagesOuts_22__0 ;
    output pagesOuts_23__15 ;
    output pagesOuts_23__14 ;
    output pagesOuts_23__13 ;
    output pagesOuts_23__12 ;
    output pagesOuts_23__11 ;
    output pagesOuts_23__10 ;
    output pagesOuts_23__9 ;
    output pagesOuts_23__8 ;
    output pagesOuts_23__7 ;
    output pagesOuts_23__6 ;
    output pagesOuts_23__5 ;
    output pagesOuts_23__4 ;
    output pagesOuts_23__3 ;
    output pagesOuts_23__2 ;
    output pagesOuts_23__1 ;
    output pagesOuts_23__0 ;
    output pagesOuts_24__15 ;
    output pagesOuts_24__14 ;
    output pagesOuts_24__13 ;
    output pagesOuts_24__12 ;
    output pagesOuts_24__11 ;
    output pagesOuts_24__10 ;
    output pagesOuts_24__9 ;
    output pagesOuts_24__8 ;
    output pagesOuts_24__7 ;
    output pagesOuts_24__6 ;
    output pagesOuts_24__5 ;
    output pagesOuts_24__4 ;
    output pagesOuts_24__3 ;
    output pagesOuts_24__2 ;
    output pagesOuts_24__1 ;
    output pagesOuts_24__0 ;
    output filtersOuts_0__7 ;
    output filtersOuts_0__6 ;
    output filtersOuts_0__5 ;
    output filtersOuts_0__4 ;
    output filtersOuts_0__3 ;
    output filtersOuts_0__2 ;
    output filtersOuts_0__1 ;
    output filtersOuts_0__0 ;
    output filtersOuts_1__7 ;
    output filtersOuts_1__6 ;
    output filtersOuts_1__5 ;
    output filtersOuts_1__4 ;
    output filtersOuts_1__3 ;
    output filtersOuts_1__2 ;
    output filtersOuts_1__1 ;
    output filtersOuts_1__0 ;
    output filtersOuts_2__7 ;
    output filtersOuts_2__6 ;
    output filtersOuts_2__5 ;
    output filtersOuts_2__4 ;
    output filtersOuts_2__3 ;
    output filtersOuts_2__2 ;
    output filtersOuts_2__1 ;
    output filtersOuts_2__0 ;
    output filtersOuts_3__7 ;
    output filtersOuts_3__6 ;
    output filtersOuts_3__5 ;
    output filtersOuts_3__4 ;
    output filtersOuts_3__3 ;
    output filtersOuts_3__2 ;
    output filtersOuts_3__1 ;
    output filtersOuts_3__0 ;
    output filtersOuts_4__7 ;
    output filtersOuts_4__6 ;
    output filtersOuts_4__5 ;
    output filtersOuts_4__4 ;
    output filtersOuts_4__3 ;
    output filtersOuts_4__2 ;
    output filtersOuts_4__1 ;
    output filtersOuts_4__0 ;
    output filtersOuts_5__7 ;
    output filtersOuts_5__6 ;
    output filtersOuts_5__5 ;
    output filtersOuts_5__4 ;
    output filtersOuts_5__3 ;
    output filtersOuts_5__2 ;
    output filtersOuts_5__1 ;
    output filtersOuts_5__0 ;
    output filtersOuts_6__7 ;
    output filtersOuts_6__6 ;
    output filtersOuts_6__5 ;
    output filtersOuts_6__4 ;
    output filtersOuts_6__3 ;
    output filtersOuts_6__2 ;
    output filtersOuts_6__1 ;
    output filtersOuts_6__0 ;
    output filtersOuts_7__7 ;
    output filtersOuts_7__6 ;
    output filtersOuts_7__5 ;
    output filtersOuts_7__4 ;
    output filtersOuts_7__3 ;
    output filtersOuts_7__2 ;
    output filtersOuts_7__1 ;
    output filtersOuts_7__0 ;
    output filtersOuts_8__7 ;
    output filtersOuts_8__6 ;
    output filtersOuts_8__5 ;
    output filtersOuts_8__4 ;
    output filtersOuts_8__3 ;
    output filtersOuts_8__2 ;
    output filtersOuts_8__1 ;
    output filtersOuts_8__0 ;
    output filtersOuts_9__7 ;
    output filtersOuts_9__6 ;
    output filtersOuts_9__5 ;
    output filtersOuts_9__4 ;
    output filtersOuts_9__3 ;
    output filtersOuts_9__2 ;
    output filtersOuts_9__1 ;
    output filtersOuts_9__0 ;
    output filtersOuts_10__7 ;
    output filtersOuts_10__6 ;
    output filtersOuts_10__5 ;
    output filtersOuts_10__4 ;
    output filtersOuts_10__3 ;
    output filtersOuts_10__2 ;
    output filtersOuts_10__1 ;
    output filtersOuts_10__0 ;
    output filtersOuts_11__7 ;
    output filtersOuts_11__6 ;
    output filtersOuts_11__5 ;
    output filtersOuts_11__4 ;
    output filtersOuts_11__3 ;
    output filtersOuts_11__2 ;
    output filtersOuts_11__1 ;
    output filtersOuts_11__0 ;
    output filtersOuts_12__7 ;
    output filtersOuts_12__6 ;
    output filtersOuts_12__5 ;
    output filtersOuts_12__4 ;
    output filtersOuts_12__3 ;
    output filtersOuts_12__2 ;
    output filtersOuts_12__1 ;
    output filtersOuts_12__0 ;
    output filtersOuts_13__7 ;
    output filtersOuts_13__6 ;
    output filtersOuts_13__5 ;
    output filtersOuts_13__4 ;
    output filtersOuts_13__3 ;
    output filtersOuts_13__2 ;
    output filtersOuts_13__1 ;
    output filtersOuts_13__0 ;
    output filtersOuts_14__7 ;
    output filtersOuts_14__6 ;
    output filtersOuts_14__5 ;
    output filtersOuts_14__4 ;
    output filtersOuts_14__3 ;
    output filtersOuts_14__2 ;
    output filtersOuts_14__1 ;
    output filtersOuts_14__0 ;
    output filtersOuts_15__7 ;
    output filtersOuts_15__6 ;
    output filtersOuts_15__5 ;
    output filtersOuts_15__4 ;
    output filtersOuts_15__3 ;
    output filtersOuts_15__2 ;
    output filtersOuts_15__1 ;
    output filtersOuts_15__0 ;
    output filtersOuts_16__7 ;
    output filtersOuts_16__6 ;
    output filtersOuts_16__5 ;
    output filtersOuts_16__4 ;
    output filtersOuts_16__3 ;
    output filtersOuts_16__2 ;
    output filtersOuts_16__1 ;
    output filtersOuts_16__0 ;
    output filtersOuts_17__7 ;
    output filtersOuts_17__6 ;
    output filtersOuts_17__5 ;
    output filtersOuts_17__4 ;
    output filtersOuts_17__3 ;
    output filtersOuts_17__2 ;
    output filtersOuts_17__1 ;
    output filtersOuts_17__0 ;
    output filtersOuts_18__7 ;
    output filtersOuts_18__6 ;
    output filtersOuts_18__5 ;
    output filtersOuts_18__4 ;
    output filtersOuts_18__3 ;
    output filtersOuts_18__2 ;
    output filtersOuts_18__1 ;
    output filtersOuts_18__0 ;
    output filtersOuts_19__7 ;
    output filtersOuts_19__6 ;
    output filtersOuts_19__5 ;
    output filtersOuts_19__4 ;
    output filtersOuts_19__3 ;
    output filtersOuts_19__2 ;
    output filtersOuts_19__1 ;
    output filtersOuts_19__0 ;
    output filtersOuts_20__7 ;
    output filtersOuts_20__6 ;
    output filtersOuts_20__5 ;
    output filtersOuts_20__4 ;
    output filtersOuts_20__3 ;
    output filtersOuts_20__2 ;
    output filtersOuts_20__1 ;
    output filtersOuts_20__0 ;
    output filtersOuts_21__7 ;
    output filtersOuts_21__6 ;
    output filtersOuts_21__5 ;
    output filtersOuts_21__4 ;
    output filtersOuts_21__3 ;
    output filtersOuts_21__2 ;
    output filtersOuts_21__1 ;
    output filtersOuts_21__0 ;
    output filtersOuts_22__7 ;
    output filtersOuts_22__6 ;
    output filtersOuts_22__5 ;
    output filtersOuts_22__4 ;
    output filtersOuts_22__3 ;
    output filtersOuts_22__2 ;
    output filtersOuts_22__1 ;
    output filtersOuts_22__0 ;
    output filtersOuts_23__7 ;
    output filtersOuts_23__6 ;
    output filtersOuts_23__5 ;
    output filtersOuts_23__4 ;
    output filtersOuts_23__3 ;
    output filtersOuts_23__2 ;
    output filtersOuts_23__1 ;
    output filtersOuts_23__0 ;
    output filtersOuts_24__7 ;
    output filtersOuts_24__6 ;
    output filtersOuts_24__5 ;
    output filtersOuts_24__4 ;
    output filtersOuts_24__3 ;
    output filtersOuts_24__2 ;
    output filtersOuts_24__1 ;
    output filtersOuts_24__0 ;

    wire page1Out_5__15, page1Out_5__14, page1Out_5__13, page1Out_5__12, 
         page1Out_5__11, page1Out_5__10, page1Out_5__9, page1Out_5__8, 
         page1Out_5__7, page1Out_5__6, page1Out_5__5, page1Out_5__4, 
         page1Out_5__3, page1Out_5__2, page1Out_5__1, page1Out_5__0, 
         page1Out_6__15, page1Out_6__14, page1Out_6__13, page1Out_6__12, 
         page1Out_6__11, page1Out_6__10, page1Out_6__9, page1Out_6__8, 
         page1Out_6__7, page1Out_6__6, page1Out_6__5, page1Out_6__4, 
         page1Out_6__3, page1Out_6__2, page1Out_6__1, page1Out_6__0, 
         page1Out_7__15, page1Out_7__14, page1Out_7__13, page1Out_7__12, 
         page1Out_7__11, page1Out_7__10, page1Out_7__9, page1Out_7__8, 
         page1Out_7__7, page1Out_7__6, page1Out_7__5, page1Out_7__4, 
         page1Out_7__3, page1Out_7__2, page1Out_7__1, page1Out_7__0, 
         page1Out_8__15, page1Out_8__14, page1Out_8__13, page1Out_8__12, 
         page1Out_8__11, page1Out_8__10, page1Out_8__9, page1Out_8__8, 
         page1Out_8__7, page1Out_8__6, page1Out_8__5, page1Out_8__4, 
         page1Out_8__3, page1Out_8__2, page1Out_8__1, page1Out_8__0, 
         page1Out_9__15, page1Out_9__14, page1Out_9__13, page1Out_9__12, 
         page1Out_9__11, page1Out_9__10, page1Out_9__9, page1Out_9__8, 
         page1Out_9__7, page1Out_9__6, page1Out_9__5, page1Out_9__4, 
         page1Out_9__3, page1Out_9__2, page1Out_9__1, page1Out_9__0, 
         page1Out_10__15, page1Out_10__14, page1Out_10__13, page1Out_10__12, 
         page1Out_10__11, page1Out_10__10, page1Out_10__9, page1Out_10__8, 
         page1Out_10__7, page1Out_10__6, page1Out_10__5, page1Out_10__4, 
         page1Out_10__3, page1Out_10__2, page1Out_10__1, page1Out_10__0, 
         page1Out_11__15, page1Out_11__14, page1Out_11__13, page1Out_11__12, 
         page1Out_11__11, page1Out_11__10, page1Out_11__9, page1Out_11__8, 
         page1Out_11__7, page1Out_11__6, page1Out_11__5, page1Out_11__4, 
         page1Out_11__3, page1Out_11__2, page1Out_11__1, page1Out_11__0, 
         page1Out_12__15, page1Out_12__14, page1Out_12__13, page1Out_12__12, 
         page1Out_12__11, page1Out_12__10, page1Out_12__9, page1Out_12__8, 
         page1Out_12__7, page1Out_12__6, page1Out_12__5, page1Out_12__4, 
         page1Out_12__3, page1Out_12__2, page1Out_12__1, page1Out_12__0, 
         page1Out_13__15, page1Out_13__14, page1Out_13__13, page1Out_13__12, 
         page1Out_13__11, page1Out_13__10, page1Out_13__9, page1Out_13__8, 
         page1Out_13__7, page1Out_13__6, page1Out_13__5, page1Out_13__4, 
         page1Out_13__3, page1Out_13__2, page1Out_13__1, page1Out_13__0, 
         page1Out_14__15, page1Out_14__14, page1Out_14__13, page1Out_14__12, 
         page1Out_14__11, page1Out_14__10, page1Out_14__9, page1Out_14__8, 
         page1Out_14__7, page1Out_14__6, page1Out_14__5, page1Out_14__4, 
         page1Out_14__3, page1Out_14__2, page1Out_14__1, page1Out_14__0, 
         page1Out_15__15, page1Out_15__14, page1Out_15__13, page1Out_15__12, 
         page1Out_15__11, page1Out_15__10, page1Out_15__9, page1Out_15__8, 
         page1Out_15__7, page1Out_15__6, page1Out_15__5, page1Out_15__4, 
         page1Out_15__3, page1Out_15__2, page1Out_15__1, page1Out_15__0, 
         page1Out_16__15, page1Out_16__14, page1Out_16__13, page1Out_16__12, 
         page1Out_16__11, page1Out_16__10, page1Out_16__9, page1Out_16__8, 
         page1Out_16__7, page1Out_16__6, page1Out_16__5, page1Out_16__4, 
         page1Out_16__3, page1Out_16__2, page1Out_16__1, page1Out_16__0, 
         page1Out_17__15, page1Out_17__14, page1Out_17__13, page1Out_17__12, 
         page1Out_17__11, page1Out_17__10, page1Out_17__9, page1Out_17__8, 
         page1Out_17__7, page1Out_17__6, page1Out_17__5, page1Out_17__4, 
         page1Out_17__3, page1Out_17__2, page1Out_17__1, page1Out_17__0, 
         page1Out_18__15, page1Out_18__14, page1Out_18__13, page1Out_18__12, 
         page1Out_18__11, page1Out_18__10, page1Out_18__9, page1Out_18__8, 
         page1Out_18__7, page1Out_18__6, page1Out_18__5, page1Out_18__4, 
         page1Out_18__3, page1Out_18__2, page1Out_18__1, page1Out_18__0, 
         page1Out_19__15, page1Out_19__14, page1Out_19__13, page1Out_19__12, 
         page1Out_19__11, page1Out_19__10, page1Out_19__9, page1Out_19__8, 
         page1Out_19__7, page1Out_19__6, page1Out_19__5, page1Out_19__4, 
         page1Out_19__3, page1Out_19__2, page1Out_19__1, page1Out_19__0, 
         page1Out_20__15, page1Out_20__14, page1Out_20__13, page1Out_20__12, 
         page1Out_20__11, page1Out_20__10, page1Out_20__9, page1Out_20__8, 
         page1Out_20__7, page1Out_20__6, page1Out_20__5, page1Out_20__4, 
         page1Out_20__3, page1Out_20__2, page1Out_20__1, page1Out_20__0, 
         page1Out_21__15, page1Out_21__14, page1Out_21__13, page1Out_21__12, 
         page1Out_21__11, page1Out_21__10, page1Out_21__9, page1Out_21__8, 
         page1Out_21__7, page1Out_21__6, page1Out_21__5, page1Out_21__4, 
         page1Out_21__3, page1Out_21__2, page1Out_21__1, page1Out_21__0, 
         page1Out_22__15, page1Out_22__14, page1Out_22__13, page1Out_22__12, 
         page1Out_22__11, page1Out_22__10, page1Out_22__9, page1Out_22__8, 
         page1Out_22__7, page1Out_22__6, page1Out_22__5, page1Out_22__4, 
         page1Out_22__3, page1Out_22__2, page1Out_22__1, page1Out_22__0, 
         page1Out_23__15, page1Out_23__14, page1Out_23__13, page1Out_23__12, 
         page1Out_23__11, page1Out_23__10, page1Out_23__9, page1Out_23__8, 
         page1Out_23__7, page1Out_23__6, page1Out_23__5, page1Out_23__4, 
         page1Out_23__3, page1Out_23__2, page1Out_23__1, page1Out_23__0, 
         page1Out_24__15, page1Out_24__14, page1Out_24__13, page1Out_24__12, 
         page1Out_24__11, page1Out_24__10, page1Out_24__9, page1Out_24__8, 
         page1Out_24__7, page1Out_24__6, page1Out_24__5, page1Out_24__4, 
         page1Out_24__3, page1Out_24__2, page1Out_24__1, page1Out_24__0, 
         page2Out_5__15, page2Out_5__14, page2Out_5__13, page2Out_5__12, 
         page2Out_5__11, page2Out_5__10, page2Out_5__9, page2Out_5__8, 
         page2Out_5__7, page2Out_5__6, page2Out_5__5, page2Out_5__4, 
         page2Out_5__3, page2Out_5__2, page2Out_5__1, page2Out_5__0, 
         page2Out_6__15, page2Out_6__14, page2Out_6__13, page2Out_6__12, 
         page2Out_6__11, page2Out_6__10, page2Out_6__9, page2Out_6__8, 
         page2Out_6__7, page2Out_6__6, page2Out_6__5, page2Out_6__4, 
         page2Out_6__3, page2Out_6__2, page2Out_6__1, page2Out_6__0, 
         page2Out_7__15, page2Out_7__14, page2Out_7__13, page2Out_7__12, 
         page2Out_7__11, page2Out_7__10, page2Out_7__9, page2Out_7__8, 
         page2Out_7__7, page2Out_7__6, page2Out_7__5, page2Out_7__4, 
         page2Out_7__3, page2Out_7__2, page2Out_7__1, page2Out_7__0, 
         page2Out_8__15, page2Out_8__14, page2Out_8__13, page2Out_8__12, 
         page2Out_8__11, page2Out_8__10, page2Out_8__9, page2Out_8__8, 
         page2Out_8__7, page2Out_8__6, page2Out_8__5, page2Out_8__4, 
         page2Out_8__3, page2Out_8__2, page2Out_8__1, page2Out_8__0, 
         page2Out_9__15, page2Out_9__14, page2Out_9__13, page2Out_9__12, 
         page2Out_9__11, page2Out_9__10, page2Out_9__9, page2Out_9__8, 
         page2Out_9__7, page2Out_9__6, page2Out_9__5, page2Out_9__4, 
         page2Out_9__3, page2Out_9__2, page2Out_9__1, page2Out_9__0, 
         page2Out_10__15, page2Out_10__14, page2Out_10__13, page2Out_10__12, 
         page2Out_10__11, page2Out_10__10, page2Out_10__9, page2Out_10__8, 
         page2Out_10__7, page2Out_10__6, page2Out_10__5, page2Out_10__4, 
         page2Out_10__3, page2Out_10__2, page2Out_10__1, page2Out_10__0, 
         page2Out_11__15, page2Out_11__14, page2Out_11__13, page2Out_11__12, 
         page2Out_11__11, page2Out_11__10, page2Out_11__9, page2Out_11__8, 
         page2Out_11__7, page2Out_11__6, page2Out_11__5, page2Out_11__4, 
         page2Out_11__3, page2Out_11__2, page2Out_11__1, page2Out_11__0, 
         page2Out_12__15, page2Out_12__14, page2Out_12__13, page2Out_12__12, 
         page2Out_12__11, page2Out_12__10, page2Out_12__9, page2Out_12__8, 
         page2Out_12__7, page2Out_12__6, page2Out_12__5, page2Out_12__4, 
         page2Out_12__3, page2Out_12__2, page2Out_12__1, page2Out_12__0, 
         page2Out_13__15, page2Out_13__14, page2Out_13__13, page2Out_13__12, 
         page2Out_13__11, page2Out_13__10, page2Out_13__9, page2Out_13__8, 
         page2Out_13__7, page2Out_13__6, page2Out_13__5, page2Out_13__4, 
         page2Out_13__3, page2Out_13__2, page2Out_13__1, page2Out_13__0, 
         page2Out_14__15, page2Out_14__14, page2Out_14__13, page2Out_14__12, 
         page2Out_14__11, page2Out_14__10, page2Out_14__9, page2Out_14__8, 
         page2Out_14__7, page2Out_14__6, page2Out_14__5, page2Out_14__4, 
         page2Out_14__3, page2Out_14__2, page2Out_14__1, page2Out_14__0, 
         page2Out_15__15, page2Out_15__14, page2Out_15__13, page2Out_15__12, 
         page2Out_15__11, page2Out_15__10, page2Out_15__9, page2Out_15__8, 
         page2Out_15__7, page2Out_15__6, page2Out_15__5, page2Out_15__4, 
         page2Out_15__3, page2Out_15__2, page2Out_15__1, page2Out_15__0, 
         page2Out_16__15, page2Out_16__14, page2Out_16__13, page2Out_16__12, 
         page2Out_16__11, page2Out_16__10, page2Out_16__9, page2Out_16__8, 
         page2Out_16__7, page2Out_16__6, page2Out_16__5, page2Out_16__4, 
         page2Out_16__3, page2Out_16__2, page2Out_16__1, page2Out_16__0, 
         page2Out_17__15, page2Out_17__14, page2Out_17__13, page2Out_17__12, 
         page2Out_17__11, page2Out_17__10, page2Out_17__9, page2Out_17__8, 
         page2Out_17__7, page2Out_17__6, page2Out_17__5, page2Out_17__4, 
         page2Out_17__3, page2Out_17__2, page2Out_17__1, page2Out_17__0, 
         page2Out_18__15, page2Out_18__14, page2Out_18__13, page2Out_18__12, 
         page2Out_18__11, page2Out_18__10, page2Out_18__9, page2Out_18__8, 
         page2Out_18__7, page2Out_18__6, page2Out_18__5, page2Out_18__4, 
         page2Out_18__3, page2Out_18__2, page2Out_18__1, page2Out_18__0, 
         page2Out_19__15, page2Out_19__14, page2Out_19__13, page2Out_19__12, 
         page2Out_19__11, page2Out_19__10, page2Out_19__9, page2Out_19__8, 
         page2Out_19__7, page2Out_19__6, page2Out_19__5, page2Out_19__4, 
         page2Out_19__3, page2Out_19__2, page2Out_19__1, page2Out_19__0, 
         page2Out_20__15, page2Out_20__14, page2Out_20__13, page2Out_20__12, 
         page2Out_20__11, page2Out_20__10, page2Out_20__9, page2Out_20__8, 
         page2Out_20__7, page2Out_20__6, page2Out_20__5, page2Out_20__4, 
         page2Out_20__3, page2Out_20__2, page2Out_20__1, page2Out_20__0, 
         page2Out_21__15, page2Out_21__14, page2Out_21__13, page2Out_21__12, 
         page2Out_21__11, page2Out_21__10, page2Out_21__9, page2Out_21__8, 
         page2Out_21__7, page2Out_21__6, page2Out_21__5, page2Out_21__4, 
         page2Out_21__3, page2Out_21__2, page2Out_21__1, page2Out_21__0, 
         page2Out_22__15, page2Out_22__14, page2Out_22__13, page2Out_22__12, 
         page2Out_22__11, page2Out_22__10, page2Out_22__9, page2Out_22__8, 
         page2Out_22__7, page2Out_22__6, page2Out_22__5, page2Out_22__4, 
         page2Out_22__3, page2Out_22__2, page2Out_22__1, page2Out_22__0, 
         page2Out_23__15, page2Out_23__14, page2Out_23__13, page2Out_23__12, 
         page2Out_23__11, page2Out_23__10, page2Out_23__9, page2Out_23__8, 
         page2Out_23__7, page2Out_23__6, page2Out_23__5, page2Out_23__4, 
         page2Out_23__3, page2Out_23__2, page2Out_23__1, page2Out_23__0, 
         page2Out_24__15, page2Out_24__14, page2Out_24__13, page2Out_24__12, 
         page2Out_24__11, page2Out_24__10, page2Out_24__9, page2Out_24__8, 
         page2Out_24__7, page2Out_24__6, page2Out_24__5, page2Out_24__4, 
         page2Out_24__3, page2Out_24__2, page2Out_24__1, page2Out_24__0, 
         page1Enables_0, page1Enables_1, page1Enables_2, page1Enables_3, 
         page1Enables_4, page2Enables_0, page2Enables_1, page2Enables_2, 
         page2Enables_3, page2Enables_4, filterEnables_0, filterEnables_1, 
         filterEnables_2, filterEnables_3, page1Out_25__15, nx4, nx62, nx3429, 
         nx3433, nx3435, nx3438, nx3440, nx3443, nx3445, nx3448, nx3452, nx3455, 
         nx3461, nx3464, nx3478, nx3480, nx3482, nx3484, nx3486, nx3488, nx3490, 
         nx3492, nx3494, nx3496;
    wire [159:0] \$dummy ;




    RegUnit_8_16 loop1_0_regRowMap_loop1_0_regUnitMap (.filterBus ({filterBus[7]
                 ,filterBus[6],filterBus[5],filterBus[4],filterBus[3],
                 filterBus[2],filterBus[1],filterBus[0]}), .windowBus ({
                 windowBus[15],windowBus[14],windowBus[13],windowBus[12],
                 windowBus[11],windowBus[10],windowBus[9],windowBus[8],
                 windowBus[7],windowBus[6],windowBus[5],windowBus[4],
                 windowBus[3],windowBus[2],windowBus[1],windowBus[0]}), .regPage1NextUnit (
                 {page1Out_5__15,page1Out_5__14,page1Out_5__13,page1Out_5__12,
                 page1Out_5__11,page1Out_5__10,page1Out_5__9,page1Out_5__8,
                 page1Out_5__7,page1Out_5__6,page1Out_5__5,page1Out_5__4,
                 page1Out_5__3,page1Out_5__2,page1Out_5__1,page1Out_5__0}), .regPage2NextUnit (
                 {page2Out_5__15,page2Out_5__14,page2Out_5__13,page2Out_5__12,
                 page2Out_5__11,page2Out_5__10,page2Out_5__9,page2Out_5__8,
                 page2Out_5__7,page2Out_5__6,page2Out_5__5,page2Out_5__4,
                 page2Out_5__3,page2Out_5__2,page2Out_5__1,page2Out_5__0}), .clk (
                 clk), .rst (rst), .enableRegPage1 (page1Enables_0), .enableRegPage2 (
                 page2Enables_0), .enableRegFilter (nx3478), .page1ReadBusOrPage2 (
                 shift2To1), .page2ReadBusOrPage1 (shift1To2), .pageTurn (
                 pageTurn), .outRegPage ({pagesOuts_0__15,pagesOuts_0__14,
                 pagesOuts_0__13,pagesOuts_0__12,pagesOuts_0__11,pagesOuts_0__10
                 ,pagesOuts_0__9,pagesOuts_0__8,pagesOuts_0__7,pagesOuts_0__6,
                 pagesOuts_0__5,pagesOuts_0__4,pagesOuts_0__3,pagesOuts_0__2,
                 pagesOuts_0__1,pagesOuts_0__0}), .outputRegPage1 ({\$dummy [0],
                 \$dummy [1],\$dummy [2],\$dummy [3],\$dummy [4],\$dummy [5],
                 \$dummy [6],\$dummy [7],\$dummy [8],\$dummy [9],\$dummy [10],
                 \$dummy [11],\$dummy [12],\$dummy [13],\$dummy [14],
                 \$dummy [15]}), .outputRegPage2 ({\$dummy [16],\$dummy [17],
                 \$dummy [18],\$dummy [19],\$dummy [20],\$dummy [21],
                 \$dummy [22],\$dummy [23],\$dummy [24],\$dummy [25],
                 \$dummy [26],\$dummy [27],\$dummy [28],\$dummy [29],
                 \$dummy [30],\$dummy [31]}), .outFilter ({filtersOuts_0__7,
                 filtersOuts_0__6,filtersOuts_0__5,filtersOuts_0__4,
                 filtersOuts_0__3,filtersOuts_0__2,filtersOuts_0__1,
                 filtersOuts_0__0})) ;
    RegUnit_8_16 loop1_0_regRowMap_loop1_1_regUnitMap (.filterBus ({
                 filterBus[15],filterBus[14],filterBus[13],filterBus[12],
                 filterBus[11],filterBus[10],filterBus[9],filterBus[8]}), .windowBus (
                 {windowBus[31],windowBus[30],windowBus[29],windowBus[28],
                 windowBus[27],windowBus[26],windowBus[25],windowBus[24],
                 windowBus[23],windowBus[22],windowBus[21],windowBus[20],
                 windowBus[19],windowBus[18],windowBus[17],windowBus[16]}), .regPage1NextUnit (
                 {page1Out_6__15,page1Out_6__14,page1Out_6__13,page1Out_6__12,
                 page1Out_6__11,page1Out_6__10,page1Out_6__9,page1Out_6__8,
                 page1Out_6__7,page1Out_6__6,page1Out_6__5,page1Out_6__4,
                 page1Out_6__3,page1Out_6__2,page1Out_6__1,page1Out_6__0}), .regPage2NextUnit (
                 {page2Out_6__15,page2Out_6__14,page2Out_6__13,page2Out_6__12,
                 page2Out_6__11,page2Out_6__10,page2Out_6__9,page2Out_6__8,
                 page2Out_6__7,page2Out_6__6,page2Out_6__5,page2Out_6__4,
                 page2Out_6__3,page2Out_6__2,page2Out_6__1,page2Out_6__0}), .clk (
                 clk), .rst (rst), .enableRegPage1 (page1Enables_0), .enableRegPage2 (
                 page2Enables_0), .enableRegFilter (nx3478), .page1ReadBusOrPage2 (
                 shift2To1), .page2ReadBusOrPage1 (shift1To2), .pageTurn (
                 pageTurn), .outRegPage ({pagesOuts_1__15,pagesOuts_1__14,
                 pagesOuts_1__13,pagesOuts_1__12,pagesOuts_1__11,pagesOuts_1__10
                 ,pagesOuts_1__9,pagesOuts_1__8,pagesOuts_1__7,pagesOuts_1__6,
                 pagesOuts_1__5,pagesOuts_1__4,pagesOuts_1__3,pagesOuts_1__2,
                 pagesOuts_1__1,pagesOuts_1__0}), .outputRegPage1 ({\$dummy [32]
                 ,\$dummy [33],\$dummy [34],\$dummy [35],\$dummy [36],
                 \$dummy [37],\$dummy [38],\$dummy [39],\$dummy [40],
                 \$dummy [41],\$dummy [42],\$dummy [43],\$dummy [44],
                 \$dummy [45],\$dummy [46],\$dummy [47]}), .outputRegPage2 ({
                 \$dummy [48],\$dummy [49],\$dummy [50],\$dummy [51],
                 \$dummy [52],\$dummy [53],\$dummy [54],\$dummy [55],
                 \$dummy [56],\$dummy [57],\$dummy [58],\$dummy [59],
                 \$dummy [60],\$dummy [61],\$dummy [62],\$dummy [63]}), .outFilter (
                 {filtersOuts_1__7,filtersOuts_1__6,filtersOuts_1__5,
                 filtersOuts_1__4,filtersOuts_1__3,filtersOuts_1__2,
                 filtersOuts_1__1,filtersOuts_1__0})) ;
    RegUnit_8_16 loop1_0_regRowMap_loop1_2_regUnitMap (.filterBus ({
                 filterBus[23],filterBus[22],filterBus[21],filterBus[20],
                 filterBus[19],filterBus[18],filterBus[17],filterBus[16]}), .windowBus (
                 {windowBus[47],windowBus[46],windowBus[45],windowBus[44],
                 windowBus[43],windowBus[42],windowBus[41],windowBus[40],
                 windowBus[39],windowBus[38],windowBus[37],windowBus[36],
                 windowBus[35],windowBus[34],windowBus[33],windowBus[32]}), .regPage1NextUnit (
                 {page1Out_7__15,page1Out_7__14,page1Out_7__13,page1Out_7__12,
                 page1Out_7__11,page1Out_7__10,page1Out_7__9,page1Out_7__8,
                 page1Out_7__7,page1Out_7__6,page1Out_7__5,page1Out_7__4,
                 page1Out_7__3,page1Out_7__2,page1Out_7__1,page1Out_7__0}), .regPage2NextUnit (
                 {page2Out_7__15,page2Out_7__14,page2Out_7__13,page2Out_7__12,
                 page2Out_7__11,page2Out_7__10,page2Out_7__9,page2Out_7__8,
                 page2Out_7__7,page2Out_7__6,page2Out_7__5,page2Out_7__4,
                 page2Out_7__3,page2Out_7__2,page2Out_7__1,page2Out_7__0}), .clk (
                 clk), .rst (rst), .enableRegPage1 (page1Enables_0), .enableRegPage2 (
                 page2Enables_0), .enableRegFilter (nx3478), .page1ReadBusOrPage2 (
                 shift2To1), .page2ReadBusOrPage1 (shift1To2), .pageTurn (
                 pageTurn), .outRegPage ({pagesOuts_2__15,pagesOuts_2__14,
                 pagesOuts_2__13,pagesOuts_2__12,pagesOuts_2__11,pagesOuts_2__10
                 ,pagesOuts_2__9,pagesOuts_2__8,pagesOuts_2__7,pagesOuts_2__6,
                 pagesOuts_2__5,pagesOuts_2__4,pagesOuts_2__3,pagesOuts_2__2,
                 pagesOuts_2__1,pagesOuts_2__0}), .outputRegPage1 ({\$dummy [64]
                 ,\$dummy [65],\$dummy [66],\$dummy [67],\$dummy [68],
                 \$dummy [69],\$dummy [70],\$dummy [71],\$dummy [72],
                 \$dummy [73],\$dummy [74],\$dummy [75],\$dummy [76],
                 \$dummy [77],\$dummy [78],\$dummy [79]}), .outputRegPage2 ({
                 \$dummy [80],\$dummy [81],\$dummy [82],\$dummy [83],
                 \$dummy [84],\$dummy [85],\$dummy [86],\$dummy [87],
                 \$dummy [88],\$dummy [89],\$dummy [90],\$dummy [91],
                 \$dummy [92],\$dummy [93],\$dummy [94],\$dummy [95]}), .outFilter (
                 {filtersOuts_2__7,filtersOuts_2__6,filtersOuts_2__5,
                 filtersOuts_2__4,filtersOuts_2__3,filtersOuts_2__2,
                 filtersOuts_2__1,filtersOuts_2__0})) ;
    RegUnit_8_16 loop1_0_regRowMap_loop1_3_regUnitMap (.filterBus ({
                 filterBus[31],filterBus[30],filterBus[29],filterBus[28],
                 filterBus[27],filterBus[26],filterBus[25],filterBus[24]}), .windowBus (
                 {windowBus[63],windowBus[62],windowBus[61],windowBus[60],
                 windowBus[59],windowBus[58],windowBus[57],windowBus[56],
                 windowBus[55],windowBus[54],windowBus[53],windowBus[52],
                 windowBus[51],windowBus[50],windowBus[49],windowBus[48]}), .regPage1NextUnit (
                 {page1Out_8__15,page1Out_8__14,page1Out_8__13,page1Out_8__12,
                 page1Out_8__11,page1Out_8__10,page1Out_8__9,page1Out_8__8,
                 page1Out_8__7,page1Out_8__6,page1Out_8__5,page1Out_8__4,
                 page1Out_8__3,page1Out_8__2,page1Out_8__1,page1Out_8__0}), .regPage2NextUnit (
                 {page2Out_8__15,page2Out_8__14,page2Out_8__13,page2Out_8__12,
                 page2Out_8__11,page2Out_8__10,page2Out_8__9,page2Out_8__8,
                 page2Out_8__7,page2Out_8__6,page2Out_8__5,page2Out_8__4,
                 page2Out_8__3,page2Out_8__2,page2Out_8__1,page2Out_8__0}), .clk (
                 clk), .rst (rst), .enableRegPage1 (page1Enables_0), .enableRegPage2 (
                 page2Enables_0), .enableRegFilter (nx3480), .page1ReadBusOrPage2 (
                 shift2To1), .page2ReadBusOrPage1 (shift1To2), .pageTurn (
                 pageTurn), .outRegPage ({pagesOuts_15__15,pagesOuts_15__14,
                 pagesOuts_15__13,pagesOuts_15__12,pagesOuts_15__11,
                 pagesOuts_15__10,pagesOuts_15__9,pagesOuts_15__8,
                 pagesOuts_15__7,pagesOuts_15__6,pagesOuts_15__5,pagesOuts_15__4
                 ,pagesOuts_15__3,pagesOuts_15__2,pagesOuts_15__1,
                 pagesOuts_15__0}), .outputRegPage1 ({\$dummy [96],\$dummy [97],
                 \$dummy [98],\$dummy [99],\$dummy [100],\$dummy [101],
                 \$dummy [102],\$dummy [103],\$dummy [104],\$dummy [105],
                 \$dummy [106],\$dummy [107],\$dummy [108],\$dummy [109],
                 \$dummy [110],\$dummy [111]}), .outputRegPage2 ({\$dummy [112],
                 \$dummy [113],\$dummy [114],\$dummy [115],\$dummy [116],
                 \$dummy [117],\$dummy [118],\$dummy [119],\$dummy [120],
                 \$dummy [121],\$dummy [122],\$dummy [123],\$dummy [124],
                 \$dummy [125],\$dummy [126],\$dummy [127]}), .outFilter ({
                 filtersOuts_15__7,filtersOuts_15__6,filtersOuts_15__5,
                 filtersOuts_15__4,filtersOuts_15__3,filtersOuts_15__2,
                 filtersOuts_15__1,filtersOuts_15__0})) ;
    RegUnit_8_16 loop1_0_regRowMap_loop1_4_regUnitMap (.filterBus ({
                 filterBus[39],filterBus[38],filterBus[37],filterBus[36],
                 filterBus[35],filterBus[34],filterBus[33],filterBus[32]}), .windowBus (
                 {windowBus[79],windowBus[78],windowBus[77],windowBus[76],
                 windowBus[75],windowBus[74],windowBus[73],windowBus[72],
                 windowBus[71],windowBus[70],windowBus[69],windowBus[68],
                 windowBus[67],windowBus[66],windowBus[65],windowBus[64]}), .regPage1NextUnit (
                 {page1Out_9__15,page1Out_9__14,page1Out_9__13,page1Out_9__12,
                 page1Out_9__11,page1Out_9__10,page1Out_9__9,page1Out_9__8,
                 page1Out_9__7,page1Out_9__6,page1Out_9__5,page1Out_9__4,
                 page1Out_9__3,page1Out_9__2,page1Out_9__1,page1Out_9__0}), .regPage2NextUnit (
                 {page2Out_9__15,page2Out_9__14,page2Out_9__13,page2Out_9__12,
                 page2Out_9__11,page2Out_9__10,page2Out_9__9,page2Out_9__8,
                 page2Out_9__7,page2Out_9__6,page2Out_9__5,page2Out_9__4,
                 page2Out_9__3,page2Out_9__2,page2Out_9__1,page2Out_9__0}), .clk (
                 clk), .rst (rst), .enableRegPage1 (page1Enables_0), .enableRegPage2 (
                 page2Enables_0), .enableRegFilter (nx3480), .page1ReadBusOrPage2 (
                 shift2To1), .page2ReadBusOrPage1 (shift1To2), .pageTurn (
                 pageTurn), .outRegPage ({pagesOuts_16__15,pagesOuts_16__14,
                 pagesOuts_16__13,pagesOuts_16__12,pagesOuts_16__11,
                 pagesOuts_16__10,pagesOuts_16__9,pagesOuts_16__8,
                 pagesOuts_16__7,pagesOuts_16__6,pagesOuts_16__5,pagesOuts_16__4
                 ,pagesOuts_16__3,pagesOuts_16__2,pagesOuts_16__1,
                 pagesOuts_16__0}), .outputRegPage1 ({\$dummy [128],
                 \$dummy [129],\$dummy [130],\$dummy [131],\$dummy [132],
                 \$dummy [133],\$dummy [134],\$dummy [135],\$dummy [136],
                 \$dummy [137],\$dummy [138],\$dummy [139],\$dummy [140],
                 \$dummy [141],\$dummy [142],\$dummy [143]}), .outputRegPage2 ({
                 \$dummy [144],\$dummy [145],\$dummy [146],\$dummy [147],
                 \$dummy [148],\$dummy [149],\$dummy [150],\$dummy [151],
                 \$dummy [152],\$dummy [153],\$dummy [154],\$dummy [155],
                 \$dummy [156],\$dummy [157],\$dummy [158],\$dummy [159]}), .outFilter (
                 {filtersOuts_16__7,filtersOuts_16__6,filtersOuts_16__5,
                 filtersOuts_16__4,filtersOuts_16__3,filtersOuts_16__2,
                 filtersOuts_16__1,filtersOuts_16__0})) ;
    RegUnit_8_16_unfolded0 loop1_1_regRowMap_loop1_0_regUnitMap (.filterBus ({
                           filterBus[7],filterBus[6],filterBus[5],filterBus[4],
                           filterBus[3],filterBus[2],filterBus[1],filterBus[0]})
                           , .windowBus ({windowBus[15],windowBus[14],
                           windowBus[13],windowBus[12],windowBus[11],
                           windowBus[10],windowBus[9],windowBus[8],windowBus[7],
                           windowBus[6],windowBus[5],windowBus[4],windowBus[3],
                           windowBus[2],windowBus[1],windowBus[0]}), .regPage1NextUnit (
                           {page1Out_10__15,page1Out_10__14,page1Out_10__13,
                           page1Out_10__12,page1Out_10__11,page1Out_10__10,
                           page1Out_10__9,page1Out_10__8,page1Out_10__7,
                           page1Out_10__6,page1Out_10__5,page1Out_10__4,
                           page1Out_10__3,page1Out_10__2,page1Out_10__1,
                           page1Out_10__0}), .regPage2NextUnit ({page2Out_10__15
                           ,page2Out_10__14,page2Out_10__13,page2Out_10__12,
                           page2Out_10__11,page2Out_10__10,page2Out_10__9,
                           page2Out_10__8,page2Out_10__7,page2Out_10__6,
                           page2Out_10__5,page2Out_10__4,page2Out_10__3,
                           page2Out_10__2,page2Out_10__1,page2Out_10__0}), .clk (
                           clk), .rst (rst), .enableRegPage1 (page1Enables_1), .enableRegPage2 (
                           page2Enables_1), .enableRegFilter (nx3482), .page1ReadBusOrPage2 (
                           shift2To1), .page2ReadBusOrPage1 (shift1To2), .pageTurn (
                           pageTurn), .outRegPage ({pagesOuts_3__15,
                           pagesOuts_3__14,pagesOuts_3__13,pagesOuts_3__12,
                           pagesOuts_3__11,pagesOuts_3__10,pagesOuts_3__9,
                           pagesOuts_3__8,pagesOuts_3__7,pagesOuts_3__6,
                           pagesOuts_3__5,pagesOuts_3__4,pagesOuts_3__3,
                           pagesOuts_3__2,pagesOuts_3__1,pagesOuts_3__0}), .outputRegPage1 (
                           {page1Out_5__15,page1Out_5__14,page1Out_5__13,
                           page1Out_5__12,page1Out_5__11,page1Out_5__10,
                           page1Out_5__9,page1Out_5__8,page1Out_5__7,
                           page1Out_5__6,page1Out_5__5,page1Out_5__4,
                           page1Out_5__3,page1Out_5__2,page1Out_5__1,
                           page1Out_5__0}), .outputRegPage2 ({page2Out_5__15,
                           page2Out_5__14,page2Out_5__13,page2Out_5__12,
                           page2Out_5__11,page2Out_5__10,page2Out_5__9,
                           page2Out_5__8,page2Out_5__7,page2Out_5__6,
                           page2Out_5__5,page2Out_5__4,page2Out_5__3,
                           page2Out_5__2,page2Out_5__1,page2Out_5__0}), .outFilter (
                           {filtersOuts_3__7,filtersOuts_3__6,filtersOuts_3__5,
                           filtersOuts_3__4,filtersOuts_3__3,filtersOuts_3__2,
                           filtersOuts_3__1,filtersOuts_3__0})) ;
    RegUnit_8_16_unfolded0 loop1_1_regRowMap_loop1_1_regUnitMap (.filterBus ({
                           filterBus[15],filterBus[14],filterBus[13],
                           filterBus[12],filterBus[11],filterBus[10],
                           filterBus[9],filterBus[8]}), .windowBus ({
                           windowBus[31],windowBus[30],windowBus[29],
                           windowBus[28],windowBus[27],windowBus[26],
                           windowBus[25],windowBus[24],windowBus[23],
                           windowBus[22],windowBus[21],windowBus[20],
                           windowBus[19],windowBus[18],windowBus[17],
                           windowBus[16]}), .regPage1NextUnit ({page1Out_11__15,
                           page1Out_11__14,page1Out_11__13,page1Out_11__12,
                           page1Out_11__11,page1Out_11__10,page1Out_11__9,
                           page1Out_11__8,page1Out_11__7,page1Out_11__6,
                           page1Out_11__5,page1Out_11__4,page1Out_11__3,
                           page1Out_11__2,page1Out_11__1,page1Out_11__0}), .regPage2NextUnit (
                           {page2Out_11__15,page2Out_11__14,page2Out_11__13,
                           page2Out_11__12,page2Out_11__11,page2Out_11__10,
                           page2Out_11__9,page2Out_11__8,page2Out_11__7,
                           page2Out_11__6,page2Out_11__5,page2Out_11__4,
                           page2Out_11__3,page2Out_11__2,page2Out_11__1,
                           page2Out_11__0}), .clk (clk), .rst (rst), .enableRegPage1 (
                           page1Enables_1), .enableRegPage2 (page2Enables_1), .enableRegFilter (
                           nx3482), .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           pagesOuts_4__15,pagesOuts_4__14,pagesOuts_4__13,
                           pagesOuts_4__12,pagesOuts_4__11,pagesOuts_4__10,
                           pagesOuts_4__9,pagesOuts_4__8,pagesOuts_4__7,
                           pagesOuts_4__6,pagesOuts_4__5,pagesOuts_4__4,
                           pagesOuts_4__3,pagesOuts_4__2,pagesOuts_4__1,
                           pagesOuts_4__0}), .outputRegPage1 ({page1Out_6__15,
                           page1Out_6__14,page1Out_6__13,page1Out_6__12,
                           page1Out_6__11,page1Out_6__10,page1Out_6__9,
                           page1Out_6__8,page1Out_6__7,page1Out_6__6,
                           page1Out_6__5,page1Out_6__4,page1Out_6__3,
                           page1Out_6__2,page1Out_6__1,page1Out_6__0}), .outputRegPage2 (
                           {page2Out_6__15,page2Out_6__14,page2Out_6__13,
                           page2Out_6__12,page2Out_6__11,page2Out_6__10,
                           page2Out_6__9,page2Out_6__8,page2Out_6__7,
                           page2Out_6__6,page2Out_6__5,page2Out_6__4,
                           page2Out_6__3,page2Out_6__2,page2Out_6__1,
                           page2Out_6__0}), .outFilter ({filtersOuts_4__7,
                           filtersOuts_4__6,filtersOuts_4__5,filtersOuts_4__4,
                           filtersOuts_4__3,filtersOuts_4__2,filtersOuts_4__1,
                           filtersOuts_4__0})) ;
    RegUnit_8_16_unfolded0 loop1_1_regRowMap_loop1_2_regUnitMap (.filterBus ({
                           filterBus[23],filterBus[22],filterBus[21],
                           filterBus[20],filterBus[19],filterBus[18],
                           filterBus[17],filterBus[16]}), .windowBus ({
                           windowBus[47],windowBus[46],windowBus[45],
                           windowBus[44],windowBus[43],windowBus[42],
                           windowBus[41],windowBus[40],windowBus[39],
                           windowBus[38],windowBus[37],windowBus[36],
                           windowBus[35],windowBus[34],windowBus[33],
                           windowBus[32]}), .regPage1NextUnit ({page1Out_12__15,
                           page1Out_12__14,page1Out_12__13,page1Out_12__12,
                           page1Out_12__11,page1Out_12__10,page1Out_12__9,
                           page1Out_12__8,page1Out_12__7,page1Out_12__6,
                           page1Out_12__5,page1Out_12__4,page1Out_12__3,
                           page1Out_12__2,page1Out_12__1,page1Out_12__0}), .regPage2NextUnit (
                           {page2Out_12__15,page2Out_12__14,page2Out_12__13,
                           page2Out_12__12,page2Out_12__11,page2Out_12__10,
                           page2Out_12__9,page2Out_12__8,page2Out_12__7,
                           page2Out_12__6,page2Out_12__5,page2Out_12__4,
                           page2Out_12__3,page2Out_12__2,page2Out_12__1,
                           page2Out_12__0}), .clk (clk), .rst (rst), .enableRegPage1 (
                           page1Enables_1), .enableRegPage2 (page2Enables_1), .enableRegFilter (
                           nx3482), .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           pagesOuts_5__15,pagesOuts_5__14,pagesOuts_5__13,
                           pagesOuts_5__12,pagesOuts_5__11,pagesOuts_5__10,
                           pagesOuts_5__9,pagesOuts_5__8,pagesOuts_5__7,
                           pagesOuts_5__6,pagesOuts_5__5,pagesOuts_5__4,
                           pagesOuts_5__3,pagesOuts_5__2,pagesOuts_5__1,
                           pagesOuts_5__0}), .outputRegPage1 ({page1Out_7__15,
                           page1Out_7__14,page1Out_7__13,page1Out_7__12,
                           page1Out_7__11,page1Out_7__10,page1Out_7__9,
                           page1Out_7__8,page1Out_7__7,page1Out_7__6,
                           page1Out_7__5,page1Out_7__4,page1Out_7__3,
                           page1Out_7__2,page1Out_7__1,page1Out_7__0}), .outputRegPage2 (
                           {page2Out_7__15,page2Out_7__14,page2Out_7__13,
                           page2Out_7__12,page2Out_7__11,page2Out_7__10,
                           page2Out_7__9,page2Out_7__8,page2Out_7__7,
                           page2Out_7__6,page2Out_7__5,page2Out_7__4,
                           page2Out_7__3,page2Out_7__2,page2Out_7__1,
                           page2Out_7__0}), .outFilter ({filtersOuts_5__7,
                           filtersOuts_5__6,filtersOuts_5__5,filtersOuts_5__4,
                           filtersOuts_5__3,filtersOuts_5__2,filtersOuts_5__1,
                           filtersOuts_5__0})) ;
    RegUnit_8_16_unfolded0 loop1_1_regRowMap_loop1_3_regUnitMap (.filterBus ({
                           filterBus[31],filterBus[30],filterBus[29],
                           filterBus[28],filterBus[27],filterBus[26],
                           filterBus[25],filterBus[24]}), .windowBus ({
                           windowBus[63],windowBus[62],windowBus[61],
                           windowBus[60],windowBus[59],windowBus[58],
                           windowBus[57],windowBus[56],windowBus[55],
                           windowBus[54],windowBus[53],windowBus[52],
                           windowBus[51],windowBus[50],windowBus[49],
                           windowBus[48]}), .regPage1NextUnit ({page1Out_13__15,
                           page1Out_13__14,page1Out_13__13,page1Out_13__12,
                           page1Out_13__11,page1Out_13__10,page1Out_13__9,
                           page1Out_13__8,page1Out_13__7,page1Out_13__6,
                           page1Out_13__5,page1Out_13__4,page1Out_13__3,
                           page1Out_13__2,page1Out_13__1,page1Out_13__0}), .regPage2NextUnit (
                           {page2Out_13__15,page2Out_13__14,page2Out_13__13,
                           page2Out_13__12,page2Out_13__11,page2Out_13__10,
                           page2Out_13__9,page2Out_13__8,page2Out_13__7,
                           page2Out_13__6,page2Out_13__5,page2Out_13__4,
                           page2Out_13__3,page2Out_13__2,page2Out_13__1,
                           page2Out_13__0}), .clk (clk), .rst (rst), .enableRegPage1 (
                           page1Enables_1), .enableRegPage2 (page2Enables_1), .enableRegFilter (
                           nx3484), .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           pagesOuts_17__15,pagesOuts_17__14,pagesOuts_17__13,
                           pagesOuts_17__12,pagesOuts_17__11,pagesOuts_17__10,
                           pagesOuts_17__9,pagesOuts_17__8,pagesOuts_17__7,
                           pagesOuts_17__6,pagesOuts_17__5,pagesOuts_17__4,
                           pagesOuts_17__3,pagesOuts_17__2,pagesOuts_17__1,
                           pagesOuts_17__0}), .outputRegPage1 ({page1Out_8__15,
                           page1Out_8__14,page1Out_8__13,page1Out_8__12,
                           page1Out_8__11,page1Out_8__10,page1Out_8__9,
                           page1Out_8__8,page1Out_8__7,page1Out_8__6,
                           page1Out_8__5,page1Out_8__4,page1Out_8__3,
                           page1Out_8__2,page1Out_8__1,page1Out_8__0}), .outputRegPage2 (
                           {page2Out_8__15,page2Out_8__14,page2Out_8__13,
                           page2Out_8__12,page2Out_8__11,page2Out_8__10,
                           page2Out_8__9,page2Out_8__8,page2Out_8__7,
                           page2Out_8__6,page2Out_8__5,page2Out_8__4,
                           page2Out_8__3,page2Out_8__2,page2Out_8__1,
                           page2Out_8__0}), .outFilter ({filtersOuts_17__7,
                           filtersOuts_17__6,filtersOuts_17__5,filtersOuts_17__4
                           ,filtersOuts_17__3,filtersOuts_17__2,
                           filtersOuts_17__1,filtersOuts_17__0})) ;
    RegUnit_8_16_unfolded0 loop1_1_regRowMap_loop1_4_regUnitMap (.filterBus ({
                           filterBus[39],filterBus[38],filterBus[37],
                           filterBus[36],filterBus[35],filterBus[34],
                           filterBus[33],filterBus[32]}), .windowBus ({
                           windowBus[79],windowBus[78],windowBus[77],
                           windowBus[76],windowBus[75],windowBus[74],
                           windowBus[73],windowBus[72],windowBus[71],
                           windowBus[70],windowBus[69],windowBus[68],
                           windowBus[67],windowBus[66],windowBus[65],
                           windowBus[64]}), .regPage1NextUnit ({page1Out_14__15,
                           page1Out_14__14,page1Out_14__13,page1Out_14__12,
                           page1Out_14__11,page1Out_14__10,page1Out_14__9,
                           page1Out_14__8,page1Out_14__7,page1Out_14__6,
                           page1Out_14__5,page1Out_14__4,page1Out_14__3,
                           page1Out_14__2,page1Out_14__1,page1Out_14__0}), .regPage2NextUnit (
                           {page2Out_14__15,page2Out_14__14,page2Out_14__13,
                           page2Out_14__12,page2Out_14__11,page2Out_14__10,
                           page2Out_14__9,page2Out_14__8,page2Out_14__7,
                           page2Out_14__6,page2Out_14__5,page2Out_14__4,
                           page2Out_14__3,page2Out_14__2,page2Out_14__1,
                           page2Out_14__0}), .clk (clk), .rst (rst), .enableRegPage1 (
                           page1Enables_1), .enableRegPage2 (page2Enables_1), .enableRegFilter (
                           nx3484), .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           pagesOuts_18__15,pagesOuts_18__14,pagesOuts_18__13,
                           pagesOuts_18__12,pagesOuts_18__11,pagesOuts_18__10,
                           pagesOuts_18__9,pagesOuts_18__8,pagesOuts_18__7,
                           pagesOuts_18__6,pagesOuts_18__5,pagesOuts_18__4,
                           pagesOuts_18__3,pagesOuts_18__2,pagesOuts_18__1,
                           pagesOuts_18__0}), .outputRegPage1 ({page1Out_9__15,
                           page1Out_9__14,page1Out_9__13,page1Out_9__12,
                           page1Out_9__11,page1Out_9__10,page1Out_9__9,
                           page1Out_9__8,page1Out_9__7,page1Out_9__6,
                           page1Out_9__5,page1Out_9__4,page1Out_9__3,
                           page1Out_9__2,page1Out_9__1,page1Out_9__0}), .outputRegPage2 (
                           {page2Out_9__15,page2Out_9__14,page2Out_9__13,
                           page2Out_9__12,page2Out_9__11,page2Out_9__10,
                           page2Out_9__9,page2Out_9__8,page2Out_9__7,
                           page2Out_9__6,page2Out_9__5,page2Out_9__4,
                           page2Out_9__3,page2Out_9__2,page2Out_9__1,
                           page2Out_9__0}), .outFilter ({filtersOuts_18__7,
                           filtersOuts_18__6,filtersOuts_18__5,filtersOuts_18__4
                           ,filtersOuts_18__3,filtersOuts_18__2,
                           filtersOuts_18__1,filtersOuts_18__0})) ;
    RegUnit_8_16_unfolded0 loop1_2_regRowMap_loop1_0_regUnitMap (.filterBus ({
                           filterBus[7],filterBus[6],filterBus[5],filterBus[4],
                           filterBus[3],filterBus[2],filterBus[1],filterBus[0]})
                           , .windowBus ({windowBus[15],windowBus[14],
                           windowBus[13],windowBus[12],windowBus[11],
                           windowBus[10],windowBus[9],windowBus[8],windowBus[7],
                           windowBus[6],windowBus[5],windowBus[4],windowBus[3],
                           windowBus[2],windowBus[1],windowBus[0]}), .regPage1NextUnit (
                           {page1Out_15__15,page1Out_15__14,page1Out_15__13,
                           page1Out_15__12,page1Out_15__11,page1Out_15__10,
                           page1Out_15__9,page1Out_15__8,page1Out_15__7,
                           page1Out_15__6,page1Out_15__5,page1Out_15__4,
                           page1Out_15__3,page1Out_15__2,page1Out_15__1,
                           page1Out_15__0}), .regPage2NextUnit ({page2Out_15__15
                           ,page2Out_15__14,page2Out_15__13,page2Out_15__12,
                           page2Out_15__11,page2Out_15__10,page2Out_15__9,
                           page2Out_15__8,page2Out_15__7,page2Out_15__6,
                           page2Out_15__5,page2Out_15__4,page2Out_15__3,
                           page2Out_15__2,page2Out_15__1,page2Out_15__0}), .clk (
                           clk), .rst (rst), .enableRegPage1 (page1Enables_2), .enableRegPage2 (
                           page2Enables_2), .enableRegFilter (nx3486), .page1ReadBusOrPage2 (
                           shift2To1), .page2ReadBusOrPage1 (shift1To2), .pageTurn (
                           pageTurn), .outRegPage ({pagesOuts_6__15,
                           pagesOuts_6__14,pagesOuts_6__13,pagesOuts_6__12,
                           pagesOuts_6__11,pagesOuts_6__10,pagesOuts_6__9,
                           pagesOuts_6__8,pagesOuts_6__7,pagesOuts_6__6,
                           pagesOuts_6__5,pagesOuts_6__4,pagesOuts_6__3,
                           pagesOuts_6__2,pagesOuts_6__1,pagesOuts_6__0}), .outputRegPage1 (
                           {page1Out_10__15,page1Out_10__14,page1Out_10__13,
                           page1Out_10__12,page1Out_10__11,page1Out_10__10,
                           page1Out_10__9,page1Out_10__8,page1Out_10__7,
                           page1Out_10__6,page1Out_10__5,page1Out_10__4,
                           page1Out_10__3,page1Out_10__2,page1Out_10__1,
                           page1Out_10__0}), .outputRegPage2 ({page2Out_10__15,
                           page2Out_10__14,page2Out_10__13,page2Out_10__12,
                           page2Out_10__11,page2Out_10__10,page2Out_10__9,
                           page2Out_10__8,page2Out_10__7,page2Out_10__6,
                           page2Out_10__5,page2Out_10__4,page2Out_10__3,
                           page2Out_10__2,page2Out_10__1,page2Out_10__0}), .outFilter (
                           {filtersOuts_6__7,filtersOuts_6__6,filtersOuts_6__5,
                           filtersOuts_6__4,filtersOuts_6__3,filtersOuts_6__2,
                           filtersOuts_6__1,filtersOuts_6__0})) ;
    RegUnit_8_16_unfolded0 loop1_2_regRowMap_loop1_1_regUnitMap (.filterBus ({
                           filterBus[15],filterBus[14],filterBus[13],
                           filterBus[12],filterBus[11],filterBus[10],
                           filterBus[9],filterBus[8]}), .windowBus ({
                           windowBus[31],windowBus[30],windowBus[29],
                           windowBus[28],windowBus[27],windowBus[26],
                           windowBus[25],windowBus[24],windowBus[23],
                           windowBus[22],windowBus[21],windowBus[20],
                           windowBus[19],windowBus[18],windowBus[17],
                           windowBus[16]}), .regPage1NextUnit ({page1Out_16__15,
                           page1Out_16__14,page1Out_16__13,page1Out_16__12,
                           page1Out_16__11,page1Out_16__10,page1Out_16__9,
                           page1Out_16__8,page1Out_16__7,page1Out_16__6,
                           page1Out_16__5,page1Out_16__4,page1Out_16__3,
                           page1Out_16__2,page1Out_16__1,page1Out_16__0}), .regPage2NextUnit (
                           {page2Out_16__15,page2Out_16__14,page2Out_16__13,
                           page2Out_16__12,page2Out_16__11,page2Out_16__10,
                           page2Out_16__9,page2Out_16__8,page2Out_16__7,
                           page2Out_16__6,page2Out_16__5,page2Out_16__4,
                           page2Out_16__3,page2Out_16__2,page2Out_16__1,
                           page2Out_16__0}), .clk (clk), .rst (rst), .enableRegPage1 (
                           page1Enables_2), .enableRegPage2 (page2Enables_2), .enableRegFilter (
                           nx3486), .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           pagesOuts_7__15,pagesOuts_7__14,pagesOuts_7__13,
                           pagesOuts_7__12,pagesOuts_7__11,pagesOuts_7__10,
                           pagesOuts_7__9,pagesOuts_7__8,pagesOuts_7__7,
                           pagesOuts_7__6,pagesOuts_7__5,pagesOuts_7__4,
                           pagesOuts_7__3,pagesOuts_7__2,pagesOuts_7__1,
                           pagesOuts_7__0}), .outputRegPage1 ({page1Out_11__15,
                           page1Out_11__14,page1Out_11__13,page1Out_11__12,
                           page1Out_11__11,page1Out_11__10,page1Out_11__9,
                           page1Out_11__8,page1Out_11__7,page1Out_11__6,
                           page1Out_11__5,page1Out_11__4,page1Out_11__3,
                           page1Out_11__2,page1Out_11__1,page1Out_11__0}), .outputRegPage2 (
                           {page2Out_11__15,page2Out_11__14,page2Out_11__13,
                           page2Out_11__12,page2Out_11__11,page2Out_11__10,
                           page2Out_11__9,page2Out_11__8,page2Out_11__7,
                           page2Out_11__6,page2Out_11__5,page2Out_11__4,
                           page2Out_11__3,page2Out_11__2,page2Out_11__1,
                           page2Out_11__0}), .outFilter ({filtersOuts_7__7,
                           filtersOuts_7__6,filtersOuts_7__5,filtersOuts_7__4,
                           filtersOuts_7__3,filtersOuts_7__2,filtersOuts_7__1,
                           filtersOuts_7__0})) ;
    RegUnit_8_16_unfolded0 loop1_2_regRowMap_loop1_2_regUnitMap (.filterBus ({
                           filterBus[23],filterBus[22],filterBus[21],
                           filterBus[20],filterBus[19],filterBus[18],
                           filterBus[17],filterBus[16]}), .windowBus ({
                           windowBus[47],windowBus[46],windowBus[45],
                           windowBus[44],windowBus[43],windowBus[42],
                           windowBus[41],windowBus[40],windowBus[39],
                           windowBus[38],windowBus[37],windowBus[36],
                           windowBus[35],windowBus[34],windowBus[33],
                           windowBus[32]}), .regPage1NextUnit ({page1Out_17__15,
                           page1Out_17__14,page1Out_17__13,page1Out_17__12,
                           page1Out_17__11,page1Out_17__10,page1Out_17__9,
                           page1Out_17__8,page1Out_17__7,page1Out_17__6,
                           page1Out_17__5,page1Out_17__4,page1Out_17__3,
                           page1Out_17__2,page1Out_17__1,page1Out_17__0}), .regPage2NextUnit (
                           {page2Out_17__15,page2Out_17__14,page2Out_17__13,
                           page2Out_17__12,page2Out_17__11,page2Out_17__10,
                           page2Out_17__9,page2Out_17__8,page2Out_17__7,
                           page2Out_17__6,page2Out_17__5,page2Out_17__4,
                           page2Out_17__3,page2Out_17__2,page2Out_17__1,
                           page2Out_17__0}), .clk (clk), .rst (rst), .enableRegPage1 (
                           page1Enables_2), .enableRegPage2 (page2Enables_2), .enableRegFilter (
                           nx3486), .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           pagesOuts_8__15,pagesOuts_8__14,pagesOuts_8__13,
                           pagesOuts_8__12,pagesOuts_8__11,pagesOuts_8__10,
                           pagesOuts_8__9,pagesOuts_8__8,pagesOuts_8__7,
                           pagesOuts_8__6,pagesOuts_8__5,pagesOuts_8__4,
                           pagesOuts_8__3,pagesOuts_8__2,pagesOuts_8__1,
                           pagesOuts_8__0}), .outputRegPage1 ({page1Out_12__15,
                           page1Out_12__14,page1Out_12__13,page1Out_12__12,
                           page1Out_12__11,page1Out_12__10,page1Out_12__9,
                           page1Out_12__8,page1Out_12__7,page1Out_12__6,
                           page1Out_12__5,page1Out_12__4,page1Out_12__3,
                           page1Out_12__2,page1Out_12__1,page1Out_12__0}), .outputRegPage2 (
                           {page2Out_12__15,page2Out_12__14,page2Out_12__13,
                           page2Out_12__12,page2Out_12__11,page2Out_12__10,
                           page2Out_12__9,page2Out_12__8,page2Out_12__7,
                           page2Out_12__6,page2Out_12__5,page2Out_12__4,
                           page2Out_12__3,page2Out_12__2,page2Out_12__1,
                           page2Out_12__0}), .outFilter ({filtersOuts_8__7,
                           filtersOuts_8__6,filtersOuts_8__5,filtersOuts_8__4,
                           filtersOuts_8__3,filtersOuts_8__2,filtersOuts_8__1,
                           filtersOuts_8__0})) ;
    RegUnit_8_16_unfolded0 loop1_2_regRowMap_loop1_3_regUnitMap (.filterBus ({
                           filterBus[31],filterBus[30],filterBus[29],
                           filterBus[28],filterBus[27],filterBus[26],
                           filterBus[25],filterBus[24]}), .windowBus ({
                           windowBus[63],windowBus[62],windowBus[61],
                           windowBus[60],windowBus[59],windowBus[58],
                           windowBus[57],windowBus[56],windowBus[55],
                           windowBus[54],windowBus[53],windowBus[52],
                           windowBus[51],windowBus[50],windowBus[49],
                           windowBus[48]}), .regPage1NextUnit ({page1Out_18__15,
                           page1Out_18__14,page1Out_18__13,page1Out_18__12,
                           page1Out_18__11,page1Out_18__10,page1Out_18__9,
                           page1Out_18__8,page1Out_18__7,page1Out_18__6,
                           page1Out_18__5,page1Out_18__4,page1Out_18__3,
                           page1Out_18__2,page1Out_18__1,page1Out_18__0}), .regPage2NextUnit (
                           {page2Out_18__15,page2Out_18__14,page2Out_18__13,
                           page2Out_18__12,page2Out_18__11,page2Out_18__10,
                           page2Out_18__9,page2Out_18__8,page2Out_18__7,
                           page2Out_18__6,page2Out_18__5,page2Out_18__4,
                           page2Out_18__3,page2Out_18__2,page2Out_18__1,
                           page2Out_18__0}), .clk (clk), .rst (rst), .enableRegPage1 (
                           page1Enables_2), .enableRegPage2 (page2Enables_2), .enableRegFilter (
                           nx3488), .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           pagesOuts_19__15,pagesOuts_19__14,pagesOuts_19__13,
                           pagesOuts_19__12,pagesOuts_19__11,pagesOuts_19__10,
                           pagesOuts_19__9,pagesOuts_19__8,pagesOuts_19__7,
                           pagesOuts_19__6,pagesOuts_19__5,pagesOuts_19__4,
                           pagesOuts_19__3,pagesOuts_19__2,pagesOuts_19__1,
                           pagesOuts_19__0}), .outputRegPage1 ({page1Out_13__15,
                           page1Out_13__14,page1Out_13__13,page1Out_13__12,
                           page1Out_13__11,page1Out_13__10,page1Out_13__9,
                           page1Out_13__8,page1Out_13__7,page1Out_13__6,
                           page1Out_13__5,page1Out_13__4,page1Out_13__3,
                           page1Out_13__2,page1Out_13__1,page1Out_13__0}), .outputRegPage2 (
                           {page2Out_13__15,page2Out_13__14,page2Out_13__13,
                           page2Out_13__12,page2Out_13__11,page2Out_13__10,
                           page2Out_13__9,page2Out_13__8,page2Out_13__7,
                           page2Out_13__6,page2Out_13__5,page2Out_13__4,
                           page2Out_13__3,page2Out_13__2,page2Out_13__1,
                           page2Out_13__0}), .outFilter ({filtersOuts_19__7,
                           filtersOuts_19__6,filtersOuts_19__5,filtersOuts_19__4
                           ,filtersOuts_19__3,filtersOuts_19__2,
                           filtersOuts_19__1,filtersOuts_19__0})) ;
    RegUnit_8_16_unfolded0 loop1_2_regRowMap_loop1_4_regUnitMap (.filterBus ({
                           filterBus[39],filterBus[38],filterBus[37],
                           filterBus[36],filterBus[35],filterBus[34],
                           filterBus[33],filterBus[32]}), .windowBus ({
                           windowBus[79],windowBus[78],windowBus[77],
                           windowBus[76],windowBus[75],windowBus[74],
                           windowBus[73],windowBus[72],windowBus[71],
                           windowBus[70],windowBus[69],windowBus[68],
                           windowBus[67],windowBus[66],windowBus[65],
                           windowBus[64]}), .regPage1NextUnit ({page1Out_19__15,
                           page1Out_19__14,page1Out_19__13,page1Out_19__12,
                           page1Out_19__11,page1Out_19__10,page1Out_19__9,
                           page1Out_19__8,page1Out_19__7,page1Out_19__6,
                           page1Out_19__5,page1Out_19__4,page1Out_19__3,
                           page1Out_19__2,page1Out_19__1,page1Out_19__0}), .regPage2NextUnit (
                           {page2Out_19__15,page2Out_19__14,page2Out_19__13,
                           page2Out_19__12,page2Out_19__11,page2Out_19__10,
                           page2Out_19__9,page2Out_19__8,page2Out_19__7,
                           page2Out_19__6,page2Out_19__5,page2Out_19__4,
                           page2Out_19__3,page2Out_19__2,page2Out_19__1,
                           page2Out_19__0}), .clk (clk), .rst (rst), .enableRegPage1 (
                           page1Enables_2), .enableRegPage2 (page2Enables_2), .enableRegFilter (
                           nx3488), .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           pagesOuts_20__15,pagesOuts_20__14,pagesOuts_20__13,
                           pagesOuts_20__12,pagesOuts_20__11,pagesOuts_20__10,
                           pagesOuts_20__9,pagesOuts_20__8,pagesOuts_20__7,
                           pagesOuts_20__6,pagesOuts_20__5,pagesOuts_20__4,
                           pagesOuts_20__3,pagesOuts_20__2,pagesOuts_20__1,
                           pagesOuts_20__0}), .outputRegPage1 ({page1Out_14__15,
                           page1Out_14__14,page1Out_14__13,page1Out_14__12,
                           page1Out_14__11,page1Out_14__10,page1Out_14__9,
                           page1Out_14__8,page1Out_14__7,page1Out_14__6,
                           page1Out_14__5,page1Out_14__4,page1Out_14__3,
                           page1Out_14__2,page1Out_14__1,page1Out_14__0}), .outputRegPage2 (
                           {page2Out_14__15,page2Out_14__14,page2Out_14__13,
                           page2Out_14__12,page2Out_14__11,page2Out_14__10,
                           page2Out_14__9,page2Out_14__8,page2Out_14__7,
                           page2Out_14__6,page2Out_14__5,page2Out_14__4,
                           page2Out_14__3,page2Out_14__2,page2Out_14__1,
                           page2Out_14__0}), .outFilter ({filtersOuts_20__7,
                           filtersOuts_20__6,filtersOuts_20__5,filtersOuts_20__4
                           ,filtersOuts_20__3,filtersOuts_20__2,
                           filtersOuts_20__1,filtersOuts_20__0})) ;
    RegUnit_8_16_unfolded0 loop1_3_regRowMap_loop1_0_regUnitMap (.filterBus ({
                           filterBus[7],filterBus[6],filterBus[5],filterBus[4],
                           filterBus[3],filterBus[2],filterBus[1],filterBus[0]})
                           , .windowBus ({windowBus[15],windowBus[14],
                           windowBus[13],windowBus[12],windowBus[11],
                           windowBus[10],windowBus[9],windowBus[8],windowBus[7],
                           windowBus[6],windowBus[5],windowBus[4],windowBus[3],
                           windowBus[2],windowBus[1],windowBus[0]}), .regPage1NextUnit (
                           {page1Out_20__15,page1Out_20__14,page1Out_20__13,
                           page1Out_20__12,page1Out_20__11,page1Out_20__10,
                           page1Out_20__9,page1Out_20__8,page1Out_20__7,
                           page1Out_20__6,page1Out_20__5,page1Out_20__4,
                           page1Out_20__3,page1Out_20__2,page1Out_20__1,
                           page1Out_20__0}), .regPage2NextUnit ({page2Out_20__15
                           ,page2Out_20__14,page2Out_20__13,page2Out_20__12,
                           page2Out_20__11,page2Out_20__10,page2Out_20__9,
                           page2Out_20__8,page2Out_20__7,page2Out_20__6,
                           page2Out_20__5,page2Out_20__4,page2Out_20__3,
                           page2Out_20__2,page2Out_20__1,page2Out_20__0}), .clk (
                           clk), .rst (rst), .enableRegPage1 (page1Enables_3), .enableRegPage2 (
                           page2Enables_3), .enableRegFilter (nx3490), .page1ReadBusOrPage2 (
                           shift2To1), .page2ReadBusOrPage1 (shift1To2), .pageTurn (
                           pageTurn), .outRegPage ({pagesOuts_9__15,
                           pagesOuts_9__14,pagesOuts_9__13,pagesOuts_9__12,
                           pagesOuts_9__11,pagesOuts_9__10,pagesOuts_9__9,
                           pagesOuts_9__8,pagesOuts_9__7,pagesOuts_9__6,
                           pagesOuts_9__5,pagesOuts_9__4,pagesOuts_9__3,
                           pagesOuts_9__2,pagesOuts_9__1,pagesOuts_9__0}), .outputRegPage1 (
                           {page1Out_15__15,page1Out_15__14,page1Out_15__13,
                           page1Out_15__12,page1Out_15__11,page1Out_15__10,
                           page1Out_15__9,page1Out_15__8,page1Out_15__7,
                           page1Out_15__6,page1Out_15__5,page1Out_15__4,
                           page1Out_15__3,page1Out_15__2,page1Out_15__1,
                           page1Out_15__0}), .outputRegPage2 ({page2Out_15__15,
                           page2Out_15__14,page2Out_15__13,page2Out_15__12,
                           page2Out_15__11,page2Out_15__10,page2Out_15__9,
                           page2Out_15__8,page2Out_15__7,page2Out_15__6,
                           page2Out_15__5,page2Out_15__4,page2Out_15__3,
                           page2Out_15__2,page2Out_15__1,page2Out_15__0}), .outFilter (
                           {filtersOuts_9__7,filtersOuts_9__6,filtersOuts_9__5,
                           filtersOuts_9__4,filtersOuts_9__3,filtersOuts_9__2,
                           filtersOuts_9__1,filtersOuts_9__0})) ;
    RegUnit_8_16_unfolded0 loop1_3_regRowMap_loop1_1_regUnitMap (.filterBus ({
                           filterBus[15],filterBus[14],filterBus[13],
                           filterBus[12],filterBus[11],filterBus[10],
                           filterBus[9],filterBus[8]}), .windowBus ({
                           windowBus[31],windowBus[30],windowBus[29],
                           windowBus[28],windowBus[27],windowBus[26],
                           windowBus[25],windowBus[24],windowBus[23],
                           windowBus[22],windowBus[21],windowBus[20],
                           windowBus[19],windowBus[18],windowBus[17],
                           windowBus[16]}), .regPage1NextUnit ({page1Out_21__15,
                           page1Out_21__14,page1Out_21__13,page1Out_21__12,
                           page1Out_21__11,page1Out_21__10,page1Out_21__9,
                           page1Out_21__8,page1Out_21__7,page1Out_21__6,
                           page1Out_21__5,page1Out_21__4,page1Out_21__3,
                           page1Out_21__2,page1Out_21__1,page1Out_21__0}), .regPage2NextUnit (
                           {page2Out_21__15,page2Out_21__14,page2Out_21__13,
                           page2Out_21__12,page2Out_21__11,page2Out_21__10,
                           page2Out_21__9,page2Out_21__8,page2Out_21__7,
                           page2Out_21__6,page2Out_21__5,page2Out_21__4,
                           page2Out_21__3,page2Out_21__2,page2Out_21__1,
                           page2Out_21__0}), .clk (clk), .rst (rst), .enableRegPage1 (
                           page1Enables_3), .enableRegPage2 (page2Enables_3), .enableRegFilter (
                           nx3490), .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           pagesOuts_10__15,pagesOuts_10__14,pagesOuts_10__13,
                           pagesOuts_10__12,pagesOuts_10__11,pagesOuts_10__10,
                           pagesOuts_10__9,pagesOuts_10__8,pagesOuts_10__7,
                           pagesOuts_10__6,pagesOuts_10__5,pagesOuts_10__4,
                           pagesOuts_10__3,pagesOuts_10__2,pagesOuts_10__1,
                           pagesOuts_10__0}), .outputRegPage1 ({page1Out_16__15,
                           page1Out_16__14,page1Out_16__13,page1Out_16__12,
                           page1Out_16__11,page1Out_16__10,page1Out_16__9,
                           page1Out_16__8,page1Out_16__7,page1Out_16__6,
                           page1Out_16__5,page1Out_16__4,page1Out_16__3,
                           page1Out_16__2,page1Out_16__1,page1Out_16__0}), .outputRegPage2 (
                           {page2Out_16__15,page2Out_16__14,page2Out_16__13,
                           page2Out_16__12,page2Out_16__11,page2Out_16__10,
                           page2Out_16__9,page2Out_16__8,page2Out_16__7,
                           page2Out_16__6,page2Out_16__5,page2Out_16__4,
                           page2Out_16__3,page2Out_16__2,page2Out_16__1,
                           page2Out_16__0}), .outFilter ({filtersOuts_10__7,
                           filtersOuts_10__6,filtersOuts_10__5,filtersOuts_10__4
                           ,filtersOuts_10__3,filtersOuts_10__2,
                           filtersOuts_10__1,filtersOuts_10__0})) ;
    RegUnit_8_16_unfolded0 loop1_3_regRowMap_loop1_2_regUnitMap (.filterBus ({
                           filterBus[23],filterBus[22],filterBus[21],
                           filterBus[20],filterBus[19],filterBus[18],
                           filterBus[17],filterBus[16]}), .windowBus ({
                           windowBus[47],windowBus[46],windowBus[45],
                           windowBus[44],windowBus[43],windowBus[42],
                           windowBus[41],windowBus[40],windowBus[39],
                           windowBus[38],windowBus[37],windowBus[36],
                           windowBus[35],windowBus[34],windowBus[33],
                           windowBus[32]}), .regPage1NextUnit ({page1Out_22__15,
                           page1Out_22__14,page1Out_22__13,page1Out_22__12,
                           page1Out_22__11,page1Out_22__10,page1Out_22__9,
                           page1Out_22__8,page1Out_22__7,page1Out_22__6,
                           page1Out_22__5,page1Out_22__4,page1Out_22__3,
                           page1Out_22__2,page1Out_22__1,page1Out_22__0}), .regPage2NextUnit (
                           {page2Out_22__15,page2Out_22__14,page2Out_22__13,
                           page2Out_22__12,page2Out_22__11,page2Out_22__10,
                           page2Out_22__9,page2Out_22__8,page2Out_22__7,
                           page2Out_22__6,page2Out_22__5,page2Out_22__4,
                           page2Out_22__3,page2Out_22__2,page2Out_22__1,
                           page2Out_22__0}), .clk (clk), .rst (rst), .enableRegPage1 (
                           page1Enables_3), .enableRegPage2 (page2Enables_3), .enableRegFilter (
                           nx3490), .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           pagesOuts_11__15,pagesOuts_11__14,pagesOuts_11__13,
                           pagesOuts_11__12,pagesOuts_11__11,pagesOuts_11__10,
                           pagesOuts_11__9,pagesOuts_11__8,pagesOuts_11__7,
                           pagesOuts_11__6,pagesOuts_11__5,pagesOuts_11__4,
                           pagesOuts_11__3,pagesOuts_11__2,pagesOuts_11__1,
                           pagesOuts_11__0}), .outputRegPage1 ({page1Out_17__15,
                           page1Out_17__14,page1Out_17__13,page1Out_17__12,
                           page1Out_17__11,page1Out_17__10,page1Out_17__9,
                           page1Out_17__8,page1Out_17__7,page1Out_17__6,
                           page1Out_17__5,page1Out_17__4,page1Out_17__3,
                           page1Out_17__2,page1Out_17__1,page1Out_17__0}), .outputRegPage2 (
                           {page2Out_17__15,page2Out_17__14,page2Out_17__13,
                           page2Out_17__12,page2Out_17__11,page2Out_17__10,
                           page2Out_17__9,page2Out_17__8,page2Out_17__7,
                           page2Out_17__6,page2Out_17__5,page2Out_17__4,
                           page2Out_17__3,page2Out_17__2,page2Out_17__1,
                           page2Out_17__0}), .outFilter ({filtersOuts_11__7,
                           filtersOuts_11__6,filtersOuts_11__5,filtersOuts_11__4
                           ,filtersOuts_11__3,filtersOuts_11__2,
                           filtersOuts_11__1,filtersOuts_11__0})) ;
    RegUnit_8_16_unfolded0 loop1_3_regRowMap_loop1_3_regUnitMap (.filterBus ({
                           filterBus[31],filterBus[30],filterBus[29],
                           filterBus[28],filterBus[27],filterBus[26],
                           filterBus[25],filterBus[24]}), .windowBus ({
                           windowBus[63],windowBus[62],windowBus[61],
                           windowBus[60],windowBus[59],windowBus[58],
                           windowBus[57],windowBus[56],windowBus[55],
                           windowBus[54],windowBus[53],windowBus[52],
                           windowBus[51],windowBus[50],windowBus[49],
                           windowBus[48]}), .regPage1NextUnit ({page1Out_23__15,
                           page1Out_23__14,page1Out_23__13,page1Out_23__12,
                           page1Out_23__11,page1Out_23__10,page1Out_23__9,
                           page1Out_23__8,page1Out_23__7,page1Out_23__6,
                           page1Out_23__5,page1Out_23__4,page1Out_23__3,
                           page1Out_23__2,page1Out_23__1,page1Out_23__0}), .regPage2NextUnit (
                           {page2Out_23__15,page2Out_23__14,page2Out_23__13,
                           page2Out_23__12,page2Out_23__11,page2Out_23__10,
                           page2Out_23__9,page2Out_23__8,page2Out_23__7,
                           page2Out_23__6,page2Out_23__5,page2Out_23__4,
                           page2Out_23__3,page2Out_23__2,page2Out_23__1,
                           page2Out_23__0}), .clk (clk), .rst (rst), .enableRegPage1 (
                           page1Enables_3), .enableRegPage2 (page2Enables_3), .enableRegFilter (
                           nx3492), .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           pagesOuts_21__15,pagesOuts_21__14,pagesOuts_21__13,
                           pagesOuts_21__12,pagesOuts_21__11,pagesOuts_21__10,
                           pagesOuts_21__9,pagesOuts_21__8,pagesOuts_21__7,
                           pagesOuts_21__6,pagesOuts_21__5,pagesOuts_21__4,
                           pagesOuts_21__3,pagesOuts_21__2,pagesOuts_21__1,
                           pagesOuts_21__0}), .outputRegPage1 ({page1Out_18__15,
                           page1Out_18__14,page1Out_18__13,page1Out_18__12,
                           page1Out_18__11,page1Out_18__10,page1Out_18__9,
                           page1Out_18__8,page1Out_18__7,page1Out_18__6,
                           page1Out_18__5,page1Out_18__4,page1Out_18__3,
                           page1Out_18__2,page1Out_18__1,page1Out_18__0}), .outputRegPage2 (
                           {page2Out_18__15,page2Out_18__14,page2Out_18__13,
                           page2Out_18__12,page2Out_18__11,page2Out_18__10,
                           page2Out_18__9,page2Out_18__8,page2Out_18__7,
                           page2Out_18__6,page2Out_18__5,page2Out_18__4,
                           page2Out_18__3,page2Out_18__2,page2Out_18__1,
                           page2Out_18__0}), .outFilter ({filtersOuts_21__7,
                           filtersOuts_21__6,filtersOuts_21__5,filtersOuts_21__4
                           ,filtersOuts_21__3,filtersOuts_21__2,
                           filtersOuts_21__1,filtersOuts_21__0})) ;
    RegUnit_8_16_unfolded0 loop1_3_regRowMap_loop1_4_regUnitMap (.filterBus ({
                           filterBus[39],filterBus[38],filterBus[37],
                           filterBus[36],filterBus[35],filterBus[34],
                           filterBus[33],filterBus[32]}), .windowBus ({
                           windowBus[79],windowBus[78],windowBus[77],
                           windowBus[76],windowBus[75],windowBus[74],
                           windowBus[73],windowBus[72],windowBus[71],
                           windowBus[70],windowBus[69],windowBus[68],
                           windowBus[67],windowBus[66],windowBus[65],
                           windowBus[64]}), .regPage1NextUnit ({page1Out_24__15,
                           page1Out_24__14,page1Out_24__13,page1Out_24__12,
                           page1Out_24__11,page1Out_24__10,page1Out_24__9,
                           page1Out_24__8,page1Out_24__7,page1Out_24__6,
                           page1Out_24__5,page1Out_24__4,page1Out_24__3,
                           page1Out_24__2,page1Out_24__1,page1Out_24__0}), .regPage2NextUnit (
                           {page2Out_24__15,page2Out_24__14,page2Out_24__13,
                           page2Out_24__12,page2Out_24__11,page2Out_24__10,
                           page2Out_24__9,page2Out_24__8,page2Out_24__7,
                           page2Out_24__6,page2Out_24__5,page2Out_24__4,
                           page2Out_24__3,page2Out_24__2,page2Out_24__1,
                           page2Out_24__0}), .clk (clk), .rst (rst), .enableRegPage1 (
                           page1Enables_3), .enableRegPage2 (page2Enables_3), .enableRegFilter (
                           nx3492), .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           pagesOuts_22__15,pagesOuts_22__14,pagesOuts_22__13,
                           pagesOuts_22__12,pagesOuts_22__11,pagesOuts_22__10,
                           pagesOuts_22__9,pagesOuts_22__8,pagesOuts_22__7,
                           pagesOuts_22__6,pagesOuts_22__5,pagesOuts_22__4,
                           pagesOuts_22__3,pagesOuts_22__2,pagesOuts_22__1,
                           pagesOuts_22__0}), .outputRegPage1 ({page1Out_19__15,
                           page1Out_19__14,page1Out_19__13,page1Out_19__12,
                           page1Out_19__11,page1Out_19__10,page1Out_19__9,
                           page1Out_19__8,page1Out_19__7,page1Out_19__6,
                           page1Out_19__5,page1Out_19__4,page1Out_19__3,
                           page1Out_19__2,page1Out_19__1,page1Out_19__0}), .outputRegPage2 (
                           {page2Out_19__15,page2Out_19__14,page2Out_19__13,
                           page2Out_19__12,page2Out_19__11,page2Out_19__10,
                           page2Out_19__9,page2Out_19__8,page2Out_19__7,
                           page2Out_19__6,page2Out_19__5,page2Out_19__4,
                           page2Out_19__3,page2Out_19__2,page2Out_19__1,
                           page2Out_19__0}), .outFilter ({filtersOuts_22__7,
                           filtersOuts_22__6,filtersOuts_22__5,filtersOuts_22__4
                           ,filtersOuts_22__3,filtersOuts_22__2,
                           filtersOuts_22__1,filtersOuts_22__0})) ;
    RegUnit_8_16_unfolded1 loop1_4_regRowMap_loop1_0_regUnitMap (.filterBus ({
                           filterBus[7],filterBus[6],filterBus[5],filterBus[4],
                           filterBus[3],filterBus[2],filterBus[1],filterBus[0]})
                           , .windowBus ({windowBus[15],windowBus[14],
                           windowBus[13],windowBus[12],windowBus[11],
                           windowBus[10],windowBus[9],windowBus[8],windowBus[7],
                           windowBus[6],windowBus[5],windowBus[4],windowBus[3],
                           windowBus[2],windowBus[1],windowBus[0]}), .regPage1NextUnit (
                           {page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15}), .regPage2NextUnit ({
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15}), .clk (clk), .rst (rst), .enableRegPage1 (
                           page1Enables_4), .enableRegPage2 (page2Enables_4), .enableRegFilter (
                           nx3494), .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           pagesOuts_12__15,pagesOuts_12__14,pagesOuts_12__13,
                           pagesOuts_12__12,pagesOuts_12__11,pagesOuts_12__10,
                           pagesOuts_12__9,pagesOuts_12__8,pagesOuts_12__7,
                           pagesOuts_12__6,pagesOuts_12__5,pagesOuts_12__4,
                           pagesOuts_12__3,pagesOuts_12__2,pagesOuts_12__1,
                           pagesOuts_12__0}), .outputRegPage1 ({page1Out_20__15,
                           page1Out_20__14,page1Out_20__13,page1Out_20__12,
                           page1Out_20__11,page1Out_20__10,page1Out_20__9,
                           page1Out_20__8,page1Out_20__7,page1Out_20__6,
                           page1Out_20__5,page1Out_20__4,page1Out_20__3,
                           page1Out_20__2,page1Out_20__1,page1Out_20__0}), .outputRegPage2 (
                           {page2Out_20__15,page2Out_20__14,page2Out_20__13,
                           page2Out_20__12,page2Out_20__11,page2Out_20__10,
                           page2Out_20__9,page2Out_20__8,page2Out_20__7,
                           page2Out_20__6,page2Out_20__5,page2Out_20__4,
                           page2Out_20__3,page2Out_20__2,page2Out_20__1,
                           page2Out_20__0}), .outFilter ({filtersOuts_12__7,
                           filtersOuts_12__6,filtersOuts_12__5,filtersOuts_12__4
                           ,filtersOuts_12__3,filtersOuts_12__2,
                           filtersOuts_12__1,filtersOuts_12__0})) ;
    RegUnit_8_16_unfolded1 loop1_4_regRowMap_loop1_1_regUnitMap (.filterBus ({
                           filterBus[15],filterBus[14],filterBus[13],
                           filterBus[12],filterBus[11],filterBus[10],
                           filterBus[9],filterBus[8]}), .windowBus ({
                           windowBus[31],windowBus[30],windowBus[29],
                           windowBus[28],windowBus[27],windowBus[26],
                           windowBus[25],windowBus[24],windowBus[23],
                           windowBus[22],windowBus[21],windowBus[20],
                           windowBus[19],windowBus[18],windowBus[17],
                           windowBus[16]}), .regPage1NextUnit ({page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15}), .regPage2NextUnit (
                           {page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15}), .clk (clk), .rst (rst), .enableRegPage1 (
                           page1Enables_4), .enableRegPage2 (page2Enables_4), .enableRegFilter (
                           nx3494), .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           pagesOuts_13__15,pagesOuts_13__14,pagesOuts_13__13,
                           pagesOuts_13__12,pagesOuts_13__11,pagesOuts_13__10,
                           pagesOuts_13__9,pagesOuts_13__8,pagesOuts_13__7,
                           pagesOuts_13__6,pagesOuts_13__5,pagesOuts_13__4,
                           pagesOuts_13__3,pagesOuts_13__2,pagesOuts_13__1,
                           pagesOuts_13__0}), .outputRegPage1 ({page1Out_21__15,
                           page1Out_21__14,page1Out_21__13,page1Out_21__12,
                           page1Out_21__11,page1Out_21__10,page1Out_21__9,
                           page1Out_21__8,page1Out_21__7,page1Out_21__6,
                           page1Out_21__5,page1Out_21__4,page1Out_21__3,
                           page1Out_21__2,page1Out_21__1,page1Out_21__0}), .outputRegPage2 (
                           {page2Out_21__15,page2Out_21__14,page2Out_21__13,
                           page2Out_21__12,page2Out_21__11,page2Out_21__10,
                           page2Out_21__9,page2Out_21__8,page2Out_21__7,
                           page2Out_21__6,page2Out_21__5,page2Out_21__4,
                           page2Out_21__3,page2Out_21__2,page2Out_21__1,
                           page2Out_21__0}), .outFilter ({filtersOuts_13__7,
                           filtersOuts_13__6,filtersOuts_13__5,filtersOuts_13__4
                           ,filtersOuts_13__3,filtersOuts_13__2,
                           filtersOuts_13__1,filtersOuts_13__0})) ;
    RegUnit_8_16_unfolded1 loop1_4_regRowMap_loop1_2_regUnitMap (.filterBus ({
                           filterBus[23],filterBus[22],filterBus[21],
                           filterBus[20],filterBus[19],filterBus[18],
                           filterBus[17],filterBus[16]}), .windowBus ({
                           windowBus[47],windowBus[46],windowBus[45],
                           windowBus[44],windowBus[43],windowBus[42],
                           windowBus[41],windowBus[40],windowBus[39],
                           windowBus[38],windowBus[37],windowBus[36],
                           windowBus[35],windowBus[34],windowBus[33],
                           windowBus[32]}), .regPage1NextUnit ({page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15}), .regPage2NextUnit (
                           {page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15}), .clk (clk), .rst (rst), .enableRegPage1 (
                           page1Enables_4), .enableRegPage2 (page2Enables_4), .enableRegFilter (
                           nx3494), .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           pagesOuts_14__15,pagesOuts_14__14,pagesOuts_14__13,
                           pagesOuts_14__12,pagesOuts_14__11,pagesOuts_14__10,
                           pagesOuts_14__9,pagesOuts_14__8,pagesOuts_14__7,
                           pagesOuts_14__6,pagesOuts_14__5,pagesOuts_14__4,
                           pagesOuts_14__3,pagesOuts_14__2,pagesOuts_14__1,
                           pagesOuts_14__0}), .outputRegPage1 ({page1Out_22__15,
                           page1Out_22__14,page1Out_22__13,page1Out_22__12,
                           page1Out_22__11,page1Out_22__10,page1Out_22__9,
                           page1Out_22__8,page1Out_22__7,page1Out_22__6,
                           page1Out_22__5,page1Out_22__4,page1Out_22__3,
                           page1Out_22__2,page1Out_22__1,page1Out_22__0}), .outputRegPage2 (
                           {page2Out_22__15,page2Out_22__14,page2Out_22__13,
                           page2Out_22__12,page2Out_22__11,page2Out_22__10,
                           page2Out_22__9,page2Out_22__8,page2Out_22__7,
                           page2Out_22__6,page2Out_22__5,page2Out_22__4,
                           page2Out_22__3,page2Out_22__2,page2Out_22__1,
                           page2Out_22__0}), .outFilter ({filtersOuts_14__7,
                           filtersOuts_14__6,filtersOuts_14__5,filtersOuts_14__4
                           ,filtersOuts_14__3,filtersOuts_14__2,
                           filtersOuts_14__1,filtersOuts_14__0})) ;
    RegUnit_8_16_unfolded1 loop1_4_regRowMap_loop1_3_regUnitMap (.filterBus ({
                           filterBus[31],filterBus[30],filterBus[29],
                           filterBus[28],filterBus[27],filterBus[26],
                           filterBus[25],filterBus[24]}), .windowBus ({
                           windowBus[63],windowBus[62],windowBus[61],
                           windowBus[60],windowBus[59],windowBus[58],
                           windowBus[57],windowBus[56],windowBus[55],
                           windowBus[54],windowBus[53],windowBus[52],
                           windowBus[51],windowBus[50],windowBus[49],
                           windowBus[48]}), .regPage1NextUnit ({page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15}), .regPage2NextUnit (
                           {page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15}), .clk (clk), .rst (rst), .enableRegPage1 (
                           page1Enables_4), .enableRegPage2 (page2Enables_4), .enableRegFilter (
                           nx3496), .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           pagesOuts_23__15,pagesOuts_23__14,pagesOuts_23__13,
                           pagesOuts_23__12,pagesOuts_23__11,pagesOuts_23__10,
                           pagesOuts_23__9,pagesOuts_23__8,pagesOuts_23__7,
                           pagesOuts_23__6,pagesOuts_23__5,pagesOuts_23__4,
                           pagesOuts_23__3,pagesOuts_23__2,pagesOuts_23__1,
                           pagesOuts_23__0}), .outputRegPage1 ({page1Out_23__15,
                           page1Out_23__14,page1Out_23__13,page1Out_23__12,
                           page1Out_23__11,page1Out_23__10,page1Out_23__9,
                           page1Out_23__8,page1Out_23__7,page1Out_23__6,
                           page1Out_23__5,page1Out_23__4,page1Out_23__3,
                           page1Out_23__2,page1Out_23__1,page1Out_23__0}), .outputRegPage2 (
                           {page2Out_23__15,page2Out_23__14,page2Out_23__13,
                           page2Out_23__12,page2Out_23__11,page2Out_23__10,
                           page2Out_23__9,page2Out_23__8,page2Out_23__7,
                           page2Out_23__6,page2Out_23__5,page2Out_23__4,
                           page2Out_23__3,page2Out_23__2,page2Out_23__1,
                           page2Out_23__0}), .outFilter ({filtersOuts_23__7,
                           filtersOuts_23__6,filtersOuts_23__5,filtersOuts_23__4
                           ,filtersOuts_23__3,filtersOuts_23__2,
                           filtersOuts_23__1,filtersOuts_23__0})) ;
    RegUnit_8_16_unfolded1 loop1_4_regRowMap_loop1_4_regUnitMap (.filterBus ({
                           filterBus[39],filterBus[38],filterBus[37],
                           filterBus[36],filterBus[35],filterBus[34],
                           filterBus[33],filterBus[32]}), .windowBus ({
                           windowBus[79],windowBus[78],windowBus[77],
                           windowBus[76],windowBus[75],windowBus[74],
                           windowBus[73],windowBus[72],windowBus[71],
                           windowBus[70],windowBus[69],windowBus[68],
                           windowBus[67],windowBus[66],windowBus[65],
                           windowBus[64]}), .regPage1NextUnit ({page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15}), .regPage2NextUnit (
                           {page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15,page1Out_25__15,page1Out_25__15,
                           page1Out_25__15}), .clk (clk), .rst (rst), .enableRegPage1 (
                           page1Enables_4), .enableRegPage2 (page2Enables_4), .enableRegFilter (
                           nx3496), .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           pagesOuts_24__15,pagesOuts_24__14,pagesOuts_24__13,
                           pagesOuts_24__12,pagesOuts_24__11,pagesOuts_24__10,
                           pagesOuts_24__9,pagesOuts_24__8,pagesOuts_24__7,
                           pagesOuts_24__6,pagesOuts_24__5,pagesOuts_24__4,
                           pagesOuts_24__3,pagesOuts_24__2,pagesOuts_24__1,
                           pagesOuts_24__0}), .outputRegPage1 ({page1Out_24__15,
                           page1Out_24__14,page1Out_24__13,page1Out_24__12,
                           page1Out_24__11,page1Out_24__10,page1Out_24__9,
                           page1Out_24__8,page1Out_24__7,page1Out_24__6,
                           page1Out_24__5,page1Out_24__4,page1Out_24__3,
                           page1Out_24__2,page1Out_24__1,page1Out_24__0}), .outputRegPage2 (
                           {page2Out_24__15,page2Out_24__14,page2Out_24__13,
                           page2Out_24__12,page2Out_24__11,page2Out_24__10,
                           page2Out_24__9,page2Out_24__8,page2Out_24__7,
                           page2Out_24__6,page2Out_24__5,page2Out_24__4,
                           page2Out_24__3,page2Out_24__2,page2Out_24__1,
                           page2Out_24__0}), .outFilter ({filtersOuts_24__7,
                           filtersOuts_24__6,filtersOuts_24__5,filtersOuts_24__4
                           ,filtersOuts_24__3,filtersOuts_24__2,
                           filtersOuts_24__1,filtersOuts_24__0})) ;
    fake_gnd ix3415 (.Y (page1Out_25__15)) ;
    nand03 ix3430 (.Y (nx3429), .A0 (enableFilterRead), .A1 (nx4), .A2 (
           decoderRow[2])) ;
    nor02_2x ix5 (.Y (nx4), .A0 (decoderRow[1]), .A1 (decoderRow[0])) ;
    nor03_2x ix29 (.Y (filterEnables_3), .A0 (nx3433), .A1 (decoderRow[2]), .A2 (
             nx3435)) ;
    inv02 ix3434 (.Y (nx3433), .A (enableFilterRead)) ;
    nand02 ix3436 (.Y (nx3435), .A0 (decoderRow[1]), .A1 (decoderRow[0])) ;
    nor03_2x ix41 (.Y (filterEnables_2), .A0 (nx3433), .A1 (decoderRow[2]), .A2 (
             nx3438)) ;
    nand02 ix3439 (.Y (nx3438), .A0 (decoderRow[1]), .A1 (nx3440)) ;
    inv01 ix3441 (.Y (nx3440), .A (decoderRow[0])) ;
    nor03_2x ix53 (.Y (filterEnables_1), .A0 (nx3433), .A1 (decoderRow[2]), .A2 (
             nx3443)) ;
    nand02 ix3444 (.Y (nx3443), .A0 (nx3445), .A1 (decoderRow[0])) ;
    inv01 ix3446 (.Y (nx3445), .A (decoderRow[1])) ;
    nor03_2x ix67 (.Y (filterEnables_0), .A0 (nx3433), .A1 (decoderRow[2]), .A2 (
             nx3448)) ;
    inv01 ix3449 (.Y (nx3448), .A (nx62)) ;
    nor02_2x ix63 (.Y (nx62), .A0 (decoderRow[1]), .A1 (decoderRow[0])) ;
    inv01 ix17 (.Y (page2Enables_4), .A (nx3452)) ;
    nand03 ix3453 (.Y (nx3452), .A0 (enablePage2Read), .A1 (nx4), .A2 (
           decoderRow[2])) ;
    nor03_2x ix31 (.Y (page2Enables_3), .A0 (nx3455), .A1 (decoderRow[2]), .A2 (
             nx3435)) ;
    inv02 ix3456 (.Y (nx3455), .A (enablePage2Read)) ;
    nor03_2x ix43 (.Y (page2Enables_2), .A0 (nx3455), .A1 (decoderRow[2]), .A2 (
             nx3438)) ;
    nor03_2x ix55 (.Y (page2Enables_1), .A0 (nx3455), .A1 (decoderRow[2]), .A2 (
             nx3443)) ;
    nor03_2x ix69 (.Y (page2Enables_0), .A0 (nx3455), .A1 (decoderRow[2]), .A2 (
             nx3448)) ;
    inv01 ix19 (.Y (page1Enables_4), .A (nx3461)) ;
    nand03 ix3462 (.Y (nx3461), .A0 (enablePage1Read), .A1 (nx4), .A2 (
           decoderRow[2])) ;
    nor03_2x ix33 (.Y (page1Enables_3), .A0 (nx3464), .A1 (decoderRow[2]), .A2 (
             nx3435)) ;
    inv02 ix3465 (.Y (nx3464), .A (enablePage1Read)) ;
    nor03_2x ix45 (.Y (page1Enables_2), .A0 (nx3464), .A1 (decoderRow[2]), .A2 (
             nx3438)) ;
    nor03_2x ix57 (.Y (page1Enables_1), .A0 (nx3464), .A1 (decoderRow[2]), .A2 (
             nx3443)) ;
    nor03_2x ix71 (.Y (page1Enables_0), .A0 (nx3464), .A1 (decoderRow[2]), .A2 (
             nx3448)) ;
    buf02 ix3477 (.Y (nx3478), .A (filterEnables_0)) ;
    buf02 ix3479 (.Y (nx3480), .A (filterEnables_0)) ;
    buf02 ix3481 (.Y (nx3482), .A (filterEnables_1)) ;
    buf02 ix3483 (.Y (nx3484), .A (filterEnables_1)) ;
    buf02 ix3485 (.Y (nx3486), .A (filterEnables_2)) ;
    buf02 ix3487 (.Y (nx3488), .A (filterEnables_2)) ;
    buf02 ix3489 (.Y (nx3490), .A (filterEnables_3)) ;
    buf02 ix3491 (.Y (nx3492), .A (filterEnables_3)) ;
    inv02 ix3493 (.Y (nx3494), .A (nx3429)) ;
    inv02 ix3495 (.Y (nx3496), .A (nx3429)) ;
endmodule


module RegUnit_8_16_unfolded1 ( filterBus, windowBus, regPage1NextUnit, 
                                regPage2NextUnit, clk, rst, enableRegPage1, 
                                enableRegPage2, enableRegFilter, 
                                page1ReadBusOrPage2, page2ReadBusOrPage1, 
                                pageTurn, outRegPage, outputRegPage1, 
                                outputRegPage2, outFilter ) ;

    input [7:0]filterBus ;
    input [15:0]windowBus ;
    input [15:0]regPage1NextUnit ;
    input [15:0]regPage2NextUnit ;
    input clk ;
    input rst ;
    input enableRegPage1 ;
    input enableRegPage2 ;
    input enableRegFilter ;
    input page1ReadBusOrPage2 ;
    input page2ReadBusOrPage1 ;
    input pageTurn ;
    output [15:0]outRegPage ;
    output [15:0]outputRegPage1 ;
    output [15:0]outputRegPage2 ;
    output [7:0]outFilter ;

    wire nx133, nx143, nx153, nx163, nx173, nx183, nx193, nx203, nx213, nx223, 
         nx233, nx243, nx253, nx263, nx273, nx283, nx293, nx303, nx313, nx323, 
         nx333, nx343, nx353, nx363, nx373, nx383, nx393, nx403, nx413, nx423, 
         nx433, nx443, nx453, nx463, nx473, nx483, nx493, nx503, nx513, nx523, 
         nx535, nx539, nx544, nx546, nx551, nx553, nx558, nx560, nx565, nx567, 
         nx572, nx574, nx579, nx581, nx586, nx588, nx593, nx595, nx597, nx599, 
         nx601, nx604, nx606, nx608, nx611, nx613, nx615, nx618, nx620, nx622, 
         nx625, nx627, nx629, nx632, nx634, nx636, nx639, nx641, nx643, nx646, 
         nx648, nx650, nx653, nx655, nx657, nx660, nx662, nx664, nx667, nx669, 
         nx671, nx674, nx676, nx678, nx681, nx683, nx685, nx688, nx690, nx692, 
         nx695, nx697, nx699, nx702, nx704, nx706, nx709, nx711, nx713, nx715, 
         nx717, nx720, nx722, nx724, nx727, nx729, nx731, nx734, nx736, nx738, 
         nx741, nx743, nx745, nx748, nx750, nx752, nx755, nx757, nx759, nx762, 
         nx764, nx766, nx769, nx771, nx773, nx776, nx778, nx780, nx783, nx785, 
         nx787, nx790, nx792, nx794, nx797, nx799, nx801, nx804, nx806, nx808, 
         nx811, nx813, nx815, nx818, nx820, nx822, nx846, nx848, nx850, nx852, 
         nx854, nx856, nx858, nx860, nx862, nx868, nx870, nx872, nx874, nx876, 
         nx878, nx880, nx882, nx884, nx886, nx888, nx890;
    wire [7:0] \$dummy ;




    dffr regFilterMap_reg_Q_0 (.Q (outFilter[0]), .QB (\$dummy [0]), .D (nx453)
         , .CLK (clk), .R (rst)) ;
    nand02 ix454 (.Y (nx453), .A0 (nx535), .A1 (nx539)) ;
    nand02 ix536 (.Y (nx535), .A0 (outFilter[0]), .A1 (nx888)) ;
    nand02 ix540 (.Y (nx539), .A0 (filterBus[0]), .A1 (nx884)) ;
    dffr regFilterMap_reg_Q_1 (.Q (outFilter[1]), .QB (\$dummy [1]), .D (nx463)
         , .CLK (clk), .R (rst)) ;
    nand02 ix464 (.Y (nx463), .A0 (nx544), .A1 (nx546)) ;
    nand02 ix545 (.Y (nx544), .A0 (outFilter[1]), .A1 (nx888)) ;
    nand02 ix547 (.Y (nx546), .A0 (filterBus[1]), .A1 (nx884)) ;
    dffr regFilterMap_reg_Q_2 (.Q (outFilter[2]), .QB (\$dummy [2]), .D (nx473)
         , .CLK (clk), .R (rst)) ;
    nand02 ix474 (.Y (nx473), .A0 (nx551), .A1 (nx553)) ;
    nand02 ix552 (.Y (nx551), .A0 (outFilter[2]), .A1 (nx888)) ;
    nand02 ix554 (.Y (nx553), .A0 (filterBus[2]), .A1 (nx884)) ;
    dffr regFilterMap_reg_Q_3 (.Q (outFilter[3]), .QB (\$dummy [3]), .D (nx483)
         , .CLK (clk), .R (rst)) ;
    nand02 ix484 (.Y (nx483), .A0 (nx558), .A1 (nx560)) ;
    nand02 ix559 (.Y (nx558), .A0 (outFilter[3]), .A1 (nx888)) ;
    nand02 ix561 (.Y (nx560), .A0 (filterBus[3]), .A1 (nx884)) ;
    dffr regFilterMap_reg_Q_4 (.Q (outFilter[4]), .QB (\$dummy [4]), .D (nx493)
         , .CLK (clk), .R (rst)) ;
    nand02 ix494 (.Y (nx493), .A0 (nx565), .A1 (nx567)) ;
    nand02 ix566 (.Y (nx565), .A0 (outFilter[4]), .A1 (nx888)) ;
    nand02 ix568 (.Y (nx567), .A0 (filterBus[4]), .A1 (nx884)) ;
    dffr regFilterMap_reg_Q_5 (.Q (outFilter[5]), .QB (\$dummy [5]), .D (nx503)
         , .CLK (clk), .R (rst)) ;
    nand02 ix504 (.Y (nx503), .A0 (nx572), .A1 (nx574)) ;
    nand02 ix573 (.Y (nx572), .A0 (outFilter[5]), .A1 (nx888)) ;
    nand02 ix575 (.Y (nx574), .A0 (filterBus[5]), .A1 (nx884)) ;
    dffr regFilterMap_reg_Q_6 (.Q (outFilter[6]), .QB (\$dummy [6]), .D (nx513)
         , .CLK (clk), .R (rst)) ;
    nand02 ix514 (.Y (nx513), .A0 (nx579), .A1 (nx581)) ;
    nand02 ix580 (.Y (nx579), .A0 (outFilter[6]), .A1 (nx888)) ;
    nand02 ix582 (.Y (nx581), .A0 (filterBus[6]), .A1 (nx884)) ;
    dffr regFilterMap_reg_Q_7 (.Q (outFilter[7]), .QB (\$dummy [7]), .D (nx523)
         , .CLK (clk), .R (rst)) ;
    nand02 ix524 (.Y (nx523), .A0 (nx586), .A1 (nx588)) ;
    nand02 ix587 (.Y (nx586), .A0 (outFilter[7]), .A1 (nx846)) ;
    nand02 ix589 (.Y (nx588), .A0 (filterBus[7]), .A1 (nx886)) ;
    dffr regPage2Map_reg_Q_0 (.Q (outputRegPage2[0]), .QB (nx601), .D (nx143), .CLK (
         clk), .R (rst)) ;
    nand02 ix144 (.Y (nx143), .A0 (nx593), .A1 (nx597)) ;
    nand02 ix594 (.Y (nx593), .A0 (outputRegPage2[0]), .A1 (nx848)) ;
    nor02_2x ix596 (.Y (nx595), .A0 (nx878), .A1 (page2ReadBusOrPage1)) ;
    nand03 ix598 (.Y (nx597), .A0 (windowBus[0]), .A1 (nx852), .A2 (nx878)) ;
    inv01 ix600 (.Y (nx599), .A (page2ReadBusOrPage1)) ;
    dffr regPage2Map_reg_Q_1 (.Q (outputRegPage2[1]), .QB (nx608), .D (nx163), .CLK (
         clk), .R (rst)) ;
    nand02 ix164 (.Y (nx163), .A0 (nx604), .A1 (nx606)) ;
    nand02 ix605 (.Y (nx604), .A0 (outputRegPage2[1]), .A1 (nx848)) ;
    nand03 ix607 (.Y (nx606), .A0 (windowBus[1]), .A1 (nx852), .A2 (nx878)) ;
    dffr regPage2Map_reg_Q_2 (.Q (outputRegPage2[2]), .QB (nx615), .D (nx183), .CLK (
         clk), .R (rst)) ;
    nand02 ix184 (.Y (nx183), .A0 (nx611), .A1 (nx613)) ;
    nand02 ix612 (.Y (nx611), .A0 (outputRegPage2[2]), .A1 (nx848)) ;
    nand03 ix614 (.Y (nx613), .A0 (windowBus[2]), .A1 (nx852), .A2 (nx878)) ;
    dffr regPage2Map_reg_Q_3 (.Q (outputRegPage2[3]), .QB (nx622), .D (nx203), .CLK (
         clk), .R (rst)) ;
    nand02 ix204 (.Y (nx203), .A0 (nx618), .A1 (nx620)) ;
    nand02 ix619 (.Y (nx618), .A0 (outputRegPage2[3]), .A1 (nx848)) ;
    nand03 ix621 (.Y (nx620), .A0 (windowBus[3]), .A1 (nx852), .A2 (nx878)) ;
    dffr regPage2Map_reg_Q_4 (.Q (outputRegPage2[4]), .QB (nx629), .D (nx223), .CLK (
         clk), .R (rst)) ;
    nand02 ix224 (.Y (nx223), .A0 (nx625), .A1 (nx627)) ;
    nand02 ix626 (.Y (nx625), .A0 (outputRegPage2[4]), .A1 (nx848)) ;
    nand03 ix628 (.Y (nx627), .A0 (windowBus[4]), .A1 (nx852), .A2 (nx878)) ;
    dffr regPage2Map_reg_Q_5 (.Q (outputRegPage2[5]), .QB (nx636), .D (nx243), .CLK (
         clk), .R (rst)) ;
    nand02 ix244 (.Y (nx243), .A0 (nx632), .A1 (nx634)) ;
    nand02 ix633 (.Y (nx632), .A0 (outputRegPage2[5]), .A1 (nx848)) ;
    nand03 ix635 (.Y (nx634), .A0 (windowBus[5]), .A1 (nx852), .A2 (nx878)) ;
    dffr regPage2Map_reg_Q_6 (.Q (outputRegPage2[6]), .QB (nx643), .D (nx263), .CLK (
         clk), .R (rst)) ;
    nand02 ix264 (.Y (nx263), .A0 (nx639), .A1 (nx641)) ;
    nand02 ix640 (.Y (nx639), .A0 (outputRegPage2[6]), .A1 (nx848)) ;
    nand03 ix642 (.Y (nx641), .A0 (windowBus[6]), .A1 (nx854), .A2 (nx880)) ;
    dffr regPage2Map_reg_Q_7 (.Q (outputRegPage2[7]), .QB (nx650), .D (nx283), .CLK (
         clk), .R (rst)) ;
    nand02 ix284 (.Y (nx283), .A0 (nx646), .A1 (nx648)) ;
    nand02 ix647 (.Y (nx646), .A0 (outputRegPage2[7]), .A1 (nx850)) ;
    nand03 ix649 (.Y (nx648), .A0 (windowBus[7]), .A1 (nx854), .A2 (nx880)) ;
    dffr regPage2Map_reg_Q_8 (.Q (outputRegPage2[8]), .QB (nx657), .D (nx303), .CLK (
         clk), .R (rst)) ;
    nand02 ix304 (.Y (nx303), .A0 (nx653), .A1 (nx655)) ;
    nand02 ix654 (.Y (nx653), .A0 (outputRegPage2[8]), .A1 (nx850)) ;
    nand03 ix656 (.Y (nx655), .A0 (windowBus[8]), .A1 (nx854), .A2 (nx880)) ;
    dffr regPage2Map_reg_Q_9 (.Q (outputRegPage2[9]), .QB (nx664), .D (nx323), .CLK (
         clk), .R (rst)) ;
    nand02 ix324 (.Y (nx323), .A0 (nx660), .A1 (nx662)) ;
    nand02 ix661 (.Y (nx660), .A0 (outputRegPage2[9]), .A1 (nx850)) ;
    nand03 ix663 (.Y (nx662), .A0 (windowBus[9]), .A1 (nx854), .A2 (nx880)) ;
    dffr regPage2Map_reg_Q_10 (.Q (outputRegPage2[10]), .QB (nx671), .D (nx343)
         , .CLK (clk), .R (rst)) ;
    nand02 ix344 (.Y (nx343), .A0 (nx667), .A1 (nx669)) ;
    nand02 ix668 (.Y (nx667), .A0 (outputRegPage2[10]), .A1 (nx850)) ;
    nand03 ix670 (.Y (nx669), .A0 (windowBus[10]), .A1 (nx854), .A2 (nx880)) ;
    dffr regPage2Map_reg_Q_11 (.Q (outputRegPage2[11]), .QB (nx678), .D (nx363)
         , .CLK (clk), .R (rst)) ;
    nand02 ix364 (.Y (nx363), .A0 (nx674), .A1 (nx676)) ;
    nand02 ix675 (.Y (nx674), .A0 (outputRegPage2[11]), .A1 (nx850)) ;
    nand03 ix677 (.Y (nx676), .A0 (windowBus[11]), .A1 (nx854), .A2 (nx880)) ;
    dffr regPage2Map_reg_Q_12 (.Q (outputRegPage2[12]), .QB (nx685), .D (nx383)
         , .CLK (clk), .R (rst)) ;
    nand02 ix384 (.Y (nx383), .A0 (nx681), .A1 (nx683)) ;
    nand02 ix682 (.Y (nx681), .A0 (outputRegPage2[12]), .A1 (nx850)) ;
    nand03 ix684 (.Y (nx683), .A0 (windowBus[12]), .A1 (nx599), .A2 (nx880)) ;
    dffr regPage2Map_reg_Q_13 (.Q (outputRegPage2[13]), .QB (nx692), .D (nx403)
         , .CLK (clk), .R (rst)) ;
    nand02 ix404 (.Y (nx403), .A0 (nx688), .A1 (nx690)) ;
    nand02 ix689 (.Y (nx688), .A0 (outputRegPage2[13]), .A1 (nx850)) ;
    nand03 ix691 (.Y (nx690), .A0 (windowBus[13]), .A1 (nx599), .A2 (nx882)) ;
    dffr regPage2Map_reg_Q_14 (.Q (outputRegPage2[14]), .QB (nx699), .D (nx423)
         , .CLK (clk), .R (rst)) ;
    nand02 ix424 (.Y (nx423), .A0 (nx695), .A1 (nx697)) ;
    nand02 ix696 (.Y (nx695), .A0 (outputRegPage2[14]), .A1 (nx595)) ;
    nand03 ix698 (.Y (nx697), .A0 (windowBus[14]), .A1 (nx599), .A2 (nx882)) ;
    dffr regPage2Map_reg_Q_15 (.Q (outputRegPage2[15]), .QB (nx706), .D (nx443)
         , .CLK (clk), .R (rst)) ;
    nand02 ix444 (.Y (nx443), .A0 (nx702), .A1 (nx704)) ;
    nand02 ix703 (.Y (nx702), .A0 (outputRegPage2[15]), .A1 (nx595)) ;
    nand03 ix705 (.Y (nx704), .A0 (windowBus[15]), .A1 (nx599), .A2 (nx882)) ;
    dffr regPage1Map_reg_Q_0 (.Q (outputRegPage1[0]), .QB (nx717), .D (nx133), .CLK (
         clk), .R (rst)) ;
    nand02 ix134 (.Y (nx133), .A0 (nx709), .A1 (nx713)) ;
    nand02 ix710 (.Y (nx709), .A0 (outputRegPage1[0]), .A1 (nx856)) ;
    nor02_2x ix712 (.Y (nx711), .A0 (nx870), .A1 (page1ReadBusOrPage2)) ;
    nand03 ix714 (.Y (nx713), .A0 (windowBus[0]), .A1 (nx860), .A2 (nx870)) ;
    inv01 ix716 (.Y (nx715), .A (page1ReadBusOrPage2)) ;
    dffr regPage1Map_reg_Q_1 (.Q (outputRegPage1[1]), .QB (nx724), .D (nx153), .CLK (
         clk), .R (rst)) ;
    nand02 ix154 (.Y (nx153), .A0 (nx720), .A1 (nx722)) ;
    nand02 ix721 (.Y (nx720), .A0 (outputRegPage1[1]), .A1 (nx856)) ;
    nand03 ix723 (.Y (nx722), .A0 (windowBus[1]), .A1 (nx860), .A2 (nx870)) ;
    dffr regPage1Map_reg_Q_2 (.Q (outputRegPage1[2]), .QB (nx731), .D (nx173), .CLK (
         clk), .R (rst)) ;
    nand02 ix174 (.Y (nx173), .A0 (nx727), .A1 (nx729)) ;
    nand02 ix728 (.Y (nx727), .A0 (outputRegPage1[2]), .A1 (nx856)) ;
    nand03 ix730 (.Y (nx729), .A0 (windowBus[2]), .A1 (nx860), .A2 (nx870)) ;
    dffr regPage1Map_reg_Q_3 (.Q (outputRegPage1[3]), .QB (nx738), .D (nx193), .CLK (
         clk), .R (rst)) ;
    nand02 ix194 (.Y (nx193), .A0 (nx734), .A1 (nx736)) ;
    nand02 ix735 (.Y (nx734), .A0 (outputRegPage1[3]), .A1 (nx856)) ;
    nand03 ix737 (.Y (nx736), .A0 (windowBus[3]), .A1 (nx860), .A2 (nx870)) ;
    dffr regPage1Map_reg_Q_4 (.Q (outputRegPage1[4]), .QB (nx745), .D (nx213), .CLK (
         clk), .R (rst)) ;
    nand02 ix214 (.Y (nx213), .A0 (nx741), .A1 (nx743)) ;
    nand02 ix742 (.Y (nx741), .A0 (outputRegPage1[4]), .A1 (nx856)) ;
    nand03 ix744 (.Y (nx743), .A0 (windowBus[4]), .A1 (nx860), .A2 (nx870)) ;
    dffr regPage1Map_reg_Q_5 (.Q (outputRegPage1[5]), .QB (nx752), .D (nx233), .CLK (
         clk), .R (rst)) ;
    nand02 ix234 (.Y (nx233), .A0 (nx748), .A1 (nx750)) ;
    nand02 ix749 (.Y (nx748), .A0 (outputRegPage1[5]), .A1 (nx856)) ;
    nand03 ix751 (.Y (nx750), .A0 (windowBus[5]), .A1 (nx860), .A2 (nx870)) ;
    dffr regPage1Map_reg_Q_6 (.Q (outputRegPage1[6]), .QB (nx759), .D (nx253), .CLK (
         clk), .R (rst)) ;
    nand02 ix254 (.Y (nx253), .A0 (nx755), .A1 (nx757)) ;
    nand02 ix756 (.Y (nx755), .A0 (outputRegPage1[6]), .A1 (nx856)) ;
    nand03 ix758 (.Y (nx757), .A0 (windowBus[6]), .A1 (nx862), .A2 (nx872)) ;
    dffr regPage1Map_reg_Q_7 (.Q (outputRegPage1[7]), .QB (nx766), .D (nx273), .CLK (
         clk), .R (rst)) ;
    nand02 ix274 (.Y (nx273), .A0 (nx762), .A1 (nx764)) ;
    nand02 ix763 (.Y (nx762), .A0 (outputRegPage1[7]), .A1 (nx858)) ;
    nand03 ix765 (.Y (nx764), .A0 (windowBus[7]), .A1 (nx862), .A2 (nx872)) ;
    dffr regPage1Map_reg_Q_8 (.Q (outputRegPage1[8]), .QB (nx773), .D (nx293), .CLK (
         clk), .R (rst)) ;
    nand02 ix294 (.Y (nx293), .A0 (nx769), .A1 (nx771)) ;
    nand02 ix770 (.Y (nx769), .A0 (outputRegPage1[8]), .A1 (nx858)) ;
    nand03 ix772 (.Y (nx771), .A0 (windowBus[8]), .A1 (nx862), .A2 (nx872)) ;
    dffr regPage1Map_reg_Q_9 (.Q (outputRegPage1[9]), .QB (nx780), .D (nx313), .CLK (
         clk), .R (rst)) ;
    nand02 ix314 (.Y (nx313), .A0 (nx776), .A1 (nx778)) ;
    nand02 ix777 (.Y (nx776), .A0 (outputRegPage1[9]), .A1 (nx858)) ;
    nand03 ix779 (.Y (nx778), .A0 (windowBus[9]), .A1 (nx862), .A2 (nx872)) ;
    dffr regPage1Map_reg_Q_10 (.Q (outputRegPage1[10]), .QB (nx787), .D (nx333)
         , .CLK (clk), .R (rst)) ;
    nand02 ix334 (.Y (nx333), .A0 (nx783), .A1 (nx785)) ;
    nand02 ix784 (.Y (nx783), .A0 (outputRegPage1[10]), .A1 (nx858)) ;
    nand03 ix786 (.Y (nx785), .A0 (windowBus[10]), .A1 (nx862), .A2 (nx872)) ;
    dffr regPage1Map_reg_Q_11 (.Q (outputRegPage1[11]), .QB (nx794), .D (nx353)
         , .CLK (clk), .R (rst)) ;
    nand02 ix354 (.Y (nx353), .A0 (nx790), .A1 (nx792)) ;
    nand02 ix791 (.Y (nx790), .A0 (outputRegPage1[11]), .A1 (nx858)) ;
    nand03 ix793 (.Y (nx792), .A0 (windowBus[11]), .A1 (nx862), .A2 (nx872)) ;
    dffr regPage1Map_reg_Q_12 (.Q (outputRegPage1[12]), .QB (nx801), .D (nx373)
         , .CLK (clk), .R (rst)) ;
    nand02 ix374 (.Y (nx373), .A0 (nx797), .A1 (nx799)) ;
    nand02 ix798 (.Y (nx797), .A0 (outputRegPage1[12]), .A1 (nx858)) ;
    nand03 ix800 (.Y (nx799), .A0 (windowBus[12]), .A1 (nx715), .A2 (nx872)) ;
    dffr regPage1Map_reg_Q_13 (.Q (outputRegPage1[13]), .QB (nx808), .D (nx393)
         , .CLK (clk), .R (rst)) ;
    nand02 ix394 (.Y (nx393), .A0 (nx804), .A1 (nx806)) ;
    nand02 ix805 (.Y (nx804), .A0 (outputRegPage1[13]), .A1 (nx858)) ;
    nand03 ix807 (.Y (nx806), .A0 (windowBus[13]), .A1 (nx715), .A2 (nx874)) ;
    dffr regPage1Map_reg_Q_14 (.Q (outputRegPage1[14]), .QB (nx815), .D (nx413)
         , .CLK (clk), .R (rst)) ;
    nand02 ix414 (.Y (nx413), .A0 (nx811), .A1 (nx813)) ;
    nand02 ix812 (.Y (nx811), .A0 (outputRegPage1[14]), .A1 (nx711)) ;
    nand03 ix814 (.Y (nx813), .A0 (windowBus[14]), .A1 (nx715), .A2 (nx874)) ;
    dffr regPage1Map_reg_Q_15 (.Q (outputRegPage1[15]), .QB (nx822), .D (nx433)
         , .CLK (clk), .R (rst)) ;
    nand02 ix434 (.Y (nx433), .A0 (nx818), .A1 (nx820)) ;
    nand02 ix819 (.Y (nx818), .A0 (outputRegPage1[15]), .A1 (nx711)) ;
    nand03 ix821 (.Y (nx820), .A0 (windowBus[15]), .A1 (nx715), .A2 (nx874)) ;
    mux21 ix25 (.Y (outRegPage[0]), .A0 (nx717), .A1 (nx601), .S0 (pageTurn)) ;
    mux21 ix45 (.Y (outRegPage[1]), .A0 (nx724), .A1 (nx608), .S0 (pageTurn)) ;
    mux21 ix65 (.Y (outRegPage[2]), .A0 (nx731), .A1 (nx615), .S0 (pageTurn)) ;
    mux21 ix85 (.Y (outRegPage[3]), .A0 (nx738), .A1 (nx622), .S0 (pageTurn)) ;
    mux21 ix105 (.Y (outRegPage[4]), .A0 (nx745), .A1 (nx629), .S0 (pageTurn)) ;
    mux21 ix125 (.Y (outRegPage[5]), .A0 (nx752), .A1 (nx636), .S0 (pageTurn)) ;
    mux21 ix145 (.Y (outRegPage[6]), .A0 (nx759), .A1 (nx643), .S0 (pageTurn)) ;
    mux21 ix165 (.Y (outRegPage[7]), .A0 (nx766), .A1 (nx650), .S0 (pageTurn)) ;
    mux21 ix185 (.Y (outRegPage[8]), .A0 (nx773), .A1 (nx657), .S0 (pageTurn)) ;
    mux21 ix205 (.Y (outRegPage[9]), .A0 (nx780), .A1 (nx664), .S0 (pageTurn)) ;
    mux21 ix225 (.Y (outRegPage[10]), .A0 (nx787), .A1 (nx671), .S0 (pageTurn)
          ) ;
    mux21 ix245 (.Y (outRegPage[11]), .A0 (nx794), .A1 (nx678), .S0 (pageTurn)
          ) ;
    mux21 ix265 (.Y (outRegPage[12]), .A0 (nx801), .A1 (nx685), .S0 (pageTurn)
          ) ;
    mux21 ix285 (.Y (outRegPage[13]), .A0 (nx808), .A1 (nx692), .S0 (pageTurn)
          ) ;
    mux21 ix305 (.Y (outRegPage[14]), .A0 (nx815), .A1 (nx699), .S0 (pageTurn)
          ) ;
    mux21 ix325 (.Y (outRegPage[15]), .A0 (nx822), .A1 (nx706), .S0 (pageTurn)
          ) ;
    inv01 ix845 (.Y (nx846), .A (nx886)) ;
    nor02_2x ix847 (.Y (nx848), .A0 (nx882), .A1 (page2ReadBusOrPage1)) ;
    nor02_2x ix849 (.Y (nx850), .A0 (nx882), .A1 (page2ReadBusOrPage1)) ;
    inv01 ix851 (.Y (nx852), .A (page2ReadBusOrPage1)) ;
    inv01 ix853 (.Y (nx854), .A (page2ReadBusOrPage1)) ;
    nor02_2x ix855 (.Y (nx856), .A0 (nx874), .A1 (page1ReadBusOrPage2)) ;
    nor02_2x ix857 (.Y (nx858), .A0 (nx874), .A1 (page1ReadBusOrPage2)) ;
    inv01 ix859 (.Y (nx860), .A (page1ReadBusOrPage2)) ;
    inv01 ix861 (.Y (nx862), .A (page1ReadBusOrPage2)) ;
    inv01 ix867 (.Y (nx868), .A (enableRegPage1)) ;
    inv02 ix869 (.Y (nx870), .A (nx868)) ;
    inv02 ix871 (.Y (nx872), .A (nx868)) ;
    inv02 ix873 (.Y (nx874), .A (nx868)) ;
    inv01 ix875 (.Y (nx876), .A (enableRegPage2)) ;
    inv02 ix877 (.Y (nx878), .A (nx876)) ;
    inv02 ix879 (.Y (nx880), .A (nx876)) ;
    inv02 ix881 (.Y (nx882), .A (nx876)) ;
    inv02 ix883 (.Y (nx884), .A (nx890)) ;
    inv02 ix885 (.Y (nx886), .A (nx890)) ;
    inv02 ix887 (.Y (nx888), .A (enableRegFilter)) ;
    inv02 ix889 (.Y (nx890), .A (enableRegFilter)) ;
endmodule


module RegUnit_8_16_unfolded0 ( filterBus, windowBus, regPage1NextUnit, 
                                regPage2NextUnit, clk, rst, enableRegPage1, 
                                enableRegPage2, enableRegFilter, 
                                page1ReadBusOrPage2, page2ReadBusOrPage1, 
                                pageTurn, outRegPage, outputRegPage1, 
                                outputRegPage2, outFilter ) ;

    input [7:0]filterBus ;
    input [15:0]windowBus ;
    input [15:0]regPage1NextUnit ;
    input [15:0]regPage2NextUnit ;
    input clk ;
    input rst ;
    input enableRegPage1 ;
    input enableRegPage2 ;
    input enableRegFilter ;
    input page1ReadBusOrPage2 ;
    input page2ReadBusOrPage1 ;
    input pageTurn ;
    output [15:0]outRegPage ;
    output [15:0]outputRegPage1 ;
    output [15:0]outputRegPage2 ;
    output [7:0]outFilter ;

    wire nx345, nx355, nx365, nx375, nx385, nx395, nx405, nx415, nx425, nx435, 
         nx445, nx455, nx465, nx475, nx485, nx495, nx505, nx515, nx525, nx535, 
         nx545, nx555, nx565, nx575, nx585, nx595, nx605, nx615, nx625, nx635, 
         nx645, nx655, nx665, nx675, nx685, nx695, nx705, nx715, nx725, nx735, 
         nx747, nx751, nx756, nx758, nx763, nx765, nx770, nx772, nx777, nx779, 
         nx784, nx786, nx791, nx793, nx798, nx800, nx805, nx807, nx809, nx811, 
         nx814, nx816, nx818, nx821, nx823, nx825, nx828, nx830, nx832, nx835, 
         nx837, nx839, nx842, nx844, nx846, nx849, nx851, nx853, nx856, nx858, 
         nx860, nx863, nx865, nx867, nx870, nx872, nx874, nx877, nx879, nx881, 
         nx884, nx886, nx888, nx891, nx893, nx895, nx898, nx900, nx902, nx905, 
         nx907, nx909, nx912, nx914, nx916, nx919, nx921, nx923, nx925, nx928, 
         nx930, nx932, nx935, nx937, nx939, nx942, nx944, nx946, nx949, nx951, 
         nx953, nx956, nx958, nx960, nx963, nx965, nx967, nx970, nx972, nx974, 
         nx977, nx979, nx981, nx984, nx986, nx988, nx991, nx993, nx995, nx998, 
         nx1000, nx1002, nx1005, nx1007, nx1009, nx1012, nx1014, nx1016, nx1019, 
         nx1021, nx1023, nx1026, nx1028, nx1030, nx1054, nx1056, nx1058, nx1060, 
         nx1062, nx1064, nx1066, nx1068, nx1070, nx1072, nx1074, nx1076, nx1078, 
         nx1084, nx1086, nx1088, nx1090;
    wire [7:0] \$dummy ;




    dffr regFilterMap_reg_Q_0 (.Q (outFilter[0]), .QB (\$dummy [0]), .D (nx665)
         , .CLK (clk), .R (rst)) ;
    nand02 ix666 (.Y (nx665), .A0 (nx747), .A1 (nx751)) ;
    nand02 ix748 (.Y (nx747), .A0 (outFilter[0]), .A1 (nx1088)) ;
    nand02 ix752 (.Y (nx751), .A0 (filterBus[0]), .A1 (nx1084)) ;
    dffr regFilterMap_reg_Q_1 (.Q (outFilter[1]), .QB (\$dummy [1]), .D (nx675)
         , .CLK (clk), .R (rst)) ;
    nand02 ix676 (.Y (nx675), .A0 (nx756), .A1 (nx758)) ;
    nand02 ix757 (.Y (nx756), .A0 (outFilter[1]), .A1 (nx1088)) ;
    nand02 ix759 (.Y (nx758), .A0 (filterBus[1]), .A1 (nx1084)) ;
    dffr regFilterMap_reg_Q_2 (.Q (outFilter[2]), .QB (\$dummy [2]), .D (nx685)
         , .CLK (clk), .R (rst)) ;
    nand02 ix686 (.Y (nx685), .A0 (nx763), .A1 (nx765)) ;
    nand02 ix764 (.Y (nx763), .A0 (outFilter[2]), .A1 (nx1088)) ;
    nand02 ix766 (.Y (nx765), .A0 (filterBus[2]), .A1 (nx1084)) ;
    dffr regFilterMap_reg_Q_3 (.Q (outFilter[3]), .QB (\$dummy [3]), .D (nx695)
         , .CLK (clk), .R (rst)) ;
    nand02 ix696 (.Y (nx695), .A0 (nx770), .A1 (nx772)) ;
    nand02 ix771 (.Y (nx770), .A0 (outFilter[3]), .A1 (nx1088)) ;
    nand02 ix773 (.Y (nx772), .A0 (filterBus[3]), .A1 (nx1084)) ;
    dffr regFilterMap_reg_Q_4 (.Q (outFilter[4]), .QB (\$dummy [4]), .D (nx705)
         , .CLK (clk), .R (rst)) ;
    nand02 ix706 (.Y (nx705), .A0 (nx777), .A1 (nx779)) ;
    nand02 ix778 (.Y (nx777), .A0 (outFilter[4]), .A1 (nx1088)) ;
    nand02 ix780 (.Y (nx779), .A0 (filterBus[4]), .A1 (nx1084)) ;
    dffr regFilterMap_reg_Q_5 (.Q (outFilter[5]), .QB (\$dummy [5]), .D (nx715)
         , .CLK (clk), .R (rst)) ;
    nand02 ix716 (.Y (nx715), .A0 (nx784), .A1 (nx786)) ;
    nand02 ix785 (.Y (nx784), .A0 (outFilter[5]), .A1 (nx1088)) ;
    nand02 ix787 (.Y (nx786), .A0 (filterBus[5]), .A1 (nx1084)) ;
    dffr regFilterMap_reg_Q_6 (.Q (outFilter[6]), .QB (\$dummy [6]), .D (nx725)
         , .CLK (clk), .R (rst)) ;
    nand02 ix726 (.Y (nx725), .A0 (nx791), .A1 (nx793)) ;
    nand02 ix792 (.Y (nx791), .A0 (outFilter[6]), .A1 (nx1088)) ;
    nand02 ix794 (.Y (nx793), .A0 (filterBus[6]), .A1 (nx1084)) ;
    dffr regFilterMap_reg_Q_7 (.Q (outFilter[7]), .QB (\$dummy [7]), .D (nx735)
         , .CLK (clk), .R (rst)) ;
    nand02 ix736 (.Y (nx735), .A0 (nx798), .A1 (nx800)) ;
    nand02 ix799 (.Y (nx798), .A0 (outFilter[7]), .A1 (nx1054)) ;
    nand02 ix801 (.Y (nx800), .A0 (filterBus[7]), .A1 (nx1086)) ;
    dffr regPage2Map_reg_Q_0 (.Q (outputRegPage2[0]), .QB (nx811), .D (nx355), .CLK (
         clk), .R (rst)) ;
    oai21 ix356 (.Y (nx355), .A0 (nx805), .A1 (nx1058), .B0 (nx809)) ;
    mux21 ix806 (.Y (nx805), .A0 (windowBus[0]), .A1 (regPage1NextUnit[0]), .S0 (
          page2ReadBusOrPage1)) ;
    nor02_2x ix808 (.Y (nx807), .A0 (enableRegPage2), .A1 (page2ReadBusOrPage1)
             ) ;
    nand02 ix810 (.Y (nx809), .A0 (outputRegPage2[0]), .A1 (nx1058)) ;
    dffr regPage2Map_reg_Q_1 (.Q (outputRegPage2[1]), .QB (nx818), .D (nx375), .CLK (
         clk), .R (rst)) ;
    oai21 ix376 (.Y (nx375), .A0 (nx814), .A1 (nx1058), .B0 (nx816)) ;
    mux21 ix815 (.Y (nx814), .A0 (windowBus[1]), .A1 (regPage1NextUnit[1]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix817 (.Y (nx816), .A0 (outputRegPage2[1]), .A1 (nx1058)) ;
    dffr regPage2Map_reg_Q_2 (.Q (outputRegPage2[2]), .QB (nx825), .D (nx395), .CLK (
         clk), .R (rst)) ;
    oai21 ix396 (.Y (nx395), .A0 (nx821), .A1 (nx1058), .B0 (nx823)) ;
    mux21 ix822 (.Y (nx821), .A0 (windowBus[2]), .A1 (regPage1NextUnit[2]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix824 (.Y (nx823), .A0 (outputRegPage2[2]), .A1 (nx1058)) ;
    dffr regPage2Map_reg_Q_3 (.Q (outputRegPage2[3]), .QB (nx832), .D (nx415), .CLK (
         clk), .R (rst)) ;
    oai21 ix416 (.Y (nx415), .A0 (nx828), .A1 (nx1058), .B0 (nx830)) ;
    mux21 ix829 (.Y (nx828), .A0 (windowBus[3]), .A1 (regPage1NextUnit[3]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix831 (.Y (nx830), .A0 (outputRegPage2[3]), .A1 (nx1060)) ;
    dffr regPage2Map_reg_Q_4 (.Q (outputRegPage2[4]), .QB (nx839), .D (nx435), .CLK (
         clk), .R (rst)) ;
    oai21 ix436 (.Y (nx435), .A0 (nx835), .A1 (nx1060), .B0 (nx837)) ;
    mux21 ix836 (.Y (nx835), .A0 (windowBus[4]), .A1 (regPage1NextUnit[4]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix838 (.Y (nx837), .A0 (outputRegPage2[4]), .A1 (nx1060)) ;
    dffr regPage2Map_reg_Q_5 (.Q (outputRegPage2[5]), .QB (nx846), .D (nx455), .CLK (
         clk), .R (rst)) ;
    oai21 ix456 (.Y (nx455), .A0 (nx842), .A1 (nx1060), .B0 (nx844)) ;
    mux21 ix843 (.Y (nx842), .A0 (windowBus[5]), .A1 (regPage1NextUnit[5]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix845 (.Y (nx844), .A0 (outputRegPage2[5]), .A1 (nx1060)) ;
    dffr regPage2Map_reg_Q_6 (.Q (outputRegPage2[6]), .QB (nx853), .D (nx475), .CLK (
         clk), .R (rst)) ;
    oai21 ix476 (.Y (nx475), .A0 (nx849), .A1 (nx1060), .B0 (nx851)) ;
    mux21 ix850 (.Y (nx849), .A0 (windowBus[6]), .A1 (regPage1NextUnit[6]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix852 (.Y (nx851), .A0 (outputRegPage2[6]), .A1 (nx1060)) ;
    dffr regPage2Map_reg_Q_7 (.Q (outputRegPage2[7]), .QB (nx860), .D (nx495), .CLK (
         clk), .R (rst)) ;
    oai21 ix496 (.Y (nx495), .A0 (nx856), .A1 (nx1062), .B0 (nx858)) ;
    mux21 ix857 (.Y (nx856), .A0 (windowBus[7]), .A1 (regPage1NextUnit[7]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix859 (.Y (nx858), .A0 (outputRegPage2[7]), .A1 (nx1062)) ;
    dffr regPage2Map_reg_Q_8 (.Q (outputRegPage2[8]), .QB (nx867), .D (nx515), .CLK (
         clk), .R (rst)) ;
    oai21 ix516 (.Y (nx515), .A0 (nx863), .A1 (nx1062), .B0 (nx865)) ;
    mux21 ix864 (.Y (nx863), .A0 (windowBus[8]), .A1 (regPage1NextUnit[8]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix866 (.Y (nx865), .A0 (outputRegPage2[8]), .A1 (nx1062)) ;
    dffr regPage2Map_reg_Q_9 (.Q (outputRegPage2[9]), .QB (nx874), .D (nx535), .CLK (
         clk), .R (rst)) ;
    oai21 ix536 (.Y (nx535), .A0 (nx870), .A1 (nx1062), .B0 (nx872)) ;
    mux21 ix871 (.Y (nx870), .A0 (windowBus[9]), .A1 (regPage1NextUnit[9]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix873 (.Y (nx872), .A0 (outputRegPage2[9]), .A1 (nx1062)) ;
    dffr regPage2Map_reg_Q_10 (.Q (outputRegPage2[10]), .QB (nx881), .D (nx555)
         , .CLK (clk), .R (rst)) ;
    oai21 ix556 (.Y (nx555), .A0 (nx877), .A1 (nx1062), .B0 (nx879)) ;
    mux21 ix878 (.Y (nx877), .A0 (windowBus[10]), .A1 (regPage1NextUnit[10]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix880 (.Y (nx879), .A0 (outputRegPage2[10]), .A1 (nx1064)) ;
    dffr regPage2Map_reg_Q_11 (.Q (outputRegPage2[11]), .QB (nx888), .D (nx575)
         , .CLK (clk), .R (rst)) ;
    oai21 ix576 (.Y (nx575), .A0 (nx884), .A1 (nx1064), .B0 (nx886)) ;
    mux21 ix885 (.Y (nx884), .A0 (windowBus[11]), .A1 (regPage1NextUnit[11]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix887 (.Y (nx886), .A0 (outputRegPage2[11]), .A1 (nx1064)) ;
    dffr regPage2Map_reg_Q_12 (.Q (outputRegPage2[12]), .QB (nx895), .D (nx595)
         , .CLK (clk), .R (rst)) ;
    oai21 ix596 (.Y (nx595), .A0 (nx891), .A1 (nx1064), .B0 (nx893)) ;
    mux21 ix892 (.Y (nx891), .A0 (windowBus[12]), .A1 (regPage1NextUnit[12]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix894 (.Y (nx893), .A0 (outputRegPage2[12]), .A1 (nx1064)) ;
    dffr regPage2Map_reg_Q_13 (.Q (outputRegPage2[13]), .QB (nx902), .D (nx615)
         , .CLK (clk), .R (rst)) ;
    oai21 ix616 (.Y (nx615), .A0 (nx898), .A1 (nx1064), .B0 (nx900)) ;
    mux21 ix899 (.Y (nx898), .A0 (windowBus[13]), .A1 (regPage1NextUnit[13]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix901 (.Y (nx900), .A0 (outputRegPage2[13]), .A1 (nx1064)) ;
    dffr regPage2Map_reg_Q_14 (.Q (outputRegPage2[14]), .QB (nx909), .D (nx635)
         , .CLK (clk), .R (rst)) ;
    oai21 ix636 (.Y (nx635), .A0 (nx905), .A1 (nx1066), .B0 (nx907)) ;
    mux21 ix906 (.Y (nx905), .A0 (windowBus[14]), .A1 (regPage1NextUnit[14]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix908 (.Y (nx907), .A0 (outputRegPage2[14]), .A1 (nx1066)) ;
    dffr regPage2Map_reg_Q_15 (.Q (outputRegPage2[15]), .QB (nx916), .D (nx655)
         , .CLK (clk), .R (rst)) ;
    oai21 ix656 (.Y (nx655), .A0 (nx912), .A1 (nx1066), .B0 (nx914)) ;
    mux21 ix913 (.Y (nx912), .A0 (windowBus[15]), .A1 (regPage1NextUnit[15]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix915 (.Y (nx914), .A0 (outputRegPage2[15]), .A1 (nx1066)) ;
    dffr regPage1Map_reg_Q_0 (.Q (outputRegPage1[0]), .QB (nx925), .D (nx345), .CLK (
         clk), .R (rst)) ;
    oai21 ix346 (.Y (nx345), .A0 (nx919), .A1 (nx1070), .B0 (nx923)) ;
    mux21 ix920 (.Y (nx919), .A0 (windowBus[0]), .A1 (regPage2NextUnit[0]), .S0 (
          page1ReadBusOrPage2)) ;
    nor02_2x ix922 (.Y (nx921), .A0 (enableRegPage1), .A1 (page1ReadBusOrPage2)
             ) ;
    nand02 ix924 (.Y (nx923), .A0 (outputRegPage1[0]), .A1 (nx1070)) ;
    dffr regPage1Map_reg_Q_1 (.Q (outputRegPage1[1]), .QB (nx932), .D (nx365), .CLK (
         clk), .R (rst)) ;
    oai21 ix366 (.Y (nx365), .A0 (nx928), .A1 (nx1070), .B0 (nx930)) ;
    mux21 ix929 (.Y (nx928), .A0 (windowBus[1]), .A1 (regPage2NextUnit[1]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix931 (.Y (nx930), .A0 (outputRegPage1[1]), .A1 (nx1070)) ;
    dffr regPage1Map_reg_Q_2 (.Q (outputRegPage1[2]), .QB (nx939), .D (nx385), .CLK (
         clk), .R (rst)) ;
    oai21 ix386 (.Y (nx385), .A0 (nx935), .A1 (nx1070), .B0 (nx937)) ;
    mux21 ix936 (.Y (nx935), .A0 (windowBus[2]), .A1 (regPage2NextUnit[2]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix938 (.Y (nx937), .A0 (outputRegPage1[2]), .A1 (nx1070)) ;
    dffr regPage1Map_reg_Q_3 (.Q (outputRegPage1[3]), .QB (nx946), .D (nx405), .CLK (
         clk), .R (rst)) ;
    oai21 ix406 (.Y (nx405), .A0 (nx942), .A1 (nx1070), .B0 (nx944)) ;
    mux21 ix943 (.Y (nx942), .A0 (windowBus[3]), .A1 (regPage2NextUnit[3]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix945 (.Y (nx944), .A0 (outputRegPage1[3]), .A1 (nx1072)) ;
    dffr regPage1Map_reg_Q_4 (.Q (outputRegPage1[4]), .QB (nx953), .D (nx425), .CLK (
         clk), .R (rst)) ;
    oai21 ix426 (.Y (nx425), .A0 (nx949), .A1 (nx1072), .B0 (nx951)) ;
    mux21 ix950 (.Y (nx949), .A0 (windowBus[4]), .A1 (regPage2NextUnit[4]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix952 (.Y (nx951), .A0 (outputRegPage1[4]), .A1 (nx1072)) ;
    dffr regPage1Map_reg_Q_5 (.Q (outputRegPage1[5]), .QB (nx960), .D (nx445), .CLK (
         clk), .R (rst)) ;
    oai21 ix446 (.Y (nx445), .A0 (nx956), .A1 (nx1072), .B0 (nx958)) ;
    mux21 ix957 (.Y (nx956), .A0 (windowBus[5]), .A1 (regPage2NextUnit[5]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix959 (.Y (nx958), .A0 (outputRegPage1[5]), .A1 (nx1072)) ;
    dffr regPage1Map_reg_Q_6 (.Q (outputRegPage1[6]), .QB (nx967), .D (nx465), .CLK (
         clk), .R (rst)) ;
    oai21 ix466 (.Y (nx465), .A0 (nx963), .A1 (nx1072), .B0 (nx965)) ;
    mux21 ix964 (.Y (nx963), .A0 (windowBus[6]), .A1 (regPage2NextUnit[6]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix966 (.Y (nx965), .A0 (outputRegPage1[6]), .A1 (nx1072)) ;
    dffr regPage1Map_reg_Q_7 (.Q (outputRegPage1[7]), .QB (nx974), .D (nx485), .CLK (
         clk), .R (rst)) ;
    oai21 ix486 (.Y (nx485), .A0 (nx970), .A1 (nx1074), .B0 (nx972)) ;
    mux21 ix971 (.Y (nx970), .A0 (windowBus[7]), .A1 (regPage2NextUnit[7]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix973 (.Y (nx972), .A0 (outputRegPage1[7]), .A1 (nx1074)) ;
    dffr regPage1Map_reg_Q_8 (.Q (outputRegPage1[8]), .QB (nx981), .D (nx505), .CLK (
         clk), .R (rst)) ;
    oai21 ix506 (.Y (nx505), .A0 (nx977), .A1 (nx1074), .B0 (nx979)) ;
    mux21 ix978 (.Y (nx977), .A0 (windowBus[8]), .A1 (regPage2NextUnit[8]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix980 (.Y (nx979), .A0 (outputRegPage1[8]), .A1 (nx1074)) ;
    dffr regPage1Map_reg_Q_9 (.Q (outputRegPage1[9]), .QB (nx988), .D (nx525), .CLK (
         clk), .R (rst)) ;
    oai21 ix526 (.Y (nx525), .A0 (nx984), .A1 (nx1074), .B0 (nx986)) ;
    mux21 ix985 (.Y (nx984), .A0 (windowBus[9]), .A1 (regPage2NextUnit[9]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix987 (.Y (nx986), .A0 (outputRegPage1[9]), .A1 (nx1074)) ;
    dffr regPage1Map_reg_Q_10 (.Q (outputRegPage1[10]), .QB (nx995), .D (nx545)
         , .CLK (clk), .R (rst)) ;
    oai21 ix546 (.Y (nx545), .A0 (nx991), .A1 (nx1074), .B0 (nx993)) ;
    mux21 ix992 (.Y (nx991), .A0 (windowBus[10]), .A1 (regPage2NextUnit[10]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix994 (.Y (nx993), .A0 (outputRegPage1[10]), .A1 (nx1076)) ;
    dffr regPage1Map_reg_Q_11 (.Q (outputRegPage1[11]), .QB (nx1002), .D (nx565)
         , .CLK (clk), .R (rst)) ;
    oai21 ix566 (.Y (nx565), .A0 (nx998), .A1 (nx1076), .B0 (nx1000)) ;
    mux21 ix999 (.Y (nx998), .A0 (windowBus[11]), .A1 (regPage2NextUnit[11]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix1001 (.Y (nx1000), .A0 (outputRegPage1[11]), .A1 (nx1076)) ;
    dffr regPage1Map_reg_Q_12 (.Q (outputRegPage1[12]), .QB (nx1009), .D (nx585)
         , .CLK (clk), .R (rst)) ;
    oai21 ix586 (.Y (nx585), .A0 (nx1005), .A1 (nx1076), .B0 (nx1007)) ;
    mux21 ix1006 (.Y (nx1005), .A0 (windowBus[12]), .A1 (regPage2NextUnit[12]), 
          .S0 (page1ReadBusOrPage2)) ;
    nand02 ix1008 (.Y (nx1007), .A0 (outputRegPage1[12]), .A1 (nx1076)) ;
    dffr regPage1Map_reg_Q_13 (.Q (outputRegPage1[13]), .QB (nx1016), .D (nx605)
         , .CLK (clk), .R (rst)) ;
    oai21 ix606 (.Y (nx605), .A0 (nx1012), .A1 (nx1076), .B0 (nx1014)) ;
    mux21 ix1013 (.Y (nx1012), .A0 (windowBus[13]), .A1 (regPage2NextUnit[13]), 
          .S0 (page1ReadBusOrPage2)) ;
    nand02 ix1015 (.Y (nx1014), .A0 (outputRegPage1[13]), .A1 (nx1076)) ;
    dffr regPage1Map_reg_Q_14 (.Q (outputRegPage1[14]), .QB (nx1023), .D (nx625)
         , .CLK (clk), .R (rst)) ;
    oai21 ix626 (.Y (nx625), .A0 (nx1019), .A1 (nx1078), .B0 (nx1021)) ;
    mux21 ix1020 (.Y (nx1019), .A0 (windowBus[14]), .A1 (regPage2NextUnit[14]), 
          .S0 (page1ReadBusOrPage2)) ;
    nand02 ix1022 (.Y (nx1021), .A0 (outputRegPage1[14]), .A1 (nx1078)) ;
    dffr regPage1Map_reg_Q_15 (.Q (outputRegPage1[15]), .QB (nx1030), .D (nx645)
         , .CLK (clk), .R (rst)) ;
    oai21 ix646 (.Y (nx645), .A0 (nx1026), .A1 (nx1078), .B0 (nx1028)) ;
    mux21 ix1027 (.Y (nx1026), .A0 (windowBus[15]), .A1 (regPage2NextUnit[15]), 
          .S0 (page1ReadBusOrPage2)) ;
    nand02 ix1029 (.Y (nx1028), .A0 (outputRegPage1[15]), .A1 (nx1078)) ;
    mux21 ix33 (.Y (outRegPage[0]), .A0 (nx925), .A1 (nx811), .S0 (pageTurn)) ;
    mux21 ix61 (.Y (outRegPage[1]), .A0 (nx932), .A1 (nx818), .S0 (pageTurn)) ;
    mux21 ix89 (.Y (outRegPage[2]), .A0 (nx939), .A1 (nx825), .S0 (pageTurn)) ;
    mux21 ix117 (.Y (outRegPage[3]), .A0 (nx946), .A1 (nx832), .S0 (pageTurn)) ;
    mux21 ix145 (.Y (outRegPage[4]), .A0 (nx953), .A1 (nx839), .S0 (pageTurn)) ;
    mux21 ix173 (.Y (outRegPage[5]), .A0 (nx960), .A1 (nx846), .S0 (pageTurn)) ;
    mux21 ix201 (.Y (outRegPage[6]), .A0 (nx967), .A1 (nx853), .S0 (pageTurn)) ;
    mux21 ix229 (.Y (outRegPage[7]), .A0 (nx974), .A1 (nx860), .S0 (pageTurn)) ;
    mux21 ix257 (.Y (outRegPage[8]), .A0 (nx981), .A1 (nx867), .S0 (pageTurn)) ;
    mux21 ix285 (.Y (outRegPage[9]), .A0 (nx988), .A1 (nx874), .S0 (pageTurn)) ;
    mux21 ix313 (.Y (outRegPage[10]), .A0 (nx995), .A1 (nx881), .S0 (pageTurn)
          ) ;
    mux21 ix341 (.Y (outRegPage[11]), .A0 (nx1002), .A1 (nx888), .S0 (pageTurn)
          ) ;
    mux21 ix369 (.Y (outRegPage[12]), .A0 (nx1009), .A1 (nx895), .S0 (pageTurn)
          ) ;
    mux21 ix397 (.Y (outRegPage[13]), .A0 (nx1016), .A1 (nx902), .S0 (pageTurn)
          ) ;
    mux21 ix425 (.Y (outRegPage[14]), .A0 (nx1023), .A1 (nx909), .S0 (pageTurn)
          ) ;
    mux21 ix453 (.Y (outRegPage[15]), .A0 (nx1030), .A1 (nx916), .S0 (pageTurn)
          ) ;
    inv01 ix1053 (.Y (nx1054), .A (nx1086)) ;
    inv01 ix1055 (.Y (nx1056), .A (nx807)) ;
    inv02 ix1057 (.Y (nx1058), .A (nx1056)) ;
    inv02 ix1059 (.Y (nx1060), .A (nx1056)) ;
    inv02 ix1061 (.Y (nx1062), .A (nx1056)) ;
    inv02 ix1063 (.Y (nx1064), .A (nx1056)) ;
    inv02 ix1065 (.Y (nx1066), .A (nx1056)) ;
    inv01 ix1067 (.Y (nx1068), .A (nx921)) ;
    inv02 ix1069 (.Y (nx1070), .A (nx1068)) ;
    inv02 ix1071 (.Y (nx1072), .A (nx1068)) ;
    inv02 ix1073 (.Y (nx1074), .A (nx1068)) ;
    inv02 ix1075 (.Y (nx1076), .A (nx1068)) ;
    inv02 ix1077 (.Y (nx1078), .A (nx1068)) ;
    inv02 ix1083 (.Y (nx1084), .A (nx1090)) ;
    inv02 ix1085 (.Y (nx1086), .A (nx1090)) ;
    inv02 ix1087 (.Y (nx1088), .A (enableRegFilter)) ;
    inv02 ix1089 (.Y (nx1090), .A (enableRegFilter)) ;
endmodule


module RegUnit_8_16 ( filterBus, windowBus, regPage1NextUnit, regPage2NextUnit, 
                      clk, rst, enableRegPage1, enableRegPage2, enableRegFilter, 
                      page1ReadBusOrPage2, page2ReadBusOrPage1, pageTurn, 
                      outRegPage, outputRegPage1, outputRegPage2, outFilter ) ;

    input [7:0]filterBus ;
    input [15:0]windowBus ;
    input [15:0]regPage1NextUnit ;
    input [15:0]regPage2NextUnit ;
    input clk ;
    input rst ;
    input enableRegPage1 ;
    input enableRegPage2 ;
    input enableRegFilter ;
    input page1ReadBusOrPage2 ;
    input page2ReadBusOrPage1 ;
    input pageTurn ;
    output [15:0]outRegPage ;
    output [15:0]outputRegPage1 ;
    output [15:0]outputRegPage2 ;
    output [7:0]outFilter ;

    wire outputRegPage1_0_rename, outputRegPage2_0_rename, 
         outputRegPage1_1_rename, outputRegPage2_1_rename, 
         outputRegPage1_2_rename, outputRegPage2_2_rename, 
         outputRegPage1_3_rename, outputRegPage2_3_rename, 
         outputRegPage1_4_rename, outputRegPage2_4_rename, 
         outputRegPage1_5_rename, outputRegPage2_5_rename, 
         outputRegPage1_6_rename, outputRegPage2_6_rename, 
         outputRegPage1_7_rename, outputRegPage2_7_rename, 
         outputRegPage1_8_rename, outputRegPage2_8_rename, 
         outputRegPage1_9_rename, outputRegPage2_9_rename, 
         outputRegPage1_10_rename, outputRegPage2_10_rename, 
         outputRegPage1_11_rename, outputRegPage2_11_rename, 
         outputRegPage1_12_rename, outputRegPage2_12_rename, 
         outputRegPage1_13_rename, outputRegPage2_13_rename, 
         outputRegPage1_14_rename, outputRegPage2_14_rename, 
         outputRegPage1_15_rename, outputRegPage2_15_rename, nx133, nx143, nx153, 
         nx163, nx173, nx183, nx193, nx203, nx213, nx223, nx233, nx243, nx253, 
         nx263, nx273, nx283, nx293, nx303, nx313, nx323, nx333, nx343, nx353, 
         nx363, nx373, nx383, nx393, nx403, nx413, nx423, nx433, nx443, nx453, 
         nx463, nx473, nx483, nx493, nx503, nx513, nx523, nx535, nx539, nx544, 
         nx546, nx551, nx553, nx558, nx560, nx565, nx567, nx572, nx574, nx579, 
         nx581, nx586, nx588, nx592, nx595, nx597, nx599, nx602, nx605, nx607, 
         nx609, nx613, nx616, nx618, nx621, nx624, nx626, nx630, nx633, nx635, 
         nx638, nx641, nx643, nx647, nx650, nx652, nx655, nx658, nx660, nx664, 
         nx667, nx669, nx672, nx675, nx677, nx681, nx684, nx686, nx689, nx692, 
         nx694, nx698, nx701, nx703, nx706, nx709, nx711, nx715, nx718, nx720, 
         nx723, nx726, nx728, nx732, nx735, nx737, nx740, nx743, nx745, nx749, 
         nx752, nx754, nx757, nx760, nx762, nx766, nx769, nx771, nx774, nx777, 
         nx779, nx783, nx786, nx788, nx791, nx794, nx796, nx800, nx803, nx805, 
         nx808, nx811, nx813, nx817, nx820, nx822, nx825, nx828, nx830, nx834, 
         nx837, nx839, nx842, nx845, nx847, nx851, nx854, nx856, nx859, nx862, 
         nx864, nx874, nx876, nx878, nx880, nx882, nx884, nx886, nx888, nx890, 
         nx892, nx894, nx896, nx898, nx904, nx906, nx908, nx910;
    wire [7:0] \$dummy ;




    assign outputRegPage1[14] = outputRegPage1[15] ;
    assign outputRegPage1[13] = outputRegPage1[15] ;
    assign outputRegPage1[12] = outputRegPage1[15] ;
    assign outputRegPage1[11] = outputRegPage1[15] ;
    assign outputRegPage1[10] = outputRegPage1[15] ;
    assign outputRegPage1[9] = outputRegPage1[15] ;
    assign outputRegPage1[8] = outputRegPage1[15] ;
    assign outputRegPage1[7] = outputRegPage1[15] ;
    assign outputRegPage1[6] = outputRegPage1[15] ;
    assign outputRegPage1[5] = outputRegPage1[15] ;
    assign outputRegPage1[4] = outputRegPage1[15] ;
    assign outputRegPage1[3] = outputRegPage1[15] ;
    assign outputRegPage1[2] = outputRegPage1[15] ;
    assign outputRegPage1[1] = outputRegPage1[15] ;
    assign outputRegPage1[0] = outputRegPage1[15] ;
    assign outputRegPage2[15] = outputRegPage1[15] ;
    assign outputRegPage2[14] = outputRegPage1[15] ;
    assign outputRegPage2[13] = outputRegPage1[15] ;
    assign outputRegPage2[12] = outputRegPage1[15] ;
    assign outputRegPage2[11] = outputRegPage1[15] ;
    assign outputRegPage2[10] = outputRegPage1[15] ;
    assign outputRegPage2[9] = outputRegPage1[15] ;
    assign outputRegPage2[8] = outputRegPage1[15] ;
    assign outputRegPage2[7] = outputRegPage1[15] ;
    assign outputRegPage2[6] = outputRegPage1[15] ;
    assign outputRegPage2[5] = outputRegPage1[15] ;
    assign outputRegPage2[4] = outputRegPage1[15] ;
    assign outputRegPage2[3] = outputRegPage1[15] ;
    assign outputRegPage2[2] = outputRegPage1[15] ;
    assign outputRegPage2[1] = outputRegPage1[15] ;
    assign outputRegPage2[0] = outputRegPage1[15] ;
    fake_gnd ix54 (.Y (outputRegPage1[15])) ;
    dffr regFilterMap_reg_Q_0 (.Q (outFilter[0]), .QB (\$dummy [0]), .D (nx453)
         , .CLK (clk), .R (rst)) ;
    nand02 ix454 (.Y (nx453), .A0 (nx535), .A1 (nx539)) ;
    nand02 ix536 (.Y (nx535), .A0 (outFilter[0]), .A1 (nx908)) ;
    nand02 ix540 (.Y (nx539), .A0 (filterBus[0]), .A1 (nx904)) ;
    dffr regFilterMap_reg_Q_1 (.Q (outFilter[1]), .QB (\$dummy [1]), .D (nx463)
         , .CLK (clk), .R (rst)) ;
    nand02 ix464 (.Y (nx463), .A0 (nx544), .A1 (nx546)) ;
    nand02 ix545 (.Y (nx544), .A0 (outFilter[1]), .A1 (nx908)) ;
    nand02 ix547 (.Y (nx546), .A0 (filterBus[1]), .A1 (nx904)) ;
    dffr regFilterMap_reg_Q_2 (.Q (outFilter[2]), .QB (\$dummy [2]), .D (nx473)
         , .CLK (clk), .R (rst)) ;
    nand02 ix474 (.Y (nx473), .A0 (nx551), .A1 (nx553)) ;
    nand02 ix552 (.Y (nx551), .A0 (outFilter[2]), .A1 (nx908)) ;
    nand02 ix554 (.Y (nx553), .A0 (filterBus[2]), .A1 (nx904)) ;
    dffr regFilterMap_reg_Q_3 (.Q (outFilter[3]), .QB (\$dummy [3]), .D (nx483)
         , .CLK (clk), .R (rst)) ;
    nand02 ix484 (.Y (nx483), .A0 (nx558), .A1 (nx560)) ;
    nand02 ix559 (.Y (nx558), .A0 (outFilter[3]), .A1 (nx908)) ;
    nand02 ix561 (.Y (nx560), .A0 (filterBus[3]), .A1 (nx904)) ;
    dffr regFilterMap_reg_Q_4 (.Q (outFilter[4]), .QB (\$dummy [4]), .D (nx493)
         , .CLK (clk), .R (rst)) ;
    nand02 ix494 (.Y (nx493), .A0 (nx565), .A1 (nx567)) ;
    nand02 ix566 (.Y (nx565), .A0 (outFilter[4]), .A1 (nx908)) ;
    nand02 ix568 (.Y (nx567), .A0 (filterBus[4]), .A1 (nx904)) ;
    dffr regFilterMap_reg_Q_5 (.Q (outFilter[5]), .QB (\$dummy [5]), .D (nx503)
         , .CLK (clk), .R (rst)) ;
    nand02 ix504 (.Y (nx503), .A0 (nx572), .A1 (nx574)) ;
    nand02 ix573 (.Y (nx572), .A0 (outFilter[5]), .A1 (nx908)) ;
    nand02 ix575 (.Y (nx574), .A0 (filterBus[5]), .A1 (nx904)) ;
    dffr regFilterMap_reg_Q_6 (.Q (outFilter[6]), .QB (\$dummy [6]), .D (nx513)
         , .CLK (clk), .R (rst)) ;
    nand02 ix514 (.Y (nx513), .A0 (nx579), .A1 (nx581)) ;
    nand02 ix580 (.Y (nx579), .A0 (outFilter[6]), .A1 (nx908)) ;
    nand02 ix582 (.Y (nx581), .A0 (filterBus[6]), .A1 (nx904)) ;
    dffr regFilterMap_reg_Q_7 (.Q (outFilter[7]), .QB (\$dummy [7]), .D (nx523)
         , .CLK (clk), .R (rst)) ;
    nand02 ix524 (.Y (nx523), .A0 (nx586), .A1 (nx588)) ;
    nand02 ix587 (.Y (nx586), .A0 (outFilter[7]), .A1 (nx874)) ;
    nand02 ix589 (.Y (nx588), .A0 (filterBus[7]), .A1 (nx906)) ;
    mux21 ix33 (.Y (outRegPage[0]), .A0 (nx592), .A1 (nx602), .S0 (pageTurn)) ;
    oai21 ix134 (.Y (nx133), .A0 (nx595), .A1 (nx878), .B0 (nx599)) ;
    mux21 ix596 (.Y (nx595), .A0 (windowBus[0]), .A1 (regPage2NextUnit[0]), .S0 (
          page1ReadBusOrPage2)) ;
    nor02_2x ix598 (.Y (nx597), .A0 (enableRegPage1), .A1 (page1ReadBusOrPage2)
             ) ;
    nand02 ix600 (.Y (nx599), .A0 (outputRegPage1_0_rename), .A1 (nx878)) ;
    dffr regPage1Map_reg_Q_0 (.Q (outputRegPage1_0_rename), .QB (nx592), .D (
         nx133), .CLK (clk), .R (rst)) ;
    oai21 ix144 (.Y (nx143), .A0 (nx605), .A1 (nx890), .B0 (nx609)) ;
    mux21 ix606 (.Y (nx605), .A0 (windowBus[0]), .A1 (regPage1NextUnit[0]), .S0 (
          page2ReadBusOrPage1)) ;
    nor02_2x ix608 (.Y (nx607), .A0 (enableRegPage2), .A1 (page2ReadBusOrPage1)
             ) ;
    nand02 ix610 (.Y (nx609), .A0 (outputRegPage2_0_rename), .A1 (nx890)) ;
    dffr regPage2Map_reg_Q_0 (.Q (outputRegPage2_0_rename), .QB (nx602), .D (
         nx143), .CLK (clk), .R (rst)) ;
    mux21 ix61 (.Y (outRegPage[1]), .A0 (nx613), .A1 (nx621), .S0 (pageTurn)) ;
    oai21 ix154 (.Y (nx153), .A0 (nx616), .A1 (nx878), .B0 (nx618)) ;
    mux21 ix617 (.Y (nx616), .A0 (windowBus[1]), .A1 (regPage2NextUnit[1]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix619 (.Y (nx618), .A0 (outputRegPage1_1_rename), .A1 (nx878)) ;
    dffr regPage1Map_reg_Q_1 (.Q (outputRegPage1_1_rename), .QB (nx613), .D (
         nx153), .CLK (clk), .R (rst)) ;
    oai21 ix164 (.Y (nx163), .A0 (nx624), .A1 (nx890), .B0 (nx626)) ;
    mux21 ix625 (.Y (nx624), .A0 (windowBus[1]), .A1 (regPage1NextUnit[1]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix627 (.Y (nx626), .A0 (outputRegPage2_1_rename), .A1 (nx890)) ;
    dffr regPage2Map_reg_Q_1 (.Q (outputRegPage2_1_rename), .QB (nx621), .D (
         nx163), .CLK (clk), .R (rst)) ;
    mux21 ix89 (.Y (outRegPage[2]), .A0 (nx630), .A1 (nx638), .S0 (pageTurn)) ;
    oai21 ix174 (.Y (nx173), .A0 (nx633), .A1 (nx878), .B0 (nx635)) ;
    mux21 ix634 (.Y (nx633), .A0 (windowBus[2]), .A1 (regPage2NextUnit[2]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix636 (.Y (nx635), .A0 (outputRegPage1_2_rename), .A1 (nx878)) ;
    dffr regPage1Map_reg_Q_2 (.Q (outputRegPage1_2_rename), .QB (nx630), .D (
         nx173), .CLK (clk), .R (rst)) ;
    oai21 ix184 (.Y (nx183), .A0 (nx641), .A1 (nx890), .B0 (nx643)) ;
    mux21 ix642 (.Y (nx641), .A0 (windowBus[2]), .A1 (regPage1NextUnit[2]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix644 (.Y (nx643), .A0 (outputRegPage2_2_rename), .A1 (nx890)) ;
    dffr regPage2Map_reg_Q_2 (.Q (outputRegPage2_2_rename), .QB (nx638), .D (
         nx183), .CLK (clk), .R (rst)) ;
    mux21 ix117 (.Y (outRegPage[3]), .A0 (nx647), .A1 (nx655), .S0 (pageTurn)) ;
    oai21 ix194 (.Y (nx193), .A0 (nx650), .A1 (nx878), .B0 (nx652)) ;
    mux21 ix651 (.Y (nx650), .A0 (windowBus[3]), .A1 (regPage2NextUnit[3]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix653 (.Y (nx652), .A0 (outputRegPage1_3_rename), .A1 (nx880)) ;
    dffr regPage1Map_reg_Q_3 (.Q (outputRegPage1_3_rename), .QB (nx647), .D (
         nx193), .CLK (clk), .R (rst)) ;
    oai21 ix204 (.Y (nx203), .A0 (nx658), .A1 (nx890), .B0 (nx660)) ;
    mux21 ix659 (.Y (nx658), .A0 (windowBus[3]), .A1 (regPage1NextUnit[3]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix661 (.Y (nx660), .A0 (outputRegPage2_3_rename), .A1 (nx892)) ;
    dffr regPage2Map_reg_Q_3 (.Q (outputRegPage2_3_rename), .QB (nx655), .D (
         nx203), .CLK (clk), .R (rst)) ;
    mux21 ix145 (.Y (outRegPage[4]), .A0 (nx664), .A1 (nx672), .S0 (pageTurn)) ;
    oai21 ix214 (.Y (nx213), .A0 (nx667), .A1 (nx880), .B0 (nx669)) ;
    mux21 ix668 (.Y (nx667), .A0 (windowBus[4]), .A1 (regPage2NextUnit[4]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix670 (.Y (nx669), .A0 (outputRegPage1_4_rename), .A1 (nx880)) ;
    dffr regPage1Map_reg_Q_4 (.Q (outputRegPage1_4_rename), .QB (nx664), .D (
         nx213), .CLK (clk), .R (rst)) ;
    oai21 ix224 (.Y (nx223), .A0 (nx675), .A1 (nx892), .B0 (nx677)) ;
    mux21 ix676 (.Y (nx675), .A0 (windowBus[4]), .A1 (regPage1NextUnit[4]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix678 (.Y (nx677), .A0 (outputRegPage2_4_rename), .A1 (nx892)) ;
    dffr regPage2Map_reg_Q_4 (.Q (outputRegPage2_4_rename), .QB (nx672), .D (
         nx223), .CLK (clk), .R (rst)) ;
    mux21 ix173 (.Y (outRegPage[5]), .A0 (nx681), .A1 (nx689), .S0 (pageTurn)) ;
    oai21 ix234 (.Y (nx233), .A0 (nx684), .A1 (nx880), .B0 (nx686)) ;
    mux21 ix685 (.Y (nx684), .A0 (windowBus[5]), .A1 (regPage2NextUnit[5]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix687 (.Y (nx686), .A0 (outputRegPage1_5_rename), .A1 (nx880)) ;
    dffr regPage1Map_reg_Q_5 (.Q (outputRegPage1_5_rename), .QB (nx681), .D (
         nx233), .CLK (clk), .R (rst)) ;
    oai21 ix244 (.Y (nx243), .A0 (nx692), .A1 (nx892), .B0 (nx694)) ;
    mux21 ix693 (.Y (nx692), .A0 (windowBus[5]), .A1 (regPage1NextUnit[5]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix695 (.Y (nx694), .A0 (outputRegPage2_5_rename), .A1 (nx892)) ;
    dffr regPage2Map_reg_Q_5 (.Q (outputRegPage2_5_rename), .QB (nx689), .D (
         nx243), .CLK (clk), .R (rst)) ;
    mux21 ix201 (.Y (outRegPage[6]), .A0 (nx698), .A1 (nx706), .S0 (pageTurn)) ;
    oai21 ix254 (.Y (nx253), .A0 (nx701), .A1 (nx880), .B0 (nx703)) ;
    mux21 ix702 (.Y (nx701), .A0 (windowBus[6]), .A1 (regPage2NextUnit[6]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix704 (.Y (nx703), .A0 (outputRegPage1_6_rename), .A1 (nx880)) ;
    dffr regPage1Map_reg_Q_6 (.Q (outputRegPage1_6_rename), .QB (nx698), .D (
         nx253), .CLK (clk), .R (rst)) ;
    oai21 ix264 (.Y (nx263), .A0 (nx709), .A1 (nx892), .B0 (nx711)) ;
    mux21 ix710 (.Y (nx709), .A0 (windowBus[6]), .A1 (regPage1NextUnit[6]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix712 (.Y (nx711), .A0 (outputRegPage2_6_rename), .A1 (nx892)) ;
    dffr regPage2Map_reg_Q_6 (.Q (outputRegPage2_6_rename), .QB (nx706), .D (
         nx263), .CLK (clk), .R (rst)) ;
    mux21 ix229 (.Y (outRegPage[7]), .A0 (nx715), .A1 (nx723), .S0 (pageTurn)) ;
    oai21 ix274 (.Y (nx273), .A0 (nx718), .A1 (nx882), .B0 (nx720)) ;
    mux21 ix719 (.Y (nx718), .A0 (windowBus[7]), .A1 (regPage2NextUnit[7]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix721 (.Y (nx720), .A0 (outputRegPage1_7_rename), .A1 (nx882)) ;
    dffr regPage1Map_reg_Q_7 (.Q (outputRegPage1_7_rename), .QB (nx715), .D (
         nx273), .CLK (clk), .R (rst)) ;
    oai21 ix284 (.Y (nx283), .A0 (nx726), .A1 (nx894), .B0 (nx728)) ;
    mux21 ix727 (.Y (nx726), .A0 (windowBus[7]), .A1 (regPage1NextUnit[7]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix729 (.Y (nx728), .A0 (outputRegPage2_7_rename), .A1 (nx894)) ;
    dffr regPage2Map_reg_Q_7 (.Q (outputRegPage2_7_rename), .QB (nx723), .D (
         nx283), .CLK (clk), .R (rst)) ;
    mux21 ix257 (.Y (outRegPage[8]), .A0 (nx732), .A1 (nx740), .S0 (pageTurn)) ;
    oai21 ix294 (.Y (nx293), .A0 (nx735), .A1 (nx882), .B0 (nx737)) ;
    mux21 ix736 (.Y (nx735), .A0 (windowBus[8]), .A1 (regPage2NextUnit[8]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix738 (.Y (nx737), .A0 (outputRegPage1_8_rename), .A1 (nx882)) ;
    dffr regPage1Map_reg_Q_8 (.Q (outputRegPage1_8_rename), .QB (nx732), .D (
         nx293), .CLK (clk), .R (rst)) ;
    oai21 ix304 (.Y (nx303), .A0 (nx743), .A1 (nx894), .B0 (nx745)) ;
    mux21 ix744 (.Y (nx743), .A0 (windowBus[8]), .A1 (regPage1NextUnit[8]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix746 (.Y (nx745), .A0 (outputRegPage2_8_rename), .A1 (nx894)) ;
    dffr regPage2Map_reg_Q_8 (.Q (outputRegPage2_8_rename), .QB (nx740), .D (
         nx303), .CLK (clk), .R (rst)) ;
    mux21 ix285 (.Y (outRegPage[9]), .A0 (nx749), .A1 (nx757), .S0 (pageTurn)) ;
    oai21 ix314 (.Y (nx313), .A0 (nx752), .A1 (nx882), .B0 (nx754)) ;
    mux21 ix753 (.Y (nx752), .A0 (windowBus[9]), .A1 (regPage2NextUnit[9]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix755 (.Y (nx754), .A0 (outputRegPage1_9_rename), .A1 (nx882)) ;
    dffr regPage1Map_reg_Q_9 (.Q (outputRegPage1_9_rename), .QB (nx749), .D (
         nx313), .CLK (clk), .R (rst)) ;
    oai21 ix324 (.Y (nx323), .A0 (nx760), .A1 (nx894), .B0 (nx762)) ;
    mux21 ix761 (.Y (nx760), .A0 (windowBus[9]), .A1 (regPage1NextUnit[9]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix763 (.Y (nx762), .A0 (outputRegPage2_9_rename), .A1 (nx894)) ;
    dffr regPage2Map_reg_Q_9 (.Q (outputRegPage2_9_rename), .QB (nx757), .D (
         nx323), .CLK (clk), .R (rst)) ;
    mux21 ix313 (.Y (outRegPage[10]), .A0 (nx766), .A1 (nx774), .S0 (pageTurn)
          ) ;
    oai21 ix334 (.Y (nx333), .A0 (nx769), .A1 (nx882), .B0 (nx771)) ;
    mux21 ix770 (.Y (nx769), .A0 (windowBus[10]), .A1 (regPage2NextUnit[10]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix772 (.Y (nx771), .A0 (outputRegPage1_10_rename), .A1 (nx884)) ;
    dffr regPage1Map_reg_Q_10 (.Q (outputRegPage1_10_rename), .QB (nx766), .D (
         nx333), .CLK (clk), .R (rst)) ;
    oai21 ix344 (.Y (nx343), .A0 (nx777), .A1 (nx894), .B0 (nx779)) ;
    mux21 ix778 (.Y (nx777), .A0 (windowBus[10]), .A1 (regPage1NextUnit[10]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix780 (.Y (nx779), .A0 (outputRegPage2_10_rename), .A1 (nx896)) ;
    dffr regPage2Map_reg_Q_10 (.Q (outputRegPage2_10_rename), .QB (nx774), .D (
         nx343), .CLK (clk), .R (rst)) ;
    mux21 ix341 (.Y (outRegPage[11]), .A0 (nx783), .A1 (nx791), .S0 (pageTurn)
          ) ;
    oai21 ix354 (.Y (nx353), .A0 (nx786), .A1 (nx884), .B0 (nx788)) ;
    mux21 ix787 (.Y (nx786), .A0 (windowBus[11]), .A1 (regPage2NextUnit[11]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix789 (.Y (nx788), .A0 (outputRegPage1_11_rename), .A1 (nx884)) ;
    dffr regPage1Map_reg_Q_11 (.Q (outputRegPage1_11_rename), .QB (nx783), .D (
         nx353), .CLK (clk), .R (rst)) ;
    oai21 ix364 (.Y (nx363), .A0 (nx794), .A1 (nx896), .B0 (nx796)) ;
    mux21 ix795 (.Y (nx794), .A0 (windowBus[11]), .A1 (regPage1NextUnit[11]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix797 (.Y (nx796), .A0 (outputRegPage2_11_rename), .A1 (nx896)) ;
    dffr regPage2Map_reg_Q_11 (.Q (outputRegPage2_11_rename), .QB (nx791), .D (
         nx363), .CLK (clk), .R (rst)) ;
    mux21 ix369 (.Y (outRegPage[12]), .A0 (nx800), .A1 (nx808), .S0 (pageTurn)
          ) ;
    oai21 ix374 (.Y (nx373), .A0 (nx803), .A1 (nx884), .B0 (nx805)) ;
    mux21 ix804 (.Y (nx803), .A0 (windowBus[12]), .A1 (regPage2NextUnit[12]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix806 (.Y (nx805), .A0 (outputRegPage1_12_rename), .A1 (nx884)) ;
    dffr regPage1Map_reg_Q_12 (.Q (outputRegPage1_12_rename), .QB (nx800), .D (
         nx373), .CLK (clk), .R (rst)) ;
    oai21 ix384 (.Y (nx383), .A0 (nx811), .A1 (nx896), .B0 (nx813)) ;
    mux21 ix812 (.Y (nx811), .A0 (windowBus[12]), .A1 (regPage1NextUnit[12]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix814 (.Y (nx813), .A0 (outputRegPage2_12_rename), .A1 (nx896)) ;
    dffr regPage2Map_reg_Q_12 (.Q (outputRegPage2_12_rename), .QB (nx808), .D (
         nx383), .CLK (clk), .R (rst)) ;
    mux21 ix397 (.Y (outRegPage[13]), .A0 (nx817), .A1 (nx825), .S0 (pageTurn)
          ) ;
    oai21 ix394 (.Y (nx393), .A0 (nx820), .A1 (nx884), .B0 (nx822)) ;
    mux21 ix821 (.Y (nx820), .A0 (windowBus[13]), .A1 (regPage2NextUnit[13]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix823 (.Y (nx822), .A0 (outputRegPage1_13_rename), .A1 (nx884)) ;
    dffr regPage1Map_reg_Q_13 (.Q (outputRegPage1_13_rename), .QB (nx817), .D (
         nx393), .CLK (clk), .R (rst)) ;
    oai21 ix404 (.Y (nx403), .A0 (nx828), .A1 (nx896), .B0 (nx830)) ;
    mux21 ix829 (.Y (nx828), .A0 (windowBus[13]), .A1 (regPage1NextUnit[13]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix831 (.Y (nx830), .A0 (outputRegPage2_13_rename), .A1 (nx896)) ;
    dffr regPage2Map_reg_Q_13 (.Q (outputRegPage2_13_rename), .QB (nx825), .D (
         nx403), .CLK (clk), .R (rst)) ;
    mux21 ix425 (.Y (outRegPage[14]), .A0 (nx834), .A1 (nx842), .S0 (pageTurn)
          ) ;
    oai21 ix414 (.Y (nx413), .A0 (nx837), .A1 (nx886), .B0 (nx839)) ;
    mux21 ix838 (.Y (nx837), .A0 (windowBus[14]), .A1 (regPage2NextUnit[14]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix840 (.Y (nx839), .A0 (outputRegPage1_14_rename), .A1 (nx886)) ;
    dffr regPage1Map_reg_Q_14 (.Q (outputRegPage1_14_rename), .QB (nx834), .D (
         nx413), .CLK (clk), .R (rst)) ;
    oai21 ix424 (.Y (nx423), .A0 (nx845), .A1 (nx898), .B0 (nx847)) ;
    mux21 ix846 (.Y (nx845), .A0 (windowBus[14]), .A1 (regPage1NextUnit[14]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix848 (.Y (nx847), .A0 (outputRegPage2_14_rename), .A1 (nx898)) ;
    dffr regPage2Map_reg_Q_14 (.Q (outputRegPage2_14_rename), .QB (nx842), .D (
         nx423), .CLK (clk), .R (rst)) ;
    mux21 ix453 (.Y (outRegPage[15]), .A0 (nx851), .A1 (nx859), .S0 (pageTurn)
          ) ;
    oai21 ix434 (.Y (nx433), .A0 (nx854), .A1 (nx886), .B0 (nx856)) ;
    mux21 ix855 (.Y (nx854), .A0 (windowBus[15]), .A1 (regPage2NextUnit[15]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix857 (.Y (nx856), .A0 (outputRegPage1_15_rename), .A1 (nx886)) ;
    dffr regPage1Map_reg_Q_15 (.Q (outputRegPage1_15_rename), .QB (nx851), .D (
         nx433), .CLK (clk), .R (rst)) ;
    oai21 ix444 (.Y (nx443), .A0 (nx862), .A1 (nx898), .B0 (nx864)) ;
    mux21 ix863 (.Y (nx862), .A0 (windowBus[15]), .A1 (regPage1NextUnit[15]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix865 (.Y (nx864), .A0 (outputRegPage2_15_rename), .A1 (nx898)) ;
    dffr regPage2Map_reg_Q_15 (.Q (outputRegPage2_15_rename), .QB (nx859), .D (
         nx443), .CLK (clk), .R (rst)) ;
    inv01 ix873 (.Y (nx874), .A (nx906)) ;
    inv01 ix875 (.Y (nx876), .A (nx597)) ;
    inv02 ix877 (.Y (nx878), .A (nx876)) ;
    inv02 ix879 (.Y (nx880), .A (nx876)) ;
    inv02 ix881 (.Y (nx882), .A (nx876)) ;
    inv02 ix883 (.Y (nx884), .A (nx876)) ;
    inv02 ix885 (.Y (nx886), .A (nx876)) ;
    inv01 ix887 (.Y (nx888), .A (nx607)) ;
    inv02 ix889 (.Y (nx890), .A (nx888)) ;
    inv02 ix891 (.Y (nx892), .A (nx888)) ;
    inv02 ix893 (.Y (nx894), .A (nx888)) ;
    inv02 ix895 (.Y (nx896), .A (nx888)) ;
    inv02 ix897 (.Y (nx898), .A (nx888)) ;
    inv02 ix903 (.Y (nx904), .A (nx910)) ;
    inv02 ix905 (.Y (nx906), .A (nx910)) ;
    inv02 ix907 (.Y (nx908), .A (enableRegFilter)) ;
    inv02 ix909 (.Y (nx910), .A (enableRegFilter)) ;
endmodule

