
-- 
-- Definition of  CNNMuls
-- 
--      Thu Apr 11 12:57:10 2019
--      
--      LeonardoSpectrum Level 3, 2018a.2
-- 

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity Reg_33 is
   port (
      D : IN std_logic_vector (32 DOWNTO 0) ;
      en : IN std_logic ;
      clk : IN std_logic ;
      rst : IN std_logic ;
      Q : OUT std_logic_vector (32 DOWNTO 0)) ;
end Reg_33 ;

architecture RegArch_unfold_1389 of Reg_33 is
   signal Q_30_EXMPLR, Q_29_EXMPLR, Q_28_EXMPLR, Q_27_EXMPLR, Q_26_EXMPLR, 
      Q_25_EXMPLR, Q_24_EXMPLR, Q_23_EXMPLR, Q_22_EXMPLR, Q_21_EXMPLR, 
      Q_20_EXMPLR, Q_19_EXMPLR, Q_18_EXMPLR, Q_17_EXMPLR, Q_16_EXMPLR, 
      Q_15_EXMPLR, Q_14_EXMPLR, Q_13_EXMPLR, Q_12_EXMPLR, Q_11_EXMPLR, 
      Q_10_EXMPLR, Q_9_EXMPLR, Q_8_EXMPLR, Q_7_EXMPLR, Q_6_EXMPLR, 
      Q_5_EXMPLR, Q_4_EXMPLR, Q_3_EXMPLR, Q_2_EXMPLR, Q_1_EXMPLR, Q_0_EXMPLR, 
      Q_32_EXMPLR, nx115, nx125, nx135, nx145, nx155, nx165, nx175, nx185, 
      nx195, nx205, nx215, nx225, nx235, nx245, nx255, nx265, nx275, nx285, 
      nx295, nx305, nx315, nx325, nx335, nx345, nx355, nx365, nx375, nx385, 
      nx395, nx405, nx415, nx427, nx431, nx436, nx438, nx443, nx445, nx450, 
      nx452, nx457, nx459, nx464, nx466, nx471, nx473, nx478, nx480, nx485, 
      nx487, nx492, nx494, nx499, nx501, nx506, nx508, nx513, nx515, nx520, 
      nx522, nx527, nx529, nx534, nx536, nx541, nx543, nx548, nx550, nx555, 
      nx557, nx562, nx564, nx569, nx571, nx576, nx578, nx583, nx585, nx590, 
      nx592, nx597, nx599, nx604, nx606, nx611, nx613, nx618, nx620, nx625, 
      nx627, nx632, nx634, nx639, nx641, nx649, nx651, nx653, nx655, nx657, 
      nx663, nx665, nx667, nx669, nx671, nx673, nx675, nx677, nx679, nx681, 
      nx683, nx685: std_logic ;

begin
   Q(32) <= Q_32_EXMPLR ;
   Q(31) <= Q_32_EXMPLR ;
   Q(30) <= Q_30_EXMPLR ;
   Q(29) <= Q_29_EXMPLR ;
   Q(28) <= Q_28_EXMPLR ;
   Q(27) <= Q_27_EXMPLR ;
   Q(26) <= Q_26_EXMPLR ;
   Q(25) <= Q_25_EXMPLR ;
   Q(24) <= Q_24_EXMPLR ;
   Q(23) <= Q_23_EXMPLR ;
   Q(22) <= Q_22_EXMPLR ;
   Q(21) <= Q_21_EXMPLR ;
   Q(20) <= Q_20_EXMPLR ;
   Q(19) <= Q_19_EXMPLR ;
   Q(18) <= Q_18_EXMPLR ;
   Q(17) <= Q_17_EXMPLR ;
   Q(16) <= Q_16_EXMPLR ;
   Q(15) <= Q_15_EXMPLR ;
   Q(14) <= Q_14_EXMPLR ;
   Q(13) <= Q_13_EXMPLR ;
   Q(12) <= Q_12_EXMPLR ;
   Q(11) <= Q_11_EXMPLR ;
   Q(10) <= Q_10_EXMPLR ;
   Q(9) <= Q_9_EXMPLR ;
   Q(8) <= Q_8_EXMPLR ;
   Q(7) <= Q_7_EXMPLR ;
   Q(6) <= Q_6_EXMPLR ;
   Q(5) <= Q_5_EXMPLR ;
   Q(4) <= Q_4_EXMPLR ;
   Q(3) <= Q_3_EXMPLR ;
   Q(2) <= Q_2_EXMPLR ;
   Q(1) <= Q_1_EXMPLR ;
   Q(0) <= Q_0_EXMPLR ;
   ix43 : fake_gnd port map ( Y=>Q_32_EXMPLR);
   reg_Q_0 : dffr port map ( Q=>Q_0_EXMPLR, QB=>OPEN, D=>nx115, CLK=>nx665, 
      R=>rst);
   ix116 : nand02 port map ( Y=>nx115, A0=>nx427, A1=>nx431);
   ix428 : nand02 port map ( Y=>nx427, A0=>Q_0_EXMPLR, A1=>nx685);
   ix432 : nand02 port map ( Y=>nx431, A0=>D(0), A1=>nx675);
   reg_Q_1 : dffr port map ( Q=>Q_1_EXMPLR, QB=>OPEN, D=>nx125, CLK=>nx665, 
      R=>rst);
   ix126 : nand02 port map ( Y=>nx125, A0=>nx436, A1=>nx438);
   ix437 : nand02 port map ( Y=>nx436, A0=>Q_1_EXMPLR, A1=>nx685);
   ix439 : nand02 port map ( Y=>nx438, A0=>D(1), A1=>nx675);
   reg_Q_2 : dffr port map ( Q=>Q_2_EXMPLR, QB=>OPEN, D=>nx135, CLK=>nx665, 
      R=>rst);
   ix136 : nand02 port map ( Y=>nx135, A0=>nx443, A1=>nx445);
   ix444 : nand02 port map ( Y=>nx443, A0=>Q_2_EXMPLR, A1=>nx685);
   ix446 : nand02 port map ( Y=>nx445, A0=>D(2), A1=>nx675);
   reg_Q_3 : dffr port map ( Q=>Q_3_EXMPLR, QB=>OPEN, D=>nx145, CLK=>nx665, 
      R=>rst);
   ix146 : nand02 port map ( Y=>nx145, A0=>nx450, A1=>nx452);
   ix451 : nand02 port map ( Y=>nx450, A0=>Q_3_EXMPLR, A1=>nx685);
   ix453 : nand02 port map ( Y=>nx452, A0=>D(3), A1=>nx675);
   reg_Q_4 : dffr port map ( Q=>Q_4_EXMPLR, QB=>OPEN, D=>nx155, CLK=>nx665, 
      R=>rst);
   ix156 : nand02 port map ( Y=>nx155, A0=>nx457, A1=>nx459);
   ix458 : nand02 port map ( Y=>nx457, A0=>Q_4_EXMPLR, A1=>nx685);
   ix460 : nand02 port map ( Y=>nx459, A0=>D(4), A1=>nx675);
   reg_Q_5 : dffr port map ( Q=>Q_5_EXMPLR, QB=>OPEN, D=>nx165, CLK=>nx665, 
      R=>rst);
   ix166 : nand02 port map ( Y=>nx165, A0=>nx464, A1=>nx466);
   ix465 : nand02 port map ( Y=>nx464, A0=>Q_5_EXMPLR, A1=>nx685);
   ix467 : nand02 port map ( Y=>nx466, A0=>D(5), A1=>nx675);
   reg_Q_6 : dffr port map ( Q=>Q_6_EXMPLR, QB=>OPEN, D=>nx175, CLK=>nx665, 
      R=>rst);
   ix176 : nand02 port map ( Y=>nx175, A0=>nx471, A1=>nx473);
   ix472 : nand02 port map ( Y=>nx471, A0=>Q_6_EXMPLR, A1=>nx685);
   ix474 : nand02 port map ( Y=>nx473, A0=>D(6), A1=>nx675);
   reg_Q_7 : dffr port map ( Q=>Q_7_EXMPLR, QB=>OPEN, D=>nx185, CLK=>nx667, 
      R=>rst);
   ix186 : nand02 port map ( Y=>nx185, A0=>nx478, A1=>nx480);
   ix479 : nand02 port map ( Y=>nx478, A0=>Q_7_EXMPLR, A1=>nx651);
   ix481 : nand02 port map ( Y=>nx480, A0=>D(7), A1=>nx677);
   reg_Q_8 : dffr port map ( Q=>Q_8_EXMPLR, QB=>OPEN, D=>nx195, CLK=>nx667, 
      R=>rst);
   ix196 : nand02 port map ( Y=>nx195, A0=>nx485, A1=>nx487);
   ix486 : nand02 port map ( Y=>nx485, A0=>Q_8_EXMPLR, A1=>nx651);
   ix488 : nand02 port map ( Y=>nx487, A0=>D(8), A1=>nx677);
   reg_Q_9 : dffr port map ( Q=>Q_9_EXMPLR, QB=>OPEN, D=>nx205, CLK=>nx667, 
      R=>rst);
   ix206 : nand02 port map ( Y=>nx205, A0=>nx492, A1=>nx494);
   ix493 : nand02 port map ( Y=>nx492, A0=>Q_9_EXMPLR, A1=>nx651);
   ix495 : nand02 port map ( Y=>nx494, A0=>D(9), A1=>nx677);
   reg_Q_10 : dffr port map ( Q=>Q_10_EXMPLR, QB=>OPEN, D=>nx215, CLK=>nx667, 
      R=>rst);
   ix216 : nand02 port map ( Y=>nx215, A0=>nx499, A1=>nx501);
   ix500 : nand02 port map ( Y=>nx499, A0=>Q_10_EXMPLR, A1=>nx651);
   ix502 : nand02 port map ( Y=>nx501, A0=>D(10), A1=>nx677);
   reg_Q_11 : dffr port map ( Q=>Q_11_EXMPLR, QB=>OPEN, D=>nx225, CLK=>nx667, 
      R=>rst);
   ix226 : nand02 port map ( Y=>nx225, A0=>nx506, A1=>nx508);
   ix507 : nand02 port map ( Y=>nx506, A0=>Q_11_EXMPLR, A1=>nx651);
   ix509 : nand02 port map ( Y=>nx508, A0=>D(11), A1=>nx677);
   reg_Q_12 : dffr port map ( Q=>Q_12_EXMPLR, QB=>OPEN, D=>nx235, CLK=>nx667, 
      R=>rst);
   ix236 : nand02 port map ( Y=>nx235, A0=>nx513, A1=>nx515);
   ix514 : nand02 port map ( Y=>nx513, A0=>Q_12_EXMPLR, A1=>nx651);
   ix516 : nand02 port map ( Y=>nx515, A0=>D(12), A1=>nx677);
   reg_Q_13 : dffr port map ( Q=>Q_13_EXMPLR, QB=>OPEN, D=>nx245, CLK=>nx667, 
      R=>rst);
   ix246 : nand02 port map ( Y=>nx245, A0=>nx520, A1=>nx522);
   ix521 : nand02 port map ( Y=>nx520, A0=>Q_13_EXMPLR, A1=>nx651);
   ix523 : nand02 port map ( Y=>nx522, A0=>D(13), A1=>nx677);
   reg_Q_14 : dffr port map ( Q=>Q_14_EXMPLR, QB=>OPEN, D=>nx255, CLK=>nx669, 
      R=>rst);
   ix256 : nand02 port map ( Y=>nx255, A0=>nx527, A1=>nx529);
   ix528 : nand02 port map ( Y=>nx527, A0=>Q_14_EXMPLR, A1=>nx653);
   ix530 : nand02 port map ( Y=>nx529, A0=>D(14), A1=>nx679);
   reg_Q_15 : dffr port map ( Q=>Q_15_EXMPLR, QB=>OPEN, D=>nx265, CLK=>nx669, 
      R=>rst);
   ix266 : nand02 port map ( Y=>nx265, A0=>nx534, A1=>nx536);
   ix535 : nand02 port map ( Y=>nx534, A0=>Q_15_EXMPLR, A1=>nx653);
   ix537 : nand02 port map ( Y=>nx536, A0=>D(15), A1=>nx679);
   reg_Q_16 : dffr port map ( Q=>Q_16_EXMPLR, QB=>OPEN, D=>nx275, CLK=>nx669, 
      R=>rst);
   ix276 : nand02 port map ( Y=>nx275, A0=>nx541, A1=>nx543);
   ix542 : nand02 port map ( Y=>nx541, A0=>Q_16_EXMPLR, A1=>nx653);
   ix544 : nand02 port map ( Y=>nx543, A0=>D(16), A1=>nx679);
   reg_Q_17 : dffr port map ( Q=>Q_17_EXMPLR, QB=>OPEN, D=>nx285, CLK=>nx669, 
      R=>rst);
   ix286 : nand02 port map ( Y=>nx285, A0=>nx548, A1=>nx550);
   ix549 : nand02 port map ( Y=>nx548, A0=>Q_17_EXMPLR, A1=>nx653);
   ix551 : nand02 port map ( Y=>nx550, A0=>D(17), A1=>nx679);
   reg_Q_18 : dffr port map ( Q=>Q_18_EXMPLR, QB=>OPEN, D=>nx295, CLK=>nx669, 
      R=>rst);
   ix296 : nand02 port map ( Y=>nx295, A0=>nx555, A1=>nx557);
   ix556 : nand02 port map ( Y=>nx555, A0=>Q_18_EXMPLR, A1=>nx653);
   ix558 : nand02 port map ( Y=>nx557, A0=>D(18), A1=>nx679);
   reg_Q_19 : dffr port map ( Q=>Q_19_EXMPLR, QB=>OPEN, D=>nx305, CLK=>nx669, 
      R=>rst);
   ix306 : nand02 port map ( Y=>nx305, A0=>nx562, A1=>nx564);
   ix563 : nand02 port map ( Y=>nx562, A0=>Q_19_EXMPLR, A1=>nx653);
   ix565 : nand02 port map ( Y=>nx564, A0=>D(19), A1=>nx679);
   reg_Q_20 : dffr port map ( Q=>Q_20_EXMPLR, QB=>OPEN, D=>nx315, CLK=>nx669, 
      R=>rst);
   ix316 : nand02 port map ( Y=>nx315, A0=>nx569, A1=>nx571);
   ix570 : nand02 port map ( Y=>nx569, A0=>Q_20_EXMPLR, A1=>nx653);
   ix572 : nand02 port map ( Y=>nx571, A0=>D(20), A1=>nx679);
   reg_Q_21 : dffr port map ( Q=>Q_21_EXMPLR, QB=>OPEN, D=>nx325, CLK=>nx671, 
      R=>rst);
   ix326 : nand02 port map ( Y=>nx325, A0=>nx576, A1=>nx578);
   ix577 : nand02 port map ( Y=>nx576, A0=>Q_21_EXMPLR, A1=>nx655);
   ix579 : nand02 port map ( Y=>nx578, A0=>D(21), A1=>nx681);
   reg_Q_22 : dffr port map ( Q=>Q_22_EXMPLR, QB=>OPEN, D=>nx335, CLK=>nx671, 
      R=>rst);
   ix336 : nand02 port map ( Y=>nx335, A0=>nx583, A1=>nx585);
   ix584 : nand02 port map ( Y=>nx583, A0=>Q_22_EXMPLR, A1=>nx655);
   ix586 : nand02 port map ( Y=>nx585, A0=>D(22), A1=>nx681);
   reg_Q_23 : dffr port map ( Q=>Q_23_EXMPLR, QB=>OPEN, D=>nx345, CLK=>nx671, 
      R=>rst);
   ix346 : nand02 port map ( Y=>nx345, A0=>nx590, A1=>nx592);
   ix591 : nand02 port map ( Y=>nx590, A0=>Q_23_EXMPLR, A1=>nx655);
   ix593 : nand02 port map ( Y=>nx592, A0=>D(23), A1=>nx681);
   reg_Q_24 : dffr port map ( Q=>Q_24_EXMPLR, QB=>OPEN, D=>nx355, CLK=>nx671, 
      R=>rst);
   ix356 : nand02 port map ( Y=>nx355, A0=>nx597, A1=>nx599);
   ix598 : nand02 port map ( Y=>nx597, A0=>Q_24_EXMPLR, A1=>nx655);
   ix600 : nand02 port map ( Y=>nx599, A0=>D(24), A1=>nx681);
   reg_Q_25 : dffr port map ( Q=>Q_25_EXMPLR, QB=>OPEN, D=>nx365, CLK=>nx671, 
      R=>rst);
   ix366 : nand02 port map ( Y=>nx365, A0=>nx604, A1=>nx606);
   ix605 : nand02 port map ( Y=>nx604, A0=>Q_25_EXMPLR, A1=>nx655);
   ix607 : nand02 port map ( Y=>nx606, A0=>D(25), A1=>nx681);
   reg_Q_26 : dffr port map ( Q=>Q_26_EXMPLR, QB=>OPEN, D=>nx375, CLK=>nx671, 
      R=>rst);
   ix376 : nand02 port map ( Y=>nx375, A0=>nx611, A1=>nx613);
   ix612 : nand02 port map ( Y=>nx611, A0=>Q_26_EXMPLR, A1=>nx655);
   ix614 : nand02 port map ( Y=>nx613, A0=>D(26), A1=>nx681);
   reg_Q_27 : dffr port map ( Q=>Q_27_EXMPLR, QB=>OPEN, D=>nx385, CLK=>nx671, 
      R=>rst);
   ix386 : nand02 port map ( Y=>nx385, A0=>nx618, A1=>nx620);
   ix619 : nand02 port map ( Y=>nx618, A0=>Q_27_EXMPLR, A1=>nx655);
   ix621 : nand02 port map ( Y=>nx620, A0=>D(27), A1=>nx681);
   reg_Q_28 : dffr port map ( Q=>Q_28_EXMPLR, QB=>OPEN, D=>nx395, CLK=>nx673, 
      R=>rst);
   ix396 : nand02 port map ( Y=>nx395, A0=>nx625, A1=>nx627);
   ix626 : nand02 port map ( Y=>nx625, A0=>Q_28_EXMPLR, A1=>nx657);
   ix628 : nand02 port map ( Y=>nx627, A0=>D(28), A1=>nx683);
   reg_Q_29 : dffr port map ( Q=>Q_29_EXMPLR, QB=>OPEN, D=>nx405, CLK=>nx673, 
      R=>rst);
   ix406 : nand02 port map ( Y=>nx405, A0=>nx632, A1=>nx634);
   ix633 : nand02 port map ( Y=>nx632, A0=>Q_29_EXMPLR, A1=>nx657);
   ix635 : nand02 port map ( Y=>nx634, A0=>D(29), A1=>nx683);
   reg_Q_30 : dffr port map ( Q=>Q_30_EXMPLR, QB=>OPEN, D=>nx415, CLK=>nx673, 
      R=>rst);
   ix416 : nand02 port map ( Y=>nx415, A0=>nx639, A1=>nx641);
   ix640 : nand02 port map ( Y=>nx639, A0=>Q_30_EXMPLR, A1=>nx657);
   ix642 : nand02 port map ( Y=>nx641, A0=>D(30), A1=>nx683);
   ix648 : inv02 port map ( Y=>nx649, A=>en);
   ix650 : inv02 port map ( Y=>nx651, A=>nx683);
   ix652 : inv02 port map ( Y=>nx653, A=>nx683);
   ix654 : inv02 port map ( Y=>nx655, A=>nx683);
   ix656 : inv02 port map ( Y=>nx657, A=>nx683);
   ix662 : inv01 port map ( Y=>nx663, A=>clk);
   ix664 : inv02 port map ( Y=>nx665, A=>nx663);
   ix666 : inv02 port map ( Y=>nx667, A=>nx663);
   ix668 : inv02 port map ( Y=>nx669, A=>nx663);
   ix670 : inv02 port map ( Y=>nx671, A=>nx663);
   ix672 : inv02 port map ( Y=>nx673, A=>nx663);
   ix674 : inv02 port map ( Y=>nx675, A=>nx649);
   ix676 : inv02 port map ( Y=>nx677, A=>nx649);
   ix678 : inv02 port map ( Y=>nx679, A=>nx649);
   ix680 : inv02 port map ( Y=>nx681, A=>nx649);
   ix682 : inv02 port map ( Y=>nx683, A=>nx649);
   ix684 : inv02 port map ( Y=>nx685, A=>en);
end RegArch_unfold_1389 ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity BinaryMux_33 is
   port (
      a : IN std_logic_vector (32 DOWNTO 0) ;
      b : IN std_logic_vector (32 DOWNTO 0) ;
      sel : IN std_logic ;
      f : OUT std_logic_vector (32 DOWNTO 0)) ;
end BinaryMux_33 ;

architecture BinaryMuxArch_unfold_1786 of BinaryMux_33 is
   signal f_32_EXMPLR, nx93, nx97, nx99, nx105, nx107, nx111, nx113, nx117, 
      nx119, nx123, nx125, nx129, nx131, nx135, nx137, nx141, nx143, nx147, 
      nx151, nx155, nx158, nx161, nx164, nx167, nx170, nx173, nx176, nx179, 
      nx182, nx185, nx188, nx191, nx194, nx197, nx200, nx203, nx206, nx209, 
      nx212, nx219, nx221, nx223, nx225, nx227, nx229, nx231: std_logic ;

begin
   f(32) <= f_32_EXMPLR ;
   f(31) <= f_32_EXMPLR ;
   ix44 : fake_gnd port map ( Y=>f_32_EXMPLR);
   ix3 : nor02_2x port map ( Y=>f(0), A0=>nx93, A1=>nx219);
   ix94 : inv01 port map ( Y=>nx93, A=>a(0));
   ix99 : nand02_2x port map ( Y=>f(1), A0=>nx97, A1=>nx99);
   ix98 : nand02 port map ( Y=>nx97, A0=>b(1), A1=>nx219);
   ix100 : nand02 port map ( Y=>nx99, A0=>a(1), A1=>nx229);
   ix107 : nand02 port map ( Y=>f(2), A0=>nx105, A1=>nx107);
   ix106 : nand02 port map ( Y=>nx105, A0=>b(2), A1=>nx219);
   ix108 : nand02 port map ( Y=>nx107, A0=>a(2), A1=>nx229);
   ix115 : nand02 port map ( Y=>f(3), A0=>nx111, A1=>nx113);
   ix112 : nand02 port map ( Y=>nx111, A0=>b(3), A1=>nx219);
   ix114 : nand02 port map ( Y=>nx113, A0=>a(3), A1=>nx229);
   ix123 : nand02 port map ( Y=>f(4), A0=>nx117, A1=>nx119);
   ix118 : nand02 port map ( Y=>nx117, A0=>b(4), A1=>nx219);
   ix120 : nand02 port map ( Y=>nx119, A0=>a(4), A1=>nx229);
   ix131 : nand02 port map ( Y=>f(5), A0=>nx123, A1=>nx125);
   ix124 : nand02 port map ( Y=>nx123, A0=>b(5), A1=>nx219);
   ix126 : nand02 port map ( Y=>nx125, A0=>a(5), A1=>nx229);
   ix139 : nand02 port map ( Y=>f(6), A0=>nx129, A1=>nx131);
   ix130 : nand02 port map ( Y=>nx129, A0=>b(6), A1=>nx219);
   ix132 : nand02 port map ( Y=>nx131, A0=>a(6), A1=>nx229);
   ix147 : nand02 port map ( Y=>f(7), A0=>nx135, A1=>nx137);
   ix136 : nand02 port map ( Y=>nx135, A0=>b(7), A1=>nx221);
   ix138 : nand02 port map ( Y=>nx137, A0=>a(7), A1=>nx229);
   ix155 : nand02 port map ( Y=>f(8), A0=>nx141, A1=>nx143);
   ix142 : nand02 port map ( Y=>nx141, A0=>nx221, A1=>b(8));
   ix144 : nand02 port map ( Y=>nx143, A0=>nx231, A1=>a(8));
   ix7 : nor02_2x port map ( Y=>f(9), A0=>nx147, A1=>nx221);
   ix148 : inv01 port map ( Y=>nx147, A=>a(9));
   ix11 : nor02_2x port map ( Y=>f(10), A0=>nx151, A1=>nx221);
   ix152 : inv01 port map ( Y=>nx151, A=>a(10));
   ix15 : nor02_2x port map ( Y=>f(11), A0=>nx155, A1=>nx221);
   ix156 : inv01 port map ( Y=>nx155, A=>a(11));
   ix19 : nor02_2x port map ( Y=>f(12), A0=>nx158, A1=>nx221);
   ix159 : inv01 port map ( Y=>nx158, A=>a(12));
   ix23 : nor02_2x port map ( Y=>f(13), A0=>nx161, A1=>nx221);
   ix162 : inv01 port map ( Y=>nx161, A=>a(13));
   ix27 : nor02_2x port map ( Y=>f(14), A0=>nx164, A1=>nx223);
   ix165 : inv01 port map ( Y=>nx164, A=>a(14));
   ix31 : nor02_2x port map ( Y=>f(15), A0=>nx167, A1=>nx223);
   ix168 : inv01 port map ( Y=>nx167, A=>a(15));
   ix35 : nor02_2x port map ( Y=>f(16), A0=>nx170, A1=>nx223);
   ix171 : inv01 port map ( Y=>nx170, A=>a(16));
   ix39 : nor02_2x port map ( Y=>f(17), A0=>nx173, A1=>nx223);
   ix174 : inv01 port map ( Y=>nx173, A=>a(17));
   ix43 : nor02_2x port map ( Y=>f(18), A0=>nx176, A1=>nx223);
   ix177 : inv01 port map ( Y=>nx176, A=>a(18));
   ix47 : nor02_2x port map ( Y=>f(19), A0=>nx179, A1=>nx223);
   ix180 : inv01 port map ( Y=>nx179, A=>a(19));
   ix51 : nor02_2x port map ( Y=>f(20), A0=>nx182, A1=>nx223);
   ix183 : inv01 port map ( Y=>nx182, A=>a(20));
   ix55 : nor02_2x port map ( Y=>f(21), A0=>nx185, A1=>nx225);
   ix186 : inv01 port map ( Y=>nx185, A=>a(21));
   ix59 : nor02_2x port map ( Y=>f(22), A0=>nx188, A1=>nx225);
   ix189 : inv01 port map ( Y=>nx188, A=>a(22));
   ix63 : nor02_2x port map ( Y=>f(23), A0=>nx191, A1=>nx225);
   ix192 : inv01 port map ( Y=>nx191, A=>a(23));
   ix67 : nor02_2x port map ( Y=>f(24), A0=>nx194, A1=>nx225);
   ix195 : inv01 port map ( Y=>nx194, A=>a(24));
   ix71 : nor02_2x port map ( Y=>f(25), A0=>nx197, A1=>nx225);
   ix198 : inv01 port map ( Y=>nx197, A=>a(25));
   ix75 : nor02_2x port map ( Y=>f(26), A0=>nx200, A1=>nx225);
   ix201 : inv01 port map ( Y=>nx200, A=>a(26));
   ix79 : nor02_2x port map ( Y=>f(27), A0=>nx203, A1=>nx225);
   ix204 : inv01 port map ( Y=>nx203, A=>a(27));
   ix83 : nor02_2x port map ( Y=>f(28), A0=>nx206, A1=>nx227);
   ix207 : inv01 port map ( Y=>nx206, A=>a(28));
   ix87 : nor02_2x port map ( Y=>f(29), A0=>nx209, A1=>nx227);
   ix210 : inv01 port map ( Y=>nx209, A=>a(29));
   ix91 : nor02_2x port map ( Y=>f(30), A0=>nx212, A1=>nx227);
   ix213 : inv01 port map ( Y=>nx212, A=>a(30));
   ix218 : inv02 port map ( Y=>nx219, A=>nx231);
   ix220 : inv02 port map ( Y=>nx221, A=>nx231);
   ix222 : inv02 port map ( Y=>nx223, A=>nx231);
   ix224 : inv02 port map ( Y=>nx225, A=>nx231);
   ix226 : inv02 port map ( Y=>nx227, A=>nx231);
   ix228 : inv02 port map ( Y=>nx229, A=>sel);
   ix230 : inv02 port map ( Y=>nx231, A=>sel);
end BinaryMuxArch_unfold_1786 ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity NBitAdder_24 is
   port (
      a : IN std_logic_vector (23 DOWNTO 0) ;
      b : IN std_logic_vector (23 DOWNTO 0) ;
      carryIn : IN std_logic ;
      sum : OUT std_logic_vector (23 DOWNTO 0) ;
      carryOut : OUT std_logic) ;
end NBitAdder_24 ;

architecture NBitAdderArch_unfold_2081 of NBitAdder_24 is
   signal nx6, nx8, nx16, nx18, nx22, nx24, nx30, nx32, nx38, nx40, nx46, 
      nx48, nx54, nx56, nx62, nx64, nx70, nx72, nx78, nx80, nx86, nx88, nx94, 
      nx96, nx102, nx104, nx110, nx112, nx118, nx120, nx126, nx128, nx134, 
      nx136, nx142, nx144, nx150, nx152, nx158, nx160, nx166, nx168, nx170, 
      nx172, nx103, nx109, nx111, nx113, nx115, nx119, nx123, nx127, nx133, 
      nx135, nx137, nx141, nx145, nx149, nx155, nx157, nx159, nx163, nx167, 
      nx171, nx177, nx179, nx181, nx185, nx189, nx193, nx199, nx201, nx203, 
      nx207, nx211, nx215, nx221, nx223, nx225, nx229, nx232, nx235, nx239, 
      nx241, nx243, nx246, nx249, nx252, nx256, nx258, nx260, nx263, nx266, 
      nx269, nx273, nx275, nx277, nx280, nx283, nx286, nx290, nx292, nx294, 
      nx297, nx300, nx303, nx307, nx309, nx311, nx314, nx317, nx320, nx323, 
      nx326, nx329, nx332, nx335, nx338, nx341, nx344, nx347, nx350, nx353, 
      nx356, nx358, nx360, nx362, nx364, nx366, nx368, nx370, nx372: 
   std_logic ;

begin
   ix44 : fake_gnd port map ( Y=>carryOut);
   ix229 : xnor2 port map ( Y=>sum(0), A0=>carryIn, A1=>nx103);
   ix104 : xnor2 port map ( Y=>nx103, A0=>a(0), A1=>b(0));
   ix227 : xnor2 port map ( Y=>sum(1), A0=>nx6, A1=>nx115);
   ix7 : oai22 port map ( Y=>nx6, A0=>nx109, A1=>nx103, B0=>nx111, B1=>nx113
   );
   ix110 : inv01 port map ( Y=>nx109, A=>carryIn);
   ix112 : inv01 port map ( Y=>nx111, A=>b(0));
   ix114 : inv01 port map ( Y=>nx113, A=>a(0));
   ix116 : xnor2 port map ( Y=>nx115, A0=>a(1), A1=>b(1));
   ix225 : xnor2 port map ( Y=>sum(2), A0=>nx119, A1=>nx16);
   ix120 : aoi22 port map ( Y=>nx119, A0=>b(1), A1=>a(1), B0=>nx6, B1=>nx8);
   ix9 : xnor2 port map ( Y=>nx8, A0=>a(1), A1=>nx123);
   ix124 : inv01 port map ( Y=>nx123, A=>b(1));
   ix17 : xnor2 port map ( Y=>nx16, A0=>a(2), A1=>nx127);
   ix128 : inv01 port map ( Y=>nx127, A=>b(2));
   ix223 : xnor2 port map ( Y=>sum(3), A0=>nx22, A1=>nx137);
   ix23 : oai21 port map ( Y=>nx22, A0=>nx119, A1=>nx133, B0=>nx135);
   ix134 : xnor2 port map ( Y=>nx133, A0=>a(2), A1=>b(2));
   ix136 : nand02 port map ( Y=>nx135, A0=>b(2), A1=>a(2));
   ix138 : xnor2 port map ( Y=>nx137, A0=>a(3), A1=>b(3));
   ix221 : xnor2 port map ( Y=>sum(4), A0=>nx141, A1=>nx32);
   ix142 : aoi22 port map ( Y=>nx141, A0=>b(3), A1=>a(3), B0=>nx22, B1=>nx24
   );
   ix25 : xnor2 port map ( Y=>nx24, A0=>a(3), A1=>nx145);
   ix146 : inv01 port map ( Y=>nx145, A=>b(3));
   ix33 : xnor2 port map ( Y=>nx32, A0=>a(4), A1=>nx149);
   ix150 : inv01 port map ( Y=>nx149, A=>b(4));
   ix219 : xnor2 port map ( Y=>sum(5), A0=>nx38, A1=>nx159);
   ix39 : oai21 port map ( Y=>nx38, A0=>nx141, A1=>nx155, B0=>nx157);
   ix156 : xnor2 port map ( Y=>nx155, A0=>a(4), A1=>b(4));
   ix158 : nand02 port map ( Y=>nx157, A0=>b(4), A1=>a(4));
   ix160 : xnor2 port map ( Y=>nx159, A0=>a(5), A1=>b(5));
   ix217 : xnor2 port map ( Y=>sum(6), A0=>nx163, A1=>nx48);
   ix164 : aoi22 port map ( Y=>nx163, A0=>b(5), A1=>a(5), B0=>nx38, B1=>nx40
   );
   ix41 : xnor2 port map ( Y=>nx40, A0=>a(5), A1=>nx167);
   ix168 : inv01 port map ( Y=>nx167, A=>b(5));
   ix49 : xnor2 port map ( Y=>nx48, A0=>a(6), A1=>nx171);
   ix172 : inv01 port map ( Y=>nx171, A=>b(6));
   ix215 : xnor2 port map ( Y=>sum(7), A0=>nx54, A1=>nx181);
   ix55 : oai21 port map ( Y=>nx54, A0=>nx163, A1=>nx177, B0=>nx179);
   ix178 : xnor2 port map ( Y=>nx177, A0=>a(6), A1=>b(6));
   ix180 : nand02 port map ( Y=>nx179, A0=>b(6), A1=>a(6));
   ix182 : xnor2 port map ( Y=>nx181, A0=>a(7), A1=>b(7));
   ix213 : xnor2 port map ( Y=>sum(8), A0=>nx185, A1=>nx64);
   ix186 : aoi22 port map ( Y=>nx185, A0=>b(7), A1=>a(7), B0=>nx54, B1=>nx56
   );
   ix57 : xnor2 port map ( Y=>nx56, A0=>a(7), A1=>nx189);
   ix190 : inv01 port map ( Y=>nx189, A=>b(7));
   ix65 : xnor2 port map ( Y=>nx64, A0=>a(8), A1=>nx193);
   ix194 : inv01 port map ( Y=>nx193, A=>b(8));
   ix211 : xnor2 port map ( Y=>sum(9), A0=>nx70, A1=>nx203);
   ix71 : oai21 port map ( Y=>nx70, A0=>nx185, A1=>nx199, B0=>nx201);
   ix200 : xnor2 port map ( Y=>nx199, A0=>a(8), A1=>b(8));
   ix202 : nand02 port map ( Y=>nx201, A0=>b(8), A1=>a(8));
   ix204 : xnor2 port map ( Y=>nx203, A0=>a(9), A1=>b(9));
   ix209 : xnor2 port map ( Y=>sum(10), A0=>nx207, A1=>nx80);
   ix208 : aoi22 port map ( Y=>nx207, A0=>b(9), A1=>a(9), B0=>nx70, B1=>nx72
   );
   ix73 : xnor2 port map ( Y=>nx72, A0=>a(9), A1=>nx211);
   ix212 : inv01 port map ( Y=>nx211, A=>b(9));
   ix81 : xnor2 port map ( Y=>nx80, A0=>a(10), A1=>nx215);
   ix216 : inv01 port map ( Y=>nx215, A=>b(10));
   ix207 : xnor2 port map ( Y=>sum(11), A0=>nx86, A1=>nx225);
   ix87 : oai21 port map ( Y=>nx86, A0=>nx207, A1=>nx221, B0=>nx223);
   ix222 : xnor2 port map ( Y=>nx221, A0=>a(10), A1=>b(10));
   ix224 : nand02 port map ( Y=>nx223, A0=>b(10), A1=>a(10));
   ix226 : xnor2 port map ( Y=>nx225, A0=>a(11), A1=>b(11));
   ix205 : xnor2 port map ( Y=>sum(12), A0=>nx229, A1=>nx96);
   ix230 : aoi22 port map ( Y=>nx229, A0=>b(11), A1=>a(11), B0=>nx86, B1=>
      nx88);
   ix89 : xnor2 port map ( Y=>nx88, A0=>a(11), A1=>nx232);
   ix233 : inv01 port map ( Y=>nx232, A=>b(11));
   ix97 : xnor2 port map ( Y=>nx96, A0=>a(12), A1=>nx235);
   ix236 : inv01 port map ( Y=>nx235, A=>b(12));
   ix203 : xnor2 port map ( Y=>sum(13), A0=>nx102, A1=>nx243);
   ix103 : oai21 port map ( Y=>nx102, A0=>nx229, A1=>nx239, B0=>nx241);
   ix240 : xnor2 port map ( Y=>nx239, A0=>a(12), A1=>b(12));
   ix242 : nand02 port map ( Y=>nx241, A0=>b(12), A1=>a(12));
   ix244 : xnor2 port map ( Y=>nx243, A0=>a(13), A1=>b(13));
   ix201 : xnor2 port map ( Y=>sum(14), A0=>nx246, A1=>nx112);
   ix247 : aoi22 port map ( Y=>nx246, A0=>b(13), A1=>a(13), B0=>nx102, B1=>
      nx104);
   ix105 : xnor2 port map ( Y=>nx104, A0=>a(13), A1=>nx249);
   ix250 : inv01 port map ( Y=>nx249, A=>b(13));
   ix113 : xnor2 port map ( Y=>nx112, A0=>a(14), A1=>nx252);
   ix253 : inv01 port map ( Y=>nx252, A=>b(14));
   ix199 : xnor2 port map ( Y=>sum(15), A0=>nx118, A1=>nx260);
   ix119 : oai21 port map ( Y=>nx118, A0=>nx246, A1=>nx256, B0=>nx258);
   ix257 : xnor2 port map ( Y=>nx256, A0=>a(14), A1=>b(14));
   ix259 : nand02 port map ( Y=>nx258, A0=>b(14), A1=>a(14));
   ix261 : xnor2 port map ( Y=>nx260, A0=>a(15), A1=>b(15));
   ix197 : xnor2 port map ( Y=>sum(16), A0=>nx263, A1=>nx128);
   ix264 : aoi22 port map ( Y=>nx263, A0=>b(15), A1=>a(15), B0=>nx118, B1=>
      nx120);
   ix121 : xnor2 port map ( Y=>nx120, A0=>a(15), A1=>nx266);
   ix267 : inv01 port map ( Y=>nx266, A=>b(15));
   ix129 : xnor2 port map ( Y=>nx128, A0=>a(16), A1=>nx269);
   ix270 : inv01 port map ( Y=>nx269, A=>b(16));
   ix195 : xnor2 port map ( Y=>sum(17), A0=>nx134, A1=>nx277);
   ix135 : oai21 port map ( Y=>nx134, A0=>nx263, A1=>nx273, B0=>nx275);
   ix274 : xnor2 port map ( Y=>nx273, A0=>a(16), A1=>b(16));
   ix276 : nand02 port map ( Y=>nx275, A0=>b(16), A1=>a(16));
   ix278 : xnor2 port map ( Y=>nx277, A0=>a(17), A1=>b(17));
   ix193 : xnor2 port map ( Y=>sum(18), A0=>nx280, A1=>nx144);
   ix281 : aoi22 port map ( Y=>nx280, A0=>b(17), A1=>a(17), B0=>nx134, B1=>
      nx136);
   ix137 : xnor2 port map ( Y=>nx136, A0=>a(17), A1=>nx283);
   ix284 : inv01 port map ( Y=>nx283, A=>b(17));
   ix145 : xnor2 port map ( Y=>nx144, A0=>a(18), A1=>nx286);
   ix287 : inv01 port map ( Y=>nx286, A=>b(18));
   ix191 : xnor2 port map ( Y=>sum(19), A0=>nx150, A1=>nx294);
   ix151 : oai21 port map ( Y=>nx150, A0=>nx280, A1=>nx290, B0=>nx292);
   ix291 : xnor2 port map ( Y=>nx290, A0=>a(18), A1=>b(18));
   ix293 : nand02 port map ( Y=>nx292, A0=>b(18), A1=>a(18));
   ix295 : xnor2 port map ( Y=>nx294, A0=>a(19), A1=>b(19));
   ix189 : xnor2 port map ( Y=>sum(20), A0=>nx297, A1=>nx160);
   ix298 : aoi22 port map ( Y=>nx297, A0=>b(19), A1=>a(19), B0=>nx150, B1=>
      nx152);
   ix153 : xnor2 port map ( Y=>nx152, A0=>a(19), A1=>nx300);
   ix301 : inv01 port map ( Y=>nx300, A=>b(19));
   ix161 : xnor2 port map ( Y=>nx160, A0=>a(20), A1=>nx303);
   ix304 : inv01 port map ( Y=>nx303, A=>b(20));
   ix187 : xnor2 port map ( Y=>sum(21), A0=>nx166, A1=>nx311);
   ix167 : oai21 port map ( Y=>nx166, A0=>nx297, A1=>nx307, B0=>nx309);
   ix308 : xnor2 port map ( Y=>nx307, A0=>a(20), A1=>b(20));
   ix310 : nand02 port map ( Y=>nx309, A0=>b(20), A1=>a(20));
   ix312 : xnor2 port map ( Y=>nx311, A0=>a(21), A1=>b(21));
   ix185 : xnor2 port map ( Y=>sum(22), A0=>b(22), A1=>nx314);
   ix315 : aoi22 port map ( Y=>nx314, A0=>b(21), A1=>a(21), B0=>nx166, B1=>
      nx168);
   ix169 : xnor2 port map ( Y=>nx168, A0=>a(21), A1=>nx317);
   ix318 : inv01 port map ( Y=>nx317, A=>b(21));
   ix179 : xnor2 port map ( Y=>sum(23), A0=>b(23), A1=>nx320);
   ix321 : oai21 port map ( Y=>nx320, A0=>nx172, A1=>nx170, B0=>b(22));
   ix173 : nor02_2x port map ( Y=>nx172, A0=>nx317, A1=>nx323);
   ix324 : inv01 port map ( Y=>nx323, A=>a(21));
   ix171 : nor02ii port map ( Y=>nx170, A0=>nx326, A1=>nx168);
   ix327 : aoi22 port map ( Y=>nx326, A0=>b(20), A1=>a(20), B0=>nx158, B1=>
      nx160);
   ix159 : oai21 port map ( Y=>nx158, A0=>nx329, A1=>nx294, B0=>nx372);
   ix330 : aoi22 port map ( Y=>nx329, A0=>b(18), A1=>a(18), B0=>nx142, B1=>
      nx144);
   ix143 : oai21 port map ( Y=>nx142, A0=>nx332, A1=>nx277, B0=>nx370);
   ix333 : aoi22 port map ( Y=>nx332, A0=>b(16), A1=>a(16), B0=>nx126, B1=>
      nx128);
   ix127 : oai21 port map ( Y=>nx126, A0=>nx335, A1=>nx260, B0=>nx368);
   ix336 : aoi22 port map ( Y=>nx335, A0=>b(14), A1=>a(14), B0=>nx110, B1=>
      nx112);
   ix111 : oai21 port map ( Y=>nx110, A0=>nx338, A1=>nx243, B0=>nx366);
   ix339 : aoi22 port map ( Y=>nx338, A0=>b(12), A1=>a(12), B0=>nx94, B1=>
      nx96);
   ix95 : oai21 port map ( Y=>nx94, A0=>nx341, A1=>nx225, B0=>nx364);
   ix342 : aoi22 port map ( Y=>nx341, A0=>b(10), A1=>a(10), B0=>nx78, B1=>
      nx80);
   ix79 : oai21 port map ( Y=>nx78, A0=>nx344, A1=>nx203, B0=>nx362);
   ix345 : aoi22 port map ( Y=>nx344, A0=>b(8), A1=>a(8), B0=>nx62, B1=>nx64
   );
   ix63 : oai21 port map ( Y=>nx62, A0=>nx347, A1=>nx181, B0=>nx360);
   ix348 : aoi22 port map ( Y=>nx347, A0=>b(6), A1=>a(6), B0=>nx46, B1=>nx48
   );
   ix47 : oai21 port map ( Y=>nx46, A0=>nx350, A1=>nx159, B0=>nx358);
   ix351 : aoi22 port map ( Y=>nx350, A0=>b(4), A1=>a(4), B0=>nx30, B1=>nx32
   );
   ix31 : oai21 port map ( Y=>nx30, A0=>nx353, A1=>nx137, B0=>nx356);
   ix354 : aoi21 port map ( Y=>nx353, A0=>b(2), A1=>a(2), B0=>nx18);
   ix19 : nor02ii port map ( Y=>nx18, A0=>nx119, A1=>nx16);
   ix357 : nand02 port map ( Y=>nx356, A0=>b(3), A1=>a(3));
   ix359 : nand02 port map ( Y=>nx358, A0=>b(5), A1=>a(5));
   ix361 : nand02 port map ( Y=>nx360, A0=>b(7), A1=>a(7));
   ix363 : nand02 port map ( Y=>nx362, A0=>b(9), A1=>a(9));
   ix365 : nand02 port map ( Y=>nx364, A0=>b(11), A1=>a(11));
   ix367 : nand02 port map ( Y=>nx366, A0=>b(13), A1=>a(13));
   ix369 : nand02 port map ( Y=>nx368, A0=>b(15), A1=>a(15));
   ix371 : nand02 port map ( Y=>nx370, A0=>b(17), A1=>a(17));
   ix373 : nand02 port map ( Y=>nx372, A0=>b(19), A1=>a(19));
end NBitAdderArch_unfold_2081 ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity CNNMuls is
   port (
      filter_24_7 : IN std_logic ;
      filter_24_6 : IN std_logic ;
      filter_24_5 : IN std_logic ;
      filter_24_4 : IN std_logic ;
      filter_24_3 : IN std_logic ;
      filter_24_2 : IN std_logic ;
      filter_24_1 : IN std_logic ;
      filter_24_0 : IN std_logic ;
      filter_23_7 : IN std_logic ;
      filter_23_6 : IN std_logic ;
      filter_23_5 : IN std_logic ;
      filter_23_4 : IN std_logic ;
      filter_23_3 : IN std_logic ;
      filter_23_2 : IN std_logic ;
      filter_23_1 : IN std_logic ;
      filter_23_0 : IN std_logic ;
      filter_22_7 : IN std_logic ;
      filter_22_6 : IN std_logic ;
      filter_22_5 : IN std_logic ;
      filter_22_4 : IN std_logic ;
      filter_22_3 : IN std_logic ;
      filter_22_2 : IN std_logic ;
      filter_22_1 : IN std_logic ;
      filter_22_0 : IN std_logic ;
      filter_21_7 : IN std_logic ;
      filter_21_6 : IN std_logic ;
      filter_21_5 : IN std_logic ;
      filter_21_4 : IN std_logic ;
      filter_21_3 : IN std_logic ;
      filter_21_2 : IN std_logic ;
      filter_21_1 : IN std_logic ;
      filter_21_0 : IN std_logic ;
      filter_20_7 : IN std_logic ;
      filter_20_6 : IN std_logic ;
      filter_20_5 : IN std_logic ;
      filter_20_4 : IN std_logic ;
      filter_20_3 : IN std_logic ;
      filter_20_2 : IN std_logic ;
      filter_20_1 : IN std_logic ;
      filter_20_0 : IN std_logic ;
      filter_19_7 : IN std_logic ;
      filter_19_6 : IN std_logic ;
      filter_19_5 : IN std_logic ;
      filter_19_4 : IN std_logic ;
      filter_19_3 : IN std_logic ;
      filter_19_2 : IN std_logic ;
      filter_19_1 : IN std_logic ;
      filter_19_0 : IN std_logic ;
      filter_18_7 : IN std_logic ;
      filter_18_6 : IN std_logic ;
      filter_18_5 : IN std_logic ;
      filter_18_4 : IN std_logic ;
      filter_18_3 : IN std_logic ;
      filter_18_2 : IN std_logic ;
      filter_18_1 : IN std_logic ;
      filter_18_0 : IN std_logic ;
      filter_17_7 : IN std_logic ;
      filter_17_6 : IN std_logic ;
      filter_17_5 : IN std_logic ;
      filter_17_4 : IN std_logic ;
      filter_17_3 : IN std_logic ;
      filter_17_2 : IN std_logic ;
      filter_17_1 : IN std_logic ;
      filter_17_0 : IN std_logic ;
      filter_16_7 : IN std_logic ;
      filter_16_6 : IN std_logic ;
      filter_16_5 : IN std_logic ;
      filter_16_4 : IN std_logic ;
      filter_16_3 : IN std_logic ;
      filter_16_2 : IN std_logic ;
      filter_16_1 : IN std_logic ;
      filter_16_0 : IN std_logic ;
      filter_15_7 : IN std_logic ;
      filter_15_6 : IN std_logic ;
      filter_15_5 : IN std_logic ;
      filter_15_4 : IN std_logic ;
      filter_15_3 : IN std_logic ;
      filter_15_2 : IN std_logic ;
      filter_15_1 : IN std_logic ;
      filter_15_0 : IN std_logic ;
      filter_14_7 : IN std_logic ;
      filter_14_6 : IN std_logic ;
      filter_14_5 : IN std_logic ;
      filter_14_4 : IN std_logic ;
      filter_14_3 : IN std_logic ;
      filter_14_2 : IN std_logic ;
      filter_14_1 : IN std_logic ;
      filter_14_0 : IN std_logic ;
      filter_13_7 : IN std_logic ;
      filter_13_6 : IN std_logic ;
      filter_13_5 : IN std_logic ;
      filter_13_4 : IN std_logic ;
      filter_13_3 : IN std_logic ;
      filter_13_2 : IN std_logic ;
      filter_13_1 : IN std_logic ;
      filter_13_0 : IN std_logic ;
      filter_12_7 : IN std_logic ;
      filter_12_6 : IN std_logic ;
      filter_12_5 : IN std_logic ;
      filter_12_4 : IN std_logic ;
      filter_12_3 : IN std_logic ;
      filter_12_2 : IN std_logic ;
      filter_12_1 : IN std_logic ;
      filter_12_0 : IN std_logic ;
      filter_11_7 : IN std_logic ;
      filter_11_6 : IN std_logic ;
      filter_11_5 : IN std_logic ;
      filter_11_4 : IN std_logic ;
      filter_11_3 : IN std_logic ;
      filter_11_2 : IN std_logic ;
      filter_11_1 : IN std_logic ;
      filter_11_0 : IN std_logic ;
      filter_10_7 : IN std_logic ;
      filter_10_6 : IN std_logic ;
      filter_10_5 : IN std_logic ;
      filter_10_4 : IN std_logic ;
      filter_10_3 : IN std_logic ;
      filter_10_2 : IN std_logic ;
      filter_10_1 : IN std_logic ;
      filter_10_0 : IN std_logic ;
      filter_9_7 : IN std_logic ;
      filter_9_6 : IN std_logic ;
      filter_9_5 : IN std_logic ;
      filter_9_4 : IN std_logic ;
      filter_9_3 : IN std_logic ;
      filter_9_2 : IN std_logic ;
      filter_9_1 : IN std_logic ;
      filter_9_0 : IN std_logic ;
      filter_8_7 : IN std_logic ;
      filter_8_6 : IN std_logic ;
      filter_8_5 : IN std_logic ;
      filter_8_4 : IN std_logic ;
      filter_8_3 : IN std_logic ;
      filter_8_2 : IN std_logic ;
      filter_8_1 : IN std_logic ;
      filter_8_0 : IN std_logic ;
      filter_7_7 : IN std_logic ;
      filter_7_6 : IN std_logic ;
      filter_7_5 : IN std_logic ;
      filter_7_4 : IN std_logic ;
      filter_7_3 : IN std_logic ;
      filter_7_2 : IN std_logic ;
      filter_7_1 : IN std_logic ;
      filter_7_0 : IN std_logic ;
      filter_6_7 : IN std_logic ;
      filter_6_6 : IN std_logic ;
      filter_6_5 : IN std_logic ;
      filter_6_4 : IN std_logic ;
      filter_6_3 : IN std_logic ;
      filter_6_2 : IN std_logic ;
      filter_6_1 : IN std_logic ;
      filter_6_0 : IN std_logic ;
      filter_5_7 : IN std_logic ;
      filter_5_6 : IN std_logic ;
      filter_5_5 : IN std_logic ;
      filter_5_4 : IN std_logic ;
      filter_5_3 : IN std_logic ;
      filter_5_2 : IN std_logic ;
      filter_5_1 : IN std_logic ;
      filter_5_0 : IN std_logic ;
      filter_4_7 : IN std_logic ;
      filter_4_6 : IN std_logic ;
      filter_4_5 : IN std_logic ;
      filter_4_4 : IN std_logic ;
      filter_4_3 : IN std_logic ;
      filter_4_2 : IN std_logic ;
      filter_4_1 : IN std_logic ;
      filter_4_0 : IN std_logic ;
      filter_3_7 : IN std_logic ;
      filter_3_6 : IN std_logic ;
      filter_3_5 : IN std_logic ;
      filter_3_4 : IN std_logic ;
      filter_3_3 : IN std_logic ;
      filter_3_2 : IN std_logic ;
      filter_3_1 : IN std_logic ;
      filter_3_0 : IN std_logic ;
      filter_2_7 : IN std_logic ;
      filter_2_6 : IN std_logic ;
      filter_2_5 : IN std_logic ;
      filter_2_4 : IN std_logic ;
      filter_2_3 : IN std_logic ;
      filter_2_2 : IN std_logic ;
      filter_2_1 : IN std_logic ;
      filter_2_0 : IN std_logic ;
      filter_1_7 : IN std_logic ;
      filter_1_6 : IN std_logic ;
      filter_1_5 : IN std_logic ;
      filter_1_4 : IN std_logic ;
      filter_1_3 : IN std_logic ;
      filter_1_2 : IN std_logic ;
      filter_1_1 : IN std_logic ;
      filter_1_0 : IN std_logic ;
      filter_0_7 : IN std_logic ;
      filter_0_6 : IN std_logic ;
      filter_0_5 : IN std_logic ;
      filter_0_4 : IN std_logic ;
      filter_0_3 : IN std_logic ;
      filter_0_2 : IN std_logic ;
      filter_0_1 : IN std_logic ;
      filter_0_0 : IN std_logic ;
      window_24_15 : IN std_logic ;
      window_24_14 : IN std_logic ;
      window_24_13 : IN std_logic ;
      window_24_12 : IN std_logic ;
      window_24_11 : IN std_logic ;
      window_24_10 : IN std_logic ;
      window_24_9 : IN std_logic ;
      window_24_8 : IN std_logic ;
      window_24_7 : IN std_logic ;
      window_24_6 : IN std_logic ;
      window_24_5 : IN std_logic ;
      window_24_4 : IN std_logic ;
      window_24_3 : IN std_logic ;
      window_24_2 : IN std_logic ;
      window_24_1 : IN std_logic ;
      window_24_0 : IN std_logic ;
      window_23_15 : IN std_logic ;
      window_23_14 : IN std_logic ;
      window_23_13 : IN std_logic ;
      window_23_12 : IN std_logic ;
      window_23_11 : IN std_logic ;
      window_23_10 : IN std_logic ;
      window_23_9 : IN std_logic ;
      window_23_8 : IN std_logic ;
      window_23_7 : IN std_logic ;
      window_23_6 : IN std_logic ;
      window_23_5 : IN std_logic ;
      window_23_4 : IN std_logic ;
      window_23_3 : IN std_logic ;
      window_23_2 : IN std_logic ;
      window_23_1 : IN std_logic ;
      window_23_0 : IN std_logic ;
      window_22_15 : IN std_logic ;
      window_22_14 : IN std_logic ;
      window_22_13 : IN std_logic ;
      window_22_12 : IN std_logic ;
      window_22_11 : IN std_logic ;
      window_22_10 : IN std_logic ;
      window_22_9 : IN std_logic ;
      window_22_8 : IN std_logic ;
      window_22_7 : IN std_logic ;
      window_22_6 : IN std_logic ;
      window_22_5 : IN std_logic ;
      window_22_4 : IN std_logic ;
      window_22_3 : IN std_logic ;
      window_22_2 : IN std_logic ;
      window_22_1 : IN std_logic ;
      window_22_0 : IN std_logic ;
      window_21_15 : IN std_logic ;
      window_21_14 : IN std_logic ;
      window_21_13 : IN std_logic ;
      window_21_12 : IN std_logic ;
      window_21_11 : IN std_logic ;
      window_21_10 : IN std_logic ;
      window_21_9 : IN std_logic ;
      window_21_8 : IN std_logic ;
      window_21_7 : IN std_logic ;
      window_21_6 : IN std_logic ;
      window_21_5 : IN std_logic ;
      window_21_4 : IN std_logic ;
      window_21_3 : IN std_logic ;
      window_21_2 : IN std_logic ;
      window_21_1 : IN std_logic ;
      window_21_0 : IN std_logic ;
      window_20_15 : IN std_logic ;
      window_20_14 : IN std_logic ;
      window_20_13 : IN std_logic ;
      window_20_12 : IN std_logic ;
      window_20_11 : IN std_logic ;
      window_20_10 : IN std_logic ;
      window_20_9 : IN std_logic ;
      window_20_8 : IN std_logic ;
      window_20_7 : IN std_logic ;
      window_20_6 : IN std_logic ;
      window_20_5 : IN std_logic ;
      window_20_4 : IN std_logic ;
      window_20_3 : IN std_logic ;
      window_20_2 : IN std_logic ;
      window_20_1 : IN std_logic ;
      window_20_0 : IN std_logic ;
      window_19_15 : IN std_logic ;
      window_19_14 : IN std_logic ;
      window_19_13 : IN std_logic ;
      window_19_12 : IN std_logic ;
      window_19_11 : IN std_logic ;
      window_19_10 : IN std_logic ;
      window_19_9 : IN std_logic ;
      window_19_8 : IN std_logic ;
      window_19_7 : IN std_logic ;
      window_19_6 : IN std_logic ;
      window_19_5 : IN std_logic ;
      window_19_4 : IN std_logic ;
      window_19_3 : IN std_logic ;
      window_19_2 : IN std_logic ;
      window_19_1 : IN std_logic ;
      window_19_0 : IN std_logic ;
      window_18_15 : IN std_logic ;
      window_18_14 : IN std_logic ;
      window_18_13 : IN std_logic ;
      window_18_12 : IN std_logic ;
      window_18_11 : IN std_logic ;
      window_18_10 : IN std_logic ;
      window_18_9 : IN std_logic ;
      window_18_8 : IN std_logic ;
      window_18_7 : IN std_logic ;
      window_18_6 : IN std_logic ;
      window_18_5 : IN std_logic ;
      window_18_4 : IN std_logic ;
      window_18_3 : IN std_logic ;
      window_18_2 : IN std_logic ;
      window_18_1 : IN std_logic ;
      window_18_0 : IN std_logic ;
      window_17_15 : IN std_logic ;
      window_17_14 : IN std_logic ;
      window_17_13 : IN std_logic ;
      window_17_12 : IN std_logic ;
      window_17_11 : IN std_logic ;
      window_17_10 : IN std_logic ;
      window_17_9 : IN std_logic ;
      window_17_8 : IN std_logic ;
      window_17_7 : IN std_logic ;
      window_17_6 : IN std_logic ;
      window_17_5 : IN std_logic ;
      window_17_4 : IN std_logic ;
      window_17_3 : IN std_logic ;
      window_17_2 : IN std_logic ;
      window_17_1 : IN std_logic ;
      window_17_0 : IN std_logic ;
      window_16_15 : IN std_logic ;
      window_16_14 : IN std_logic ;
      window_16_13 : IN std_logic ;
      window_16_12 : IN std_logic ;
      window_16_11 : IN std_logic ;
      window_16_10 : IN std_logic ;
      window_16_9 : IN std_logic ;
      window_16_8 : IN std_logic ;
      window_16_7 : IN std_logic ;
      window_16_6 : IN std_logic ;
      window_16_5 : IN std_logic ;
      window_16_4 : IN std_logic ;
      window_16_3 : IN std_logic ;
      window_16_2 : IN std_logic ;
      window_16_1 : IN std_logic ;
      window_16_0 : IN std_logic ;
      window_15_15 : IN std_logic ;
      window_15_14 : IN std_logic ;
      window_15_13 : IN std_logic ;
      window_15_12 : IN std_logic ;
      window_15_11 : IN std_logic ;
      window_15_10 : IN std_logic ;
      window_15_9 : IN std_logic ;
      window_15_8 : IN std_logic ;
      window_15_7 : IN std_logic ;
      window_15_6 : IN std_logic ;
      window_15_5 : IN std_logic ;
      window_15_4 : IN std_logic ;
      window_15_3 : IN std_logic ;
      window_15_2 : IN std_logic ;
      window_15_1 : IN std_logic ;
      window_15_0 : IN std_logic ;
      window_14_15 : IN std_logic ;
      window_14_14 : IN std_logic ;
      window_14_13 : IN std_logic ;
      window_14_12 : IN std_logic ;
      window_14_11 : IN std_logic ;
      window_14_10 : IN std_logic ;
      window_14_9 : IN std_logic ;
      window_14_8 : IN std_logic ;
      window_14_7 : IN std_logic ;
      window_14_6 : IN std_logic ;
      window_14_5 : IN std_logic ;
      window_14_4 : IN std_logic ;
      window_14_3 : IN std_logic ;
      window_14_2 : IN std_logic ;
      window_14_1 : IN std_logic ;
      window_14_0 : IN std_logic ;
      window_13_15 : IN std_logic ;
      window_13_14 : IN std_logic ;
      window_13_13 : IN std_logic ;
      window_13_12 : IN std_logic ;
      window_13_11 : IN std_logic ;
      window_13_10 : IN std_logic ;
      window_13_9 : IN std_logic ;
      window_13_8 : IN std_logic ;
      window_13_7 : IN std_logic ;
      window_13_6 : IN std_logic ;
      window_13_5 : IN std_logic ;
      window_13_4 : IN std_logic ;
      window_13_3 : IN std_logic ;
      window_13_2 : IN std_logic ;
      window_13_1 : IN std_logic ;
      window_13_0 : IN std_logic ;
      window_12_15 : IN std_logic ;
      window_12_14 : IN std_logic ;
      window_12_13 : IN std_logic ;
      window_12_12 : IN std_logic ;
      window_12_11 : IN std_logic ;
      window_12_10 : IN std_logic ;
      window_12_9 : IN std_logic ;
      window_12_8 : IN std_logic ;
      window_12_7 : IN std_logic ;
      window_12_6 : IN std_logic ;
      window_12_5 : IN std_logic ;
      window_12_4 : IN std_logic ;
      window_12_3 : IN std_logic ;
      window_12_2 : IN std_logic ;
      window_12_1 : IN std_logic ;
      window_12_0 : IN std_logic ;
      window_11_15 : IN std_logic ;
      window_11_14 : IN std_logic ;
      window_11_13 : IN std_logic ;
      window_11_12 : IN std_logic ;
      window_11_11 : IN std_logic ;
      window_11_10 : IN std_logic ;
      window_11_9 : IN std_logic ;
      window_11_8 : IN std_logic ;
      window_11_7 : IN std_logic ;
      window_11_6 : IN std_logic ;
      window_11_5 : IN std_logic ;
      window_11_4 : IN std_logic ;
      window_11_3 : IN std_logic ;
      window_11_2 : IN std_logic ;
      window_11_1 : IN std_logic ;
      window_11_0 : IN std_logic ;
      window_10_15 : IN std_logic ;
      window_10_14 : IN std_logic ;
      window_10_13 : IN std_logic ;
      window_10_12 : IN std_logic ;
      window_10_11 : IN std_logic ;
      window_10_10 : IN std_logic ;
      window_10_9 : IN std_logic ;
      window_10_8 : IN std_logic ;
      window_10_7 : IN std_logic ;
      window_10_6 : IN std_logic ;
      window_10_5 : IN std_logic ;
      window_10_4 : IN std_logic ;
      window_10_3 : IN std_logic ;
      window_10_2 : IN std_logic ;
      window_10_1 : IN std_logic ;
      window_10_0 : IN std_logic ;
      window_9_15 : IN std_logic ;
      window_9_14 : IN std_logic ;
      window_9_13 : IN std_logic ;
      window_9_12 : IN std_logic ;
      window_9_11 : IN std_logic ;
      window_9_10 : IN std_logic ;
      window_9_9 : IN std_logic ;
      window_9_8 : IN std_logic ;
      window_9_7 : IN std_logic ;
      window_9_6 : IN std_logic ;
      window_9_5 : IN std_logic ;
      window_9_4 : IN std_logic ;
      window_9_3 : IN std_logic ;
      window_9_2 : IN std_logic ;
      window_9_1 : IN std_logic ;
      window_9_0 : IN std_logic ;
      window_8_15 : IN std_logic ;
      window_8_14 : IN std_logic ;
      window_8_13 : IN std_logic ;
      window_8_12 : IN std_logic ;
      window_8_11 : IN std_logic ;
      window_8_10 : IN std_logic ;
      window_8_9 : IN std_logic ;
      window_8_8 : IN std_logic ;
      window_8_7 : IN std_logic ;
      window_8_6 : IN std_logic ;
      window_8_5 : IN std_logic ;
      window_8_4 : IN std_logic ;
      window_8_3 : IN std_logic ;
      window_8_2 : IN std_logic ;
      window_8_1 : IN std_logic ;
      window_8_0 : IN std_logic ;
      window_7_15 : IN std_logic ;
      window_7_14 : IN std_logic ;
      window_7_13 : IN std_logic ;
      window_7_12 : IN std_logic ;
      window_7_11 : IN std_logic ;
      window_7_10 : IN std_logic ;
      window_7_9 : IN std_logic ;
      window_7_8 : IN std_logic ;
      window_7_7 : IN std_logic ;
      window_7_6 : IN std_logic ;
      window_7_5 : IN std_logic ;
      window_7_4 : IN std_logic ;
      window_7_3 : IN std_logic ;
      window_7_2 : IN std_logic ;
      window_7_1 : IN std_logic ;
      window_7_0 : IN std_logic ;
      window_6_15 : IN std_logic ;
      window_6_14 : IN std_logic ;
      window_6_13 : IN std_logic ;
      window_6_12 : IN std_logic ;
      window_6_11 : IN std_logic ;
      window_6_10 : IN std_logic ;
      window_6_9 : IN std_logic ;
      window_6_8 : IN std_logic ;
      window_6_7 : IN std_logic ;
      window_6_6 : IN std_logic ;
      window_6_5 : IN std_logic ;
      window_6_4 : IN std_logic ;
      window_6_3 : IN std_logic ;
      window_6_2 : IN std_logic ;
      window_6_1 : IN std_logic ;
      window_6_0 : IN std_logic ;
      window_5_15 : IN std_logic ;
      window_5_14 : IN std_logic ;
      window_5_13 : IN std_logic ;
      window_5_12 : IN std_logic ;
      window_5_11 : IN std_logic ;
      window_5_10 : IN std_logic ;
      window_5_9 : IN std_logic ;
      window_5_8 : IN std_logic ;
      window_5_7 : IN std_logic ;
      window_5_6 : IN std_logic ;
      window_5_5 : IN std_logic ;
      window_5_4 : IN std_logic ;
      window_5_3 : IN std_logic ;
      window_5_2 : IN std_logic ;
      window_5_1 : IN std_logic ;
      window_5_0 : IN std_logic ;
      window_4_15 : IN std_logic ;
      window_4_14 : IN std_logic ;
      window_4_13 : IN std_logic ;
      window_4_12 : IN std_logic ;
      window_4_11 : IN std_logic ;
      window_4_10 : IN std_logic ;
      window_4_9 : IN std_logic ;
      window_4_8 : IN std_logic ;
      window_4_7 : IN std_logic ;
      window_4_6 : IN std_logic ;
      window_4_5 : IN std_logic ;
      window_4_4 : IN std_logic ;
      window_4_3 : IN std_logic ;
      window_4_2 : IN std_logic ;
      window_4_1 : IN std_logic ;
      window_4_0 : IN std_logic ;
      window_3_15 : IN std_logic ;
      window_3_14 : IN std_logic ;
      window_3_13 : IN std_logic ;
      window_3_12 : IN std_logic ;
      window_3_11 : IN std_logic ;
      window_3_10 : IN std_logic ;
      window_3_9 : IN std_logic ;
      window_3_8 : IN std_logic ;
      window_3_7 : IN std_logic ;
      window_3_6 : IN std_logic ;
      window_3_5 : IN std_logic ;
      window_3_4 : IN std_logic ;
      window_3_3 : IN std_logic ;
      window_3_2 : IN std_logic ;
      window_3_1 : IN std_logic ;
      window_3_0 : IN std_logic ;
      window_2_15 : IN std_logic ;
      window_2_14 : IN std_logic ;
      window_2_13 : IN std_logic ;
      window_2_12 : IN std_logic ;
      window_2_11 : IN std_logic ;
      window_2_10 : IN std_logic ;
      window_2_9 : IN std_logic ;
      window_2_8 : IN std_logic ;
      window_2_7 : IN std_logic ;
      window_2_6 : IN std_logic ;
      window_2_5 : IN std_logic ;
      window_2_4 : IN std_logic ;
      window_2_3 : IN std_logic ;
      window_2_2 : IN std_logic ;
      window_2_1 : IN std_logic ;
      window_2_0 : IN std_logic ;
      window_1_15 : IN std_logic ;
      window_1_14 : IN std_logic ;
      window_1_13 : IN std_logic ;
      window_1_12 : IN std_logic ;
      window_1_11 : IN std_logic ;
      window_1_10 : IN std_logic ;
      window_1_9 : IN std_logic ;
      window_1_8 : IN std_logic ;
      window_1_7 : IN std_logic ;
      window_1_6 : IN std_logic ;
      window_1_5 : IN std_logic ;
      window_1_4 : IN std_logic ;
      window_1_3 : IN std_logic ;
      window_1_2 : IN std_logic ;
      window_1_1 : IN std_logic ;
      window_1_0 : IN std_logic ;
      window_0_15 : IN std_logic ;
      window_0_14 : IN std_logic ;
      window_0_13 : IN std_logic ;
      window_0_12 : IN std_logic ;
      window_0_11 : IN std_logic ;
      window_0_10 : IN std_logic ;
      window_0_9 : IN std_logic ;
      window_0_8 : IN std_logic ;
      window_0_7 : IN std_logic ;
      window_0_6 : IN std_logic ;
      window_0_5 : IN std_logic ;
      window_0_4 : IN std_logic ;
      window_0_3 : IN std_logic ;
      window_0_2 : IN std_logic ;
      window_0_1 : IN std_logic ;
      window_0_0 : IN std_logic ;
      outputs_24_15 : INOUT std_logic ;
      outputs_24_14 : INOUT std_logic ;
      outputs_24_13 : INOUT std_logic ;
      outputs_24_12 : INOUT std_logic ;
      outputs_24_11 : INOUT std_logic ;
      outputs_24_10 : INOUT std_logic ;
      outputs_24_9 : INOUT std_logic ;
      outputs_24_8 : INOUT std_logic ;
      outputs_24_7 : INOUT std_logic ;
      outputs_24_6 : INOUT std_logic ;
      outputs_24_5 : INOUT std_logic ;
      outputs_24_4 : INOUT std_logic ;
      outputs_24_3 : INOUT std_logic ;
      outputs_24_2 : INOUT std_logic ;
      outputs_24_1 : INOUT std_logic ;
      outputs_24_0 : INOUT std_logic ;
      outputs_23_15 : INOUT std_logic ;
      outputs_23_14 : INOUT std_logic ;
      outputs_23_13 : INOUT std_logic ;
      outputs_23_12 : INOUT std_logic ;
      outputs_23_11 : INOUT std_logic ;
      outputs_23_10 : INOUT std_logic ;
      outputs_23_9 : INOUT std_logic ;
      outputs_23_8 : INOUT std_logic ;
      outputs_23_7 : INOUT std_logic ;
      outputs_23_6 : INOUT std_logic ;
      outputs_23_5 : INOUT std_logic ;
      outputs_23_4 : INOUT std_logic ;
      outputs_23_3 : INOUT std_logic ;
      outputs_23_2 : INOUT std_logic ;
      outputs_23_1 : INOUT std_logic ;
      outputs_23_0 : INOUT std_logic ;
      outputs_22_15 : INOUT std_logic ;
      outputs_22_14 : INOUT std_logic ;
      outputs_22_13 : INOUT std_logic ;
      outputs_22_12 : INOUT std_logic ;
      outputs_22_11 : INOUT std_logic ;
      outputs_22_10 : INOUT std_logic ;
      outputs_22_9 : INOUT std_logic ;
      outputs_22_8 : INOUT std_logic ;
      outputs_22_7 : INOUT std_logic ;
      outputs_22_6 : INOUT std_logic ;
      outputs_22_5 : INOUT std_logic ;
      outputs_22_4 : INOUT std_logic ;
      outputs_22_3 : INOUT std_logic ;
      outputs_22_2 : INOUT std_logic ;
      outputs_22_1 : INOUT std_logic ;
      outputs_22_0 : INOUT std_logic ;
      outputs_21_15 : INOUT std_logic ;
      outputs_21_14 : INOUT std_logic ;
      outputs_21_13 : INOUT std_logic ;
      outputs_21_12 : INOUT std_logic ;
      outputs_21_11 : INOUT std_logic ;
      outputs_21_10 : INOUT std_logic ;
      outputs_21_9 : INOUT std_logic ;
      outputs_21_8 : INOUT std_logic ;
      outputs_21_7 : INOUT std_logic ;
      outputs_21_6 : INOUT std_logic ;
      outputs_21_5 : INOUT std_logic ;
      outputs_21_4 : INOUT std_logic ;
      outputs_21_3 : INOUT std_logic ;
      outputs_21_2 : INOUT std_logic ;
      outputs_21_1 : INOUT std_logic ;
      outputs_21_0 : INOUT std_logic ;
      outputs_20_15 : INOUT std_logic ;
      outputs_20_14 : INOUT std_logic ;
      outputs_20_13 : INOUT std_logic ;
      outputs_20_12 : INOUT std_logic ;
      outputs_20_11 : INOUT std_logic ;
      outputs_20_10 : INOUT std_logic ;
      outputs_20_9 : INOUT std_logic ;
      outputs_20_8 : INOUT std_logic ;
      outputs_20_7 : INOUT std_logic ;
      outputs_20_6 : INOUT std_logic ;
      outputs_20_5 : INOUT std_logic ;
      outputs_20_4 : INOUT std_logic ;
      outputs_20_3 : INOUT std_logic ;
      outputs_20_2 : INOUT std_logic ;
      outputs_20_1 : INOUT std_logic ;
      outputs_20_0 : INOUT std_logic ;
      outputs_19_15 : INOUT std_logic ;
      outputs_19_14 : INOUT std_logic ;
      outputs_19_13 : INOUT std_logic ;
      outputs_19_12 : INOUT std_logic ;
      outputs_19_11 : INOUT std_logic ;
      outputs_19_10 : INOUT std_logic ;
      outputs_19_9 : INOUT std_logic ;
      outputs_19_8 : INOUT std_logic ;
      outputs_19_7 : INOUT std_logic ;
      outputs_19_6 : INOUT std_logic ;
      outputs_19_5 : INOUT std_logic ;
      outputs_19_4 : INOUT std_logic ;
      outputs_19_3 : INOUT std_logic ;
      outputs_19_2 : INOUT std_logic ;
      outputs_19_1 : INOUT std_logic ;
      outputs_19_0 : INOUT std_logic ;
      outputs_18_15 : INOUT std_logic ;
      outputs_18_14 : INOUT std_logic ;
      outputs_18_13 : INOUT std_logic ;
      outputs_18_12 : INOUT std_logic ;
      outputs_18_11 : INOUT std_logic ;
      outputs_18_10 : INOUT std_logic ;
      outputs_18_9 : INOUT std_logic ;
      outputs_18_8 : INOUT std_logic ;
      outputs_18_7 : INOUT std_logic ;
      outputs_18_6 : INOUT std_logic ;
      outputs_18_5 : INOUT std_logic ;
      outputs_18_4 : INOUT std_logic ;
      outputs_18_3 : INOUT std_logic ;
      outputs_18_2 : INOUT std_logic ;
      outputs_18_1 : INOUT std_logic ;
      outputs_18_0 : INOUT std_logic ;
      outputs_17_15 : INOUT std_logic ;
      outputs_17_14 : INOUT std_logic ;
      outputs_17_13 : INOUT std_logic ;
      outputs_17_12 : INOUT std_logic ;
      outputs_17_11 : INOUT std_logic ;
      outputs_17_10 : INOUT std_logic ;
      outputs_17_9 : INOUT std_logic ;
      outputs_17_8 : INOUT std_logic ;
      outputs_17_7 : INOUT std_logic ;
      outputs_17_6 : INOUT std_logic ;
      outputs_17_5 : INOUT std_logic ;
      outputs_17_4 : INOUT std_logic ;
      outputs_17_3 : INOUT std_logic ;
      outputs_17_2 : INOUT std_logic ;
      outputs_17_1 : INOUT std_logic ;
      outputs_17_0 : INOUT std_logic ;
      outputs_16_15 : INOUT std_logic ;
      outputs_16_14 : INOUT std_logic ;
      outputs_16_13 : INOUT std_logic ;
      outputs_16_12 : INOUT std_logic ;
      outputs_16_11 : INOUT std_logic ;
      outputs_16_10 : INOUT std_logic ;
      outputs_16_9 : INOUT std_logic ;
      outputs_16_8 : INOUT std_logic ;
      outputs_16_7 : INOUT std_logic ;
      outputs_16_6 : INOUT std_logic ;
      outputs_16_5 : INOUT std_logic ;
      outputs_16_4 : INOUT std_logic ;
      outputs_16_3 : INOUT std_logic ;
      outputs_16_2 : INOUT std_logic ;
      outputs_16_1 : INOUT std_logic ;
      outputs_16_0 : INOUT std_logic ;
      outputs_15_15 : INOUT std_logic ;
      outputs_15_14 : INOUT std_logic ;
      outputs_15_13 : INOUT std_logic ;
      outputs_15_12 : INOUT std_logic ;
      outputs_15_11 : INOUT std_logic ;
      outputs_15_10 : INOUT std_logic ;
      outputs_15_9 : INOUT std_logic ;
      outputs_15_8 : INOUT std_logic ;
      outputs_15_7 : INOUT std_logic ;
      outputs_15_6 : INOUT std_logic ;
      outputs_15_5 : INOUT std_logic ;
      outputs_15_4 : INOUT std_logic ;
      outputs_15_3 : INOUT std_logic ;
      outputs_15_2 : INOUT std_logic ;
      outputs_15_1 : INOUT std_logic ;
      outputs_15_0 : INOUT std_logic ;
      outputs_14_15 : INOUT std_logic ;
      outputs_14_14 : INOUT std_logic ;
      outputs_14_13 : INOUT std_logic ;
      outputs_14_12 : INOUT std_logic ;
      outputs_14_11 : INOUT std_logic ;
      outputs_14_10 : INOUT std_logic ;
      outputs_14_9 : INOUT std_logic ;
      outputs_14_8 : INOUT std_logic ;
      outputs_14_7 : INOUT std_logic ;
      outputs_14_6 : INOUT std_logic ;
      outputs_14_5 : INOUT std_logic ;
      outputs_14_4 : INOUT std_logic ;
      outputs_14_3 : INOUT std_logic ;
      outputs_14_2 : INOUT std_logic ;
      outputs_14_1 : INOUT std_logic ;
      outputs_14_0 : INOUT std_logic ;
      outputs_13_15 : INOUT std_logic ;
      outputs_13_14 : INOUT std_logic ;
      outputs_13_13 : INOUT std_logic ;
      outputs_13_12 : INOUT std_logic ;
      outputs_13_11 : INOUT std_logic ;
      outputs_13_10 : INOUT std_logic ;
      outputs_13_9 : INOUT std_logic ;
      outputs_13_8 : INOUT std_logic ;
      outputs_13_7 : INOUT std_logic ;
      outputs_13_6 : INOUT std_logic ;
      outputs_13_5 : INOUT std_logic ;
      outputs_13_4 : INOUT std_logic ;
      outputs_13_3 : INOUT std_logic ;
      outputs_13_2 : INOUT std_logic ;
      outputs_13_1 : INOUT std_logic ;
      outputs_13_0 : INOUT std_logic ;
      outputs_12_15 : INOUT std_logic ;
      outputs_12_14 : INOUT std_logic ;
      outputs_12_13 : INOUT std_logic ;
      outputs_12_12 : INOUT std_logic ;
      outputs_12_11 : INOUT std_logic ;
      outputs_12_10 : INOUT std_logic ;
      outputs_12_9 : INOUT std_logic ;
      outputs_12_8 : INOUT std_logic ;
      outputs_12_7 : INOUT std_logic ;
      outputs_12_6 : INOUT std_logic ;
      outputs_12_5 : INOUT std_logic ;
      outputs_12_4 : INOUT std_logic ;
      outputs_12_3 : INOUT std_logic ;
      outputs_12_2 : INOUT std_logic ;
      outputs_12_1 : INOUT std_logic ;
      outputs_12_0 : INOUT std_logic ;
      outputs_11_15 : INOUT std_logic ;
      outputs_11_14 : INOUT std_logic ;
      outputs_11_13 : INOUT std_logic ;
      outputs_11_12 : INOUT std_logic ;
      outputs_11_11 : INOUT std_logic ;
      outputs_11_10 : INOUT std_logic ;
      outputs_11_9 : INOUT std_logic ;
      outputs_11_8 : INOUT std_logic ;
      outputs_11_7 : INOUT std_logic ;
      outputs_11_6 : INOUT std_logic ;
      outputs_11_5 : INOUT std_logic ;
      outputs_11_4 : INOUT std_logic ;
      outputs_11_3 : INOUT std_logic ;
      outputs_11_2 : INOUT std_logic ;
      outputs_11_1 : INOUT std_logic ;
      outputs_11_0 : INOUT std_logic ;
      outputs_10_15 : INOUT std_logic ;
      outputs_10_14 : INOUT std_logic ;
      outputs_10_13 : INOUT std_logic ;
      outputs_10_12 : INOUT std_logic ;
      outputs_10_11 : INOUT std_logic ;
      outputs_10_10 : INOUT std_logic ;
      outputs_10_9 : INOUT std_logic ;
      outputs_10_8 : INOUT std_logic ;
      outputs_10_7 : INOUT std_logic ;
      outputs_10_6 : INOUT std_logic ;
      outputs_10_5 : INOUT std_logic ;
      outputs_10_4 : INOUT std_logic ;
      outputs_10_3 : INOUT std_logic ;
      outputs_10_2 : INOUT std_logic ;
      outputs_10_1 : INOUT std_logic ;
      outputs_10_0 : INOUT std_logic ;
      outputs_9_15 : INOUT std_logic ;
      outputs_9_14 : INOUT std_logic ;
      outputs_9_13 : INOUT std_logic ;
      outputs_9_12 : INOUT std_logic ;
      outputs_9_11 : INOUT std_logic ;
      outputs_9_10 : INOUT std_logic ;
      outputs_9_9 : INOUT std_logic ;
      outputs_9_8 : INOUT std_logic ;
      outputs_9_7 : INOUT std_logic ;
      outputs_9_6 : INOUT std_logic ;
      outputs_9_5 : INOUT std_logic ;
      outputs_9_4 : INOUT std_logic ;
      outputs_9_3 : INOUT std_logic ;
      outputs_9_2 : INOUT std_logic ;
      outputs_9_1 : INOUT std_logic ;
      outputs_9_0 : INOUT std_logic ;
      outputs_8_15 : INOUT std_logic ;
      outputs_8_14 : INOUT std_logic ;
      outputs_8_13 : INOUT std_logic ;
      outputs_8_12 : INOUT std_logic ;
      outputs_8_11 : INOUT std_logic ;
      outputs_8_10 : INOUT std_logic ;
      outputs_8_9 : INOUT std_logic ;
      outputs_8_8 : INOUT std_logic ;
      outputs_8_7 : INOUT std_logic ;
      outputs_8_6 : INOUT std_logic ;
      outputs_8_5 : INOUT std_logic ;
      outputs_8_4 : INOUT std_logic ;
      outputs_8_3 : INOUT std_logic ;
      outputs_8_2 : INOUT std_logic ;
      outputs_8_1 : INOUT std_logic ;
      outputs_8_0 : INOUT std_logic ;
      outputs_7_15 : INOUT std_logic ;
      outputs_7_14 : INOUT std_logic ;
      outputs_7_13 : INOUT std_logic ;
      outputs_7_12 : INOUT std_logic ;
      outputs_7_11 : INOUT std_logic ;
      outputs_7_10 : INOUT std_logic ;
      outputs_7_9 : INOUT std_logic ;
      outputs_7_8 : INOUT std_logic ;
      outputs_7_7 : INOUT std_logic ;
      outputs_7_6 : INOUT std_logic ;
      outputs_7_5 : INOUT std_logic ;
      outputs_7_4 : INOUT std_logic ;
      outputs_7_3 : INOUT std_logic ;
      outputs_7_2 : INOUT std_logic ;
      outputs_7_1 : INOUT std_logic ;
      outputs_7_0 : INOUT std_logic ;
      outputs_6_15 : INOUT std_logic ;
      outputs_6_14 : INOUT std_logic ;
      outputs_6_13 : INOUT std_logic ;
      outputs_6_12 : INOUT std_logic ;
      outputs_6_11 : INOUT std_logic ;
      outputs_6_10 : INOUT std_logic ;
      outputs_6_9 : INOUT std_logic ;
      outputs_6_8 : INOUT std_logic ;
      outputs_6_7 : INOUT std_logic ;
      outputs_6_6 : INOUT std_logic ;
      outputs_6_5 : INOUT std_logic ;
      outputs_6_4 : INOUT std_logic ;
      outputs_6_3 : INOUT std_logic ;
      outputs_6_2 : INOUT std_logic ;
      outputs_6_1 : INOUT std_logic ;
      outputs_6_0 : INOUT std_logic ;
      outputs_5_15 : INOUT std_logic ;
      outputs_5_14 : INOUT std_logic ;
      outputs_5_13 : INOUT std_logic ;
      outputs_5_12 : INOUT std_logic ;
      outputs_5_11 : INOUT std_logic ;
      outputs_5_10 : INOUT std_logic ;
      outputs_5_9 : INOUT std_logic ;
      outputs_5_8 : INOUT std_logic ;
      outputs_5_7 : INOUT std_logic ;
      outputs_5_6 : INOUT std_logic ;
      outputs_5_5 : INOUT std_logic ;
      outputs_5_4 : INOUT std_logic ;
      outputs_5_3 : INOUT std_logic ;
      outputs_5_2 : INOUT std_logic ;
      outputs_5_1 : INOUT std_logic ;
      outputs_5_0 : INOUT std_logic ;
      outputs_4_15 : INOUT std_logic ;
      outputs_4_14 : INOUT std_logic ;
      outputs_4_13 : INOUT std_logic ;
      outputs_4_12 : INOUT std_logic ;
      outputs_4_11 : INOUT std_logic ;
      outputs_4_10 : INOUT std_logic ;
      outputs_4_9 : INOUT std_logic ;
      outputs_4_8 : INOUT std_logic ;
      outputs_4_7 : INOUT std_logic ;
      outputs_4_6 : INOUT std_logic ;
      outputs_4_5 : INOUT std_logic ;
      outputs_4_4 : INOUT std_logic ;
      outputs_4_3 : INOUT std_logic ;
      outputs_4_2 : INOUT std_logic ;
      outputs_4_1 : INOUT std_logic ;
      outputs_4_0 : INOUT std_logic ;
      outputs_3_15 : INOUT std_logic ;
      outputs_3_14 : INOUT std_logic ;
      outputs_3_13 : INOUT std_logic ;
      outputs_3_12 : INOUT std_logic ;
      outputs_3_11 : INOUT std_logic ;
      outputs_3_10 : INOUT std_logic ;
      outputs_3_9 : INOUT std_logic ;
      outputs_3_8 : INOUT std_logic ;
      outputs_3_7 : INOUT std_logic ;
      outputs_3_6 : INOUT std_logic ;
      outputs_3_5 : INOUT std_logic ;
      outputs_3_4 : INOUT std_logic ;
      outputs_3_3 : INOUT std_logic ;
      outputs_3_2 : INOUT std_logic ;
      outputs_3_1 : INOUT std_logic ;
      outputs_3_0 : INOUT std_logic ;
      outputs_2_15 : INOUT std_logic ;
      outputs_2_14 : INOUT std_logic ;
      outputs_2_13 : INOUT std_logic ;
      outputs_2_12 : INOUT std_logic ;
      outputs_2_11 : INOUT std_logic ;
      outputs_2_10 : INOUT std_logic ;
      outputs_2_9 : INOUT std_logic ;
      outputs_2_8 : INOUT std_logic ;
      outputs_2_7 : INOUT std_logic ;
      outputs_2_6 : INOUT std_logic ;
      outputs_2_5 : INOUT std_logic ;
      outputs_2_4 : INOUT std_logic ;
      outputs_2_3 : INOUT std_logic ;
      outputs_2_2 : INOUT std_logic ;
      outputs_2_1 : INOUT std_logic ;
      outputs_2_0 : INOUT std_logic ;
      outputs_1_15 : INOUT std_logic ;
      outputs_1_14 : INOUT std_logic ;
      outputs_1_13 : INOUT std_logic ;
      outputs_1_12 : INOUT std_logic ;
      outputs_1_11 : INOUT std_logic ;
      outputs_1_10 : INOUT std_logic ;
      outputs_1_9 : INOUT std_logic ;
      outputs_1_8 : INOUT std_logic ;
      outputs_1_7 : INOUT std_logic ;
      outputs_1_6 : INOUT std_logic ;
      outputs_1_5 : INOUT std_logic ;
      outputs_1_4 : INOUT std_logic ;
      outputs_1_3 : INOUT std_logic ;
      outputs_1_2 : INOUT std_logic ;
      outputs_1_1 : INOUT std_logic ;
      outputs_1_0 : INOUT std_logic ;
      outputs_0_15 : INOUT std_logic ;
      outputs_0_14 : INOUT std_logic ;
      outputs_0_13 : INOUT std_logic ;
      outputs_0_12 : INOUT std_logic ;
      outputs_0_11 : INOUT std_logic ;
      outputs_0_10 : INOUT std_logic ;
      outputs_0_9 : INOUT std_logic ;
      outputs_0_8 : INOUT std_logic ;
      outputs_0_7 : INOUT std_logic ;
      outputs_0_6 : INOUT std_logic ;
      outputs_0_5 : INOUT std_logic ;
      outputs_0_4 : INOUT std_logic ;
      outputs_0_3 : INOUT std_logic ;
      outputs_0_2 : INOUT std_logic ;
      outputs_0_1 : INOUT std_logic ;
      outputs_0_0 : INOUT std_logic ;
      clk : IN std_logic ;
      start : IN std_logic ;
      rst : IN std_logic ;
      done : INOUT std_logic ;
      working : INOUT std_logic) ;
end CNNMuls ;

architecture CNNMulsArch of CNNMuls is
   component Reg_33
      port (
         D : IN std_logic_vector (32 DOWNTO 0) ;
         en : IN std_logic ;
         clk : IN std_logic ;
         rst : IN std_logic ;
         Q : OUT std_logic_vector (32 DOWNTO 0)) ;
   end component ;
   component BinaryMux_33
      port (
         a : IN std_logic_vector (32 DOWNTO 0) ;
         b : IN std_logic_vector (32 DOWNTO 0) ;
         sel : IN std_logic ;
         f : OUT std_logic_vector (32 DOWNTO 0)) ;
   end component ;
   component NBitAdder_24
      port (
         a : IN std_logic_vector (23 DOWNTO 0) ;
         b : IN std_logic_vector (23 DOWNTO 0) ;
         carryIn : IN std_logic ;
         sum : OUT std_logic_vector (23 DOWNTO 0) ;
         carryOut : OUT std_logic) ;
   end component ;
   signal gen_24_cmp_pBs_30, gen_24_cmp_pBs_29, gen_24_cmp_pBs_28, 
      gen_24_cmp_pBs_27, gen_24_cmp_pBs_26, gen_24_cmp_pBs_25, 
      gen_24_cmp_pBs_24, gen_24_cmp_pBs_23, gen_24_cmp_pMux_30, 
      gen_24_cmp_pMux_29, gen_24_cmp_pMux_28, gen_24_cmp_pMux_27, 
      gen_24_cmp_pMux_26, gen_24_cmp_pMux_25, gen_24_cmp_pMux_24, 
      gen_24_cmp_pMux_23, gen_24_cmp_pMux_22, gen_24_cmp_pMux_21, 
      gen_24_cmp_pMux_20, gen_24_cmp_pMux_19, gen_24_cmp_pMux_18, 
      gen_24_cmp_pMux_17, gen_24_cmp_pMux_16, gen_24_cmp_pMux_15, 
      gen_24_cmp_pMux_14, gen_24_cmp_pMux_13, gen_24_cmp_pMux_12, 
      gen_24_cmp_pMux_11, gen_24_cmp_pMux_10, gen_24_cmp_pMux_9, 
      gen_24_cmp_pMux_8, gen_24_cmp_pMux_7, gen_24_cmp_pMux_6, 
      gen_24_cmp_pMux_5, gen_24_cmp_pMux_4, gen_24_cmp_pMux_3, 
      gen_24_cmp_pMux_2, gen_24_cmp_pMux_1, gen_24_cmp_pMux_0, 
      gen_24_cmp_pReg_30, gen_24_cmp_pReg_29, gen_24_cmp_pReg_28, 
      gen_24_cmp_pReg_27, gen_24_cmp_pReg_26, gen_24_cmp_pReg_25, 
      gen_24_cmp_pReg_24, gen_24_cmp_pReg_23, gen_24_cmp_pReg_22, 
      gen_24_cmp_pReg_21, gen_24_cmp_pReg_20, gen_24_cmp_pReg_19, 
      gen_24_cmp_pReg_18, gen_24_cmp_pReg_17, gen_24_cmp_pReg_16, 
      gen_24_cmp_pReg_15, gen_24_cmp_pReg_14, gen_24_cmp_pReg_13, 
      gen_24_cmp_pReg_12, gen_24_cmp_pReg_11, gen_24_cmp_pReg_10, 
      gen_24_cmp_pReg_9, gen_24_cmp_pReg_8, gen_24_cmp_pReg_7, 
      gen_24_cmp_pReg_6, gen_24_cmp_pReg_5, gen_24_cmp_pReg_4, 
      gen_24_cmp_pReg_3, gen_24_cmp_pReg_2, gen_24_cmp_pReg_1, 
      gen_24_cmp_pReg_0, gen_24_cmp_BSCmp_op2_0, gen_24_cmp_BSCmp_carryIn, 
      gen_23_cmp_pBs_30, gen_23_cmp_pBs_29, gen_23_cmp_pBs_28, 
      gen_23_cmp_pBs_27, gen_23_cmp_pBs_26, gen_23_cmp_pBs_25, 
      gen_23_cmp_pBs_24, gen_23_cmp_pBs_23, gen_23_cmp_pMux_30, 
      gen_23_cmp_pMux_29, gen_23_cmp_pMux_28, gen_23_cmp_pMux_27, 
      gen_23_cmp_pMux_26, gen_23_cmp_pMux_25, gen_23_cmp_pMux_24, 
      gen_23_cmp_pMux_23, gen_23_cmp_pMux_22, gen_23_cmp_pMux_21, 
      gen_23_cmp_pMux_20, gen_23_cmp_pMux_19, gen_23_cmp_pMux_18, 
      gen_23_cmp_pMux_17, gen_23_cmp_pMux_16, gen_23_cmp_pMux_15, 
      gen_23_cmp_pMux_14, gen_23_cmp_pMux_13, gen_23_cmp_pMux_12, 
      gen_23_cmp_pMux_11, gen_23_cmp_pMux_10, gen_23_cmp_pMux_9, 
      gen_23_cmp_pMux_8, gen_23_cmp_pMux_7, gen_23_cmp_pMux_6, 
      gen_23_cmp_pMux_5, gen_23_cmp_pMux_4, gen_23_cmp_pMux_3, 
      gen_23_cmp_pMux_2, gen_23_cmp_pMux_1, gen_23_cmp_pMux_0, 
      gen_23_cmp_pReg_30, gen_23_cmp_pReg_29, gen_23_cmp_pReg_28, 
      gen_23_cmp_pReg_27, gen_23_cmp_pReg_26, gen_23_cmp_pReg_25, 
      gen_23_cmp_pReg_24, gen_23_cmp_pReg_23, gen_23_cmp_pReg_22, 
      gen_23_cmp_pReg_21, gen_23_cmp_pReg_20, gen_23_cmp_pReg_19, 
      gen_23_cmp_pReg_18, gen_23_cmp_pReg_17, gen_23_cmp_pReg_16, 
      gen_23_cmp_pReg_15, gen_23_cmp_pReg_14, gen_23_cmp_pReg_13, 
      gen_23_cmp_pReg_12, gen_23_cmp_pReg_11, gen_23_cmp_pReg_10, 
      gen_23_cmp_pReg_9, gen_23_cmp_pReg_8, gen_23_cmp_pReg_7, 
      gen_23_cmp_pReg_6, gen_23_cmp_pReg_5, gen_23_cmp_pReg_4, 
      gen_23_cmp_pReg_3, gen_23_cmp_pReg_2, gen_23_cmp_pReg_1, 
      gen_23_cmp_pReg_0, gen_23_cmp_BSCmp_op2_0, gen_23_cmp_BSCmp_carryIn, 
      gen_22_cmp_pBs_30, gen_22_cmp_pBs_29, gen_22_cmp_pBs_28, 
      gen_22_cmp_pBs_27, gen_22_cmp_pBs_26, gen_22_cmp_pBs_25, 
      gen_22_cmp_pBs_24, gen_22_cmp_pBs_23, gen_22_cmp_pMux_30, 
      gen_22_cmp_pMux_29, gen_22_cmp_pMux_28, gen_22_cmp_pMux_27, 
      gen_22_cmp_pMux_26, gen_22_cmp_pMux_25, gen_22_cmp_pMux_24, 
      gen_22_cmp_pMux_23, gen_22_cmp_pMux_22, gen_22_cmp_pMux_21, 
      gen_22_cmp_pMux_20, gen_22_cmp_pMux_19, gen_22_cmp_pMux_18, 
      gen_22_cmp_pMux_17, gen_22_cmp_pMux_16, gen_22_cmp_pMux_15, 
      gen_22_cmp_pMux_14, gen_22_cmp_pMux_13, gen_22_cmp_pMux_12, 
      gen_22_cmp_pMux_11, gen_22_cmp_pMux_10, gen_22_cmp_pMux_9, 
      gen_22_cmp_pMux_8, gen_22_cmp_pMux_7, gen_22_cmp_pMux_6, 
      gen_22_cmp_pMux_5, gen_22_cmp_pMux_4, gen_22_cmp_pMux_3, 
      gen_22_cmp_pMux_2, gen_22_cmp_pMux_1, gen_22_cmp_pMux_0, 
      gen_22_cmp_pReg_30, gen_22_cmp_pReg_29, gen_22_cmp_pReg_28, 
      gen_22_cmp_pReg_27, gen_22_cmp_pReg_26, gen_22_cmp_pReg_25, 
      gen_22_cmp_pReg_24, gen_22_cmp_pReg_23, gen_22_cmp_pReg_22, 
      gen_22_cmp_pReg_21, gen_22_cmp_pReg_20, gen_22_cmp_pReg_19, 
      gen_22_cmp_pReg_18, gen_22_cmp_pReg_17, gen_22_cmp_pReg_16, 
      gen_22_cmp_pReg_15, gen_22_cmp_pReg_14, gen_22_cmp_pReg_13, 
      gen_22_cmp_pReg_12, gen_22_cmp_pReg_11, gen_22_cmp_pReg_10, 
      gen_22_cmp_pReg_9, gen_22_cmp_pReg_8, gen_22_cmp_pReg_7, 
      gen_22_cmp_pReg_6, gen_22_cmp_pReg_5, gen_22_cmp_pReg_4, 
      gen_22_cmp_pReg_3, gen_22_cmp_pReg_2, gen_22_cmp_pReg_1, 
      gen_22_cmp_pReg_0, gen_22_cmp_BSCmp_op2_0, gen_22_cmp_BSCmp_carryIn, 
      gen_21_cmp_pBs_30, gen_21_cmp_pBs_29, gen_21_cmp_pBs_28, 
      gen_21_cmp_pBs_27, gen_21_cmp_pBs_26, gen_21_cmp_pBs_25, 
      gen_21_cmp_pBs_24, gen_21_cmp_pBs_23, gen_21_cmp_pMux_30, 
      gen_21_cmp_pMux_29, gen_21_cmp_pMux_28, gen_21_cmp_pMux_27, 
      gen_21_cmp_pMux_26, gen_21_cmp_pMux_25, gen_21_cmp_pMux_24, 
      gen_21_cmp_pMux_23, gen_21_cmp_pMux_22, gen_21_cmp_pMux_21, 
      gen_21_cmp_pMux_20, gen_21_cmp_pMux_19, gen_21_cmp_pMux_18, 
      gen_21_cmp_pMux_17, gen_21_cmp_pMux_16, gen_21_cmp_pMux_15, 
      gen_21_cmp_pMux_14, gen_21_cmp_pMux_13, gen_21_cmp_pMux_12, 
      gen_21_cmp_pMux_11, gen_21_cmp_pMux_10, gen_21_cmp_pMux_9, 
      gen_21_cmp_pMux_8, gen_21_cmp_pMux_7, gen_21_cmp_pMux_6, 
      gen_21_cmp_pMux_5, gen_21_cmp_pMux_4, gen_21_cmp_pMux_3, 
      gen_21_cmp_pMux_2, gen_21_cmp_pMux_1, gen_21_cmp_pMux_0, 
      gen_21_cmp_pReg_30, gen_21_cmp_pReg_29, gen_21_cmp_pReg_28, 
      gen_21_cmp_pReg_27, gen_21_cmp_pReg_26, gen_21_cmp_pReg_25, 
      gen_21_cmp_pReg_24, gen_21_cmp_pReg_23, gen_21_cmp_pReg_22, 
      gen_21_cmp_pReg_21, gen_21_cmp_pReg_20, gen_21_cmp_pReg_19, 
      gen_21_cmp_pReg_18, gen_21_cmp_pReg_17, gen_21_cmp_pReg_16, 
      gen_21_cmp_pReg_15, gen_21_cmp_pReg_14, gen_21_cmp_pReg_13, 
      gen_21_cmp_pReg_12, gen_21_cmp_pReg_11, gen_21_cmp_pReg_10, 
      gen_21_cmp_pReg_9, gen_21_cmp_pReg_8, gen_21_cmp_pReg_7, 
      gen_21_cmp_pReg_6, gen_21_cmp_pReg_5, gen_21_cmp_pReg_4, 
      gen_21_cmp_pReg_3, gen_21_cmp_pReg_2, gen_21_cmp_pReg_1, 
      gen_21_cmp_pReg_0, gen_21_cmp_BSCmp_op2_0, gen_21_cmp_BSCmp_carryIn, 
      gen_20_cmp_pBs_30, gen_20_cmp_pBs_29, gen_20_cmp_pBs_28, 
      gen_20_cmp_pBs_27, gen_20_cmp_pBs_26, gen_20_cmp_pBs_25, 
      gen_20_cmp_pBs_24, gen_20_cmp_pBs_23, gen_20_cmp_pMux_30, 
      gen_20_cmp_pMux_29, gen_20_cmp_pMux_28, gen_20_cmp_pMux_27, 
      gen_20_cmp_pMux_26, gen_20_cmp_pMux_25, gen_20_cmp_pMux_24, 
      gen_20_cmp_pMux_23, gen_20_cmp_pMux_22, gen_20_cmp_pMux_21, 
      gen_20_cmp_pMux_20, gen_20_cmp_pMux_19, gen_20_cmp_pMux_18, 
      gen_20_cmp_pMux_17, gen_20_cmp_pMux_16, gen_20_cmp_pMux_15, 
      gen_20_cmp_pMux_14, gen_20_cmp_pMux_13, gen_20_cmp_pMux_12, 
      gen_20_cmp_pMux_11, gen_20_cmp_pMux_10, gen_20_cmp_pMux_9, 
      gen_20_cmp_pMux_8, gen_20_cmp_pMux_7, gen_20_cmp_pMux_6, 
      gen_20_cmp_pMux_5, gen_20_cmp_pMux_4, gen_20_cmp_pMux_3, 
      gen_20_cmp_pMux_2, gen_20_cmp_pMux_1, gen_20_cmp_pMux_0, 
      gen_20_cmp_pReg_30, gen_20_cmp_pReg_29, gen_20_cmp_pReg_28, 
      gen_20_cmp_pReg_27, gen_20_cmp_pReg_26, gen_20_cmp_pReg_25, 
      gen_20_cmp_pReg_24, gen_20_cmp_pReg_23, gen_20_cmp_pReg_22, 
      gen_20_cmp_pReg_21, gen_20_cmp_pReg_20, gen_20_cmp_pReg_19, 
      gen_20_cmp_pReg_18, gen_20_cmp_pReg_17, gen_20_cmp_pReg_16, 
      gen_20_cmp_pReg_15, gen_20_cmp_pReg_14, gen_20_cmp_pReg_13, 
      gen_20_cmp_pReg_12, gen_20_cmp_pReg_11, gen_20_cmp_pReg_10, 
      gen_20_cmp_pReg_9, gen_20_cmp_pReg_8, gen_20_cmp_pReg_7, 
      gen_20_cmp_pReg_6, gen_20_cmp_pReg_5, gen_20_cmp_pReg_4, 
      gen_20_cmp_pReg_3, gen_20_cmp_pReg_2, gen_20_cmp_pReg_1, 
      gen_20_cmp_pReg_0, gen_20_cmp_BSCmp_op2_0, gen_20_cmp_BSCmp_carryIn, 
      gen_19_cmp_pBs_30, gen_19_cmp_pBs_29, gen_19_cmp_pBs_28, 
      gen_19_cmp_pBs_27, gen_19_cmp_pBs_26, gen_19_cmp_pBs_25, 
      gen_19_cmp_pBs_24, gen_19_cmp_pBs_23, gen_19_cmp_pMux_30, 
      gen_19_cmp_pMux_29, gen_19_cmp_pMux_28, gen_19_cmp_pMux_27, 
      gen_19_cmp_pMux_26, gen_19_cmp_pMux_25, gen_19_cmp_pMux_24, 
      gen_19_cmp_pMux_23, gen_19_cmp_pMux_22, gen_19_cmp_pMux_21, 
      gen_19_cmp_pMux_20, gen_19_cmp_pMux_19, gen_19_cmp_pMux_18, 
      gen_19_cmp_pMux_17, gen_19_cmp_pMux_16, gen_19_cmp_pMux_15, 
      gen_19_cmp_pMux_14, gen_19_cmp_pMux_13, gen_19_cmp_pMux_12, 
      gen_19_cmp_pMux_11, gen_19_cmp_pMux_10, gen_19_cmp_pMux_9, 
      gen_19_cmp_pMux_8, gen_19_cmp_pMux_7, gen_19_cmp_pMux_6, 
      gen_19_cmp_pMux_5, gen_19_cmp_pMux_4, gen_19_cmp_pMux_3, 
      gen_19_cmp_pMux_2, gen_19_cmp_pMux_1, gen_19_cmp_pMux_0, 
      gen_19_cmp_pReg_30, gen_19_cmp_pReg_29, gen_19_cmp_pReg_28, 
      gen_19_cmp_pReg_27, gen_19_cmp_pReg_26, gen_19_cmp_pReg_25, 
      gen_19_cmp_pReg_24, gen_19_cmp_pReg_23, gen_19_cmp_pReg_22, 
      gen_19_cmp_pReg_21, gen_19_cmp_pReg_20, gen_19_cmp_pReg_19, 
      gen_19_cmp_pReg_18, gen_19_cmp_pReg_17, gen_19_cmp_pReg_16, 
      gen_19_cmp_pReg_15, gen_19_cmp_pReg_14, gen_19_cmp_pReg_13, 
      gen_19_cmp_pReg_12, gen_19_cmp_pReg_11, gen_19_cmp_pReg_10, 
      gen_19_cmp_pReg_9, gen_19_cmp_pReg_8, gen_19_cmp_pReg_7, 
      gen_19_cmp_pReg_6, gen_19_cmp_pReg_5, gen_19_cmp_pReg_4, 
      gen_19_cmp_pReg_3, gen_19_cmp_pReg_2, gen_19_cmp_pReg_1, 
      gen_19_cmp_pReg_0, gen_19_cmp_BSCmp_op2_0, gen_19_cmp_BSCmp_carryIn, 
      gen_18_cmp_pBs_30, gen_18_cmp_pBs_29, gen_18_cmp_pBs_28, 
      gen_18_cmp_pBs_27, gen_18_cmp_pBs_26, gen_18_cmp_pBs_25, 
      gen_18_cmp_pBs_24, gen_18_cmp_pBs_23, gen_18_cmp_pMux_30, 
      gen_18_cmp_pMux_29, gen_18_cmp_pMux_28, gen_18_cmp_pMux_27, 
      gen_18_cmp_pMux_26, gen_18_cmp_pMux_25, gen_18_cmp_pMux_24, 
      gen_18_cmp_pMux_23, gen_18_cmp_pMux_22, gen_18_cmp_pMux_21, 
      gen_18_cmp_pMux_20, gen_18_cmp_pMux_19, gen_18_cmp_pMux_18, 
      gen_18_cmp_pMux_17, gen_18_cmp_pMux_16, gen_18_cmp_pMux_15, 
      gen_18_cmp_pMux_14, gen_18_cmp_pMux_13, gen_18_cmp_pMux_12, 
      gen_18_cmp_pMux_11, gen_18_cmp_pMux_10, gen_18_cmp_pMux_9, 
      gen_18_cmp_pMux_8, gen_18_cmp_pMux_7, gen_18_cmp_pMux_6, 
      gen_18_cmp_pMux_5, gen_18_cmp_pMux_4, gen_18_cmp_pMux_3, 
      gen_18_cmp_pMux_2, gen_18_cmp_pMux_1, gen_18_cmp_pMux_0, 
      gen_18_cmp_pReg_30, gen_18_cmp_pReg_29, gen_18_cmp_pReg_28, 
      gen_18_cmp_pReg_27, gen_18_cmp_pReg_26, gen_18_cmp_pReg_25, 
      gen_18_cmp_pReg_24, gen_18_cmp_pReg_23, gen_18_cmp_pReg_22, 
      gen_18_cmp_pReg_21, gen_18_cmp_pReg_20, gen_18_cmp_pReg_19, 
      gen_18_cmp_pReg_18, gen_18_cmp_pReg_17, gen_18_cmp_pReg_16, 
      gen_18_cmp_pReg_15, gen_18_cmp_pReg_14, gen_18_cmp_pReg_13, 
      gen_18_cmp_pReg_12, gen_18_cmp_pReg_11, gen_18_cmp_pReg_10, 
      gen_18_cmp_pReg_9, gen_18_cmp_pReg_8, gen_18_cmp_pReg_7, 
      gen_18_cmp_pReg_6, gen_18_cmp_pReg_5, gen_18_cmp_pReg_4, 
      gen_18_cmp_pReg_3, gen_18_cmp_pReg_2, gen_18_cmp_pReg_1, 
      gen_18_cmp_pReg_0, gen_18_cmp_BSCmp_op2_0, gen_18_cmp_BSCmp_carryIn, 
      gen_17_cmp_pBs_30, gen_17_cmp_pBs_29, gen_17_cmp_pBs_28, 
      gen_17_cmp_pBs_27, gen_17_cmp_pBs_26, gen_17_cmp_pBs_25, 
      gen_17_cmp_pBs_24, gen_17_cmp_pBs_23, gen_17_cmp_pMux_30, 
      gen_17_cmp_pMux_29, gen_17_cmp_pMux_28, gen_17_cmp_pMux_27, 
      gen_17_cmp_pMux_26, gen_17_cmp_pMux_25, gen_17_cmp_pMux_24, 
      gen_17_cmp_pMux_23, gen_17_cmp_pMux_22, gen_17_cmp_pMux_21, 
      gen_17_cmp_pMux_20, gen_17_cmp_pMux_19, gen_17_cmp_pMux_18, 
      gen_17_cmp_pMux_17, gen_17_cmp_pMux_16, gen_17_cmp_pMux_15, 
      gen_17_cmp_pMux_14, gen_17_cmp_pMux_13, gen_17_cmp_pMux_12, 
      gen_17_cmp_pMux_11, gen_17_cmp_pMux_10, gen_17_cmp_pMux_9, 
      gen_17_cmp_pMux_8, gen_17_cmp_pMux_7, gen_17_cmp_pMux_6, 
      gen_17_cmp_pMux_5, gen_17_cmp_pMux_4, gen_17_cmp_pMux_3, 
      gen_17_cmp_pMux_2, gen_17_cmp_pMux_1, gen_17_cmp_pMux_0, 
      gen_17_cmp_pReg_30, gen_17_cmp_pReg_29, gen_17_cmp_pReg_28, 
      gen_17_cmp_pReg_27, gen_17_cmp_pReg_26, gen_17_cmp_pReg_25, 
      gen_17_cmp_pReg_24, gen_17_cmp_pReg_23, gen_17_cmp_pReg_22, 
      gen_17_cmp_pReg_21, gen_17_cmp_pReg_20, gen_17_cmp_pReg_19, 
      gen_17_cmp_pReg_18, gen_17_cmp_pReg_17, gen_17_cmp_pReg_16, 
      gen_17_cmp_pReg_15, gen_17_cmp_pReg_14, gen_17_cmp_pReg_13, 
      gen_17_cmp_pReg_12, gen_17_cmp_pReg_11, gen_17_cmp_pReg_10, 
      gen_17_cmp_pReg_9, gen_17_cmp_pReg_8, gen_17_cmp_pReg_7, 
      gen_17_cmp_pReg_6, gen_17_cmp_pReg_5, gen_17_cmp_pReg_4, 
      gen_17_cmp_pReg_3, gen_17_cmp_pReg_2, gen_17_cmp_pReg_1, 
      gen_17_cmp_pReg_0, gen_17_cmp_BSCmp_op2_0, gen_17_cmp_BSCmp_carryIn, 
      gen_16_cmp_pBs_30, gen_16_cmp_pBs_29, gen_16_cmp_pBs_28, 
      gen_16_cmp_pBs_27, gen_16_cmp_pBs_26, gen_16_cmp_pBs_25, 
      gen_16_cmp_pBs_24, gen_16_cmp_pBs_23, gen_16_cmp_pMux_30, 
      gen_16_cmp_pMux_29, gen_16_cmp_pMux_28, gen_16_cmp_pMux_27, 
      gen_16_cmp_pMux_26, gen_16_cmp_pMux_25, gen_16_cmp_pMux_24, 
      gen_16_cmp_pMux_23, gen_16_cmp_pMux_22, gen_16_cmp_pMux_21, 
      gen_16_cmp_pMux_20, gen_16_cmp_pMux_19, gen_16_cmp_pMux_18, 
      gen_16_cmp_pMux_17, gen_16_cmp_pMux_16, gen_16_cmp_pMux_15, 
      gen_16_cmp_pMux_14, gen_16_cmp_pMux_13, gen_16_cmp_pMux_12, 
      gen_16_cmp_pMux_11, gen_16_cmp_pMux_10, gen_16_cmp_pMux_9, 
      gen_16_cmp_pMux_8, gen_16_cmp_pMux_7, gen_16_cmp_pMux_6, 
      gen_16_cmp_pMux_5, gen_16_cmp_pMux_4, gen_16_cmp_pMux_3, 
      gen_16_cmp_pMux_2, gen_16_cmp_pMux_1, gen_16_cmp_pMux_0, 
      gen_16_cmp_pReg_30, gen_16_cmp_pReg_29, gen_16_cmp_pReg_28, 
      gen_16_cmp_pReg_27, gen_16_cmp_pReg_26, gen_16_cmp_pReg_25, 
      gen_16_cmp_pReg_24, gen_16_cmp_pReg_23, gen_16_cmp_pReg_22, 
      gen_16_cmp_pReg_21, gen_16_cmp_pReg_20, gen_16_cmp_pReg_19, 
      gen_16_cmp_pReg_18, gen_16_cmp_pReg_17, gen_16_cmp_pReg_16, 
      gen_16_cmp_pReg_15, gen_16_cmp_pReg_14, gen_16_cmp_pReg_13, 
      gen_16_cmp_pReg_12, gen_16_cmp_pReg_11, gen_16_cmp_pReg_10, 
      gen_16_cmp_pReg_9, gen_16_cmp_pReg_8, gen_16_cmp_pReg_7, 
      gen_16_cmp_pReg_6, gen_16_cmp_pReg_5, gen_16_cmp_pReg_4, 
      gen_16_cmp_pReg_3, gen_16_cmp_pReg_2, gen_16_cmp_pReg_1, 
      gen_16_cmp_pReg_0, gen_16_cmp_BSCmp_op2_0, gen_16_cmp_BSCmp_carryIn, 
      gen_15_cmp_pBs_30, gen_15_cmp_pBs_29, gen_15_cmp_pBs_28, 
      gen_15_cmp_pBs_27, gen_15_cmp_pBs_26, gen_15_cmp_pBs_25, 
      gen_15_cmp_pBs_24, gen_15_cmp_pBs_23, gen_15_cmp_pMux_30, 
      gen_15_cmp_pMux_29, gen_15_cmp_pMux_28, gen_15_cmp_pMux_27, 
      gen_15_cmp_pMux_26, gen_15_cmp_pMux_25, gen_15_cmp_pMux_24, 
      gen_15_cmp_pMux_23, gen_15_cmp_pMux_22, gen_15_cmp_pMux_21, 
      gen_15_cmp_pMux_20, gen_15_cmp_pMux_19, gen_15_cmp_pMux_18, 
      gen_15_cmp_pMux_17, gen_15_cmp_pMux_16, gen_15_cmp_pMux_15, 
      gen_15_cmp_pMux_14, gen_15_cmp_pMux_13, gen_15_cmp_pMux_12, 
      gen_15_cmp_pMux_11, gen_15_cmp_pMux_10, gen_15_cmp_pMux_9, 
      gen_15_cmp_pMux_8, gen_15_cmp_pMux_7, gen_15_cmp_pMux_6, 
      gen_15_cmp_pMux_5, gen_15_cmp_pMux_4, gen_15_cmp_pMux_3, 
      gen_15_cmp_pMux_2, gen_15_cmp_pMux_1, gen_15_cmp_pMux_0, 
      gen_15_cmp_pReg_30, gen_15_cmp_pReg_29, gen_15_cmp_pReg_28, 
      gen_15_cmp_pReg_27, gen_15_cmp_pReg_26, gen_15_cmp_pReg_25, 
      gen_15_cmp_pReg_24, gen_15_cmp_pReg_23, gen_15_cmp_pReg_22, 
      gen_15_cmp_pReg_21, gen_15_cmp_pReg_20, gen_15_cmp_pReg_19, 
      gen_15_cmp_pReg_18, gen_15_cmp_pReg_17, gen_15_cmp_pReg_16, 
      gen_15_cmp_pReg_15, gen_15_cmp_pReg_14, gen_15_cmp_pReg_13, 
      gen_15_cmp_pReg_12, gen_15_cmp_pReg_11, gen_15_cmp_pReg_10, 
      gen_15_cmp_pReg_9, gen_15_cmp_pReg_8, gen_15_cmp_pReg_7, 
      gen_15_cmp_pReg_6, gen_15_cmp_pReg_5, gen_15_cmp_pReg_4, 
      gen_15_cmp_pReg_3, gen_15_cmp_pReg_2, gen_15_cmp_pReg_1, 
      gen_15_cmp_pReg_0, gen_15_cmp_BSCmp_op2_0, gen_15_cmp_BSCmp_carryIn, 
      gen_14_cmp_pBs_30, gen_14_cmp_pBs_29, gen_14_cmp_pBs_28, 
      gen_14_cmp_pBs_27, gen_14_cmp_pBs_26, gen_14_cmp_pBs_25, 
      gen_14_cmp_pBs_24, gen_14_cmp_pBs_23, gen_14_cmp_pMux_30, 
      gen_14_cmp_pMux_29, gen_14_cmp_pMux_28, gen_14_cmp_pMux_27, 
      gen_14_cmp_pMux_26, gen_14_cmp_pMux_25, gen_14_cmp_pMux_24, 
      gen_14_cmp_pMux_23, gen_14_cmp_pMux_22, gen_14_cmp_pMux_21, 
      gen_14_cmp_pMux_20, gen_14_cmp_pMux_19, gen_14_cmp_pMux_18, 
      gen_14_cmp_pMux_17, gen_14_cmp_pMux_16, gen_14_cmp_pMux_15, 
      gen_14_cmp_pMux_14, gen_14_cmp_pMux_13, gen_14_cmp_pMux_12, 
      gen_14_cmp_pMux_11, gen_14_cmp_pMux_10, gen_14_cmp_pMux_9, 
      gen_14_cmp_pMux_8, gen_14_cmp_pMux_7, gen_14_cmp_pMux_6, 
      gen_14_cmp_pMux_5, gen_14_cmp_pMux_4, gen_14_cmp_pMux_3, 
      gen_14_cmp_pMux_2, gen_14_cmp_pMux_1, gen_14_cmp_pMux_0, 
      gen_14_cmp_pReg_30, gen_14_cmp_pReg_29, gen_14_cmp_pReg_28, 
      gen_14_cmp_pReg_27, gen_14_cmp_pReg_26, gen_14_cmp_pReg_25, 
      gen_14_cmp_pReg_24, gen_14_cmp_pReg_23, gen_14_cmp_pReg_22, 
      gen_14_cmp_pReg_21, gen_14_cmp_pReg_20, gen_14_cmp_pReg_19, 
      gen_14_cmp_pReg_18, gen_14_cmp_pReg_17, gen_14_cmp_pReg_16, 
      gen_14_cmp_pReg_15, gen_14_cmp_pReg_14, gen_14_cmp_pReg_13, 
      gen_14_cmp_pReg_12, gen_14_cmp_pReg_11, gen_14_cmp_pReg_10, 
      gen_14_cmp_pReg_9, gen_14_cmp_pReg_8, gen_14_cmp_pReg_7, 
      gen_14_cmp_pReg_6, gen_14_cmp_pReg_5, gen_14_cmp_pReg_4, 
      gen_14_cmp_pReg_3, gen_14_cmp_pReg_2, gen_14_cmp_pReg_1, 
      gen_14_cmp_pReg_0, gen_14_cmp_BSCmp_op2_0, gen_14_cmp_BSCmp_carryIn, 
      gen_13_cmp_pBs_30, gen_13_cmp_pBs_29, gen_13_cmp_pBs_28, 
      gen_13_cmp_pBs_27, gen_13_cmp_pBs_26, gen_13_cmp_pBs_25, 
      gen_13_cmp_pBs_24, gen_13_cmp_pBs_23, gen_13_cmp_pMux_30, 
      gen_13_cmp_pMux_29, gen_13_cmp_pMux_28, gen_13_cmp_pMux_27, 
      gen_13_cmp_pMux_26, gen_13_cmp_pMux_25, gen_13_cmp_pMux_24, 
      gen_13_cmp_pMux_23, gen_13_cmp_pMux_22, gen_13_cmp_pMux_21, 
      gen_13_cmp_pMux_20, gen_13_cmp_pMux_19, gen_13_cmp_pMux_18, 
      gen_13_cmp_pMux_17, gen_13_cmp_pMux_16, gen_13_cmp_pMux_15, 
      gen_13_cmp_pMux_14, gen_13_cmp_pMux_13, gen_13_cmp_pMux_12, 
      gen_13_cmp_pMux_11, gen_13_cmp_pMux_10, gen_13_cmp_pMux_9, 
      gen_13_cmp_pMux_8, gen_13_cmp_pMux_7, gen_13_cmp_pMux_6, 
      gen_13_cmp_pMux_5, gen_13_cmp_pMux_4, gen_13_cmp_pMux_3, 
      gen_13_cmp_pMux_2, gen_13_cmp_pMux_1, gen_13_cmp_pMux_0, 
      gen_13_cmp_pReg_30, gen_13_cmp_pReg_29, gen_13_cmp_pReg_28, 
      gen_13_cmp_pReg_27, gen_13_cmp_pReg_26, gen_13_cmp_pReg_25, 
      gen_13_cmp_pReg_24, gen_13_cmp_pReg_23, gen_13_cmp_pReg_22, 
      gen_13_cmp_pReg_21, gen_13_cmp_pReg_20, gen_13_cmp_pReg_19, 
      gen_13_cmp_pReg_18, gen_13_cmp_pReg_17, gen_13_cmp_pReg_16, 
      gen_13_cmp_pReg_15, gen_13_cmp_pReg_14, gen_13_cmp_pReg_13, 
      gen_13_cmp_pReg_12, gen_13_cmp_pReg_11, gen_13_cmp_pReg_10, 
      gen_13_cmp_pReg_9, gen_13_cmp_pReg_8, gen_13_cmp_pReg_7, 
      gen_13_cmp_pReg_6, gen_13_cmp_pReg_5, gen_13_cmp_pReg_4, 
      gen_13_cmp_pReg_3, gen_13_cmp_pReg_2, gen_13_cmp_pReg_1, 
      gen_13_cmp_pReg_0, gen_13_cmp_BSCmp_op2_0, gen_13_cmp_BSCmp_carryIn, 
      gen_12_cmp_pBs_30, gen_12_cmp_pBs_29, gen_12_cmp_pBs_28, 
      gen_12_cmp_pBs_27, gen_12_cmp_pBs_26, gen_12_cmp_pBs_25, 
      gen_12_cmp_pBs_24, gen_12_cmp_pBs_23, gen_12_cmp_pMux_30, 
      gen_12_cmp_pMux_29, gen_12_cmp_pMux_28, gen_12_cmp_pMux_27, 
      gen_12_cmp_pMux_26, gen_12_cmp_pMux_25, gen_12_cmp_pMux_24, 
      gen_12_cmp_pMux_23, gen_12_cmp_pMux_22, gen_12_cmp_pMux_21, 
      gen_12_cmp_pMux_20, gen_12_cmp_pMux_19, gen_12_cmp_pMux_18, 
      gen_12_cmp_pMux_17, gen_12_cmp_pMux_16, gen_12_cmp_pMux_15, 
      gen_12_cmp_pMux_14, gen_12_cmp_pMux_13, gen_12_cmp_pMux_12, 
      gen_12_cmp_pMux_11, gen_12_cmp_pMux_10, gen_12_cmp_pMux_9, 
      gen_12_cmp_pMux_8, gen_12_cmp_pMux_7, gen_12_cmp_pMux_6, 
      gen_12_cmp_pMux_5, gen_12_cmp_pMux_4, gen_12_cmp_pMux_3, 
      gen_12_cmp_pMux_2, gen_12_cmp_pMux_1, gen_12_cmp_pMux_0, 
      gen_12_cmp_pReg_30, gen_12_cmp_pReg_29, gen_12_cmp_pReg_28, 
      gen_12_cmp_pReg_27, gen_12_cmp_pReg_26, gen_12_cmp_pReg_25, 
      gen_12_cmp_pReg_24, gen_12_cmp_pReg_23, gen_12_cmp_pReg_22, 
      gen_12_cmp_pReg_21, gen_12_cmp_pReg_20, gen_12_cmp_pReg_19, 
      gen_12_cmp_pReg_18, gen_12_cmp_pReg_17, gen_12_cmp_pReg_16, 
      gen_12_cmp_pReg_15, gen_12_cmp_pReg_14, gen_12_cmp_pReg_13, 
      gen_12_cmp_pReg_12, gen_12_cmp_pReg_11, gen_12_cmp_pReg_10, 
      gen_12_cmp_pReg_9, gen_12_cmp_pReg_8, gen_12_cmp_pReg_7, 
      gen_12_cmp_pReg_6, gen_12_cmp_pReg_5, gen_12_cmp_pReg_4, 
      gen_12_cmp_pReg_3, gen_12_cmp_pReg_2, gen_12_cmp_pReg_1, 
      gen_12_cmp_pReg_0, gen_12_cmp_BSCmp_op2_0, gen_12_cmp_BSCmp_carryIn, 
      gen_11_cmp_pBs_30, gen_11_cmp_pBs_29, gen_11_cmp_pBs_28, 
      gen_11_cmp_pBs_27, gen_11_cmp_pBs_26, gen_11_cmp_pBs_25, 
      gen_11_cmp_pBs_24, gen_11_cmp_pBs_23, gen_11_cmp_pMux_30, 
      gen_11_cmp_pMux_29, gen_11_cmp_pMux_28, gen_11_cmp_pMux_27, 
      gen_11_cmp_pMux_26, gen_11_cmp_pMux_25, gen_11_cmp_pMux_24, 
      gen_11_cmp_pMux_23, gen_11_cmp_pMux_22, gen_11_cmp_pMux_21, 
      gen_11_cmp_pMux_20, gen_11_cmp_pMux_19, gen_11_cmp_pMux_18, 
      gen_11_cmp_pMux_17, gen_11_cmp_pMux_16, gen_11_cmp_pMux_15, 
      gen_11_cmp_pMux_14, gen_11_cmp_pMux_13, gen_11_cmp_pMux_12, 
      gen_11_cmp_pMux_11, gen_11_cmp_pMux_10, gen_11_cmp_pMux_9, 
      gen_11_cmp_pMux_8, gen_11_cmp_pMux_7, gen_11_cmp_pMux_6, 
      gen_11_cmp_pMux_5, gen_11_cmp_pMux_4, gen_11_cmp_pMux_3, 
      gen_11_cmp_pMux_2, gen_11_cmp_pMux_1, gen_11_cmp_pMux_0, 
      gen_11_cmp_pReg_30, gen_11_cmp_pReg_29, gen_11_cmp_pReg_28, 
      gen_11_cmp_pReg_27, gen_11_cmp_pReg_26, gen_11_cmp_pReg_25, 
      gen_11_cmp_pReg_24, gen_11_cmp_pReg_23, gen_11_cmp_pReg_22, 
      gen_11_cmp_pReg_21, gen_11_cmp_pReg_20, gen_11_cmp_pReg_19, 
      gen_11_cmp_pReg_18, gen_11_cmp_pReg_17, gen_11_cmp_pReg_16, 
      gen_11_cmp_pReg_15, gen_11_cmp_pReg_14, gen_11_cmp_pReg_13, 
      gen_11_cmp_pReg_12, gen_11_cmp_pReg_11, gen_11_cmp_pReg_10, 
      gen_11_cmp_pReg_9, gen_11_cmp_pReg_8, gen_11_cmp_pReg_7, 
      gen_11_cmp_pReg_6, gen_11_cmp_pReg_5, gen_11_cmp_pReg_4, 
      gen_11_cmp_pReg_3, gen_11_cmp_pReg_2, gen_11_cmp_pReg_1, 
      gen_11_cmp_pReg_0, gen_11_cmp_BSCmp_op2_0, gen_11_cmp_BSCmp_carryIn, 
      gen_10_cmp_pBs_30, gen_10_cmp_pBs_29, gen_10_cmp_pBs_28, 
      gen_10_cmp_pBs_27, gen_10_cmp_pBs_26, gen_10_cmp_pBs_25, 
      gen_10_cmp_pBs_24, gen_10_cmp_pBs_23, gen_10_cmp_pMux_30, 
      gen_10_cmp_pMux_29, gen_10_cmp_pMux_28, gen_10_cmp_pMux_27, 
      gen_10_cmp_pMux_26, gen_10_cmp_pMux_25, gen_10_cmp_pMux_24, 
      gen_10_cmp_pMux_23, gen_10_cmp_pMux_22, gen_10_cmp_pMux_21, 
      gen_10_cmp_pMux_20, gen_10_cmp_pMux_19, gen_10_cmp_pMux_18, 
      gen_10_cmp_pMux_17, gen_10_cmp_pMux_16, gen_10_cmp_pMux_15, 
      gen_10_cmp_pMux_14, gen_10_cmp_pMux_13, gen_10_cmp_pMux_12, 
      gen_10_cmp_pMux_11, gen_10_cmp_pMux_10, gen_10_cmp_pMux_9, 
      gen_10_cmp_pMux_8, gen_10_cmp_pMux_7, gen_10_cmp_pMux_6, 
      gen_10_cmp_pMux_5, gen_10_cmp_pMux_4, gen_10_cmp_pMux_3, 
      gen_10_cmp_pMux_2, gen_10_cmp_pMux_1, gen_10_cmp_pMux_0, 
      gen_10_cmp_pReg_30, gen_10_cmp_pReg_29, gen_10_cmp_pReg_28, 
      gen_10_cmp_pReg_27, gen_10_cmp_pReg_26, gen_10_cmp_pReg_25, 
      gen_10_cmp_pReg_24, gen_10_cmp_pReg_23, gen_10_cmp_pReg_22, 
      gen_10_cmp_pReg_21, gen_10_cmp_pReg_20, gen_10_cmp_pReg_19, 
      gen_10_cmp_pReg_18, gen_10_cmp_pReg_17, gen_10_cmp_pReg_16, 
      gen_10_cmp_pReg_15, gen_10_cmp_pReg_14, gen_10_cmp_pReg_13, 
      gen_10_cmp_pReg_12, gen_10_cmp_pReg_11, gen_10_cmp_pReg_10, 
      gen_10_cmp_pReg_9, gen_10_cmp_pReg_8, gen_10_cmp_pReg_7, 
      gen_10_cmp_pReg_6, gen_10_cmp_pReg_5, gen_10_cmp_pReg_4, 
      gen_10_cmp_pReg_3, gen_10_cmp_pReg_2, gen_10_cmp_pReg_1, 
      gen_10_cmp_pReg_0, gen_10_cmp_BSCmp_op2_0, gen_10_cmp_BSCmp_carryIn, 
      gen_9_cmp_pBs_30, gen_9_cmp_pBs_29, gen_9_cmp_pBs_28, gen_9_cmp_pBs_27, 
      gen_9_cmp_pBs_26, gen_9_cmp_pBs_25, gen_9_cmp_pBs_24, gen_9_cmp_pBs_23, 
      gen_9_cmp_pMux_30, gen_9_cmp_pMux_29, gen_9_cmp_pMux_28, 
      gen_9_cmp_pMux_27, gen_9_cmp_pMux_26, gen_9_cmp_pMux_25, 
      gen_9_cmp_pMux_24, gen_9_cmp_pMux_23, gen_9_cmp_pMux_22, 
      gen_9_cmp_pMux_21, gen_9_cmp_pMux_20, gen_9_cmp_pMux_19, 
      gen_9_cmp_pMux_18, gen_9_cmp_pMux_17, gen_9_cmp_pMux_16, 
      gen_9_cmp_pMux_15, gen_9_cmp_pMux_14, gen_9_cmp_pMux_13, 
      gen_9_cmp_pMux_12, gen_9_cmp_pMux_11, gen_9_cmp_pMux_10, 
      gen_9_cmp_pMux_9, gen_9_cmp_pMux_8, gen_9_cmp_pMux_7, gen_9_cmp_pMux_6, 
      gen_9_cmp_pMux_5, gen_9_cmp_pMux_4, gen_9_cmp_pMux_3, gen_9_cmp_pMux_2, 
      gen_9_cmp_pMux_1, gen_9_cmp_pMux_0, gen_9_cmp_pReg_30, 
      gen_9_cmp_pReg_29, gen_9_cmp_pReg_28, gen_9_cmp_pReg_27, 
      gen_9_cmp_pReg_26, gen_9_cmp_pReg_25, gen_9_cmp_pReg_24, 
      gen_9_cmp_pReg_23, gen_9_cmp_pReg_22, gen_9_cmp_pReg_21, 
      gen_9_cmp_pReg_20, gen_9_cmp_pReg_19, gen_9_cmp_pReg_18, 
      gen_9_cmp_pReg_17, gen_9_cmp_pReg_16, gen_9_cmp_pReg_15, 
      gen_9_cmp_pReg_14, gen_9_cmp_pReg_13, gen_9_cmp_pReg_12, 
      gen_9_cmp_pReg_11, gen_9_cmp_pReg_10, gen_9_cmp_pReg_9, 
      gen_9_cmp_pReg_8, gen_9_cmp_pReg_7, gen_9_cmp_pReg_6, gen_9_cmp_pReg_5, 
      gen_9_cmp_pReg_4, gen_9_cmp_pReg_3, gen_9_cmp_pReg_2, gen_9_cmp_pReg_1, 
      gen_9_cmp_pReg_0, gen_9_cmp_BSCmp_op2_0, gen_9_cmp_BSCmp_carryIn, 
      gen_8_cmp_pBs_30, gen_8_cmp_pBs_29, gen_8_cmp_pBs_28, gen_8_cmp_pBs_27, 
      gen_8_cmp_pBs_26, gen_8_cmp_pBs_25, gen_8_cmp_pBs_24, gen_8_cmp_pBs_23, 
      gen_8_cmp_pMux_30, gen_8_cmp_pMux_29, gen_8_cmp_pMux_28, 
      gen_8_cmp_pMux_27, gen_8_cmp_pMux_26, gen_8_cmp_pMux_25, 
      gen_8_cmp_pMux_24, gen_8_cmp_pMux_23, gen_8_cmp_pMux_22, 
      gen_8_cmp_pMux_21, gen_8_cmp_pMux_20, gen_8_cmp_pMux_19, 
      gen_8_cmp_pMux_18, gen_8_cmp_pMux_17, gen_8_cmp_pMux_16, 
      gen_8_cmp_pMux_15, gen_8_cmp_pMux_14, gen_8_cmp_pMux_13, 
      gen_8_cmp_pMux_12, gen_8_cmp_pMux_11, gen_8_cmp_pMux_10, 
      gen_8_cmp_pMux_9, gen_8_cmp_pMux_8, gen_8_cmp_pMux_7, gen_8_cmp_pMux_6, 
      gen_8_cmp_pMux_5, gen_8_cmp_pMux_4, gen_8_cmp_pMux_3, gen_8_cmp_pMux_2, 
      gen_8_cmp_pMux_1, gen_8_cmp_pMux_0, gen_8_cmp_pReg_30, 
      gen_8_cmp_pReg_29, gen_8_cmp_pReg_28, gen_8_cmp_pReg_27, 
      gen_8_cmp_pReg_26, gen_8_cmp_pReg_25, gen_8_cmp_pReg_24, 
      gen_8_cmp_pReg_23, gen_8_cmp_pReg_22, gen_8_cmp_pReg_21, 
      gen_8_cmp_pReg_20, gen_8_cmp_pReg_19, gen_8_cmp_pReg_18, 
      gen_8_cmp_pReg_17, gen_8_cmp_pReg_16, gen_8_cmp_pReg_15, 
      gen_8_cmp_pReg_14, gen_8_cmp_pReg_13, gen_8_cmp_pReg_12, 
      gen_8_cmp_pReg_11, gen_8_cmp_pReg_10, gen_8_cmp_pReg_9, 
      gen_8_cmp_pReg_8, gen_8_cmp_pReg_7, gen_8_cmp_pReg_6, gen_8_cmp_pReg_5, 
      gen_8_cmp_pReg_4, gen_8_cmp_pReg_3, gen_8_cmp_pReg_2, gen_8_cmp_pReg_1, 
      gen_8_cmp_pReg_0, gen_8_cmp_BSCmp_op2_0, gen_8_cmp_BSCmp_carryIn, 
      gen_7_cmp_pBs_30, gen_7_cmp_pBs_29, gen_7_cmp_pBs_28, gen_7_cmp_pBs_27, 
      gen_7_cmp_pBs_26, gen_7_cmp_pBs_25, gen_7_cmp_pBs_24, gen_7_cmp_pBs_23, 
      gen_7_cmp_pMux_30, gen_7_cmp_pMux_29, gen_7_cmp_pMux_28, 
      gen_7_cmp_pMux_27, gen_7_cmp_pMux_26, gen_7_cmp_pMux_25, 
      gen_7_cmp_pMux_24, gen_7_cmp_pMux_23, gen_7_cmp_pMux_22, 
      gen_7_cmp_pMux_21, gen_7_cmp_pMux_20, gen_7_cmp_pMux_19, 
      gen_7_cmp_pMux_18, gen_7_cmp_pMux_17, gen_7_cmp_pMux_16, 
      gen_7_cmp_pMux_15, gen_7_cmp_pMux_14, gen_7_cmp_pMux_13, 
      gen_7_cmp_pMux_12, gen_7_cmp_pMux_11, gen_7_cmp_pMux_10, 
      gen_7_cmp_pMux_9, gen_7_cmp_pMux_8, gen_7_cmp_pMux_7, gen_7_cmp_pMux_6, 
      gen_7_cmp_pMux_5, gen_7_cmp_pMux_4, gen_7_cmp_pMux_3, gen_7_cmp_pMux_2, 
      gen_7_cmp_pMux_1, gen_7_cmp_pMux_0, gen_7_cmp_pReg_30, 
      gen_7_cmp_pReg_29, gen_7_cmp_pReg_28, gen_7_cmp_pReg_27, 
      gen_7_cmp_pReg_26, gen_7_cmp_pReg_25, gen_7_cmp_pReg_24, 
      gen_7_cmp_pReg_23, gen_7_cmp_pReg_22, gen_7_cmp_pReg_21, 
      gen_7_cmp_pReg_20, gen_7_cmp_pReg_19, gen_7_cmp_pReg_18, 
      gen_7_cmp_pReg_17, gen_7_cmp_pReg_16, gen_7_cmp_pReg_15, 
      gen_7_cmp_pReg_14, gen_7_cmp_pReg_13, gen_7_cmp_pReg_12, 
      gen_7_cmp_pReg_11, gen_7_cmp_pReg_10, gen_7_cmp_pReg_9, 
      gen_7_cmp_pReg_8, gen_7_cmp_pReg_7, gen_7_cmp_pReg_6, gen_7_cmp_pReg_5, 
      gen_7_cmp_pReg_4, gen_7_cmp_pReg_3, gen_7_cmp_pReg_2, gen_7_cmp_pReg_1, 
      gen_7_cmp_pReg_0, gen_7_cmp_BSCmp_op2_0, gen_7_cmp_BSCmp_carryIn, 
      gen_6_cmp_pBs_30, gen_6_cmp_pBs_29, gen_6_cmp_pBs_28, gen_6_cmp_pBs_27, 
      gen_6_cmp_pBs_26, gen_6_cmp_pBs_25, gen_6_cmp_pBs_24, gen_6_cmp_pBs_23, 
      gen_6_cmp_pMux_30, gen_6_cmp_pMux_29, gen_6_cmp_pMux_28, 
      gen_6_cmp_pMux_27, gen_6_cmp_pMux_26, gen_6_cmp_pMux_25, 
      gen_6_cmp_pMux_24, gen_6_cmp_pMux_23, gen_6_cmp_pMux_22, 
      gen_6_cmp_pMux_21, gen_6_cmp_pMux_20, gen_6_cmp_pMux_19, 
      gen_6_cmp_pMux_18, gen_6_cmp_pMux_17, gen_6_cmp_pMux_16, 
      gen_6_cmp_pMux_15, gen_6_cmp_pMux_14, gen_6_cmp_pMux_13, 
      gen_6_cmp_pMux_12, gen_6_cmp_pMux_11, gen_6_cmp_pMux_10, 
      gen_6_cmp_pMux_9, gen_6_cmp_pMux_8, gen_6_cmp_pMux_7, gen_6_cmp_pMux_6, 
      gen_6_cmp_pMux_5, gen_6_cmp_pMux_4, gen_6_cmp_pMux_3, gen_6_cmp_pMux_2, 
      gen_6_cmp_pMux_1, gen_6_cmp_pMux_0, gen_6_cmp_pReg_30, 
      gen_6_cmp_pReg_29, gen_6_cmp_pReg_28, gen_6_cmp_pReg_27, 
      gen_6_cmp_pReg_26, gen_6_cmp_pReg_25, gen_6_cmp_pReg_24, 
      gen_6_cmp_pReg_23, gen_6_cmp_pReg_22, gen_6_cmp_pReg_21, 
      gen_6_cmp_pReg_20, gen_6_cmp_pReg_19, gen_6_cmp_pReg_18, 
      gen_6_cmp_pReg_17, gen_6_cmp_pReg_16, gen_6_cmp_pReg_15, 
      gen_6_cmp_pReg_14, gen_6_cmp_pReg_13, gen_6_cmp_pReg_12, 
      gen_6_cmp_pReg_11, gen_6_cmp_pReg_10, gen_6_cmp_pReg_9, 
      gen_6_cmp_pReg_8, gen_6_cmp_pReg_7, gen_6_cmp_pReg_6, gen_6_cmp_pReg_5, 
      gen_6_cmp_pReg_4, gen_6_cmp_pReg_3, gen_6_cmp_pReg_2, gen_6_cmp_pReg_1, 
      gen_6_cmp_pReg_0, gen_6_cmp_BSCmp_op2_0, gen_6_cmp_BSCmp_carryIn, 
      gen_5_cmp_pBs_30, gen_5_cmp_pBs_29, gen_5_cmp_pBs_28, gen_5_cmp_pBs_27, 
      gen_5_cmp_pBs_26, gen_5_cmp_pBs_25, gen_5_cmp_pBs_24, gen_5_cmp_pBs_23, 
      gen_5_cmp_pMux_30, gen_5_cmp_pMux_29, gen_5_cmp_pMux_28, 
      gen_5_cmp_pMux_27, gen_5_cmp_pMux_26, gen_5_cmp_pMux_25, 
      gen_5_cmp_pMux_24, gen_5_cmp_pMux_23, gen_5_cmp_pMux_22, 
      gen_5_cmp_pMux_21, gen_5_cmp_pMux_20, gen_5_cmp_pMux_19, 
      gen_5_cmp_pMux_18, gen_5_cmp_pMux_17, gen_5_cmp_pMux_16, 
      gen_5_cmp_pMux_15, gen_5_cmp_pMux_14, gen_5_cmp_pMux_13, 
      gen_5_cmp_pMux_12, gen_5_cmp_pMux_11, gen_5_cmp_pMux_10, 
      gen_5_cmp_pMux_9, gen_5_cmp_pMux_8, gen_5_cmp_pMux_7, gen_5_cmp_pMux_6, 
      gen_5_cmp_pMux_5, gen_5_cmp_pMux_4, gen_5_cmp_pMux_3, gen_5_cmp_pMux_2, 
      gen_5_cmp_pMux_1, gen_5_cmp_pMux_0, gen_5_cmp_pReg_30, 
      gen_5_cmp_pReg_29, gen_5_cmp_pReg_28, gen_5_cmp_pReg_27, 
      gen_5_cmp_pReg_26, gen_5_cmp_pReg_25, gen_5_cmp_pReg_24, 
      gen_5_cmp_pReg_23, gen_5_cmp_pReg_22, gen_5_cmp_pReg_21, 
      gen_5_cmp_pReg_20, gen_5_cmp_pReg_19, gen_5_cmp_pReg_18, 
      gen_5_cmp_pReg_17, gen_5_cmp_pReg_16, gen_5_cmp_pReg_15, 
      gen_5_cmp_pReg_14, gen_5_cmp_pReg_13, gen_5_cmp_pReg_12, 
      gen_5_cmp_pReg_11, gen_5_cmp_pReg_10, gen_5_cmp_pReg_9, 
      gen_5_cmp_pReg_8, gen_5_cmp_pReg_7, gen_5_cmp_pReg_6, gen_5_cmp_pReg_5, 
      gen_5_cmp_pReg_4, gen_5_cmp_pReg_3, gen_5_cmp_pReg_2, gen_5_cmp_pReg_1, 
      gen_5_cmp_pReg_0, gen_5_cmp_BSCmp_op2_0, gen_5_cmp_BSCmp_carryIn, 
      gen_4_cmp_pBs_30, gen_4_cmp_pBs_29, gen_4_cmp_pBs_28, gen_4_cmp_pBs_27, 
      gen_4_cmp_pBs_26, gen_4_cmp_pBs_25, gen_4_cmp_pBs_24, gen_4_cmp_pBs_23, 
      gen_4_cmp_pMux_30, gen_4_cmp_pMux_29, gen_4_cmp_pMux_28, 
      gen_4_cmp_pMux_27, gen_4_cmp_pMux_26, gen_4_cmp_pMux_25, 
      gen_4_cmp_pMux_24, gen_4_cmp_pMux_23, gen_4_cmp_pMux_22, 
      gen_4_cmp_pMux_21, gen_4_cmp_pMux_20, gen_4_cmp_pMux_19, 
      gen_4_cmp_pMux_18, gen_4_cmp_pMux_17, gen_4_cmp_pMux_16, 
      gen_4_cmp_pMux_15, gen_4_cmp_pMux_14, gen_4_cmp_pMux_13, 
      gen_4_cmp_pMux_12, gen_4_cmp_pMux_11, gen_4_cmp_pMux_10, 
      gen_4_cmp_pMux_9, gen_4_cmp_pMux_8, gen_4_cmp_pMux_7, gen_4_cmp_pMux_6, 
      gen_4_cmp_pMux_5, gen_4_cmp_pMux_4, gen_4_cmp_pMux_3, gen_4_cmp_pMux_2, 
      gen_4_cmp_pMux_1, gen_4_cmp_pMux_0, gen_4_cmp_pReg_30, 
      gen_4_cmp_pReg_29, gen_4_cmp_pReg_28, gen_4_cmp_pReg_27, 
      gen_4_cmp_pReg_26, gen_4_cmp_pReg_25, gen_4_cmp_pReg_24, 
      gen_4_cmp_pReg_23, gen_4_cmp_pReg_22, gen_4_cmp_pReg_21, 
      gen_4_cmp_pReg_20, gen_4_cmp_pReg_19, gen_4_cmp_pReg_18, 
      gen_4_cmp_pReg_17, gen_4_cmp_pReg_16, gen_4_cmp_pReg_15, 
      gen_4_cmp_pReg_14, gen_4_cmp_pReg_13, gen_4_cmp_pReg_12, 
      gen_4_cmp_pReg_11, gen_4_cmp_pReg_10, gen_4_cmp_pReg_9, 
      gen_4_cmp_pReg_8, gen_4_cmp_pReg_7, gen_4_cmp_pReg_6, gen_4_cmp_pReg_5, 
      gen_4_cmp_pReg_4, gen_4_cmp_pReg_3, gen_4_cmp_pReg_2, gen_4_cmp_pReg_1, 
      gen_4_cmp_pReg_0, gen_4_cmp_BSCmp_op2_0, gen_4_cmp_BSCmp_carryIn, 
      gen_3_cmp_pBs_30, gen_3_cmp_pBs_29, gen_3_cmp_pBs_28, gen_3_cmp_pBs_27, 
      gen_3_cmp_pBs_26, gen_3_cmp_pBs_25, gen_3_cmp_pBs_24, gen_3_cmp_pBs_23, 
      gen_3_cmp_pMux_30, gen_3_cmp_pMux_29, gen_3_cmp_pMux_28, 
      gen_3_cmp_pMux_27, gen_3_cmp_pMux_26, gen_3_cmp_pMux_25, 
      gen_3_cmp_pMux_24, gen_3_cmp_pMux_23, gen_3_cmp_pMux_22, 
      gen_3_cmp_pMux_21, gen_3_cmp_pMux_20, gen_3_cmp_pMux_19, 
      gen_3_cmp_pMux_18, gen_3_cmp_pMux_17, gen_3_cmp_pMux_16, 
      gen_3_cmp_pMux_15, gen_3_cmp_pMux_14, gen_3_cmp_pMux_13, 
      gen_3_cmp_pMux_12, gen_3_cmp_pMux_11, gen_3_cmp_pMux_10, 
      gen_3_cmp_pMux_9, gen_3_cmp_pMux_8, gen_3_cmp_pMux_7, gen_3_cmp_pMux_6, 
      gen_3_cmp_pMux_5, gen_3_cmp_pMux_4, gen_3_cmp_pMux_3, gen_3_cmp_pMux_2, 
      gen_3_cmp_pMux_1, gen_3_cmp_pMux_0, gen_3_cmp_pReg_30, 
      gen_3_cmp_pReg_29, gen_3_cmp_pReg_28, gen_3_cmp_pReg_27, 
      gen_3_cmp_pReg_26, gen_3_cmp_pReg_25, gen_3_cmp_pReg_24, 
      gen_3_cmp_pReg_23, gen_3_cmp_pReg_22, gen_3_cmp_pReg_21, 
      gen_3_cmp_pReg_20, gen_3_cmp_pReg_19, gen_3_cmp_pReg_18, 
      gen_3_cmp_pReg_17, gen_3_cmp_pReg_16, gen_3_cmp_pReg_15, 
      gen_3_cmp_pReg_14, gen_3_cmp_pReg_13, gen_3_cmp_pReg_12, 
      gen_3_cmp_pReg_11, gen_3_cmp_pReg_10, gen_3_cmp_pReg_9, 
      gen_3_cmp_pReg_8, gen_3_cmp_pReg_7, gen_3_cmp_pReg_6, gen_3_cmp_pReg_5, 
      gen_3_cmp_pReg_4, gen_3_cmp_pReg_3, gen_3_cmp_pReg_2, gen_3_cmp_pReg_1, 
      gen_3_cmp_pReg_0, gen_3_cmp_BSCmp_op2_0, gen_3_cmp_BSCmp_carryIn, 
      gen_2_cmp_pBs_30, gen_2_cmp_pBs_29, gen_2_cmp_pBs_28, gen_2_cmp_pBs_27, 
      gen_2_cmp_pBs_26, gen_2_cmp_pBs_25, gen_2_cmp_pBs_24, gen_2_cmp_pBs_23, 
      gen_2_cmp_pMux_30, gen_2_cmp_pMux_29, gen_2_cmp_pMux_28, 
      gen_2_cmp_pMux_27, gen_2_cmp_pMux_26, gen_2_cmp_pMux_25, 
      gen_2_cmp_pMux_24, gen_2_cmp_pMux_23, gen_2_cmp_pMux_22, 
      gen_2_cmp_pMux_21, gen_2_cmp_pMux_20, gen_2_cmp_pMux_19, 
      gen_2_cmp_pMux_18, gen_2_cmp_pMux_17, gen_2_cmp_pMux_16, 
      gen_2_cmp_pMux_15, gen_2_cmp_pMux_14, gen_2_cmp_pMux_13, 
      gen_2_cmp_pMux_12, gen_2_cmp_pMux_11, gen_2_cmp_pMux_10, 
      gen_2_cmp_pMux_9, gen_2_cmp_pMux_8, gen_2_cmp_pMux_7, gen_2_cmp_pMux_6, 
      gen_2_cmp_pMux_5, gen_2_cmp_pMux_4, gen_2_cmp_pMux_3, gen_2_cmp_pMux_2, 
      gen_2_cmp_pMux_1, gen_2_cmp_pMux_0, gen_2_cmp_pReg_30, 
      gen_2_cmp_pReg_29, gen_2_cmp_pReg_28, gen_2_cmp_pReg_27, 
      gen_2_cmp_pReg_26, gen_2_cmp_pReg_25, gen_2_cmp_pReg_24, 
      gen_2_cmp_pReg_23, gen_2_cmp_pReg_22, gen_2_cmp_pReg_21, 
      gen_2_cmp_pReg_20, gen_2_cmp_pReg_19, gen_2_cmp_pReg_18, 
      gen_2_cmp_pReg_17, gen_2_cmp_pReg_16, gen_2_cmp_pReg_15, 
      gen_2_cmp_pReg_14, gen_2_cmp_pReg_13, gen_2_cmp_pReg_12, 
      gen_2_cmp_pReg_11, gen_2_cmp_pReg_10, gen_2_cmp_pReg_9, 
      gen_2_cmp_pReg_8, gen_2_cmp_pReg_7, gen_2_cmp_pReg_6, gen_2_cmp_pReg_5, 
      gen_2_cmp_pReg_4, gen_2_cmp_pReg_3, gen_2_cmp_pReg_2, gen_2_cmp_pReg_1, 
      gen_2_cmp_pReg_0, gen_2_cmp_BSCmp_op2_0, gen_2_cmp_BSCmp_carryIn, 
      gen_1_cmp_pBs_30, gen_1_cmp_pBs_29, gen_1_cmp_pBs_28, gen_1_cmp_pBs_27, 
      gen_1_cmp_pBs_26, gen_1_cmp_pBs_25, gen_1_cmp_pBs_24, gen_1_cmp_pBs_23, 
      gen_1_cmp_pMux_30, gen_1_cmp_pMux_29, gen_1_cmp_pMux_28, 
      gen_1_cmp_pMux_27, gen_1_cmp_pMux_26, gen_1_cmp_pMux_25, 
      gen_1_cmp_pMux_24, gen_1_cmp_pMux_23, gen_1_cmp_pMux_22, 
      gen_1_cmp_pMux_21, gen_1_cmp_pMux_20, gen_1_cmp_pMux_19, 
      gen_1_cmp_pMux_18, gen_1_cmp_pMux_17, gen_1_cmp_pMux_16, 
      gen_1_cmp_pMux_15, gen_1_cmp_pMux_14, gen_1_cmp_pMux_13, 
      gen_1_cmp_pMux_12, gen_1_cmp_pMux_11, gen_1_cmp_pMux_10, 
      gen_1_cmp_pMux_9, gen_1_cmp_pMux_8, gen_1_cmp_pMux_7, gen_1_cmp_pMux_6, 
      gen_1_cmp_pMux_5, gen_1_cmp_pMux_4, gen_1_cmp_pMux_3, gen_1_cmp_pMux_2, 
      gen_1_cmp_pMux_1, gen_1_cmp_pMux_0, gen_1_cmp_pReg_30, 
      gen_1_cmp_pReg_29, gen_1_cmp_pReg_28, gen_1_cmp_pReg_27, 
      gen_1_cmp_pReg_26, gen_1_cmp_pReg_25, gen_1_cmp_pReg_24, 
      gen_1_cmp_pReg_23, gen_1_cmp_pReg_22, gen_1_cmp_pReg_21, 
      gen_1_cmp_pReg_20, gen_1_cmp_pReg_19, gen_1_cmp_pReg_18, 
      gen_1_cmp_pReg_17, gen_1_cmp_pReg_16, gen_1_cmp_pReg_15, 
      gen_1_cmp_pReg_14, gen_1_cmp_pReg_13, gen_1_cmp_pReg_12, 
      gen_1_cmp_pReg_11, gen_1_cmp_pReg_10, gen_1_cmp_pReg_9, 
      gen_1_cmp_pReg_8, gen_1_cmp_pReg_7, gen_1_cmp_pReg_6, gen_1_cmp_pReg_5, 
      gen_1_cmp_pReg_4, gen_1_cmp_pReg_3, gen_1_cmp_pReg_2, gen_1_cmp_pReg_1, 
      gen_1_cmp_pReg_0, gen_1_cmp_BSCmp_op2_0, gen_1_cmp_BSCmp_carryIn, 
      gen_0_cmp_pBs_30, gen_0_cmp_pBs_29, gen_0_cmp_pBs_28, gen_0_cmp_pBs_27, 
      gen_0_cmp_pBs_26, gen_0_cmp_pBs_25, gen_0_cmp_pBs_24, gen_0_cmp_pBs_23, 
      gen_0_cmp_pMux_30, gen_0_cmp_pMux_29, gen_0_cmp_pMux_28, 
      gen_0_cmp_pMux_27, gen_0_cmp_pMux_26, gen_0_cmp_pMux_25, 
      gen_0_cmp_pMux_24, gen_0_cmp_pMux_23, gen_0_cmp_pMux_22, 
      gen_0_cmp_pMux_21, gen_0_cmp_pMux_20, gen_0_cmp_pMux_19, 
      gen_0_cmp_pMux_18, gen_0_cmp_pMux_17, gen_0_cmp_pMux_16, 
      gen_0_cmp_pMux_15, gen_0_cmp_pMux_14, gen_0_cmp_pMux_13, 
      gen_0_cmp_pMux_12, gen_0_cmp_pMux_11, gen_0_cmp_pMux_10, 
      gen_0_cmp_pMux_9, gen_0_cmp_pMux_8, gen_0_cmp_pMux_7, gen_0_cmp_pMux_6, 
      gen_0_cmp_pMux_5, gen_0_cmp_pMux_4, gen_0_cmp_pMux_3, gen_0_cmp_pMux_2, 
      gen_0_cmp_pMux_1, gen_0_cmp_pMux_0, gen_0_cmp_pReg_30, 
      gen_0_cmp_pReg_29, gen_0_cmp_pReg_28, gen_0_cmp_pReg_27, 
      gen_0_cmp_pReg_26, gen_0_cmp_pReg_25, gen_0_cmp_pReg_24, 
      gen_0_cmp_pReg_23, gen_0_cmp_pReg_22, gen_0_cmp_pReg_21, 
      gen_0_cmp_pReg_20, gen_0_cmp_pReg_19, gen_0_cmp_pReg_18, 
      gen_0_cmp_pReg_17, gen_0_cmp_pReg_16, gen_0_cmp_pReg_15, 
      gen_0_cmp_pReg_14, gen_0_cmp_pReg_13, gen_0_cmp_pReg_12, 
      gen_0_cmp_pReg_11, gen_0_cmp_pReg_10, gen_0_cmp_pReg_9, 
      gen_0_cmp_pReg_8, gen_0_cmp_pReg_7, gen_0_cmp_pReg_6, gen_0_cmp_pReg_5, 
      gen_0_cmp_pReg_4, gen_0_cmp_pReg_3, gen_0_cmp_pReg_2, gen_0_cmp_pReg_1, 
      gen_0_cmp_pReg_0, gen_0_cmp_BSCmp_op2_0, gen_0_cmp_BSCmp_carryIn, 
      gen_24_cmp_BSCmp_op2_16, gen_24_cmp_BSCmp_op2_15, 
      gen_24_cmp_BSCmp_op2_14, gen_24_cmp_BSCmp_op2_13, 
      gen_24_cmp_BSCmp_op2_12, gen_24_cmp_BSCmp_op2_11, 
      gen_24_cmp_BSCmp_op2_10, gen_24_cmp_BSCmp_op2_9, 
      gen_24_cmp_BSCmp_op2_8, gen_24_cmp_BSCmp_op2_7, gen_24_cmp_BSCmp_op2_6, 
      gen_24_cmp_BSCmp_op2_5, gen_24_cmp_BSCmp_op2_4, gen_24_cmp_BSCmp_op2_3, 
      gen_24_cmp_BSCmp_op2_2, gen_24_cmp_BSCmp_op2_1, 
      gen_23_cmp_BSCmp_op2_16, gen_23_cmp_BSCmp_op2_15, 
      gen_23_cmp_BSCmp_op2_14, gen_23_cmp_BSCmp_op2_13, 
      gen_23_cmp_BSCmp_op2_12, gen_23_cmp_BSCmp_op2_11, 
      gen_23_cmp_BSCmp_op2_10, gen_23_cmp_BSCmp_op2_9, 
      gen_23_cmp_BSCmp_op2_8, gen_23_cmp_BSCmp_op2_7, gen_23_cmp_BSCmp_op2_6, 
      gen_23_cmp_BSCmp_op2_5, gen_23_cmp_BSCmp_op2_4, gen_23_cmp_BSCmp_op2_3, 
      gen_23_cmp_BSCmp_op2_2, gen_23_cmp_BSCmp_op2_1, 
      gen_22_cmp_BSCmp_op2_16, gen_22_cmp_BSCmp_op2_15, 
      gen_22_cmp_BSCmp_op2_14, gen_22_cmp_BSCmp_op2_13, 
      gen_22_cmp_BSCmp_op2_12, gen_22_cmp_BSCmp_op2_11, 
      gen_22_cmp_BSCmp_op2_10, gen_22_cmp_BSCmp_op2_9, 
      gen_22_cmp_BSCmp_op2_8, gen_22_cmp_BSCmp_op2_7, gen_22_cmp_BSCmp_op2_6, 
      gen_22_cmp_BSCmp_op2_5, gen_22_cmp_BSCmp_op2_4, gen_22_cmp_BSCmp_op2_3, 
      gen_22_cmp_BSCmp_op2_2, gen_22_cmp_BSCmp_op2_1, 
      gen_21_cmp_BSCmp_op2_16, gen_21_cmp_BSCmp_op2_15, 
      gen_21_cmp_BSCmp_op2_14, gen_21_cmp_BSCmp_op2_13, 
      gen_21_cmp_BSCmp_op2_12, gen_21_cmp_BSCmp_op2_11, 
      gen_21_cmp_BSCmp_op2_10, gen_21_cmp_BSCmp_op2_9, 
      gen_21_cmp_BSCmp_op2_8, gen_21_cmp_BSCmp_op2_7, gen_21_cmp_BSCmp_op2_6, 
      gen_21_cmp_BSCmp_op2_5, gen_21_cmp_BSCmp_op2_4, gen_21_cmp_BSCmp_op2_3, 
      gen_21_cmp_BSCmp_op2_2, gen_21_cmp_BSCmp_op2_1, 
      gen_20_cmp_BSCmp_op2_16, gen_20_cmp_BSCmp_op2_15, 
      gen_20_cmp_BSCmp_op2_14, gen_20_cmp_BSCmp_op2_13, 
      gen_20_cmp_BSCmp_op2_12, gen_20_cmp_BSCmp_op2_11, 
      gen_20_cmp_BSCmp_op2_10, gen_20_cmp_BSCmp_op2_9, 
      gen_20_cmp_BSCmp_op2_8, gen_20_cmp_BSCmp_op2_7, gen_20_cmp_BSCmp_op2_6, 
      gen_20_cmp_BSCmp_op2_5, gen_20_cmp_BSCmp_op2_4, gen_20_cmp_BSCmp_op2_3, 
      gen_20_cmp_BSCmp_op2_2, gen_20_cmp_BSCmp_op2_1, 
      gen_19_cmp_BSCmp_op2_16, gen_19_cmp_BSCmp_op2_15, 
      gen_19_cmp_BSCmp_op2_14, gen_19_cmp_BSCmp_op2_13, 
      gen_19_cmp_BSCmp_op2_12, gen_19_cmp_BSCmp_op2_11, 
      gen_19_cmp_BSCmp_op2_10, gen_19_cmp_BSCmp_op2_9, 
      gen_19_cmp_BSCmp_op2_8, gen_19_cmp_BSCmp_op2_7, gen_19_cmp_BSCmp_op2_6, 
      gen_19_cmp_BSCmp_op2_5, gen_19_cmp_BSCmp_op2_4, gen_19_cmp_BSCmp_op2_3, 
      gen_19_cmp_BSCmp_op2_2, gen_19_cmp_BSCmp_op2_1, 
      gen_18_cmp_BSCmp_op2_16, gen_18_cmp_BSCmp_op2_15, 
      gen_18_cmp_BSCmp_op2_14, gen_18_cmp_BSCmp_op2_13, 
      gen_18_cmp_BSCmp_op2_12, gen_18_cmp_BSCmp_op2_11, 
      gen_18_cmp_BSCmp_op2_10, gen_18_cmp_BSCmp_op2_9, 
      gen_18_cmp_BSCmp_op2_8, gen_18_cmp_BSCmp_op2_7, gen_18_cmp_BSCmp_op2_6, 
      gen_18_cmp_BSCmp_op2_5, gen_18_cmp_BSCmp_op2_4, gen_18_cmp_BSCmp_op2_3, 
      gen_18_cmp_BSCmp_op2_2, gen_18_cmp_BSCmp_op2_1, 
      gen_17_cmp_BSCmp_op2_16, gen_17_cmp_BSCmp_op2_15, 
      gen_17_cmp_BSCmp_op2_14, gen_17_cmp_BSCmp_op2_13, 
      gen_17_cmp_BSCmp_op2_12, gen_17_cmp_BSCmp_op2_11, 
      gen_17_cmp_BSCmp_op2_10, gen_17_cmp_BSCmp_op2_9, 
      gen_17_cmp_BSCmp_op2_8, gen_17_cmp_BSCmp_op2_7, gen_17_cmp_BSCmp_op2_6, 
      gen_17_cmp_BSCmp_op2_5, gen_17_cmp_BSCmp_op2_4, gen_17_cmp_BSCmp_op2_3, 
      gen_17_cmp_BSCmp_op2_2, gen_17_cmp_BSCmp_op2_1, 
      gen_16_cmp_BSCmp_op2_16, gen_16_cmp_BSCmp_op2_15, 
      gen_16_cmp_BSCmp_op2_14, gen_16_cmp_BSCmp_op2_13, 
      gen_16_cmp_BSCmp_op2_12, gen_16_cmp_BSCmp_op2_11, 
      gen_16_cmp_BSCmp_op2_10, gen_16_cmp_BSCmp_op2_9, 
      gen_16_cmp_BSCmp_op2_8, gen_16_cmp_BSCmp_op2_7, gen_16_cmp_BSCmp_op2_6, 
      gen_16_cmp_BSCmp_op2_5, gen_16_cmp_BSCmp_op2_4, gen_16_cmp_BSCmp_op2_3, 
      gen_16_cmp_BSCmp_op2_2, gen_16_cmp_BSCmp_op2_1, 
      gen_15_cmp_BSCmp_op2_16, gen_15_cmp_BSCmp_op2_15, 
      gen_15_cmp_BSCmp_op2_14, gen_15_cmp_BSCmp_op2_13, 
      gen_15_cmp_BSCmp_op2_12, gen_15_cmp_BSCmp_op2_11, 
      gen_15_cmp_BSCmp_op2_10, gen_15_cmp_BSCmp_op2_9, 
      gen_15_cmp_BSCmp_op2_8, gen_15_cmp_BSCmp_op2_7, gen_15_cmp_BSCmp_op2_6, 
      gen_15_cmp_BSCmp_op2_5, gen_15_cmp_BSCmp_op2_4, gen_15_cmp_BSCmp_op2_3, 
      gen_15_cmp_BSCmp_op2_2, gen_15_cmp_BSCmp_op2_1, 
      gen_14_cmp_BSCmp_op2_16, gen_14_cmp_BSCmp_op2_15, 
      gen_14_cmp_BSCmp_op2_14, gen_14_cmp_BSCmp_op2_13, 
      gen_14_cmp_BSCmp_op2_12, gen_14_cmp_BSCmp_op2_11, 
      gen_14_cmp_BSCmp_op2_10, gen_14_cmp_BSCmp_op2_9, 
      gen_14_cmp_BSCmp_op2_8, gen_14_cmp_BSCmp_op2_7, gen_14_cmp_BSCmp_op2_6, 
      gen_14_cmp_BSCmp_op2_5, gen_14_cmp_BSCmp_op2_4, gen_14_cmp_BSCmp_op2_3, 
      gen_14_cmp_BSCmp_op2_2, gen_14_cmp_BSCmp_op2_1, 
      gen_13_cmp_BSCmp_op2_16, gen_13_cmp_BSCmp_op2_15, 
      gen_13_cmp_BSCmp_op2_14, gen_13_cmp_BSCmp_op2_13, 
      gen_13_cmp_BSCmp_op2_12, gen_13_cmp_BSCmp_op2_11, 
      gen_13_cmp_BSCmp_op2_10, gen_13_cmp_BSCmp_op2_9, 
      gen_13_cmp_BSCmp_op2_8, gen_13_cmp_BSCmp_op2_7, gen_13_cmp_BSCmp_op2_6, 
      gen_13_cmp_BSCmp_op2_5, gen_13_cmp_BSCmp_op2_4, gen_13_cmp_BSCmp_op2_3, 
      gen_13_cmp_BSCmp_op2_2, gen_13_cmp_BSCmp_op2_1, 
      gen_12_cmp_BSCmp_op2_16, gen_12_cmp_BSCmp_op2_15, 
      gen_12_cmp_BSCmp_op2_14, gen_12_cmp_BSCmp_op2_13, 
      gen_12_cmp_BSCmp_op2_12, gen_12_cmp_BSCmp_op2_11, 
      gen_12_cmp_BSCmp_op2_10, gen_12_cmp_BSCmp_op2_9, 
      gen_12_cmp_BSCmp_op2_8, gen_12_cmp_BSCmp_op2_7, gen_12_cmp_BSCmp_op2_6, 
      gen_12_cmp_BSCmp_op2_5, gen_12_cmp_BSCmp_op2_4, gen_12_cmp_BSCmp_op2_3, 
      gen_12_cmp_BSCmp_op2_2, gen_12_cmp_BSCmp_op2_1, 
      gen_11_cmp_BSCmp_op2_16, gen_11_cmp_BSCmp_op2_15, 
      gen_11_cmp_BSCmp_op2_14, gen_11_cmp_BSCmp_op2_13, 
      gen_11_cmp_BSCmp_op2_12, gen_11_cmp_BSCmp_op2_11, 
      gen_11_cmp_BSCmp_op2_10, gen_11_cmp_BSCmp_op2_9, 
      gen_11_cmp_BSCmp_op2_8, gen_11_cmp_BSCmp_op2_7, gen_11_cmp_BSCmp_op2_6, 
      gen_11_cmp_BSCmp_op2_5, gen_11_cmp_BSCmp_op2_4, gen_11_cmp_BSCmp_op2_3, 
      gen_11_cmp_BSCmp_op2_2, gen_11_cmp_BSCmp_op2_1, 
      gen_10_cmp_BSCmp_op2_16, gen_10_cmp_BSCmp_op2_15, 
      gen_10_cmp_BSCmp_op2_14, gen_10_cmp_BSCmp_op2_13, 
      gen_10_cmp_BSCmp_op2_12, gen_10_cmp_BSCmp_op2_11, 
      gen_10_cmp_BSCmp_op2_10, gen_10_cmp_BSCmp_op2_9, 
      gen_10_cmp_BSCmp_op2_8, gen_10_cmp_BSCmp_op2_7, gen_10_cmp_BSCmp_op2_6, 
      gen_10_cmp_BSCmp_op2_5, gen_10_cmp_BSCmp_op2_4, gen_10_cmp_BSCmp_op2_3, 
      gen_10_cmp_BSCmp_op2_2, gen_10_cmp_BSCmp_op2_1, gen_9_cmp_BSCmp_op2_16, 
      gen_9_cmp_BSCmp_op2_15, gen_9_cmp_BSCmp_op2_14, gen_9_cmp_BSCmp_op2_13, 
      gen_9_cmp_BSCmp_op2_12, gen_9_cmp_BSCmp_op2_11, gen_9_cmp_BSCmp_op2_10, 
      gen_9_cmp_BSCmp_op2_9, gen_9_cmp_BSCmp_op2_8, gen_9_cmp_BSCmp_op2_7, 
      gen_9_cmp_BSCmp_op2_6, gen_9_cmp_BSCmp_op2_5, gen_9_cmp_BSCmp_op2_4, 
      gen_9_cmp_BSCmp_op2_3, gen_9_cmp_BSCmp_op2_2, gen_9_cmp_BSCmp_op2_1, 
      gen_8_cmp_BSCmp_op2_16, gen_8_cmp_BSCmp_op2_15, gen_8_cmp_BSCmp_op2_14, 
      gen_8_cmp_BSCmp_op2_13, gen_8_cmp_BSCmp_op2_12, gen_8_cmp_BSCmp_op2_11, 
      gen_8_cmp_BSCmp_op2_10, gen_8_cmp_BSCmp_op2_9, gen_8_cmp_BSCmp_op2_8, 
      gen_8_cmp_BSCmp_op2_7, gen_8_cmp_BSCmp_op2_6, gen_8_cmp_BSCmp_op2_5, 
      gen_8_cmp_BSCmp_op2_4, gen_8_cmp_BSCmp_op2_3, gen_8_cmp_BSCmp_op2_2, 
      gen_8_cmp_BSCmp_op2_1, gen_7_cmp_BSCmp_op2_16, gen_7_cmp_BSCmp_op2_15, 
      gen_7_cmp_BSCmp_op2_14, gen_7_cmp_BSCmp_op2_13, gen_7_cmp_BSCmp_op2_12, 
      gen_7_cmp_BSCmp_op2_11, gen_7_cmp_BSCmp_op2_10, gen_7_cmp_BSCmp_op2_9, 
      gen_7_cmp_BSCmp_op2_8, gen_7_cmp_BSCmp_op2_7, gen_7_cmp_BSCmp_op2_6, 
      gen_7_cmp_BSCmp_op2_5, gen_7_cmp_BSCmp_op2_4, gen_7_cmp_BSCmp_op2_3, 
      gen_7_cmp_BSCmp_op2_2, gen_7_cmp_BSCmp_op2_1, gen_6_cmp_BSCmp_op2_16, 
      gen_6_cmp_BSCmp_op2_15, gen_6_cmp_BSCmp_op2_14, gen_6_cmp_BSCmp_op2_13, 
      gen_6_cmp_BSCmp_op2_12, gen_6_cmp_BSCmp_op2_11, gen_6_cmp_BSCmp_op2_10, 
      gen_6_cmp_BSCmp_op2_9, gen_6_cmp_BSCmp_op2_8, gen_6_cmp_BSCmp_op2_7, 
      gen_6_cmp_BSCmp_op2_6, gen_6_cmp_BSCmp_op2_5, gen_6_cmp_BSCmp_op2_4, 
      gen_6_cmp_BSCmp_op2_3, gen_6_cmp_BSCmp_op2_2, gen_6_cmp_BSCmp_op2_1, 
      gen_5_cmp_BSCmp_op2_16, gen_5_cmp_BSCmp_op2_15, gen_5_cmp_BSCmp_op2_14, 
      gen_5_cmp_BSCmp_op2_13, gen_5_cmp_BSCmp_op2_12, gen_5_cmp_BSCmp_op2_11, 
      gen_5_cmp_BSCmp_op2_10, gen_5_cmp_BSCmp_op2_9, gen_5_cmp_BSCmp_op2_8, 
      gen_5_cmp_BSCmp_op2_7, gen_5_cmp_BSCmp_op2_6, gen_5_cmp_BSCmp_op2_5, 
      gen_5_cmp_BSCmp_op2_4, gen_5_cmp_BSCmp_op2_3, gen_5_cmp_BSCmp_op2_2, 
      gen_5_cmp_BSCmp_op2_1, gen_4_cmp_BSCmp_op2_16, gen_4_cmp_BSCmp_op2_15, 
      gen_4_cmp_BSCmp_op2_14, gen_4_cmp_BSCmp_op2_13, gen_4_cmp_BSCmp_op2_12, 
      gen_4_cmp_BSCmp_op2_11, gen_4_cmp_BSCmp_op2_10, gen_4_cmp_BSCmp_op2_9, 
      gen_4_cmp_BSCmp_op2_8, gen_4_cmp_BSCmp_op2_7, gen_4_cmp_BSCmp_op2_6, 
      gen_4_cmp_BSCmp_op2_5, gen_4_cmp_BSCmp_op2_4, gen_4_cmp_BSCmp_op2_3, 
      gen_4_cmp_BSCmp_op2_2, gen_4_cmp_BSCmp_op2_1, gen_3_cmp_BSCmp_op2_16, 
      gen_3_cmp_BSCmp_op2_15, gen_3_cmp_BSCmp_op2_14, gen_3_cmp_BSCmp_op2_13, 
      gen_3_cmp_BSCmp_op2_12, gen_3_cmp_BSCmp_op2_11, gen_3_cmp_BSCmp_op2_10, 
      gen_3_cmp_BSCmp_op2_9, gen_3_cmp_BSCmp_op2_8, gen_3_cmp_BSCmp_op2_7, 
      gen_3_cmp_BSCmp_op2_6, gen_3_cmp_BSCmp_op2_5, gen_3_cmp_BSCmp_op2_4, 
      gen_3_cmp_BSCmp_op2_3, gen_3_cmp_BSCmp_op2_2, gen_3_cmp_BSCmp_op2_1, 
      gen_2_cmp_BSCmp_op2_16, gen_2_cmp_BSCmp_op2_15, gen_2_cmp_BSCmp_op2_14, 
      gen_2_cmp_BSCmp_op2_13, gen_2_cmp_BSCmp_op2_12, gen_2_cmp_BSCmp_op2_11, 
      gen_2_cmp_BSCmp_op2_10, gen_2_cmp_BSCmp_op2_9, gen_2_cmp_BSCmp_op2_8, 
      gen_2_cmp_BSCmp_op2_7, gen_2_cmp_BSCmp_op2_6, gen_2_cmp_BSCmp_op2_5, 
      gen_2_cmp_BSCmp_op2_4, gen_2_cmp_BSCmp_op2_3, gen_2_cmp_BSCmp_op2_2, 
      gen_2_cmp_BSCmp_op2_1, gen_1_cmp_BSCmp_op2_16, gen_1_cmp_BSCmp_op2_15, 
      gen_1_cmp_BSCmp_op2_14, gen_1_cmp_BSCmp_op2_13, gen_1_cmp_BSCmp_op2_12, 
      gen_1_cmp_BSCmp_op2_11, gen_1_cmp_BSCmp_op2_10, gen_1_cmp_BSCmp_op2_9, 
      gen_1_cmp_BSCmp_op2_8, gen_1_cmp_BSCmp_op2_7, gen_1_cmp_BSCmp_op2_6, 
      gen_1_cmp_BSCmp_op2_5, gen_1_cmp_BSCmp_op2_4, gen_1_cmp_BSCmp_op2_3, 
      gen_1_cmp_BSCmp_op2_2, gen_1_cmp_BSCmp_op2_1, gen_0_cmp_BSCmp_op2_16, 
      gen_0_cmp_BSCmp_op2_15, gen_0_cmp_BSCmp_op2_14, gen_0_cmp_BSCmp_op2_13, 
      gen_0_cmp_BSCmp_op2_12, gen_0_cmp_BSCmp_op2_11, gen_0_cmp_BSCmp_op2_10, 
      gen_0_cmp_BSCmp_op2_9, gen_0_cmp_BSCmp_op2_8, gen_0_cmp_BSCmp_op2_7, 
      gen_0_cmp_BSCmp_op2_6, gen_0_cmp_BSCmp_op2_5, gen_0_cmp_BSCmp_op2_4, 
      gen_0_cmp_BSCmp_op2_3, gen_0_cmp_BSCmp_op2_2, gen_0_cmp_BSCmp_op2_1, 
      gen_24_cmp_pInit_32, nx6, gen_0_cmp_mReg_0, nx26, nx34, 
      gen_0_cmp_mReg_1, nx46, nx48, nx58, nx62, gen_0_cmp_mReg_2, nx74, nx76, 
      nx80, nx84, gen_0_cmp_mReg_3, nx96, nx98, nx102, nx106, 
      gen_0_cmp_mReg_4, nx118, nx120, nx124, nx128, gen_0_cmp_mReg_5, nx140, 
      nx142, nx146, nx150, gen_0_cmp_mReg_6, nx162, nx164, nx168, nx172, 
      gen_0_cmp_mReg_7, nx184, nx186, nx190, nx194, gen_0_cmp_mReg_8, nx206, 
      nx208, nx212, nx216, gen_0_cmp_mReg_9, nx228, nx230, nx234, nx238, 
      gen_0_cmp_mReg_10, nx250, nx252, nx256, nx260, gen_0_cmp_mReg_11, 
      nx272, nx274, nx278, nx282, gen_0_cmp_mReg_12, nx294, nx296, nx300, 
      nx304, gen_0_cmp_mReg_13, nx316, nx318, nx322, nx326, 
      gen_0_cmp_mReg_14, nx338, nx340, nx344, nx348, gen_0_cmp_mReg_15, 
      nx360, nx362, nx366, nx370, nx376, nx380, nx392, gen_1_cmp_mReg_0, 
      nx412, nx420, gen_1_cmp_mReg_1, nx432, nx434, nx444, nx448, 
      gen_1_cmp_mReg_2, nx460, nx462, nx466, nx470, gen_1_cmp_mReg_3, nx482, 
      nx484, nx488, nx492, gen_1_cmp_mReg_4, nx504, nx506, nx510, nx514, 
      gen_1_cmp_mReg_5, nx526, nx528, nx532, nx536, gen_1_cmp_mReg_6, nx548, 
      nx550, nx554, nx558, gen_1_cmp_mReg_7, nx570, nx572, nx576, nx580, 
      gen_1_cmp_mReg_8, nx592, nx594, nx598, nx602, gen_1_cmp_mReg_9, nx614, 
      nx616, nx620, nx624, gen_1_cmp_mReg_10, nx636, nx638, nx642, nx646, 
      gen_1_cmp_mReg_11, nx658, nx660, nx664, nx668, gen_1_cmp_mReg_12, 
      nx680, nx682, nx686, nx690, gen_1_cmp_mReg_13, nx702, nx704, nx708, 
      nx712, gen_1_cmp_mReg_14, nx724, nx726, nx730, nx734, 
      gen_1_cmp_mReg_15, nx746, nx748, nx752, nx756, nx762, nx766, nx778, 
      gen_2_cmp_mReg_0, nx798, nx806, gen_2_cmp_mReg_1, nx818, nx820, nx830, 
      nx834, gen_2_cmp_mReg_2, nx846, nx848, nx852, nx856, gen_2_cmp_mReg_3, 
      nx868, nx870, nx874, nx878, gen_2_cmp_mReg_4, nx890, nx892, nx896, 
      nx900, gen_2_cmp_mReg_5, nx912, nx914, nx918, nx922, gen_2_cmp_mReg_6, 
      nx934, nx936, nx940, nx944, gen_2_cmp_mReg_7, nx956, nx958, nx962, 
      nx966, gen_2_cmp_mReg_8, nx978, nx980, nx984, nx988, gen_2_cmp_mReg_9, 
      nx1000, nx1002, nx1006, nx1010, gen_2_cmp_mReg_10, nx1022, nx1024, 
      nx1028, nx1032, gen_2_cmp_mReg_11, nx1044, nx1046, nx1050, nx1054, 
      gen_2_cmp_mReg_12, nx1066, nx1068, nx1072, nx1076, gen_2_cmp_mReg_13, 
      nx1088, nx1090, nx1094, nx1098, gen_2_cmp_mReg_14, nx1110, nx1112, 
      nx1116, nx1120, gen_2_cmp_mReg_15, nx1132, nx1134, nx1138, nx1142, 
      nx1148, nx1152, nx1164, gen_3_cmp_mReg_0, nx1184, nx1192, 
      gen_3_cmp_mReg_1, nx1204, nx1206, nx1216, nx1220, gen_3_cmp_mReg_2, 
      nx1232, nx1234, nx1238, nx1242, gen_3_cmp_mReg_3, nx1254, nx1256, 
      nx1260, nx1264, gen_3_cmp_mReg_4, nx1276, nx1278, nx1282, nx1286, 
      gen_3_cmp_mReg_5, nx1298, nx1300, nx1304, nx1308, gen_3_cmp_mReg_6, 
      nx1320, nx1322, nx1326, nx1330, gen_3_cmp_mReg_7, nx1342, nx1344, 
      nx1348, nx1352, gen_3_cmp_mReg_8, nx1364, nx1366, nx1370, nx1374, 
      gen_3_cmp_mReg_9, nx1386, nx1388, nx1392, nx1396, gen_3_cmp_mReg_10, 
      nx1408, nx1410, nx1414, nx1418, gen_3_cmp_mReg_11, nx1430, nx1432, 
      nx1436, nx1440, gen_3_cmp_mReg_12, nx1452, nx1454, nx1458, nx1462, 
      gen_3_cmp_mReg_13, nx1474, nx1476, nx1480, nx1484, gen_3_cmp_mReg_14, 
      nx1496, nx1498, nx1502, nx1506, gen_3_cmp_mReg_15, nx1518, nx1520, 
      nx1524, nx1528, nx1534, nx1538, nx1550, gen_4_cmp_mReg_0, nx1570, 
      nx1578, gen_4_cmp_mReg_1, nx1590, nx1592, nx1602, nx1606, 
      gen_4_cmp_mReg_2, nx1618, nx1620, nx1624, nx1628, gen_4_cmp_mReg_3, 
      nx1640, nx1642, nx1646, nx1650, gen_4_cmp_mReg_4, nx1662, nx1664, 
      nx1668, nx1672, gen_4_cmp_mReg_5, nx1684, nx1686, nx1690, nx1694, 
      gen_4_cmp_mReg_6, nx1706, nx1708, nx1712, nx1716, gen_4_cmp_mReg_7, 
      nx1728, nx1730, nx1734, nx1738, gen_4_cmp_mReg_8, nx1750, nx1752, 
      nx1756, nx1760, gen_4_cmp_mReg_9, nx1772, nx1774, nx1778, nx1782, 
      gen_4_cmp_mReg_10, nx1794, nx1796, nx1800, nx1804, gen_4_cmp_mReg_11, 
      nx1816, nx1818, nx1822, nx1826, gen_4_cmp_mReg_12, nx1838, nx1840, 
      nx1844, nx1848, gen_4_cmp_mReg_13, nx1860, nx1862, nx1866, nx1870, 
      gen_4_cmp_mReg_14, nx1882, nx1884, nx1888, nx1892, gen_4_cmp_mReg_15, 
      nx1904, nx1906, nx1910, nx1914, nx1920, nx1924, nx1936, 
      gen_5_cmp_mReg_0, nx1956, nx1964, gen_5_cmp_mReg_1, nx1976, nx1978, 
      nx1988, nx1992, gen_5_cmp_mReg_2, nx2004, nx2006, nx2010, nx2014, 
      gen_5_cmp_mReg_3, nx2026, nx2028, nx2032, nx2036, gen_5_cmp_mReg_4, 
      nx2048, nx2050, nx2054, nx2058, gen_5_cmp_mReg_5, nx2070, nx2072, 
      nx2076, nx2080, gen_5_cmp_mReg_6, nx2092, nx2094, nx2098, nx2102, 
      gen_5_cmp_mReg_7, nx2114, nx2116, nx2120, nx2124, gen_5_cmp_mReg_8, 
      nx2136, nx2138, nx2142, nx2146, gen_5_cmp_mReg_9, nx2158, nx2160, 
      nx2164, nx2168, gen_5_cmp_mReg_10, nx2180, nx2182, nx2186, nx2190, 
      gen_5_cmp_mReg_11, nx2202, nx2204, nx2208, nx2212, gen_5_cmp_mReg_12, 
      nx2224, nx2226, nx2230, nx2234, gen_5_cmp_mReg_13, nx2246, nx2248, 
      nx2252, nx2256, gen_5_cmp_mReg_14, nx2268, nx2270, nx2274, nx2278, 
      gen_5_cmp_mReg_15, nx2290, nx2292, nx2296, nx2300, nx2306, nx2310, 
      nx2322, gen_6_cmp_mReg_0, nx2342, nx2350, gen_6_cmp_mReg_1, nx2362, 
      nx2364, nx2374, nx2378, gen_6_cmp_mReg_2, nx2390, nx2392, nx2396, 
      nx2400, gen_6_cmp_mReg_3, nx2412, nx2414, nx2418, nx2422, 
      gen_6_cmp_mReg_4, nx2434, nx2436, nx2440, nx2444, gen_6_cmp_mReg_5, 
      nx2456, nx2458, nx2462, nx2466, gen_6_cmp_mReg_6, nx2478, nx2480, 
      nx2484, nx2488, gen_6_cmp_mReg_7, nx2500, nx2502, nx2506, nx2510, 
      gen_6_cmp_mReg_8, nx2522, nx2524, nx2528, nx2532, gen_6_cmp_mReg_9, 
      nx2544, nx2546, nx2550, nx2554, gen_6_cmp_mReg_10, nx2566, nx2568, 
      nx2572, nx2576, gen_6_cmp_mReg_11, nx2588, nx2590, nx2594, nx2598, 
      gen_6_cmp_mReg_12, nx2610, nx2612, nx2616, nx2620, gen_6_cmp_mReg_13, 
      nx2632, nx2634, nx2638, nx2642, gen_6_cmp_mReg_14, nx2654, nx2656, 
      nx2660, nx2664, gen_6_cmp_mReg_15, nx2676, nx2678, nx2682, nx2686, 
      nx2692, nx2696, nx2708, gen_7_cmp_mReg_0, nx2728, nx2736, 
      gen_7_cmp_mReg_1, nx2748, nx2750, nx2760, nx2764, gen_7_cmp_mReg_2, 
      nx2776, nx2778, nx2782, nx2786, gen_7_cmp_mReg_3, nx2798, nx2800, 
      nx2804, nx2808, gen_7_cmp_mReg_4, nx2820, nx2822, nx2826, nx2830, 
      gen_7_cmp_mReg_5, nx2842, nx2844, nx2848, nx2852, gen_7_cmp_mReg_6, 
      nx2864, nx2866, nx2870, nx2874, gen_7_cmp_mReg_7, nx2886, nx2888, 
      nx2892, nx2896, gen_7_cmp_mReg_8, nx2908, nx2910, nx2914, nx2918, 
      gen_7_cmp_mReg_9, nx2930, nx2932, nx2936, nx2940, gen_7_cmp_mReg_10, 
      nx2952, nx2954, nx2958, nx2962, gen_7_cmp_mReg_11, nx2974, nx2976, 
      nx2980, nx2984, gen_7_cmp_mReg_12, nx2996, nx2998, nx3002, nx3006, 
      gen_7_cmp_mReg_13, nx3018, nx3020, nx3024, nx3028, gen_7_cmp_mReg_14, 
      nx3040, nx3042, nx3046, nx3050, gen_7_cmp_mReg_15, nx3062, nx3064, 
      nx3068, nx3072, nx3078, nx3082, nx3094, gen_8_cmp_mReg_0, nx3114, 
      nx3122, gen_8_cmp_mReg_1, nx3134, nx3136, nx3146, nx3150, 
      gen_8_cmp_mReg_2, nx3162, nx3164, nx3168, nx3172, gen_8_cmp_mReg_3, 
      nx3184, nx3186, nx3190, nx3194, gen_8_cmp_mReg_4, nx3206, nx3208, 
      nx3212, nx3216, gen_8_cmp_mReg_5, nx3228, nx3230, nx3234, nx3238, 
      gen_8_cmp_mReg_6, nx3250, nx3252, nx3256, nx3260, gen_8_cmp_mReg_7, 
      nx3272, nx3274, nx3278, nx3282, gen_8_cmp_mReg_8, nx3294, nx3296, 
      nx3300, nx3304, gen_8_cmp_mReg_9, nx3316, nx3318, nx3322, nx3326, 
      gen_8_cmp_mReg_10, nx3338, nx3340, nx3344, nx3348, gen_8_cmp_mReg_11, 
      nx3360, nx3362, nx3366, nx3370, gen_8_cmp_mReg_12, nx3382, nx3384, 
      nx3388, nx3392, gen_8_cmp_mReg_13, nx3404, nx3406, nx3410, nx3414, 
      gen_8_cmp_mReg_14, nx3426, nx3428, nx3432, nx3436, gen_8_cmp_mReg_15, 
      nx3448, nx3450, nx3454, nx3458, nx3464, nx3468, nx3480, 
      gen_9_cmp_mReg_0, nx3500, nx3508, gen_9_cmp_mReg_1, nx3520, nx3522, 
      nx3532, nx3536, gen_9_cmp_mReg_2, nx3548, nx3550, nx3554, nx3558, 
      gen_9_cmp_mReg_3, nx3570, nx3572, nx3576, nx3580, gen_9_cmp_mReg_4, 
      nx3592, nx3594, nx3598, nx3602, gen_9_cmp_mReg_5, nx3614, nx3616, 
      nx3620, nx3624, gen_9_cmp_mReg_6, nx3636, nx3638, nx3642, nx3646, 
      gen_9_cmp_mReg_7, nx3658, nx3660, nx3664, nx3668, gen_9_cmp_mReg_8, 
      nx3680, nx3682, nx3686, nx3690, gen_9_cmp_mReg_9, nx3702, nx3704, 
      nx3708, nx3712, gen_9_cmp_mReg_10, nx3724, nx3726, nx3730, nx3734, 
      gen_9_cmp_mReg_11, nx3746, nx3748, nx3752, nx3756, gen_9_cmp_mReg_12, 
      nx3768, nx3770, nx3774, nx3778, gen_9_cmp_mReg_13, nx3790, nx3792, 
      nx3796, nx3800, gen_9_cmp_mReg_14, nx3812, nx3814, nx3818, nx3822, 
      gen_9_cmp_mReg_15, nx3834, nx3836, nx3840, nx3844, nx3850, nx3854, 
      nx3866, gen_10_cmp_mReg_0, nx3886, nx3894, gen_10_cmp_mReg_1, nx3906, 
      nx3908, nx3918, nx3922, gen_10_cmp_mReg_2, nx3934, nx3936, nx3940, 
      nx3944, gen_10_cmp_mReg_3, nx3956, nx3958, nx3962, nx3966, 
      gen_10_cmp_mReg_4, nx3978, nx3980, nx3984, nx3988, gen_10_cmp_mReg_5, 
      nx4000, nx4002, nx4006, nx4010, gen_10_cmp_mReg_6, nx4022, nx4024, 
      nx4028, nx4032, gen_10_cmp_mReg_7, nx4044, nx4046, nx4050, nx4054, 
      gen_10_cmp_mReg_8, nx4066, nx4068, nx4072, nx4076, gen_10_cmp_mReg_9, 
      nx4088, nx4090, nx4094, nx4098, gen_10_cmp_mReg_10, nx4110, nx4112, 
      nx4116, nx4120, gen_10_cmp_mReg_11, nx4132, nx4134, nx4138, nx4142, 
      gen_10_cmp_mReg_12, nx4154, nx4156, nx4160, nx4164, gen_10_cmp_mReg_13, 
      nx4176, nx4178, nx4182, nx4186, gen_10_cmp_mReg_14, nx4198, nx4200, 
      nx4204, nx4208, gen_10_cmp_mReg_15, nx4220, nx4222, nx4226, nx4230, 
      nx4236, nx4240, nx4252, gen_11_cmp_mReg_0, nx4272, nx4280, 
      gen_11_cmp_mReg_1, nx4292, nx4294, nx4304, nx4308, gen_11_cmp_mReg_2, 
      nx4320, nx4322, nx4326, nx4330, gen_11_cmp_mReg_3, nx4342, nx4344, 
      nx4348, nx4352, gen_11_cmp_mReg_4, nx4364, nx4366, nx4370, nx4374, 
      gen_11_cmp_mReg_5, nx4386, nx4388, nx4392, nx4396, gen_11_cmp_mReg_6, 
      nx4408, nx4410, nx4414, nx4418, gen_11_cmp_mReg_7, nx4430, nx4432, 
      nx4436, nx4440, gen_11_cmp_mReg_8, nx4452, nx4454, nx4458, nx4462, 
      gen_11_cmp_mReg_9, nx4474, nx4476, nx4480, nx4484, gen_11_cmp_mReg_10, 
      nx4496, nx4498, nx4502, nx4506, gen_11_cmp_mReg_11, nx4518, nx4520, 
      nx4524, nx4528, gen_11_cmp_mReg_12, nx4540, nx4542, nx4546, nx4550, 
      gen_11_cmp_mReg_13, nx4562, nx4564, nx4568, nx4572, gen_11_cmp_mReg_14, 
      nx4584, nx4586, nx4590, nx4594, gen_11_cmp_mReg_15, nx4606, nx4608, 
      nx4612, nx4616, nx4622, nx4626, nx4638, gen_12_cmp_mReg_0, nx4658, 
      nx4666, gen_12_cmp_mReg_1, nx4678, nx4680, nx4690, nx4694, 
      gen_12_cmp_mReg_2, nx4706, nx4708, nx4712, nx4716, gen_12_cmp_mReg_3, 
      nx4728, nx4730, nx4734, nx4738, gen_12_cmp_mReg_4, nx4750, nx4752, 
      nx4756, nx4760, gen_12_cmp_mReg_5, nx4772, nx4774, nx4778, nx4782, 
      gen_12_cmp_mReg_6, nx4794, nx4796, nx4800, nx4804, gen_12_cmp_mReg_7, 
      nx4816, nx4818, nx4822, nx4826, gen_12_cmp_mReg_8, nx4838, nx4840, 
      nx4844, nx4848, gen_12_cmp_mReg_9, nx4860, nx4862, nx4866, nx4870, 
      gen_12_cmp_mReg_10, nx4882, nx4884, nx4888, nx4892, gen_12_cmp_mReg_11, 
      nx4904, nx4906, nx4910, nx4914, gen_12_cmp_mReg_12, nx4926, nx4928, 
      nx4932, nx4936, gen_12_cmp_mReg_13, nx4948, nx4950, nx4954, nx4958, 
      gen_12_cmp_mReg_14, nx4970, nx4972, nx4976, nx4980, gen_12_cmp_mReg_15, 
      nx4992, nx4994, nx4998, nx5002, nx5008, nx5012, nx5024, 
      gen_13_cmp_mReg_0, nx5044, nx5052, gen_13_cmp_mReg_1, nx5064, nx5066, 
      nx5076, nx5080, gen_13_cmp_mReg_2, nx5092, nx5094, nx5098, nx5102, 
      gen_13_cmp_mReg_3, nx5114, nx5116, nx5120, nx5124, gen_13_cmp_mReg_4, 
      nx5136, nx5138, nx5142, nx5146, gen_13_cmp_mReg_5, nx5158, nx5160, 
      nx5164, nx5168, gen_13_cmp_mReg_6, nx5180, nx5182, nx5186, nx5190, 
      gen_13_cmp_mReg_7, nx5202, nx5204, nx5208, nx5212, gen_13_cmp_mReg_8, 
      nx5224, nx5226, nx5230, nx5234, gen_13_cmp_mReg_9, nx5246, nx5248, 
      nx5252, nx5256, gen_13_cmp_mReg_10, nx5268, nx5270, nx5274, nx5278, 
      gen_13_cmp_mReg_11, nx5290, nx5292, nx5296, nx5300, gen_13_cmp_mReg_12, 
      nx5312, nx5314, nx5318, nx5322, gen_13_cmp_mReg_13, nx5334, nx5336, 
      nx5340, nx5344, gen_13_cmp_mReg_14, nx5356, nx5358, nx5362, nx5366, 
      gen_13_cmp_mReg_15, nx5378, nx5380, nx5384, nx5388, nx5394, nx5398, 
      nx5410, gen_14_cmp_mReg_0, nx5430, nx5438, gen_14_cmp_mReg_1, nx5450, 
      nx5452, nx5462, nx5466, gen_14_cmp_mReg_2, nx5478, nx5480, nx5484, 
      nx5488, gen_14_cmp_mReg_3, nx5500, nx5502, nx5506, nx5510, 
      gen_14_cmp_mReg_4, nx5522, nx5524, nx5528, nx5532, gen_14_cmp_mReg_5, 
      nx5544, nx5546, nx5550, nx5554, gen_14_cmp_mReg_6, nx5566, nx5568, 
      nx5572, nx5576, gen_14_cmp_mReg_7, nx5588, nx5590, nx5594, nx5598, 
      gen_14_cmp_mReg_8, nx5610, nx5612, nx5616, nx5620, gen_14_cmp_mReg_9, 
      nx5632, nx5634, nx5638, nx5642, gen_14_cmp_mReg_10, nx5654, nx5656, 
      nx5660, nx5664, gen_14_cmp_mReg_11, nx5676, nx5678, nx5682, nx5686, 
      gen_14_cmp_mReg_12, nx5698, nx5700, nx5704, nx5708, gen_14_cmp_mReg_13, 
      nx5720, nx5722, nx5726, nx5730, gen_14_cmp_mReg_14, nx5742, nx5744, 
      nx5748, nx5752, gen_14_cmp_mReg_15, nx5764, nx5766, nx5770, nx5774, 
      nx5780, nx5784, nx5796, gen_15_cmp_mReg_0, nx5816, nx5824, 
      gen_15_cmp_mReg_1, nx5836, nx5838, nx5848, nx5852, gen_15_cmp_mReg_2, 
      nx5864, nx5866, nx5870, nx5874, gen_15_cmp_mReg_3, nx5886, nx5888, 
      nx5892, nx5896, gen_15_cmp_mReg_4, nx5908, nx5910, nx5914, nx5918, 
      gen_15_cmp_mReg_5, nx5930, nx5932, nx5936, nx5940, gen_15_cmp_mReg_6, 
      nx5952, nx5954, nx5958, nx5962, gen_15_cmp_mReg_7, nx5974, nx5976, 
      nx5980, nx5984, gen_15_cmp_mReg_8, nx5996, nx5998, nx6002, nx6006, 
      gen_15_cmp_mReg_9, nx6018, nx6020, nx6024, nx6028, gen_15_cmp_mReg_10, 
      nx6040, nx6042, nx6046, nx6050, gen_15_cmp_mReg_11, nx6062, nx6064, 
      nx6068, nx6072, gen_15_cmp_mReg_12, nx6084, nx6086, nx6090, nx6094, 
      gen_15_cmp_mReg_13, nx6106, nx6108, nx6112, nx6116, gen_15_cmp_mReg_14, 
      nx6128, nx6130, nx6134, nx6138, gen_15_cmp_mReg_15, nx6150, nx6152, 
      nx6156, nx6160, nx6166, nx6170, nx6182, gen_16_cmp_mReg_0, nx6202, 
      nx6210, gen_16_cmp_mReg_1, nx6222, nx6224, nx6234, nx6238, 
      gen_16_cmp_mReg_2, nx6250, nx6252, nx6256, nx6260, gen_16_cmp_mReg_3, 
      nx6272, nx6274, nx6278, nx6282, gen_16_cmp_mReg_4, nx6294, nx6296, 
      nx6300, nx6304, gen_16_cmp_mReg_5, nx6316, nx6318, nx6322, nx6326, 
      gen_16_cmp_mReg_6, nx6338, nx6340, nx6344, nx6348, gen_16_cmp_mReg_7, 
      nx6360, nx6362, nx6366, nx6370, gen_16_cmp_mReg_8, nx6382, nx6384, 
      nx6388, nx6392, gen_16_cmp_mReg_9, nx6404, nx6406, nx6410, nx6414, 
      gen_16_cmp_mReg_10, nx6426, nx6428, nx6432, nx6436, gen_16_cmp_mReg_11, 
      nx6448, nx6450, nx6454, nx6458, gen_16_cmp_mReg_12, nx6470, nx6472, 
      nx6476, nx6480, gen_16_cmp_mReg_13, nx6492, nx6494, nx6498, nx6502, 
      gen_16_cmp_mReg_14, nx6514, nx6516, nx6520, nx6524, gen_16_cmp_mReg_15, 
      nx6536, nx6538, nx6542, nx6546, nx6552, nx6556, nx6568, 
      gen_17_cmp_mReg_0, nx6588, nx6596, gen_17_cmp_mReg_1, nx6608, nx6610, 
      nx6620, nx6624, gen_17_cmp_mReg_2, nx6636, nx6638, nx6642, nx6646, 
      gen_17_cmp_mReg_3, nx6658, nx6660, nx6664, nx6668, gen_17_cmp_mReg_4, 
      nx6680, nx6682, nx6686, nx6690, gen_17_cmp_mReg_5, nx6702, nx6704, 
      nx6708, nx6712, gen_17_cmp_mReg_6, nx6724, nx6726, nx6730, nx6734, 
      gen_17_cmp_mReg_7, nx6746, nx6748, nx6752, nx6756, gen_17_cmp_mReg_8, 
      nx6768, nx6770, nx6774, nx6778, gen_17_cmp_mReg_9, nx6790, nx6792, 
      nx6796, nx6800, gen_17_cmp_mReg_10, nx6812, nx6814, nx6818, nx6822, 
      gen_17_cmp_mReg_11, nx6834, nx6836, nx6840, nx6844, gen_17_cmp_mReg_12, 
      nx6856, nx6858, nx6862, nx6866, gen_17_cmp_mReg_13, nx6878, nx6880, 
      nx6884, nx6888, gen_17_cmp_mReg_14, nx6900, nx6902, nx6906, nx6910, 
      gen_17_cmp_mReg_15, nx6922, nx6924, nx6928, nx6932, nx6938, nx6942, 
      nx6954, gen_18_cmp_mReg_0, nx6974, nx6982, gen_18_cmp_mReg_1, nx6994, 
      nx6996, nx7006, nx7010, gen_18_cmp_mReg_2, nx7022, nx7024, nx7028, 
      nx7032, gen_18_cmp_mReg_3, nx7044, nx7046, nx7050, nx7054, 
      gen_18_cmp_mReg_4, nx7066, nx7068, nx7072, nx7076, gen_18_cmp_mReg_5, 
      nx7088, nx7090, nx7094, nx7098, gen_18_cmp_mReg_6, nx7110, nx7112, 
      nx7116, nx7120, gen_18_cmp_mReg_7, nx7132, nx7134, nx7138, nx7142, 
      gen_18_cmp_mReg_8, nx7154, nx7156, nx7160, nx7164, gen_18_cmp_mReg_9, 
      nx7176, nx7178, nx7182, nx7186, gen_18_cmp_mReg_10, nx7198, nx7200, 
      nx7204, nx7208, gen_18_cmp_mReg_11, nx7220, nx7222, nx7226, nx7230, 
      gen_18_cmp_mReg_12, nx7242, nx7244, nx7248, nx7252, gen_18_cmp_mReg_13, 
      nx7264, nx7266, nx7270, nx7274, gen_18_cmp_mReg_14, nx7286, nx7288, 
      nx7292, nx7296, gen_18_cmp_mReg_15, nx7308, nx7310, nx7314, nx7318, 
      nx7324, nx7328, nx7340, gen_19_cmp_mReg_0, nx7360, nx7368, 
      gen_19_cmp_mReg_1, nx7380, nx7382, nx7392, nx7396, gen_19_cmp_mReg_2, 
      nx7408, nx7410, nx7414, nx7418, gen_19_cmp_mReg_3, nx7430, nx7432, 
      nx7436, nx7440, gen_19_cmp_mReg_4, nx7452, nx7454, nx7458, nx7462, 
      gen_19_cmp_mReg_5, nx7474, nx7476, nx7480, nx7484, gen_19_cmp_mReg_6, 
      nx7496, nx7498, nx7502, nx7506, gen_19_cmp_mReg_7, nx7518, nx7520, 
      nx7524, nx7528, gen_19_cmp_mReg_8, nx7540, nx7542, nx7546, nx7550, 
      gen_19_cmp_mReg_9, nx7562, nx7564, nx7568, nx7572, gen_19_cmp_mReg_10, 
      nx7584, nx7586, nx7590, nx7594, gen_19_cmp_mReg_11, nx7606, nx7608, 
      nx7612, nx7616, gen_19_cmp_mReg_12, nx7628, nx7630, nx7634, nx7638, 
      gen_19_cmp_mReg_13, nx7650, nx7652, nx7656, nx7660, gen_19_cmp_mReg_14, 
      nx7672, nx7674, nx7678, nx7682, gen_19_cmp_mReg_15, nx7694, nx7696, 
      nx7700, nx7704, nx7710, nx7714, nx7726, gen_20_cmp_mReg_0, nx7746, 
      nx7754, gen_20_cmp_mReg_1, nx7766, nx7768, nx7778, nx7782, 
      gen_20_cmp_mReg_2, nx7794, nx7796, nx7800, nx7804, gen_20_cmp_mReg_3, 
      nx7816, nx7818, nx7822, nx7826, gen_20_cmp_mReg_4, nx7838, nx7840, 
      nx7844, nx7848, gen_20_cmp_mReg_5, nx7860, nx7862, nx7866, nx7870, 
      gen_20_cmp_mReg_6, nx7882, nx7884, nx7888, nx7892, gen_20_cmp_mReg_7, 
      nx7904, nx7906, nx7910, nx7914, gen_20_cmp_mReg_8, nx7926, nx7928, 
      nx7932, nx7936, gen_20_cmp_mReg_9, nx7948, nx7950, nx7954, nx7958, 
      gen_20_cmp_mReg_10, nx7970, nx7972, nx7976, nx7980, gen_20_cmp_mReg_11, 
      nx7992, nx7994, nx7998, nx8002, gen_20_cmp_mReg_12, nx8014, nx8016, 
      nx8020, nx8024, gen_20_cmp_mReg_13, nx8036, nx8038, nx8042, nx8046, 
      gen_20_cmp_mReg_14, nx8058, nx8060, nx8064, nx8068, gen_20_cmp_mReg_15, 
      nx8080, nx8082, nx8086, nx8090, nx8096, nx8100, nx8112, 
      gen_21_cmp_mReg_0, nx8132, nx8140, gen_21_cmp_mReg_1, nx8152, nx8154, 
      nx8164, nx8168, gen_21_cmp_mReg_2, nx8180, nx8182, nx8186, nx8190, 
      gen_21_cmp_mReg_3, nx8202, nx8204, nx8208, nx8212, gen_21_cmp_mReg_4, 
      nx8224, nx8226, nx8230, nx8234, gen_21_cmp_mReg_5, nx8246, nx8248, 
      nx8252, nx8256, gen_21_cmp_mReg_6, nx8268, nx8270, nx8274, nx8278, 
      gen_21_cmp_mReg_7, nx8290, nx8292, nx8296, nx8300, gen_21_cmp_mReg_8, 
      nx8312, nx8314, nx8318, nx8322, gen_21_cmp_mReg_9, nx8334, nx8336, 
      nx8340, nx8344, gen_21_cmp_mReg_10, nx8356, nx8358, nx8362, nx8366, 
      gen_21_cmp_mReg_11, nx8378, nx8380, nx8384, nx8388, gen_21_cmp_mReg_12, 
      nx8400, nx8402, nx8406, nx8410, gen_21_cmp_mReg_13, nx8422, nx8424, 
      nx8428, nx8432, gen_21_cmp_mReg_14, nx8444, nx8446, nx8450, nx8454, 
      gen_21_cmp_mReg_15, nx8466, nx8468, nx8472, nx8476, nx8482, nx8486, 
      nx8498, gen_22_cmp_mReg_0, nx8518, nx8526, gen_22_cmp_mReg_1, nx8538, 
      nx8540, nx8550, nx8554, gen_22_cmp_mReg_2, nx8566, nx8568, nx8572, 
      nx8576, gen_22_cmp_mReg_3, nx8588, nx8590, nx8594, nx8598, 
      gen_22_cmp_mReg_4, nx8610, nx8612, nx8616, nx8620, gen_22_cmp_mReg_5, 
      nx8632, nx8634, nx8638, nx8642, gen_22_cmp_mReg_6, nx8654, nx8656, 
      nx8660, nx8664, gen_22_cmp_mReg_7, nx8676, nx8678, nx8682, nx8686, 
      gen_22_cmp_mReg_8, nx8698, nx8700, nx8704, nx8708, gen_22_cmp_mReg_9, 
      nx8720, nx8722, nx8726, nx8730, gen_22_cmp_mReg_10, nx8742, nx8744, 
      nx8748, nx8752, gen_22_cmp_mReg_11, nx8764, nx8766, nx8770, nx8774, 
      gen_22_cmp_mReg_12, nx8786, nx8788, nx8792, nx8796, gen_22_cmp_mReg_13, 
      nx8808, nx8810, nx8814, nx8818, gen_22_cmp_mReg_14, nx8830, nx8832, 
      nx8836, nx8840, gen_22_cmp_mReg_15, nx8852, nx8854, nx8858, nx8862, 
      nx8868, nx8872, nx8884, gen_23_cmp_mReg_0, nx8904, nx8912, 
      gen_23_cmp_mReg_1, nx8924, nx8926, nx8936, nx8940, gen_23_cmp_mReg_2, 
      nx8952, nx8954, nx8958, nx8962, gen_23_cmp_mReg_3, nx8974, nx8976, 
      nx8980, nx8984, gen_23_cmp_mReg_4, nx8996, nx8998, nx9002, nx9006, 
      gen_23_cmp_mReg_5, nx9018, nx9020, nx9024, nx9028, gen_23_cmp_mReg_6, 
      nx9040, nx9042, nx9046, nx9050, gen_23_cmp_mReg_7, nx9062, nx9064, 
      nx9068, nx9072, gen_23_cmp_mReg_8, nx9084, nx9086, nx9090, nx9094, 
      gen_23_cmp_mReg_9, nx9106, nx9108, nx9112, nx9116, gen_23_cmp_mReg_10, 
      nx9128, nx9130, nx9134, nx9138, gen_23_cmp_mReg_11, nx9150, nx9152, 
      nx9156, nx9160, gen_23_cmp_mReg_12, nx9172, nx9174, nx9178, nx9182, 
      gen_23_cmp_mReg_13, nx9194, nx9196, nx9200, nx9204, gen_23_cmp_mReg_14, 
      nx9216, nx9218, nx9222, nx9226, gen_23_cmp_mReg_15, nx9238, nx9240, 
      nx9244, nx9248, nx9254, nx9258, nx9270, gen_24_cmp_mReg_0, nx9290, 
      nx9298, gen_24_cmp_mReg_1, nx9310, nx9312, nx9322, nx9326, 
      gen_24_cmp_mReg_2, nx9338, nx9340, nx9344, nx9348, gen_24_cmp_mReg_3, 
      nx9360, nx9362, nx9366, nx9370, gen_24_cmp_mReg_4, nx9382, nx9384, 
      nx9388, nx9392, gen_24_cmp_mReg_5, nx9404, nx9406, nx9410, nx9414, 
      gen_24_cmp_mReg_6, nx9426, nx9428, nx9432, nx9436, gen_24_cmp_mReg_7, 
      nx9448, nx9450, nx9454, nx9458, gen_24_cmp_mReg_8, nx9470, nx9472, 
      nx9476, nx9480, gen_24_cmp_mReg_9, nx9492, nx9494, nx9498, nx9502, 
      gen_24_cmp_mReg_10, nx9514, nx9516, nx9520, nx9524, gen_24_cmp_mReg_11, 
      nx9536, nx9538, nx9542, nx9546, gen_24_cmp_mReg_12, nx9558, nx9560, 
      nx9564, nx9568, gen_24_cmp_mReg_13, nx9580, nx9582, nx9586, nx9590, 
      gen_24_cmp_mReg_14, nx9602, nx9604, nx9608, nx9612, gen_24_cmp_mReg_15, 
      nx9624, nx9626, nx9630, nx9634, nx9640, nx9644, CounterCmp_outp_1, 
      restartDetection, nx9650, StartCaptuerCmp_d, nx9660, nx9666, nx3671, 
      nx3681, nx3691, nx3697, nx3713, nx3720, nx3729, nx3733, nx3737, nx3741, 
      nx3745, nx3751, nx3757, nx3761, nx3769, nx3771, nx3775, nx3786, nx3791, 
      nx3795, nx3801, nx3807, nx3810, nx3817, nx3823, nx3827, nx3831, nx3837, 
      nx3841, nx3845, nx3851, nx3855, nx3861, nx3867, nx3870, nx3874, nx3879, 
      nx3883, nx3889, nx3895, nx3899, nx3903, nx3909, nx3913, nx3919, nx3923, 
      nx3927, nx3931, nx3937, nx3941, nx3945, nx3951, nx3954, nx3961, nx3967, 
      nx3971, nx3975, nx3981, nx3985, nx3989, nx3996, nx4001, nx4005, nx4013, 
      nx4015, nx4018, nx4031, nx4037, nx4040, nx4045, nx4051, nx4055, nx4061, 
      nx4065, nx4069, nx4075, nx4081, nx4084, nx4089, nx4095, nx4099, nx4105, 
      nx4109, nx4113, nx4119, nx4125, nx4128, nx4133, nx4139, nx4143, nx4149, 
      nx4153, nx4157, nx4163, nx4169, nx4172, nx4177, nx4183, nx4187, nx4193, 
      nx4197, nx4201, nx4207, nx4213, nx4216, nx4221, nx4227, nx4231, nx4237, 
      nx4243, nx4249, nx4253, nx4260, nx4263, nx4267, nx4279, nx4285, nx4288, 
      nx4293, nx4299, nx4303, nx4309, nx4315, nx4318, nx4325, nx4331, nx4335, 
      nx4339, nx4345, nx4349, nx4353, nx4359, nx4362, nx4369, nx4375, nx4379, 
      nx4383, nx4389, nx4393, nx4397, nx4403, nx4406, nx4413, nx4419, nx4423, 
      nx4427, nx4433, nx4437, nx4441, nx4447, nx4450, nx4457, nx4463, nx4467, 
      nx4471, nx4477, nx4481, nx4485, nx4492, nx4497, nx4501, nx4509, nx4511, 
      nx4514, nx4527, nx4533, nx4536, nx4541, nx4547, nx4551, nx4557, nx4561, 
      nx4565, nx4571, nx4577, nx4580, nx4585, nx4591, nx4595, nx4601, nx4605, 
      nx4609, nx4615, nx4621, nx4625, nx4631, nx4637, nx4641, nx4645, nx4649, 
      nx4653, nx4659, nx4665, nx4669, nx4674, nx4679, nx4683, nx4687, nx4693, 
      nx4697, nx4702, nx4707, nx4711, nx4717, nx4723, nx4726, nx4733, nx4739, 
      nx4745, nx4748, nx4757, nx4759, nx4763, nx4773, nx4779, nx4783, nx4789, 
      nx4793, nx4797, nx4803, nx4809, nx4812, nx4817, nx4823, nx4827, nx4833, 
      nx4837, nx4841, nx4847, nx4853, nx4856, nx4861, nx4867, nx4871, nx4877, 
      nx4881, nx4885, nx4891, nx4897, nx4900, nx4905, nx4911, nx4915, nx4921, 
      nx4925, nx4929, nx4935, nx4941, nx4944, nx4949, nx4955, nx4959, nx4965, 
      nx4969, nx4973, nx4979, nx4987, nx4991, nx4995, nx5003, nx5005, nx5009, 
      nx5021, nx5027, nx5030, nx5035, nx5041, nx5045, nx5051, nx5057, nx5060, 
      nx5065, nx5071, nx5075, nx5081, nx5087, nx5090, nx5097, nx5103, nx5107, 
      nx5111, nx5117, nx5121, nx5125, nx5131, nx5134, nx5141, nx5147, nx5151, 
      nx5155, nx5161, nx5165, nx5169, nx5175, nx5178, nx5185, nx5191, nx5195, 
      nx5199, nx5205, nx5209, nx5213, nx5219, nx5222, nx5229, nx5235, nx5241, 
      nx5244, nx5253, nx5255, nx5259, nx5269, nx5275, nx5279, nx5285, nx5289, 
      nx5293, nx5299, nx5305, nx5308, nx5313, nx5319, nx5323, nx5329, nx5333, 
      nx5337, nx5343, nx5349, nx5352, nx5357, nx5363, nx5367, nx5373, nx5377, 
      nx5381, nx5387, nx5393, nx5397, nx5403, nx5409, nx5413, nx5417, nx5421, 
      nx5425, nx5431, nx5437, nx5441, nx5446, nx5451, nx5455, nx5459, nx5465, 
      nx5469, nx5474, nx5481, nx5487, nx5491, nx5499, nx5501, nx5505, nx5515, 
      nx5519, nx5523, nx5529, nx5533, nx5537, nx5541, nx5547, nx5551, nx5555, 
      nx5561, nx5564, nx5571, nx5577, nx5581, nx5585, nx5591, nx5595, nx5599, 
      nx5605, nx5608, nx5615, nx5621, nx5625, nx5629, nx5635, nx5639, nx5643, 
      nx5649, nx5652, nx5659, nx5665, nx5669, nx5673, nx5679, nx5683, nx5687, 
      nx5693, nx5696, nx5703, nx5709, nx5713, nx5717, nx5725, nx5731, nx5735, 
      nx5743, nx5745, nx5749, nx5760, nx5765, nx5769, nx5775, nx5781, nx5785, 
      nx5791, nx5797, nx5800, nx5804, nx5809, nx5813, nx5819, nx5825, nx5829, 
      nx5833, nx5839, nx5843, nx5849, nx5853, nx5857, nx5861, nx5867, nx5871, 
      nx5875, nx5881, nx5884, nx5891, nx5897, nx5901, nx5905, nx5911, nx5915, 
      nx5919, nx5925, nx5928, nx5935, nx5941, nx5945, nx5949, nx5955, nx5959, 
      nx5963, nx5970, nx5975, nx5979, nx5987, nx5989, nx5992, nx6005, nx6011, 
      nx6014, nx6019, nx6025, nx6029, nx6035, nx6039, nx6043, nx6049, nx6055, 
      nx6058, nx6063, nx6069, nx6073, nx6079, nx6083, nx6087, nx6093, nx6099, 
      nx6102, nx6107, nx6113, nx6117, nx6123, nx6127, nx6131, nx6137, nx6143, 
      nx6146, nx6151, nx6157, nx6161, nx6167, nx6171, nx6175, nx6181, nx6186, 
      nx6189, nx6193, nx6199, nx6203, nx6209, nx6217, nx6221, nx6225, nx6233, 
      nx6235, nx6239, nx6249, nx6255, nx6259, nx6265, nx6269, nx6273, nx6279, 
      nx6283, nx6287, nx6291, nx6297, nx6301, nx6305, nx6311, nx6314, nx6321, 
      nx6327, nx6331, nx6335, nx6341, nx6345, nx6349, nx6355, nx6358, nx6365, 
      nx6371, nx6375, nx6379, nx6385, nx6389, nx6393, nx6399, nx6402, nx6409, 
      nx6415, nx6419, nx6423, nx6429, nx6433, nx6437, nx6443, nx6446, nx6453, 
      nx6459, nx6465, nx6468, nx6477, nx6479, nx6483, nx6493, nx6499, nx6503, 
      nx6509, nx6513, nx6517, nx6523, nx6529, nx6532, nx6537, nx6543, nx6547, 
      nx6553, nx6557, nx6561, nx6567, nx6572, nx6575, nx6579, nx6585, nx6589, 
      nx6595, nx6601, nx6604, nx6609, nx6615, nx6619, nx6625, nx6631, nx6634, 
      nx6641, nx6647, nx6651, nx6655, nx6661, nx6665, nx6669, nx6675, nx6678, 
      nx6685, nx6691, nx6695, nx6699, nx6707, nx6713, nx6717, nx6725, nx6727, 
      nx6731, nx6742, nx6747, nx6751, nx6757, nx6763, nx6766, nx6773, nx6779, 
      nx6783, nx6787, nx6793, nx6797, nx6801, nx6807, nx6810, nx6817, nx6823, 
      nx6827, nx6831, nx6837, nx6841, nx6845, nx6851, nx6854, nx6861, nx6867, 
      nx6871, nx6875, nx6881, nx6885, nx6889, nx6895, nx6898, nx6905, nx6911, 
      nx6915, nx6919, nx6925, nx6929, nx6933, nx6939, nx6943, nx6949, nx6957, 
      nx6961, nx6965, nx6973, nx6975, nx6979, nx6990, nx6995, nx6999, nx7003, 
      nx7009, nx7013, nx7018, nx7023, nx7027, nx7033, nx7039, nx7042, nx7049, 
      nx7055, nx7059, nx7063, nx7069, nx7073, nx7077, nx7083, nx7086, nx7093, 
      nx7099, nx7103, nx7107, nx7113, nx7117, nx7121, nx7127, nx7130, nx7137, 
      nx7143, nx7147, nx7151, nx7157, nx7161, nx7165, nx7171, nx7174, nx7181, 
      nx7187, nx7191, nx7195, nx7203, nx7209, nx7213, nx7221, nx7223, nx7227, 
      nx7238, nx7243, nx7247, nx7253, nx7259, nx7262, nx7269, nx7275, nx7279, 
      nx7283, nx7289, nx7293, nx7297, nx7303, nx7306, nx7313, nx7319, nx7323, 
      nx7329, nx7335, nx7339, nx7344, nx7348, nx7351, nx7357, nx7363, nx7367, 
      nx7373, nx7377, nx7381, nx7387, nx7393, nx7397, nx7403, nx7407, nx7411, 
      nx7417, nx7423, nx7426, nx7431, nx7437, nx7441, nx7447, nx7453, nx7459, 
      nx7463, nx7471, nx7473, nx7477, nx7489, nx7493, nx7497, nx7503, nx7507, 
      nx7511, nx7515, nx7521, nx7525, nx7529, nx7535, nx7538, nx7545, nx7551, 
      nx7555, nx7559, nx7565, nx7569, nx7573, nx7579, nx7582, nx7589, nx7595, 
      nx7599, nx7603, nx7609, nx7613, nx7617, nx7623, nx7626, nx7633, nx7639, 
      nx7643, nx7647, nx7653, nx7657, nx7661, nx7667, nx7670, nx7677, nx7683, 
      nx7687, nx7691, nx7699, nx7705, nx7709, nx7717, nx7719, nx7723, nx7733, 
      nx7737, nx7741, nx7747, nx7753, nx7757, nx7762, nx7767, nx7771, nx7775, 
      nx7781, nx7785, nx7790, nx7795, nx7799, nx7805, nx7811, nx7814, nx7821, 
      nx7827, nx7831, nx7835, nx7841, nx7845, nx7849, nx7855, nx7858, nx7865, 
      nx7871, nx7875, nx7879, nx7885, nx7889, nx7893, nx7899, nx7902, nx7909, 
      nx7915, nx7919, nx7923, nx7929, nx7933, nx7937, nx7944, nx7949, nx7953, 
      nx7961, nx7963, nx7966, nx7979, nx7985, nx7988, nx7993, nx7999, nx8003, 
      nx8009, nx8013, nx8017, nx8023, nx8029, nx8032, nx8037, nx8043, nx8047, 
      nx8053, nx8057, nx8061, nx8067, nx8073, nx8076, nx8081, nx8087, nx8091, 
      nx8097, nx8101, nx8105, nx8111, nx8116, nx8119, nx8123, nx8129, nx8133, 
      nx8139, nx8145, nx8148, nx8153, nx8159, nx8163, nx8169, nx8175, nx8178, 
      nx8185, nx8191, nx8197, nx8200, nx8209, nx8211, nx8215, nx8225, nx8231, 
      nx8235, nx8241, nx8245, nx8249, nx8255, nx8261, nx8264, nx8269, nx8275, 
      nx8279, nx8285, nx8289, nx8293, nx8299, nx8305, nx8308, nx8313, nx8319, 
      nx8323, nx8329, nx8333, nx8337, nx8343, nx8349, nx8352, nx8357, nx8363, 
      nx8367, nx8373, nx8377, nx8381, nx8387, nx8393, nx8396, nx8401, nx8407, 
      nx8411, nx8417, nx8421, nx8425, nx8431, nx8439, nx8443, nx8447, nx8455, 
      nx8457, nx8461, nx8473, nx8477, nx8481, nx8487, nx8493, nx8497, nx8502, 
      nx8506, nx8509, nx8515, nx8521, nx8525, nx8531, nx8535, nx8539, nx8545, 
      nx8551, nx8555, nx8561, nx8565, nx8569, nx8575, nx8581, nx8584, nx8589, 
      nx8595, nx8599, nx8605, nx8609, nx8613, nx8619, nx8625, nx8628, nx8633, 
      nx8639, nx8643, nx8649, nx8653, nx8657, nx8663, nx8669, nx8672, nx8677, 
      nx8685, nx8691, nx8694, nx8701, nx8703, nx8707, nx8718, nx8725, nx8729, 
      nx8735, nx8739, nx8743, nx8749, nx8753, nx8757, nx8761, nx8767, nx8771, 
      nx8775, nx8781, nx8784, nx8791, nx8797, nx8801, nx8805, nx8811, nx8815, 
      nx8819, nx8825, nx8828, nx8835, nx8841, nx8845, nx8849, nx8855, nx8859, 
      nx8863, nx8869, nx8873, nx8879, nx8885, nx8888, nx8892, nx8897, nx8901, 
      nx8907, nx8913, nx8917, nx8921, nx8929, nx8933, nx8937, nx8945, nx8947, 
      nx8950, nx8963, nx8969, nx8972, nx8979, nx8985, nx8989, nx8993, nx8999, 
      nx9003, nx9007, nx9013, nx9016, nx9023, nx9029, nx9033, nx9037, nx9043, 
      nx9047, nx9051, nx9057, nx9060, nx9067, nx9073, nx9077, nx9081, nx9087, 
      nx9091, nx9095, nx9101, nx9104, nx9111, nx9117, nx9121, nx9125, nx9131, 
      nx9135, nx9139, nx9145, nx9148, nx9155, nx9161, nx9165, nx9169, nx9177, 
      nx9183, nx9187, nx9195, nx9197, nx9201, nx9212, nx9217, nx9221, nx9227, 
      nx9233, nx9236, nx9243, nx9249, nx9253, nx9259, nx9265, nx9269, nx9274, 
      nx9278, nx9281, nx9287, nx9293, nx9297, nx9303, nx9307, nx9311, nx9317, 
      nx9323, nx9327, nx9333, nx9337, nx9341, nx9347, nx9353, nx9356, nx9361, 
      nx9367, nx9371, nx9377, nx9381, nx9385, nx9391, nx9397, nx9400, nx9405, 
      nx9411, nx9415, nx9421, nx9427, nx9433, nx9437, nx9445, nx9447, nx9451, 
      nx9463, nx9467, nx9471, nx9477, nx9481, nx9485, nx9489, nx9495, nx9499, 
      nx9503, nx9509, nx9512, nx9519, nx9525, nx9529, nx9533, nx9539, nx9543, 
      nx9547, nx9553, nx9556, nx9563, nx9569, nx9573, nx9577, nx9583, nx9587, 
      nx9591, nx9597, nx9600, nx9607, nx9613, nx9617, nx9621, nx9627, nx9631, 
      nx9635, nx9641, nx9645, nx9651, nx9655, nx9658, nx9663, nx9669, nx9673, 
      nx9676, nx9683, nx9685, nx9688, nx9698, nx9702, nx9705, nx9709, nx9713, 
      nx9716, nx9720, nx9724, nx9727, nx9731, nx9735, nx9738, nx9742, nx9746, 
      nx9749, nx9753, nx9757, nx9760, nx9764, nx9768, nx9771, nx9775, nx9779, 
      nx9782, nx9786, nx9790, nx9793, nx9797, nx9801, nx9804, nx9808, nx9812, 
      nx9815, nx9819, nx9823, nx9826, nx9830, nx9834, nx9837, nx9841, nx9845, 
      nx9848, nx9852, nx9857, nx9860, nx9864, nx9867, nx9870, nx9874, nx9877, 
      nx9880, nx9884, nx9887, nx9890, nx9894, nx9897, nx9900, nx9904, nx9907, 
      nx9910, nx9914, nx9917, nx9920, nx9924, nx9927, nx9930, nx9934, nx9937, 
      nx9940, nx9944, nx9947, nx9950, nx9954, nx9957, nx9960, nx9964, nx9967, 
      nx9970, nx9974, nx9977, nx9980, nx9984, nx9987, nx9990, nx9994, nx9997, 
      nx10000, nx10004, nx10007, nx10010, nx10014, nx10017, nx10020, nx10024, 
      nx10027, nx10030, nx10034, nx10037, nx10040, nx10044, nx10047, nx10050, 
      nx10054, nx10057, nx10060, nx10064, nx10067, nx10070, nx10074, nx10077, 
      nx10080, nx10084, nx10087, nx10090, nx10094, nx10097, nx10100, nx10104, 
      nx10107, nx10120, nx10122, nx10124, nx10126, nx10128, nx10130, nx10132, 
      nx10134, nx10136, nx10138, nx10140, nx10142, nx10144, nx10146, nx10148, 
      nx10150, nx10152, nx10154, nx10156, nx10158, nx10160, nx10162, nx10164, 
      nx10166, nx10168, nx10170, nx10172, nx10174, nx10176, nx10178, nx10180, 
      nx10182, nx10184, nx10186, nx10188, nx10190, nx10192, nx10194, nx10196, 
      nx10198, nx10200, nx10202, nx10204, nx10206, nx10208, nx10210, nx10212, 
      nx10214, nx10216, nx10218, nx10220, nx10222, nx10224, nx10226, nx10228, 
      nx10230, nx10232, nx10234, nx10236, nx10238, nx10240, nx10242, nx10244, 
      nx10246, nx10248, nx10250, nx10252, nx10254, nx10256, nx10258, nx10260, 
      nx10262, nx10264, nx10266, nx10268, nx10270, nx10272, nx10274, nx10276, 
      nx10278, nx10280, nx10282, nx10284, nx10286, nx10288, nx10290, nx10292, 
      nx10294, nx10296, nx10298, nx10300, nx10302, nx10304, nx10306, nx10308, 
      nx10310, nx10312, nx10314, nx10316, nx10318, nx10320, nx10322, nx10324, 
      nx10326, nx10328, nx10330, nx10332, nx10334, nx10336, nx10338, nx10340, 
      nx10342, nx10344, nx10346, nx10348, nx10350, nx10352, nx10354, nx10356, 
      nx10358, nx10360, nx10362, nx10364, nx10366, nx10368, nx10370, nx10372, 
      nx10374, nx10376, nx10378, nx10380, nx10382, nx10384, nx10386, nx10388, 
      nx10390, nx10392, nx10394, nx10396, nx10398, nx10400, nx10402, nx10404, 
      nx10406, nx10408, nx10410, nx10412, nx10414, nx10416, nx10418, nx10420, 
      nx10422, nx10424, nx10426, nx10428, nx10430, nx10432, nx10434, nx10436, 
      nx10438, nx10440, nx10442, nx10444, nx10446, nx10448, nx10450, nx10452, 
      nx10454, nx10456, nx10458, nx10460, nx10462, nx10464, nx10466, nx10468, 
      nx10470, nx10472, nx10474, nx10476, nx10478, nx10480, nx10482, nx10484, 
      nx10486, nx10488, nx10490, nx10492, nx10494, nx10496, nx10498, nx10500, 
      nx10502, nx10504, nx10506, nx10508, nx10510, nx10512, nx10514, nx10516, 
      nx10518, nx10520, nx10522, nx10524, nx10526, nx10528, nx10530, nx10532, 
      nx10534, nx10536, nx10538, nx10540, nx10542, nx10544, nx10546, nx10548, 
      nx10550, nx10552, nx10554, nx10556, nx10558, nx10560, nx10562, nx10564, 
      nx10566, nx10568, nx10570, nx10572, nx10574, nx10576, nx10578, nx10580, 
      nx10582, nx10584, nx10586, nx10588, nx10590, nx10592, nx10594, nx10596, 
      nx10598, nx10600, nx10602, nx10604, nx10606, nx10608, nx10610, nx10612, 
      nx10614, nx10616, nx10618, nx10620, nx10622, nx10624, nx10626, nx10628, 
      nx10630, nx10632, nx10634, nx10636, nx10638, nx10640, nx10642, nx10644, 
      nx10646, nx10648, nx10650, nx10652, nx10654, nx10656, nx10658, nx10660, 
      nx10662, nx10664, nx10666, nx10668, nx10670, nx10672, nx10674, nx10676, 
      nx10678, nx10680, nx10682, nx10684, nx10686, nx10688, nx10690, nx10692, 
      nx10694, nx10696, nx10698, nx10700, nx10702, nx10704, nx10706, nx10708, 
      nx10710, nx10712, nx10714, nx10716, nx10718, nx10720, nx10722, nx10724, 
      nx10726, nx10728, nx10730, nx10732, nx10734, nx10736, nx10738, nx10740, 
      nx10742, nx10744, nx10746, nx10748, nx10750, nx10752, nx10754, nx10756, 
      nx10758, nx10760, nx10762, nx10764, nx10766, nx10768, nx10770, nx10772, 
      nx10774, nx10776, nx10778, nx10780, nx10782, nx10784, nx10786, nx10788, 
      nx10790, nx10792, nx10794, nx10796, nx10798, nx10800, nx10802, nx10804, 
      nx10806, nx10808, nx10810, nx10812, nx10814, nx10816, nx10818, nx10820, 
      nx10822, nx10824, nx10826, nx10828, nx10830, nx10832, nx10834, nx10836, 
      nx10838, nx10840, nx10842, nx10844, nx10846, nx10848, nx10850, nx10852, 
      nx10854, nx10856, nx10858, nx10860, nx10862, nx10864, nx10866, nx10868, 
      nx10870, nx10872, nx10874, nx10876, nx10878, nx10880, nx10882, nx10884, 
      nx10886, nx10888, nx10890, nx10892, nx10894, nx10896, nx10898, nx10900, 
      nx10902, nx10904, nx10906, nx10908, nx10910, nx10912, nx10914, nx10916, 
      nx10918, nx10920, nx10922, nx10924, nx10926, nx10928, nx10930, nx10932, 
      nx10934, nx10936, nx10938, nx10940, nx10942, nx10944, nx10946, nx10948, 
      nx10950, nx10952, nx10954, nx10956, nx10958, nx10960, nx10962, nx10964, 
      nx10966, nx10968, nx10970, nx10972, nx10974, nx10976, nx10978, nx10980, 
      nx10982, nx10984, nx10986, nx10988, nx10990, nx10992, nx10994, nx10996, 
      nx10998, nx11000, nx11002, nx11004, nx11006, nx11008, nx11010, nx11012, 
      nx11014, nx11016, nx11018, nx11020, nx11022, nx11024, nx11026, nx11028, 
      nx11030, nx11032, nx11034, nx11036, nx11038, nx11040, nx11042, nx11044, 
      nx11046, nx11048, nx11050, nx11052, nx11054, nx11056, nx11058, nx11060, 
      nx11062, nx11064, nx11066, nx11068, nx11070, nx11072, nx11074, nx11076, 
      nx11078, nx11080, nx11082, nx11084, nx11086, nx11088, nx11090, nx11092, 
      nx11094, nx11096, nx11098, nx11100, nx11102, nx11104, nx11106, nx11108, 
      nx11110, nx11112, nx11114, nx11116, nx11118, nx11120, nx11122, nx11124, 
      nx11126, nx11128, nx11130, nx11132, nx11134, nx11136, nx11138, nx11140, 
      nx11142, nx11144, nx11146, nx11148, nx11150, nx11152, nx11154, nx11156, 
      nx11158, nx11160, nx11162, nx11164, nx11166, nx11168, nx11170, nx11172, 
      nx11174, nx11176, nx11178, nx11180, nx11182, nx11184, nx11186, nx11188, 
      nx11190, nx11192, nx11194, nx11196, nx11198, nx11200, nx11202, nx11204, 
      nx11206, nx11208, nx11210, nx11212, nx11214, nx11216, nx11218, nx11220, 
      nx11222, nx11224, nx11226, nx11228, nx11230, nx11232, nx11234, nx11236, 
      nx11238, nx11240, nx11242, nx11244, nx11246, nx11248, nx11250, nx11252, 
      nx11254, nx11256, nx11258, nx11260, nx11262, nx11264, nx11266, nx11268, 
      nx11270, nx11272, nx11274, nx11276, nx11278, nx11280, nx11282, nx11284, 
      nx11286, nx11288, nx11290, nx11292, nx11294, nx11296, nx11298, nx11300, 
      nx11302, nx11304, nx11306, nx11308, nx11310, nx11312, nx11314, nx11316, 
      nx11318, nx11320, nx11322, nx11324, nx11326, nx11328, nx11330, nx11332, 
      nx11334, nx11336, nx11338, nx11340, nx11342, nx11344, nx11346, nx11348, 
      nx11350, nx11352, nx11354, nx11356, nx11358, nx11360, nx11362, nx11364, 
      nx11366, nx11368, nx11370, nx11372, nx11374, nx11376, nx11378, nx11380, 
      nx11382, nx11384, nx11386, nx11388, nx11390, nx11392, nx11394, nx11396, 
      nx11398, nx11400, nx11402, nx11404, nx11406, nx11408, nx11410, nx11412, 
      nx11414, nx11416, nx11418, nx11420, nx11422, nx11424, nx11426, nx11428, 
      nx11430, nx11432, nx11434, nx11436, nx11438, nx11440, nx11442, nx11444, 
      nx11446, nx11448, nx11450, nx11452, nx11454, nx11456, nx11458, nx11460, 
      nx11462, nx11464, nx11466, nx11468, nx11470, nx11472, nx11474, nx11476, 
      nx11478, nx11480, nx11482, nx11484, nx11486, nx11488, nx11490, nx11492, 
      nx11494, nx11496, nx11498, nx11500, nx11502, nx11504, nx11506, nx11508, 
      nx11510, nx11512, nx11514, nx11516, nx11518, nx11520, nx11522, nx11524, 
      nx11526, nx11528, nx11530, nx11532, nx11534, nx11536, nx11538, nx11540, 
      nx11542, nx11544, nx11546, nx11548, nx11550, nx11552, nx11554, nx11556, 
      nx11558, nx11560, nx11562, nx11564, nx11566, nx11568, nx11570, nx11572, 
      nx11574, nx11576, nx11578, nx11580, nx11582, nx11584, nx11586, nx11588, 
      nx11590, nx11592, nx11594, nx11596, nx11598, nx11600, nx11602, nx11604, 
      nx11606, nx11608, nx11610, nx11612, nx11614, nx11616, nx11618, nx11620, 
      nx11622, nx11624, nx11626, nx11628, nx11630, nx11632, nx11634, nx11636, 
      nx11638, nx11640, nx11642, nx11644, nx11646, nx11648, nx11650, nx11652, 
      nx11654, nx11656, nx11658, nx11660, nx11662, nx11664, nx11666, nx11668, 
      nx11670, nx11672, nx11674, nx11676, nx11678, nx11680, nx11682, nx11684, 
      nx11686, nx11688, nx11690, nx11692, nx11694, nx11696, nx11698, nx11700, 
      nx11702, nx11704, nx11706, nx11708, nx11710, nx11712, nx11714, nx11716, 
      nx11718, nx11720, nx11722, nx11724, nx11726, nx11728, nx11730, nx11732, 
      nx11734, nx11736, nx11738, nx11740, nx11742, nx11744, nx11746, nx11748, 
      nx11750, nx11752, nx11754, nx11756, nx11758, nx11760, nx11762, nx11764, 
      nx11766, nx11768, nx11770, nx11772, nx11774, nx11776, nx11778, nx11780, 
      nx11782, nx11784, nx11786, nx11788, nx11790, nx11792, nx11794, nx11796, 
      nx11798, nx11800, nx11802, nx11804, nx11806, nx11808, nx11810, nx11812, 
      nx11814, nx11816, nx11818, nx11820, nx11822, nx11824, nx11826, nx11828, 
      nx11830, nx11832, nx11834, nx11836, nx11838, nx11840, nx11842, nx11844, 
      nx11846, nx11848, nx11850, nx11852, nx11854, nx11856, nx11858, nx11860, 
      nx11862, nx11864, nx11866, nx11868, nx11870, nx11872, nx11874, nx11876, 
      nx11878, nx11880, nx11882, nx11884, nx11886, nx11896, nx11898, nx11900, 
      nx11902, nx11904, nx11906, nx11908, nx11910, nx11912, nx11914, nx11916, 
      nx11918, nx11920, nx11922, nx11924, nx11926, nx11928, nx11934, nx11936, 
      nx11938, nx11940: std_logic ;
   
   signal DANGLING : std_logic_vector (124 downto 0 );

begin
   gen_24_cmp_pRegCmp : Reg_33 port map ( D(32)=>gen_24_cmp_pInit_32, D(31)
      =>gen_24_cmp_pInit_32, D(30)=>gen_24_cmp_pBs_30, D(29)=>
      gen_24_cmp_pBs_29, D(28)=>gen_24_cmp_pBs_28, D(27)=>gen_24_cmp_pBs_27, 
      D(26)=>gen_24_cmp_pBs_26, D(25)=>gen_24_cmp_pBs_25, D(24)=>
      gen_24_cmp_pBs_24, D(23)=>gen_24_cmp_pBs_23, D(22)=>outputs_24_15, 
      D(21)=>outputs_24_14, D(20)=>outputs_24_13, D(19)=>outputs_24_12, 
      D(18)=>outputs_24_11, D(17)=>outputs_24_10, D(16)=>outputs_24_9, D(15)
      =>outputs_24_8, D(14)=>outputs_24_7, D(13)=>outputs_24_6, D(12)=>
      outputs_24_5, D(11)=>outputs_24_4, D(10)=>outputs_24_3, D(9)=>
      outputs_24_2, D(8)=>outputs_24_1, D(7)=>outputs_24_0, D(6)=>
      gen_24_cmp_pMux_8, D(5)=>gen_24_cmp_pMux_7, D(4)=>gen_24_cmp_pMux_6, 
      D(3)=>gen_24_cmp_pMux_5, D(2)=>gen_24_cmp_pMux_4, D(1)=>
      gen_24_cmp_pMux_3, D(0)=>nx10130, en=>nx11916, clk=>nx10122, rst=>rst, 
      Q(32)=>DANGLING(0), Q(31)=>DANGLING(1), Q(30)=>gen_24_cmp_pReg_30, 
      Q(29)=>gen_24_cmp_pReg_29, Q(28)=>gen_24_cmp_pReg_28, Q(27)=>
      gen_24_cmp_pReg_27, Q(26)=>gen_24_cmp_pReg_26, Q(25)=>
      gen_24_cmp_pReg_25, Q(24)=>gen_24_cmp_pReg_24, Q(23)=>
      gen_24_cmp_pReg_23, Q(22)=>gen_24_cmp_pReg_22, Q(21)=>
      gen_24_cmp_pReg_21, Q(20)=>gen_24_cmp_pReg_20, Q(19)=>
      gen_24_cmp_pReg_19, Q(18)=>gen_24_cmp_pReg_18, Q(17)=>
      gen_24_cmp_pReg_17, Q(16)=>gen_24_cmp_pReg_16, Q(15)=>
      gen_24_cmp_pReg_15, Q(14)=>gen_24_cmp_pReg_14, Q(13)=>
      gen_24_cmp_pReg_13, Q(12)=>gen_24_cmp_pReg_12, Q(11)=>
      gen_24_cmp_pReg_11, Q(10)=>gen_24_cmp_pReg_10, Q(9)=>gen_24_cmp_pReg_9, 
      Q(8)=>gen_24_cmp_pReg_8, Q(7)=>gen_24_cmp_pReg_7, Q(6)=>
      gen_24_cmp_pReg_6, Q(5)=>gen_24_cmp_pReg_5, Q(4)=>gen_24_cmp_pReg_4, 
      Q(3)=>gen_24_cmp_pReg_3, Q(2)=>gen_24_cmp_pReg_2, Q(1)=>
      gen_24_cmp_pReg_1, Q(0)=>gen_24_cmp_pReg_0);
   gen_24_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>gen_24_cmp_pInit_32, 
      a(31)=>gen_24_cmp_pInit_32, a(30)=>gen_24_cmp_pReg_30, a(29)=>
      gen_24_cmp_pReg_29, a(28)=>gen_24_cmp_pReg_28, a(27)=>
      gen_24_cmp_pReg_27, a(26)=>gen_24_cmp_pReg_26, a(25)=>
      gen_24_cmp_pReg_25, a(24)=>gen_24_cmp_pReg_24, a(23)=>
      gen_24_cmp_pReg_23, a(22)=>gen_24_cmp_pReg_22, a(21)=>
      gen_24_cmp_pReg_21, a(20)=>gen_24_cmp_pReg_20, a(19)=>
      gen_24_cmp_pReg_19, a(18)=>gen_24_cmp_pReg_18, a(17)=>
      gen_24_cmp_pReg_17, a(16)=>gen_24_cmp_pReg_16, a(15)=>
      gen_24_cmp_pReg_15, a(14)=>gen_24_cmp_pReg_14, a(13)=>
      gen_24_cmp_pReg_13, a(12)=>gen_24_cmp_pReg_12, a(11)=>
      gen_24_cmp_pReg_11, a(10)=>gen_24_cmp_pReg_10, a(9)=>gen_24_cmp_pReg_9, 
      a(8)=>gen_24_cmp_pReg_8, a(7)=>gen_24_cmp_pReg_7, a(6)=>
      gen_24_cmp_pReg_6, a(5)=>gen_24_cmp_pReg_5, a(4)=>gen_24_cmp_pReg_4, 
      a(3)=>gen_24_cmp_pReg_3, a(2)=>gen_24_cmp_pReg_2, a(1)=>
      gen_24_cmp_pReg_1, a(0)=>gen_24_cmp_pReg_0, b(32)=>gen_24_cmp_pInit_32, 
      b(31)=>gen_24_cmp_pInit_32, b(30)=>gen_24_cmp_pInit_32, b(29)=>
      gen_24_cmp_pInit_32, b(28)=>gen_24_cmp_pInit_32, b(27)=>
      gen_24_cmp_pInit_32, b(26)=>gen_24_cmp_pInit_32, b(25)=>
      gen_24_cmp_pInit_32, b(24)=>gen_24_cmp_pInit_32, b(23)=>
      gen_24_cmp_pInit_32, b(22)=>gen_24_cmp_pInit_32, b(21)=>
      gen_24_cmp_pInit_32, b(20)=>gen_24_cmp_pInit_32, b(19)=>
      gen_24_cmp_pInit_32, b(18)=>gen_24_cmp_pInit_32, b(17)=>
      gen_24_cmp_pInit_32, b(16)=>gen_24_cmp_pInit_32, b(15)=>
      gen_24_cmp_pInit_32, b(14)=>gen_24_cmp_pInit_32, b(13)=>
      gen_24_cmp_pInit_32, b(12)=>gen_24_cmp_pInit_32, b(11)=>
      gen_24_cmp_pInit_32, b(10)=>gen_24_cmp_pInit_32, b(9)=>
      gen_24_cmp_pInit_32, b(8)=>filter_24_7, b(7)=>filter_24_6, b(6)=>
      filter_24_5, b(5)=>filter_24_4, b(4)=>filter_24_3, b(3)=>filter_24_2, 
      b(2)=>filter_24_1, b(1)=>filter_24_0, b(0)=>gen_24_cmp_pInit_32, sel=>
      nx11896, f(32)=>DANGLING(2), f(31)=>DANGLING(3), f(30)=>
      gen_24_cmp_pMux_30, f(29)=>gen_24_cmp_pMux_29, f(28)=>
      gen_24_cmp_pMux_28, f(27)=>gen_24_cmp_pMux_27, f(26)=>
      gen_24_cmp_pMux_26, f(25)=>gen_24_cmp_pMux_25, f(24)=>
      gen_24_cmp_pMux_24, f(23)=>gen_24_cmp_pMux_23, f(22)=>
      gen_24_cmp_pMux_22, f(21)=>gen_24_cmp_pMux_21, f(20)=>
      gen_24_cmp_pMux_20, f(19)=>gen_24_cmp_pMux_19, f(18)=>
      gen_24_cmp_pMux_18, f(17)=>gen_24_cmp_pMux_17, f(16)=>
      gen_24_cmp_pMux_16, f(15)=>gen_24_cmp_pMux_15, f(14)=>
      gen_24_cmp_pMux_14, f(13)=>gen_24_cmp_pMux_13, f(12)=>
      gen_24_cmp_pMux_12, f(11)=>gen_24_cmp_pMux_11, f(10)=>
      gen_24_cmp_pMux_10, f(9)=>gen_24_cmp_pMux_9, f(8)=>gen_24_cmp_pMux_8, 
      f(7)=>gen_24_cmp_pMux_7, f(6)=>gen_24_cmp_pMux_6, f(5)=>
      gen_24_cmp_pMux_5, f(4)=>gen_24_cmp_pMux_4, f(3)=>gen_24_cmp_pMux_3, 
      f(2)=>gen_24_cmp_pMux_2, f(1)=>gen_24_cmp_pMux_1, f(0)=>
      gen_24_cmp_pMux_0);
   gen_24_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>
      gen_24_cmp_pInit_32, a(22)=>gen_24_cmp_pInit_32, a(21)=>
      gen_24_cmp_pMux_30, a(20)=>gen_24_cmp_pMux_29, a(19)=>
      gen_24_cmp_pMux_28, a(18)=>gen_24_cmp_pMux_27, a(17)=>
      gen_24_cmp_pMux_26, a(16)=>gen_24_cmp_pMux_25, a(15)=>
      gen_24_cmp_pMux_24, a(14)=>gen_24_cmp_pMux_23, a(13)=>
      gen_24_cmp_pMux_22, a(12)=>gen_24_cmp_pMux_21, a(11)=>
      gen_24_cmp_pMux_20, a(10)=>gen_24_cmp_pMux_19, a(9)=>
      gen_24_cmp_pMux_18, a(8)=>gen_24_cmp_pMux_17, a(7)=>gen_24_cmp_pMux_16, 
      a(6)=>gen_24_cmp_pMux_15, a(5)=>gen_24_cmp_pMux_14, a(4)=>
      gen_24_cmp_pMux_13, a(3)=>gen_24_cmp_pMux_12, a(2)=>gen_24_cmp_pMux_11, 
      a(1)=>gen_24_cmp_pMux_10, a(0)=>gen_24_cmp_pMux_9, b(23)=>nx10434, 
      b(22)=>nx10434, b(21)=>nx10432, b(20)=>nx10440, b(19)=>nx10438, b(18)
      =>nx10436, b(17)=>nx10434, b(16)=>nx10432, b(15)=>
      gen_24_cmp_BSCmp_op2_15, b(14)=>gen_24_cmp_BSCmp_op2_14, b(13)=>
      gen_24_cmp_BSCmp_op2_13, b(12)=>gen_24_cmp_BSCmp_op2_12, b(11)=>
      gen_24_cmp_BSCmp_op2_11, b(10)=>gen_24_cmp_BSCmp_op2_10, b(9)=>
      gen_24_cmp_BSCmp_op2_9, b(8)=>gen_24_cmp_BSCmp_op2_8, b(7)=>
      gen_24_cmp_BSCmp_op2_7, b(6)=>gen_24_cmp_BSCmp_op2_6, b(5)=>
      gen_24_cmp_BSCmp_op2_5, b(4)=>gen_24_cmp_BSCmp_op2_4, b(3)=>
      gen_24_cmp_BSCmp_op2_3, b(2)=>gen_24_cmp_BSCmp_op2_2, b(1)=>
      gen_24_cmp_BSCmp_op2_1, b(0)=>gen_24_cmp_BSCmp_op2_0, carryIn=>
      gen_24_cmp_BSCmp_carryIn, sum(23)=>gen_24_cmp_pBs_30, sum(22)=>
      gen_24_cmp_pBs_29, sum(21)=>gen_24_cmp_pBs_28, sum(20)=>
      gen_24_cmp_pBs_27, sum(19)=>gen_24_cmp_pBs_26, sum(18)=>
      gen_24_cmp_pBs_25, sum(17)=>gen_24_cmp_pBs_24, sum(16)=>
      gen_24_cmp_pBs_23, sum(15)=>outputs_24_15, sum(14)=>outputs_24_14, 
      sum(13)=>outputs_24_13, sum(12)=>outputs_24_12, sum(11)=>outputs_24_11, 
      sum(10)=>outputs_24_10, sum(9)=>outputs_24_9, sum(8)=>outputs_24_8, 
      sum(7)=>outputs_24_7, sum(6)=>outputs_24_6, sum(5)=>outputs_24_5, 
      sum(4)=>outputs_24_4, sum(3)=>outputs_24_3, sum(2)=>outputs_24_2, 
      sum(1)=>outputs_24_1, sum(0)=>outputs_24_0, carryOut=>DANGLING(4));
   gen_23_cmp_pRegCmp : Reg_33 port map ( D(32)=>gen_24_cmp_pInit_32, D(31)
      =>gen_24_cmp_pInit_32, D(30)=>gen_23_cmp_pBs_30, D(29)=>
      gen_23_cmp_pBs_29, D(28)=>gen_23_cmp_pBs_28, D(27)=>gen_23_cmp_pBs_27, 
      D(26)=>gen_23_cmp_pBs_26, D(25)=>gen_23_cmp_pBs_25, D(24)=>
      gen_23_cmp_pBs_24, D(23)=>gen_23_cmp_pBs_23, D(22)=>outputs_23_15, 
      D(21)=>outputs_23_14, D(20)=>outputs_23_13, D(19)=>outputs_23_12, 
      D(18)=>outputs_23_11, D(17)=>outputs_23_10, D(16)=>outputs_23_9, D(15)
      =>outputs_23_8, D(14)=>outputs_23_7, D(13)=>outputs_23_6, D(12)=>
      outputs_23_5, D(11)=>outputs_23_4, D(10)=>outputs_23_3, D(9)=>
      outputs_23_2, D(8)=>outputs_23_1, D(7)=>outputs_23_0, D(6)=>
      gen_23_cmp_pMux_8, D(5)=>gen_23_cmp_pMux_7, D(4)=>gen_23_cmp_pMux_6, 
      D(3)=>gen_23_cmp_pMux_5, D(2)=>gen_23_cmp_pMux_4, D(1)=>
      gen_23_cmp_pMux_3, D(0)=>nx10142, en=>nx11916, clk=>nx10122, rst=>rst, 
      Q(32)=>DANGLING(5), Q(31)=>DANGLING(6), Q(30)=>gen_23_cmp_pReg_30, 
      Q(29)=>gen_23_cmp_pReg_29, Q(28)=>gen_23_cmp_pReg_28, Q(27)=>
      gen_23_cmp_pReg_27, Q(26)=>gen_23_cmp_pReg_26, Q(25)=>
      gen_23_cmp_pReg_25, Q(24)=>gen_23_cmp_pReg_24, Q(23)=>
      gen_23_cmp_pReg_23, Q(22)=>gen_23_cmp_pReg_22, Q(21)=>
      gen_23_cmp_pReg_21, Q(20)=>gen_23_cmp_pReg_20, Q(19)=>
      gen_23_cmp_pReg_19, Q(18)=>gen_23_cmp_pReg_18, Q(17)=>
      gen_23_cmp_pReg_17, Q(16)=>gen_23_cmp_pReg_16, Q(15)=>
      gen_23_cmp_pReg_15, Q(14)=>gen_23_cmp_pReg_14, Q(13)=>
      gen_23_cmp_pReg_13, Q(12)=>gen_23_cmp_pReg_12, Q(11)=>
      gen_23_cmp_pReg_11, Q(10)=>gen_23_cmp_pReg_10, Q(9)=>gen_23_cmp_pReg_9, 
      Q(8)=>gen_23_cmp_pReg_8, Q(7)=>gen_23_cmp_pReg_7, Q(6)=>
      gen_23_cmp_pReg_6, Q(5)=>gen_23_cmp_pReg_5, Q(4)=>gen_23_cmp_pReg_4, 
      Q(3)=>gen_23_cmp_pReg_3, Q(2)=>gen_23_cmp_pReg_2, Q(1)=>
      gen_23_cmp_pReg_1, Q(0)=>gen_23_cmp_pReg_0);
   gen_23_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>gen_24_cmp_pInit_32, 
      a(31)=>gen_24_cmp_pInit_32, a(30)=>gen_23_cmp_pReg_30, a(29)=>
      gen_23_cmp_pReg_29, a(28)=>gen_23_cmp_pReg_28, a(27)=>
      gen_23_cmp_pReg_27, a(26)=>gen_23_cmp_pReg_26, a(25)=>
      gen_23_cmp_pReg_25, a(24)=>gen_23_cmp_pReg_24, a(23)=>
      gen_23_cmp_pReg_23, a(22)=>gen_23_cmp_pReg_22, a(21)=>
      gen_23_cmp_pReg_21, a(20)=>gen_23_cmp_pReg_20, a(19)=>
      gen_23_cmp_pReg_19, a(18)=>gen_23_cmp_pReg_18, a(17)=>
      gen_23_cmp_pReg_17, a(16)=>gen_23_cmp_pReg_16, a(15)=>
      gen_23_cmp_pReg_15, a(14)=>gen_23_cmp_pReg_14, a(13)=>
      gen_23_cmp_pReg_13, a(12)=>gen_23_cmp_pReg_12, a(11)=>
      gen_23_cmp_pReg_11, a(10)=>gen_23_cmp_pReg_10, a(9)=>gen_23_cmp_pReg_9, 
      a(8)=>gen_23_cmp_pReg_8, a(7)=>gen_23_cmp_pReg_7, a(6)=>
      gen_23_cmp_pReg_6, a(5)=>gen_23_cmp_pReg_5, a(4)=>gen_23_cmp_pReg_4, 
      a(3)=>gen_23_cmp_pReg_3, a(2)=>gen_23_cmp_pReg_2, a(1)=>
      gen_23_cmp_pReg_1, a(0)=>gen_23_cmp_pReg_0, b(32)=>gen_24_cmp_pInit_32, 
      b(31)=>gen_24_cmp_pInit_32, b(30)=>gen_24_cmp_pInit_32, b(29)=>
      gen_24_cmp_pInit_32, b(28)=>gen_24_cmp_pInit_32, b(27)=>
      gen_24_cmp_pInit_32, b(26)=>gen_24_cmp_pInit_32, b(25)=>
      gen_24_cmp_pInit_32, b(24)=>gen_24_cmp_pInit_32, b(23)=>
      gen_24_cmp_pInit_32, b(22)=>gen_24_cmp_pInit_32, b(21)=>
      gen_24_cmp_pInit_32, b(20)=>gen_24_cmp_pInit_32, b(19)=>
      gen_24_cmp_pInit_32, b(18)=>gen_24_cmp_pInit_32, b(17)=>
      gen_24_cmp_pInit_32, b(16)=>gen_24_cmp_pInit_32, b(15)=>
      gen_24_cmp_pInit_32, b(14)=>gen_24_cmp_pInit_32, b(13)=>
      gen_24_cmp_pInit_32, b(12)=>gen_24_cmp_pInit_32, b(11)=>
      gen_24_cmp_pInit_32, b(10)=>gen_24_cmp_pInit_32, b(9)=>
      gen_24_cmp_pInit_32, b(8)=>filter_23_7, b(7)=>filter_23_6, b(6)=>
      filter_23_5, b(5)=>filter_23_4, b(4)=>filter_23_3, b(3)=>filter_23_2, 
      b(2)=>filter_23_1, b(1)=>filter_23_0, b(0)=>gen_24_cmp_pInit_32, sel=>
      nx11896, f(32)=>DANGLING(7), f(31)=>DANGLING(8), f(30)=>
      gen_23_cmp_pMux_30, f(29)=>gen_23_cmp_pMux_29, f(28)=>
      gen_23_cmp_pMux_28, f(27)=>gen_23_cmp_pMux_27, f(26)=>
      gen_23_cmp_pMux_26, f(25)=>gen_23_cmp_pMux_25, f(24)=>
      gen_23_cmp_pMux_24, f(23)=>gen_23_cmp_pMux_23, f(22)=>
      gen_23_cmp_pMux_22, f(21)=>gen_23_cmp_pMux_21, f(20)=>
      gen_23_cmp_pMux_20, f(19)=>gen_23_cmp_pMux_19, f(18)=>
      gen_23_cmp_pMux_18, f(17)=>gen_23_cmp_pMux_17, f(16)=>
      gen_23_cmp_pMux_16, f(15)=>gen_23_cmp_pMux_15, f(14)=>
      gen_23_cmp_pMux_14, f(13)=>gen_23_cmp_pMux_13, f(12)=>
      gen_23_cmp_pMux_12, f(11)=>gen_23_cmp_pMux_11, f(10)=>
      gen_23_cmp_pMux_10, f(9)=>gen_23_cmp_pMux_9, f(8)=>gen_23_cmp_pMux_8, 
      f(7)=>gen_23_cmp_pMux_7, f(6)=>gen_23_cmp_pMux_6, f(5)=>
      gen_23_cmp_pMux_5, f(4)=>gen_23_cmp_pMux_4, f(3)=>gen_23_cmp_pMux_3, 
      f(2)=>gen_23_cmp_pMux_2, f(1)=>gen_23_cmp_pMux_1, f(0)=>
      gen_23_cmp_pMux_0);
   gen_23_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>
      gen_24_cmp_pInit_32, a(22)=>gen_24_cmp_pInit_32, a(21)=>
      gen_23_cmp_pMux_30, a(20)=>gen_23_cmp_pMux_29, a(19)=>
      gen_23_cmp_pMux_28, a(18)=>gen_23_cmp_pMux_27, a(17)=>
      gen_23_cmp_pMux_26, a(16)=>gen_23_cmp_pMux_25, a(15)=>
      gen_23_cmp_pMux_24, a(14)=>gen_23_cmp_pMux_23, a(13)=>
      gen_23_cmp_pMux_22, a(12)=>gen_23_cmp_pMux_21, a(11)=>
      gen_23_cmp_pMux_20, a(10)=>gen_23_cmp_pMux_19, a(9)=>
      gen_23_cmp_pMux_18, a(8)=>gen_23_cmp_pMux_17, a(7)=>gen_23_cmp_pMux_16, 
      a(6)=>gen_23_cmp_pMux_15, a(5)=>gen_23_cmp_pMux_14, a(4)=>
      gen_23_cmp_pMux_13, a(3)=>gen_23_cmp_pMux_12, a(2)=>gen_23_cmp_pMux_11, 
      a(1)=>gen_23_cmp_pMux_10, a(0)=>gen_23_cmp_pMux_9, b(23)=>nx10446, 
      b(22)=>nx10446, b(21)=>nx10444, b(20)=>nx10452, b(19)=>nx10450, b(18)
      =>nx10448, b(17)=>nx10446, b(16)=>nx10444, b(15)=>
      gen_23_cmp_BSCmp_op2_15, b(14)=>gen_23_cmp_BSCmp_op2_14, b(13)=>
      gen_23_cmp_BSCmp_op2_13, b(12)=>gen_23_cmp_BSCmp_op2_12, b(11)=>
      gen_23_cmp_BSCmp_op2_11, b(10)=>gen_23_cmp_BSCmp_op2_10, b(9)=>
      gen_23_cmp_BSCmp_op2_9, b(8)=>gen_23_cmp_BSCmp_op2_8, b(7)=>
      gen_23_cmp_BSCmp_op2_7, b(6)=>gen_23_cmp_BSCmp_op2_6, b(5)=>
      gen_23_cmp_BSCmp_op2_5, b(4)=>gen_23_cmp_BSCmp_op2_4, b(3)=>
      gen_23_cmp_BSCmp_op2_3, b(2)=>gen_23_cmp_BSCmp_op2_2, b(1)=>
      gen_23_cmp_BSCmp_op2_1, b(0)=>gen_23_cmp_BSCmp_op2_0, carryIn=>
      gen_23_cmp_BSCmp_carryIn, sum(23)=>gen_23_cmp_pBs_30, sum(22)=>
      gen_23_cmp_pBs_29, sum(21)=>gen_23_cmp_pBs_28, sum(20)=>
      gen_23_cmp_pBs_27, sum(19)=>gen_23_cmp_pBs_26, sum(18)=>
      gen_23_cmp_pBs_25, sum(17)=>gen_23_cmp_pBs_24, sum(16)=>
      gen_23_cmp_pBs_23, sum(15)=>outputs_23_15, sum(14)=>outputs_23_14, 
      sum(13)=>outputs_23_13, sum(12)=>outputs_23_12, sum(11)=>outputs_23_11, 
      sum(10)=>outputs_23_10, sum(9)=>outputs_23_9, sum(8)=>outputs_23_8, 
      sum(7)=>outputs_23_7, sum(6)=>outputs_23_6, sum(5)=>outputs_23_5, 
      sum(4)=>outputs_23_4, sum(3)=>outputs_23_3, sum(2)=>outputs_23_2, 
      sum(1)=>outputs_23_1, sum(0)=>outputs_23_0, carryOut=>DANGLING(9));
   gen_22_cmp_pRegCmp : Reg_33 port map ( D(32)=>gen_24_cmp_pInit_32, D(31)
      =>gen_24_cmp_pInit_32, D(30)=>gen_22_cmp_pBs_30, D(29)=>
      gen_22_cmp_pBs_29, D(28)=>gen_22_cmp_pBs_28, D(27)=>gen_22_cmp_pBs_27, 
      D(26)=>gen_22_cmp_pBs_26, D(25)=>gen_22_cmp_pBs_25, D(24)=>
      gen_22_cmp_pBs_24, D(23)=>gen_22_cmp_pBs_23, D(22)=>outputs_22_15, 
      D(21)=>outputs_22_14, D(20)=>outputs_22_13, D(19)=>outputs_22_12, 
      D(18)=>outputs_22_11, D(17)=>outputs_22_10, D(16)=>outputs_22_9, D(15)
      =>outputs_22_8, D(14)=>outputs_22_7, D(13)=>outputs_22_6, D(12)=>
      outputs_22_5, D(11)=>outputs_22_4, D(10)=>outputs_22_3, D(9)=>
      outputs_22_2, D(8)=>outputs_22_1, D(7)=>outputs_22_0, D(6)=>
      gen_22_cmp_pMux_8, D(5)=>gen_22_cmp_pMux_7, D(4)=>gen_22_cmp_pMux_6, 
      D(3)=>gen_22_cmp_pMux_5, D(2)=>gen_22_cmp_pMux_4, D(1)=>
      gen_22_cmp_pMux_3, D(0)=>nx10154, en=>nx11916, clk=>nx10122, rst=>rst, 
      Q(32)=>DANGLING(10), Q(31)=>DANGLING(11), Q(30)=>gen_22_cmp_pReg_30, 
      Q(29)=>gen_22_cmp_pReg_29, Q(28)=>gen_22_cmp_pReg_28, Q(27)=>
      gen_22_cmp_pReg_27, Q(26)=>gen_22_cmp_pReg_26, Q(25)=>
      gen_22_cmp_pReg_25, Q(24)=>gen_22_cmp_pReg_24, Q(23)=>
      gen_22_cmp_pReg_23, Q(22)=>gen_22_cmp_pReg_22, Q(21)=>
      gen_22_cmp_pReg_21, Q(20)=>gen_22_cmp_pReg_20, Q(19)=>
      gen_22_cmp_pReg_19, Q(18)=>gen_22_cmp_pReg_18, Q(17)=>
      gen_22_cmp_pReg_17, Q(16)=>gen_22_cmp_pReg_16, Q(15)=>
      gen_22_cmp_pReg_15, Q(14)=>gen_22_cmp_pReg_14, Q(13)=>
      gen_22_cmp_pReg_13, Q(12)=>gen_22_cmp_pReg_12, Q(11)=>
      gen_22_cmp_pReg_11, Q(10)=>gen_22_cmp_pReg_10, Q(9)=>gen_22_cmp_pReg_9, 
      Q(8)=>gen_22_cmp_pReg_8, Q(7)=>gen_22_cmp_pReg_7, Q(6)=>
      gen_22_cmp_pReg_6, Q(5)=>gen_22_cmp_pReg_5, Q(4)=>gen_22_cmp_pReg_4, 
      Q(3)=>gen_22_cmp_pReg_3, Q(2)=>gen_22_cmp_pReg_2, Q(1)=>
      gen_22_cmp_pReg_1, Q(0)=>gen_22_cmp_pReg_0);
   gen_22_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>gen_24_cmp_pInit_32, 
      a(31)=>gen_24_cmp_pInit_32, a(30)=>gen_22_cmp_pReg_30, a(29)=>
      gen_22_cmp_pReg_29, a(28)=>gen_22_cmp_pReg_28, a(27)=>
      gen_22_cmp_pReg_27, a(26)=>gen_22_cmp_pReg_26, a(25)=>
      gen_22_cmp_pReg_25, a(24)=>gen_22_cmp_pReg_24, a(23)=>
      gen_22_cmp_pReg_23, a(22)=>gen_22_cmp_pReg_22, a(21)=>
      gen_22_cmp_pReg_21, a(20)=>gen_22_cmp_pReg_20, a(19)=>
      gen_22_cmp_pReg_19, a(18)=>gen_22_cmp_pReg_18, a(17)=>
      gen_22_cmp_pReg_17, a(16)=>gen_22_cmp_pReg_16, a(15)=>
      gen_22_cmp_pReg_15, a(14)=>gen_22_cmp_pReg_14, a(13)=>
      gen_22_cmp_pReg_13, a(12)=>gen_22_cmp_pReg_12, a(11)=>
      gen_22_cmp_pReg_11, a(10)=>gen_22_cmp_pReg_10, a(9)=>gen_22_cmp_pReg_9, 
      a(8)=>gen_22_cmp_pReg_8, a(7)=>gen_22_cmp_pReg_7, a(6)=>
      gen_22_cmp_pReg_6, a(5)=>gen_22_cmp_pReg_5, a(4)=>gen_22_cmp_pReg_4, 
      a(3)=>gen_22_cmp_pReg_3, a(2)=>gen_22_cmp_pReg_2, a(1)=>
      gen_22_cmp_pReg_1, a(0)=>gen_22_cmp_pReg_0, b(32)=>gen_24_cmp_pInit_32, 
      b(31)=>gen_24_cmp_pInit_32, b(30)=>gen_24_cmp_pInit_32, b(29)=>
      gen_24_cmp_pInit_32, b(28)=>gen_24_cmp_pInit_32, b(27)=>
      gen_24_cmp_pInit_32, b(26)=>gen_24_cmp_pInit_32, b(25)=>
      gen_24_cmp_pInit_32, b(24)=>gen_24_cmp_pInit_32, b(23)=>
      gen_24_cmp_pInit_32, b(22)=>gen_24_cmp_pInit_32, b(21)=>
      gen_24_cmp_pInit_32, b(20)=>gen_24_cmp_pInit_32, b(19)=>
      gen_24_cmp_pInit_32, b(18)=>gen_24_cmp_pInit_32, b(17)=>
      gen_24_cmp_pInit_32, b(16)=>gen_24_cmp_pInit_32, b(15)=>
      gen_24_cmp_pInit_32, b(14)=>gen_24_cmp_pInit_32, b(13)=>
      gen_24_cmp_pInit_32, b(12)=>gen_24_cmp_pInit_32, b(11)=>
      gen_24_cmp_pInit_32, b(10)=>gen_24_cmp_pInit_32, b(9)=>
      gen_24_cmp_pInit_32, b(8)=>filter_22_7, b(7)=>filter_22_6, b(6)=>
      filter_22_5, b(5)=>filter_22_4, b(4)=>filter_22_3, b(3)=>filter_22_2, 
      b(2)=>filter_22_1, b(1)=>filter_22_0, b(0)=>gen_24_cmp_pInit_32, sel=>
      nx11896, f(32)=>DANGLING(12), f(31)=>DANGLING(13), f(30)=>
      gen_22_cmp_pMux_30, f(29)=>gen_22_cmp_pMux_29, f(28)=>
      gen_22_cmp_pMux_28, f(27)=>gen_22_cmp_pMux_27, f(26)=>
      gen_22_cmp_pMux_26, f(25)=>gen_22_cmp_pMux_25, f(24)=>
      gen_22_cmp_pMux_24, f(23)=>gen_22_cmp_pMux_23, f(22)=>
      gen_22_cmp_pMux_22, f(21)=>gen_22_cmp_pMux_21, f(20)=>
      gen_22_cmp_pMux_20, f(19)=>gen_22_cmp_pMux_19, f(18)=>
      gen_22_cmp_pMux_18, f(17)=>gen_22_cmp_pMux_17, f(16)=>
      gen_22_cmp_pMux_16, f(15)=>gen_22_cmp_pMux_15, f(14)=>
      gen_22_cmp_pMux_14, f(13)=>gen_22_cmp_pMux_13, f(12)=>
      gen_22_cmp_pMux_12, f(11)=>gen_22_cmp_pMux_11, f(10)=>
      gen_22_cmp_pMux_10, f(9)=>gen_22_cmp_pMux_9, f(8)=>gen_22_cmp_pMux_8, 
      f(7)=>gen_22_cmp_pMux_7, f(6)=>gen_22_cmp_pMux_6, f(5)=>
      gen_22_cmp_pMux_5, f(4)=>gen_22_cmp_pMux_4, f(3)=>gen_22_cmp_pMux_3, 
      f(2)=>gen_22_cmp_pMux_2, f(1)=>gen_22_cmp_pMux_1, f(0)=>
      gen_22_cmp_pMux_0);
   gen_22_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>
      gen_24_cmp_pInit_32, a(22)=>gen_24_cmp_pInit_32, a(21)=>
      gen_22_cmp_pMux_30, a(20)=>gen_22_cmp_pMux_29, a(19)=>
      gen_22_cmp_pMux_28, a(18)=>gen_22_cmp_pMux_27, a(17)=>
      gen_22_cmp_pMux_26, a(16)=>gen_22_cmp_pMux_25, a(15)=>
      gen_22_cmp_pMux_24, a(14)=>gen_22_cmp_pMux_23, a(13)=>
      gen_22_cmp_pMux_22, a(12)=>gen_22_cmp_pMux_21, a(11)=>
      gen_22_cmp_pMux_20, a(10)=>gen_22_cmp_pMux_19, a(9)=>
      gen_22_cmp_pMux_18, a(8)=>gen_22_cmp_pMux_17, a(7)=>gen_22_cmp_pMux_16, 
      a(6)=>gen_22_cmp_pMux_15, a(5)=>gen_22_cmp_pMux_14, a(4)=>
      gen_22_cmp_pMux_13, a(3)=>gen_22_cmp_pMux_12, a(2)=>gen_22_cmp_pMux_11, 
      a(1)=>gen_22_cmp_pMux_10, a(0)=>gen_22_cmp_pMux_9, b(23)=>nx10458, 
      b(22)=>nx10458, b(21)=>nx10456, b(20)=>nx10464, b(19)=>nx10462, b(18)
      =>nx10460, b(17)=>nx10458, b(16)=>nx10456, b(15)=>
      gen_22_cmp_BSCmp_op2_15, b(14)=>gen_22_cmp_BSCmp_op2_14, b(13)=>
      gen_22_cmp_BSCmp_op2_13, b(12)=>gen_22_cmp_BSCmp_op2_12, b(11)=>
      gen_22_cmp_BSCmp_op2_11, b(10)=>gen_22_cmp_BSCmp_op2_10, b(9)=>
      gen_22_cmp_BSCmp_op2_9, b(8)=>gen_22_cmp_BSCmp_op2_8, b(7)=>
      gen_22_cmp_BSCmp_op2_7, b(6)=>gen_22_cmp_BSCmp_op2_6, b(5)=>
      gen_22_cmp_BSCmp_op2_5, b(4)=>gen_22_cmp_BSCmp_op2_4, b(3)=>
      gen_22_cmp_BSCmp_op2_3, b(2)=>gen_22_cmp_BSCmp_op2_2, b(1)=>
      gen_22_cmp_BSCmp_op2_1, b(0)=>gen_22_cmp_BSCmp_op2_0, carryIn=>
      gen_22_cmp_BSCmp_carryIn, sum(23)=>gen_22_cmp_pBs_30, sum(22)=>
      gen_22_cmp_pBs_29, sum(21)=>gen_22_cmp_pBs_28, sum(20)=>
      gen_22_cmp_pBs_27, sum(19)=>gen_22_cmp_pBs_26, sum(18)=>
      gen_22_cmp_pBs_25, sum(17)=>gen_22_cmp_pBs_24, sum(16)=>
      gen_22_cmp_pBs_23, sum(15)=>outputs_22_15, sum(14)=>outputs_22_14, 
      sum(13)=>outputs_22_13, sum(12)=>outputs_22_12, sum(11)=>outputs_22_11, 
      sum(10)=>outputs_22_10, sum(9)=>outputs_22_9, sum(8)=>outputs_22_8, 
      sum(7)=>outputs_22_7, sum(6)=>outputs_22_6, sum(5)=>outputs_22_5, 
      sum(4)=>outputs_22_4, sum(3)=>outputs_22_3, sum(2)=>outputs_22_2, 
      sum(1)=>outputs_22_1, sum(0)=>outputs_22_0, carryOut=>DANGLING(14));
   gen_21_cmp_pRegCmp : Reg_33 port map ( D(32)=>gen_24_cmp_pInit_32, D(31)
      =>gen_24_cmp_pInit_32, D(30)=>gen_21_cmp_pBs_30, D(29)=>
      gen_21_cmp_pBs_29, D(28)=>gen_21_cmp_pBs_28, D(27)=>gen_21_cmp_pBs_27, 
      D(26)=>gen_21_cmp_pBs_26, D(25)=>gen_21_cmp_pBs_25, D(24)=>
      gen_21_cmp_pBs_24, D(23)=>gen_21_cmp_pBs_23, D(22)=>outputs_21_15, 
      D(21)=>outputs_21_14, D(20)=>outputs_21_13, D(19)=>outputs_21_12, 
      D(18)=>outputs_21_11, D(17)=>outputs_21_10, D(16)=>outputs_21_9, D(15)
      =>outputs_21_8, D(14)=>outputs_21_7, D(13)=>outputs_21_6, D(12)=>
      outputs_21_5, D(11)=>outputs_21_4, D(10)=>outputs_21_3, D(9)=>
      outputs_21_2, D(8)=>outputs_21_1, D(7)=>outputs_21_0, D(6)=>
      gen_21_cmp_pMux_8, D(5)=>gen_21_cmp_pMux_7, D(4)=>gen_21_cmp_pMux_6, 
      D(3)=>gen_21_cmp_pMux_5, D(2)=>gen_21_cmp_pMux_4, D(1)=>
      gen_21_cmp_pMux_3, D(0)=>nx10166, en=>nx11918, clk=>nx10122, rst=>rst, 
      Q(32)=>DANGLING(15), Q(31)=>DANGLING(16), Q(30)=>gen_21_cmp_pReg_30, 
      Q(29)=>gen_21_cmp_pReg_29, Q(28)=>gen_21_cmp_pReg_28, Q(27)=>
      gen_21_cmp_pReg_27, Q(26)=>gen_21_cmp_pReg_26, Q(25)=>
      gen_21_cmp_pReg_25, Q(24)=>gen_21_cmp_pReg_24, Q(23)=>
      gen_21_cmp_pReg_23, Q(22)=>gen_21_cmp_pReg_22, Q(21)=>
      gen_21_cmp_pReg_21, Q(20)=>gen_21_cmp_pReg_20, Q(19)=>
      gen_21_cmp_pReg_19, Q(18)=>gen_21_cmp_pReg_18, Q(17)=>
      gen_21_cmp_pReg_17, Q(16)=>gen_21_cmp_pReg_16, Q(15)=>
      gen_21_cmp_pReg_15, Q(14)=>gen_21_cmp_pReg_14, Q(13)=>
      gen_21_cmp_pReg_13, Q(12)=>gen_21_cmp_pReg_12, Q(11)=>
      gen_21_cmp_pReg_11, Q(10)=>gen_21_cmp_pReg_10, Q(9)=>gen_21_cmp_pReg_9, 
      Q(8)=>gen_21_cmp_pReg_8, Q(7)=>gen_21_cmp_pReg_7, Q(6)=>
      gen_21_cmp_pReg_6, Q(5)=>gen_21_cmp_pReg_5, Q(4)=>gen_21_cmp_pReg_4, 
      Q(3)=>gen_21_cmp_pReg_3, Q(2)=>gen_21_cmp_pReg_2, Q(1)=>
      gen_21_cmp_pReg_1, Q(0)=>gen_21_cmp_pReg_0);
   gen_21_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>gen_24_cmp_pInit_32, 
      a(31)=>gen_24_cmp_pInit_32, a(30)=>gen_21_cmp_pReg_30, a(29)=>
      gen_21_cmp_pReg_29, a(28)=>gen_21_cmp_pReg_28, a(27)=>
      gen_21_cmp_pReg_27, a(26)=>gen_21_cmp_pReg_26, a(25)=>
      gen_21_cmp_pReg_25, a(24)=>gen_21_cmp_pReg_24, a(23)=>
      gen_21_cmp_pReg_23, a(22)=>gen_21_cmp_pReg_22, a(21)=>
      gen_21_cmp_pReg_21, a(20)=>gen_21_cmp_pReg_20, a(19)=>
      gen_21_cmp_pReg_19, a(18)=>gen_21_cmp_pReg_18, a(17)=>
      gen_21_cmp_pReg_17, a(16)=>gen_21_cmp_pReg_16, a(15)=>
      gen_21_cmp_pReg_15, a(14)=>gen_21_cmp_pReg_14, a(13)=>
      gen_21_cmp_pReg_13, a(12)=>gen_21_cmp_pReg_12, a(11)=>
      gen_21_cmp_pReg_11, a(10)=>gen_21_cmp_pReg_10, a(9)=>gen_21_cmp_pReg_9, 
      a(8)=>gen_21_cmp_pReg_8, a(7)=>gen_21_cmp_pReg_7, a(6)=>
      gen_21_cmp_pReg_6, a(5)=>gen_21_cmp_pReg_5, a(4)=>gen_21_cmp_pReg_4, 
      a(3)=>gen_21_cmp_pReg_3, a(2)=>gen_21_cmp_pReg_2, a(1)=>
      gen_21_cmp_pReg_1, a(0)=>gen_21_cmp_pReg_0, b(32)=>gen_24_cmp_pInit_32, 
      b(31)=>gen_24_cmp_pInit_32, b(30)=>gen_24_cmp_pInit_32, b(29)=>
      gen_24_cmp_pInit_32, b(28)=>gen_24_cmp_pInit_32, b(27)=>
      gen_24_cmp_pInit_32, b(26)=>gen_24_cmp_pInit_32, b(25)=>
      gen_24_cmp_pInit_32, b(24)=>gen_24_cmp_pInit_32, b(23)=>
      gen_24_cmp_pInit_32, b(22)=>gen_24_cmp_pInit_32, b(21)=>
      gen_24_cmp_pInit_32, b(20)=>gen_24_cmp_pInit_32, b(19)=>
      gen_24_cmp_pInit_32, b(18)=>gen_24_cmp_pInit_32, b(17)=>
      gen_24_cmp_pInit_32, b(16)=>gen_24_cmp_pInit_32, b(15)=>
      gen_24_cmp_pInit_32, b(14)=>gen_24_cmp_pInit_32, b(13)=>
      gen_24_cmp_pInit_32, b(12)=>gen_24_cmp_pInit_32, b(11)=>
      gen_24_cmp_pInit_32, b(10)=>gen_24_cmp_pInit_32, b(9)=>
      gen_24_cmp_pInit_32, b(8)=>filter_21_7, b(7)=>filter_21_6, b(6)=>
      filter_21_5, b(5)=>filter_21_4, b(4)=>filter_21_3, b(3)=>filter_21_2, 
      b(2)=>filter_21_1, b(1)=>filter_21_0, b(0)=>gen_24_cmp_pInit_32, sel=>
      nx11898, f(32)=>DANGLING(17), f(31)=>DANGLING(18), f(30)=>
      gen_21_cmp_pMux_30, f(29)=>gen_21_cmp_pMux_29, f(28)=>
      gen_21_cmp_pMux_28, f(27)=>gen_21_cmp_pMux_27, f(26)=>
      gen_21_cmp_pMux_26, f(25)=>gen_21_cmp_pMux_25, f(24)=>
      gen_21_cmp_pMux_24, f(23)=>gen_21_cmp_pMux_23, f(22)=>
      gen_21_cmp_pMux_22, f(21)=>gen_21_cmp_pMux_21, f(20)=>
      gen_21_cmp_pMux_20, f(19)=>gen_21_cmp_pMux_19, f(18)=>
      gen_21_cmp_pMux_18, f(17)=>gen_21_cmp_pMux_17, f(16)=>
      gen_21_cmp_pMux_16, f(15)=>gen_21_cmp_pMux_15, f(14)=>
      gen_21_cmp_pMux_14, f(13)=>gen_21_cmp_pMux_13, f(12)=>
      gen_21_cmp_pMux_12, f(11)=>gen_21_cmp_pMux_11, f(10)=>
      gen_21_cmp_pMux_10, f(9)=>gen_21_cmp_pMux_9, f(8)=>gen_21_cmp_pMux_8, 
      f(7)=>gen_21_cmp_pMux_7, f(6)=>gen_21_cmp_pMux_6, f(5)=>
      gen_21_cmp_pMux_5, f(4)=>gen_21_cmp_pMux_4, f(3)=>gen_21_cmp_pMux_3, 
      f(2)=>gen_21_cmp_pMux_2, f(1)=>gen_21_cmp_pMux_1, f(0)=>
      gen_21_cmp_pMux_0);
   gen_21_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>
      gen_24_cmp_pInit_32, a(22)=>gen_24_cmp_pInit_32, a(21)=>
      gen_21_cmp_pMux_30, a(20)=>gen_21_cmp_pMux_29, a(19)=>
      gen_21_cmp_pMux_28, a(18)=>gen_21_cmp_pMux_27, a(17)=>
      gen_21_cmp_pMux_26, a(16)=>gen_21_cmp_pMux_25, a(15)=>
      gen_21_cmp_pMux_24, a(14)=>gen_21_cmp_pMux_23, a(13)=>
      gen_21_cmp_pMux_22, a(12)=>gen_21_cmp_pMux_21, a(11)=>
      gen_21_cmp_pMux_20, a(10)=>gen_21_cmp_pMux_19, a(9)=>
      gen_21_cmp_pMux_18, a(8)=>gen_21_cmp_pMux_17, a(7)=>gen_21_cmp_pMux_16, 
      a(6)=>gen_21_cmp_pMux_15, a(5)=>gen_21_cmp_pMux_14, a(4)=>
      gen_21_cmp_pMux_13, a(3)=>gen_21_cmp_pMux_12, a(2)=>gen_21_cmp_pMux_11, 
      a(1)=>gen_21_cmp_pMux_10, a(0)=>gen_21_cmp_pMux_9, b(23)=>nx10470, 
      b(22)=>nx10470, b(21)=>nx10468, b(20)=>nx10476, b(19)=>nx10474, b(18)
      =>nx10472, b(17)=>nx10470, b(16)=>nx10468, b(15)=>
      gen_21_cmp_BSCmp_op2_15, b(14)=>gen_21_cmp_BSCmp_op2_14, b(13)=>
      gen_21_cmp_BSCmp_op2_13, b(12)=>gen_21_cmp_BSCmp_op2_12, b(11)=>
      gen_21_cmp_BSCmp_op2_11, b(10)=>gen_21_cmp_BSCmp_op2_10, b(9)=>
      gen_21_cmp_BSCmp_op2_9, b(8)=>gen_21_cmp_BSCmp_op2_8, b(7)=>
      gen_21_cmp_BSCmp_op2_7, b(6)=>gen_21_cmp_BSCmp_op2_6, b(5)=>
      gen_21_cmp_BSCmp_op2_5, b(4)=>gen_21_cmp_BSCmp_op2_4, b(3)=>
      gen_21_cmp_BSCmp_op2_3, b(2)=>gen_21_cmp_BSCmp_op2_2, b(1)=>
      gen_21_cmp_BSCmp_op2_1, b(0)=>gen_21_cmp_BSCmp_op2_0, carryIn=>
      gen_21_cmp_BSCmp_carryIn, sum(23)=>gen_21_cmp_pBs_30, sum(22)=>
      gen_21_cmp_pBs_29, sum(21)=>gen_21_cmp_pBs_28, sum(20)=>
      gen_21_cmp_pBs_27, sum(19)=>gen_21_cmp_pBs_26, sum(18)=>
      gen_21_cmp_pBs_25, sum(17)=>gen_21_cmp_pBs_24, sum(16)=>
      gen_21_cmp_pBs_23, sum(15)=>outputs_21_15, sum(14)=>outputs_21_14, 
      sum(13)=>outputs_21_13, sum(12)=>outputs_21_12, sum(11)=>outputs_21_11, 
      sum(10)=>outputs_21_10, sum(9)=>outputs_21_9, sum(8)=>outputs_21_8, 
      sum(7)=>outputs_21_7, sum(6)=>outputs_21_6, sum(5)=>outputs_21_5, 
      sum(4)=>outputs_21_4, sum(3)=>outputs_21_3, sum(2)=>outputs_21_2, 
      sum(1)=>outputs_21_1, sum(0)=>outputs_21_0, carryOut=>DANGLING(19));
   gen_20_cmp_pRegCmp : Reg_33 port map ( D(32)=>gen_24_cmp_pInit_32, D(31)
      =>gen_24_cmp_pInit_32, D(30)=>gen_20_cmp_pBs_30, D(29)=>
      gen_20_cmp_pBs_29, D(28)=>gen_20_cmp_pBs_28, D(27)=>gen_20_cmp_pBs_27, 
      D(26)=>gen_20_cmp_pBs_26, D(25)=>gen_20_cmp_pBs_25, D(24)=>
      gen_20_cmp_pBs_24, D(23)=>gen_20_cmp_pBs_23, D(22)=>outputs_20_15, 
      D(21)=>outputs_20_14, D(20)=>outputs_20_13, D(19)=>outputs_20_12, 
      D(18)=>outputs_20_11, D(17)=>outputs_20_10, D(16)=>outputs_20_9, D(15)
      =>outputs_20_8, D(14)=>outputs_20_7, D(13)=>outputs_20_6, D(12)=>
      outputs_20_5, D(11)=>outputs_20_4, D(10)=>outputs_20_3, D(9)=>
      outputs_20_2, D(8)=>outputs_20_1, D(7)=>outputs_20_0, D(6)=>
      gen_20_cmp_pMux_8, D(5)=>gen_20_cmp_pMux_7, D(4)=>gen_20_cmp_pMux_6, 
      D(3)=>gen_20_cmp_pMux_5, D(2)=>gen_20_cmp_pMux_4, D(1)=>
      gen_20_cmp_pMux_3, D(0)=>nx10178, en=>nx11918, clk=>nx10122, rst=>rst, 
      Q(32)=>DANGLING(20), Q(31)=>DANGLING(21), Q(30)=>gen_20_cmp_pReg_30, 
      Q(29)=>gen_20_cmp_pReg_29, Q(28)=>gen_20_cmp_pReg_28, Q(27)=>
      gen_20_cmp_pReg_27, Q(26)=>gen_20_cmp_pReg_26, Q(25)=>
      gen_20_cmp_pReg_25, Q(24)=>gen_20_cmp_pReg_24, Q(23)=>
      gen_20_cmp_pReg_23, Q(22)=>gen_20_cmp_pReg_22, Q(21)=>
      gen_20_cmp_pReg_21, Q(20)=>gen_20_cmp_pReg_20, Q(19)=>
      gen_20_cmp_pReg_19, Q(18)=>gen_20_cmp_pReg_18, Q(17)=>
      gen_20_cmp_pReg_17, Q(16)=>gen_20_cmp_pReg_16, Q(15)=>
      gen_20_cmp_pReg_15, Q(14)=>gen_20_cmp_pReg_14, Q(13)=>
      gen_20_cmp_pReg_13, Q(12)=>gen_20_cmp_pReg_12, Q(11)=>
      gen_20_cmp_pReg_11, Q(10)=>gen_20_cmp_pReg_10, Q(9)=>gen_20_cmp_pReg_9, 
      Q(8)=>gen_20_cmp_pReg_8, Q(7)=>gen_20_cmp_pReg_7, Q(6)=>
      gen_20_cmp_pReg_6, Q(5)=>gen_20_cmp_pReg_5, Q(4)=>gen_20_cmp_pReg_4, 
      Q(3)=>gen_20_cmp_pReg_3, Q(2)=>gen_20_cmp_pReg_2, Q(1)=>
      gen_20_cmp_pReg_1, Q(0)=>gen_20_cmp_pReg_0);
   gen_20_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>gen_24_cmp_pInit_32, 
      a(31)=>gen_24_cmp_pInit_32, a(30)=>gen_20_cmp_pReg_30, a(29)=>
      gen_20_cmp_pReg_29, a(28)=>gen_20_cmp_pReg_28, a(27)=>
      gen_20_cmp_pReg_27, a(26)=>gen_20_cmp_pReg_26, a(25)=>
      gen_20_cmp_pReg_25, a(24)=>gen_20_cmp_pReg_24, a(23)=>
      gen_20_cmp_pReg_23, a(22)=>gen_20_cmp_pReg_22, a(21)=>
      gen_20_cmp_pReg_21, a(20)=>gen_20_cmp_pReg_20, a(19)=>
      gen_20_cmp_pReg_19, a(18)=>gen_20_cmp_pReg_18, a(17)=>
      gen_20_cmp_pReg_17, a(16)=>gen_20_cmp_pReg_16, a(15)=>
      gen_20_cmp_pReg_15, a(14)=>gen_20_cmp_pReg_14, a(13)=>
      gen_20_cmp_pReg_13, a(12)=>gen_20_cmp_pReg_12, a(11)=>
      gen_20_cmp_pReg_11, a(10)=>gen_20_cmp_pReg_10, a(9)=>gen_20_cmp_pReg_9, 
      a(8)=>gen_20_cmp_pReg_8, a(7)=>gen_20_cmp_pReg_7, a(6)=>
      gen_20_cmp_pReg_6, a(5)=>gen_20_cmp_pReg_5, a(4)=>gen_20_cmp_pReg_4, 
      a(3)=>gen_20_cmp_pReg_3, a(2)=>gen_20_cmp_pReg_2, a(1)=>
      gen_20_cmp_pReg_1, a(0)=>gen_20_cmp_pReg_0, b(32)=>gen_24_cmp_pInit_32, 
      b(31)=>gen_24_cmp_pInit_32, b(30)=>gen_24_cmp_pInit_32, b(29)=>
      gen_24_cmp_pInit_32, b(28)=>gen_24_cmp_pInit_32, b(27)=>
      gen_24_cmp_pInit_32, b(26)=>gen_24_cmp_pInit_32, b(25)=>
      gen_24_cmp_pInit_32, b(24)=>gen_24_cmp_pInit_32, b(23)=>
      gen_24_cmp_pInit_32, b(22)=>gen_24_cmp_pInit_32, b(21)=>
      gen_24_cmp_pInit_32, b(20)=>gen_24_cmp_pInit_32, b(19)=>
      gen_24_cmp_pInit_32, b(18)=>gen_24_cmp_pInit_32, b(17)=>
      gen_24_cmp_pInit_32, b(16)=>gen_24_cmp_pInit_32, b(15)=>
      gen_24_cmp_pInit_32, b(14)=>gen_24_cmp_pInit_32, b(13)=>
      gen_24_cmp_pInit_32, b(12)=>gen_24_cmp_pInit_32, b(11)=>
      gen_24_cmp_pInit_32, b(10)=>gen_24_cmp_pInit_32, b(9)=>
      gen_24_cmp_pInit_32, b(8)=>filter_20_7, b(7)=>filter_20_6, b(6)=>
      filter_20_5, b(5)=>filter_20_4, b(4)=>filter_20_3, b(3)=>filter_20_2, 
      b(2)=>filter_20_1, b(1)=>filter_20_0, b(0)=>gen_24_cmp_pInit_32, sel=>
      nx11898, f(32)=>DANGLING(22), f(31)=>DANGLING(23), f(30)=>
      gen_20_cmp_pMux_30, f(29)=>gen_20_cmp_pMux_29, f(28)=>
      gen_20_cmp_pMux_28, f(27)=>gen_20_cmp_pMux_27, f(26)=>
      gen_20_cmp_pMux_26, f(25)=>gen_20_cmp_pMux_25, f(24)=>
      gen_20_cmp_pMux_24, f(23)=>gen_20_cmp_pMux_23, f(22)=>
      gen_20_cmp_pMux_22, f(21)=>gen_20_cmp_pMux_21, f(20)=>
      gen_20_cmp_pMux_20, f(19)=>gen_20_cmp_pMux_19, f(18)=>
      gen_20_cmp_pMux_18, f(17)=>gen_20_cmp_pMux_17, f(16)=>
      gen_20_cmp_pMux_16, f(15)=>gen_20_cmp_pMux_15, f(14)=>
      gen_20_cmp_pMux_14, f(13)=>gen_20_cmp_pMux_13, f(12)=>
      gen_20_cmp_pMux_12, f(11)=>gen_20_cmp_pMux_11, f(10)=>
      gen_20_cmp_pMux_10, f(9)=>gen_20_cmp_pMux_9, f(8)=>gen_20_cmp_pMux_8, 
      f(7)=>gen_20_cmp_pMux_7, f(6)=>gen_20_cmp_pMux_6, f(5)=>
      gen_20_cmp_pMux_5, f(4)=>gen_20_cmp_pMux_4, f(3)=>gen_20_cmp_pMux_3, 
      f(2)=>gen_20_cmp_pMux_2, f(1)=>gen_20_cmp_pMux_1, f(0)=>
      gen_20_cmp_pMux_0);
   gen_20_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>
      gen_24_cmp_pInit_32, a(22)=>gen_24_cmp_pInit_32, a(21)=>
      gen_20_cmp_pMux_30, a(20)=>gen_20_cmp_pMux_29, a(19)=>
      gen_20_cmp_pMux_28, a(18)=>gen_20_cmp_pMux_27, a(17)=>
      gen_20_cmp_pMux_26, a(16)=>gen_20_cmp_pMux_25, a(15)=>
      gen_20_cmp_pMux_24, a(14)=>gen_20_cmp_pMux_23, a(13)=>
      gen_20_cmp_pMux_22, a(12)=>gen_20_cmp_pMux_21, a(11)=>
      gen_20_cmp_pMux_20, a(10)=>gen_20_cmp_pMux_19, a(9)=>
      gen_20_cmp_pMux_18, a(8)=>gen_20_cmp_pMux_17, a(7)=>gen_20_cmp_pMux_16, 
      a(6)=>gen_20_cmp_pMux_15, a(5)=>gen_20_cmp_pMux_14, a(4)=>
      gen_20_cmp_pMux_13, a(3)=>gen_20_cmp_pMux_12, a(2)=>gen_20_cmp_pMux_11, 
      a(1)=>gen_20_cmp_pMux_10, a(0)=>gen_20_cmp_pMux_9, b(23)=>nx10482, 
      b(22)=>nx10482, b(21)=>nx10480, b(20)=>nx10488, b(19)=>nx10486, b(18)
      =>nx10484, b(17)=>nx10482, b(16)=>nx10480, b(15)=>
      gen_20_cmp_BSCmp_op2_15, b(14)=>gen_20_cmp_BSCmp_op2_14, b(13)=>
      gen_20_cmp_BSCmp_op2_13, b(12)=>gen_20_cmp_BSCmp_op2_12, b(11)=>
      gen_20_cmp_BSCmp_op2_11, b(10)=>gen_20_cmp_BSCmp_op2_10, b(9)=>
      gen_20_cmp_BSCmp_op2_9, b(8)=>gen_20_cmp_BSCmp_op2_8, b(7)=>
      gen_20_cmp_BSCmp_op2_7, b(6)=>gen_20_cmp_BSCmp_op2_6, b(5)=>
      gen_20_cmp_BSCmp_op2_5, b(4)=>gen_20_cmp_BSCmp_op2_4, b(3)=>
      gen_20_cmp_BSCmp_op2_3, b(2)=>gen_20_cmp_BSCmp_op2_2, b(1)=>
      gen_20_cmp_BSCmp_op2_1, b(0)=>gen_20_cmp_BSCmp_op2_0, carryIn=>
      gen_20_cmp_BSCmp_carryIn, sum(23)=>gen_20_cmp_pBs_30, sum(22)=>
      gen_20_cmp_pBs_29, sum(21)=>gen_20_cmp_pBs_28, sum(20)=>
      gen_20_cmp_pBs_27, sum(19)=>gen_20_cmp_pBs_26, sum(18)=>
      gen_20_cmp_pBs_25, sum(17)=>gen_20_cmp_pBs_24, sum(16)=>
      gen_20_cmp_pBs_23, sum(15)=>outputs_20_15, sum(14)=>outputs_20_14, 
      sum(13)=>outputs_20_13, sum(12)=>outputs_20_12, sum(11)=>outputs_20_11, 
      sum(10)=>outputs_20_10, sum(9)=>outputs_20_9, sum(8)=>outputs_20_8, 
      sum(7)=>outputs_20_7, sum(6)=>outputs_20_6, sum(5)=>outputs_20_5, 
      sum(4)=>outputs_20_4, sum(3)=>outputs_20_3, sum(2)=>outputs_20_2, 
      sum(1)=>outputs_20_1, sum(0)=>outputs_20_0, carryOut=>DANGLING(24));
   gen_19_cmp_pRegCmp : Reg_33 port map ( D(32)=>gen_24_cmp_pInit_32, D(31)
      =>gen_24_cmp_pInit_32, D(30)=>gen_19_cmp_pBs_30, D(29)=>
      gen_19_cmp_pBs_29, D(28)=>gen_19_cmp_pBs_28, D(27)=>gen_19_cmp_pBs_27, 
      D(26)=>gen_19_cmp_pBs_26, D(25)=>gen_19_cmp_pBs_25, D(24)=>
      gen_19_cmp_pBs_24, D(23)=>gen_19_cmp_pBs_23, D(22)=>outputs_19_15, 
      D(21)=>outputs_19_14, D(20)=>outputs_19_13, D(19)=>outputs_19_12, 
      D(18)=>outputs_19_11, D(17)=>outputs_19_10, D(16)=>outputs_19_9, D(15)
      =>outputs_19_8, D(14)=>outputs_19_7, D(13)=>outputs_19_6, D(12)=>
      outputs_19_5, D(11)=>outputs_19_4, D(10)=>outputs_19_3, D(9)=>
      outputs_19_2, D(8)=>outputs_19_1, D(7)=>outputs_19_0, D(6)=>
      gen_19_cmp_pMux_8, D(5)=>gen_19_cmp_pMux_7, D(4)=>gen_19_cmp_pMux_6, 
      D(3)=>gen_19_cmp_pMux_5, D(2)=>gen_19_cmp_pMux_4, D(1)=>
      gen_19_cmp_pMux_3, D(0)=>nx10190, en=>nx11918, clk=>nx10122, rst=>rst, 
      Q(32)=>DANGLING(25), Q(31)=>DANGLING(26), Q(30)=>gen_19_cmp_pReg_30, 
      Q(29)=>gen_19_cmp_pReg_29, Q(28)=>gen_19_cmp_pReg_28, Q(27)=>
      gen_19_cmp_pReg_27, Q(26)=>gen_19_cmp_pReg_26, Q(25)=>
      gen_19_cmp_pReg_25, Q(24)=>gen_19_cmp_pReg_24, Q(23)=>
      gen_19_cmp_pReg_23, Q(22)=>gen_19_cmp_pReg_22, Q(21)=>
      gen_19_cmp_pReg_21, Q(20)=>gen_19_cmp_pReg_20, Q(19)=>
      gen_19_cmp_pReg_19, Q(18)=>gen_19_cmp_pReg_18, Q(17)=>
      gen_19_cmp_pReg_17, Q(16)=>gen_19_cmp_pReg_16, Q(15)=>
      gen_19_cmp_pReg_15, Q(14)=>gen_19_cmp_pReg_14, Q(13)=>
      gen_19_cmp_pReg_13, Q(12)=>gen_19_cmp_pReg_12, Q(11)=>
      gen_19_cmp_pReg_11, Q(10)=>gen_19_cmp_pReg_10, Q(9)=>gen_19_cmp_pReg_9, 
      Q(8)=>gen_19_cmp_pReg_8, Q(7)=>gen_19_cmp_pReg_7, Q(6)=>
      gen_19_cmp_pReg_6, Q(5)=>gen_19_cmp_pReg_5, Q(4)=>gen_19_cmp_pReg_4, 
      Q(3)=>gen_19_cmp_pReg_3, Q(2)=>gen_19_cmp_pReg_2, Q(1)=>
      gen_19_cmp_pReg_1, Q(0)=>gen_19_cmp_pReg_0);
   gen_19_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>gen_24_cmp_pInit_32, 
      a(31)=>gen_24_cmp_pInit_32, a(30)=>gen_19_cmp_pReg_30, a(29)=>
      gen_19_cmp_pReg_29, a(28)=>gen_19_cmp_pReg_28, a(27)=>
      gen_19_cmp_pReg_27, a(26)=>gen_19_cmp_pReg_26, a(25)=>
      gen_19_cmp_pReg_25, a(24)=>gen_19_cmp_pReg_24, a(23)=>
      gen_19_cmp_pReg_23, a(22)=>gen_19_cmp_pReg_22, a(21)=>
      gen_19_cmp_pReg_21, a(20)=>gen_19_cmp_pReg_20, a(19)=>
      gen_19_cmp_pReg_19, a(18)=>gen_19_cmp_pReg_18, a(17)=>
      gen_19_cmp_pReg_17, a(16)=>gen_19_cmp_pReg_16, a(15)=>
      gen_19_cmp_pReg_15, a(14)=>gen_19_cmp_pReg_14, a(13)=>
      gen_19_cmp_pReg_13, a(12)=>gen_19_cmp_pReg_12, a(11)=>
      gen_19_cmp_pReg_11, a(10)=>gen_19_cmp_pReg_10, a(9)=>gen_19_cmp_pReg_9, 
      a(8)=>gen_19_cmp_pReg_8, a(7)=>gen_19_cmp_pReg_7, a(6)=>
      gen_19_cmp_pReg_6, a(5)=>gen_19_cmp_pReg_5, a(4)=>gen_19_cmp_pReg_4, 
      a(3)=>gen_19_cmp_pReg_3, a(2)=>gen_19_cmp_pReg_2, a(1)=>
      gen_19_cmp_pReg_1, a(0)=>gen_19_cmp_pReg_0, b(32)=>gen_24_cmp_pInit_32, 
      b(31)=>gen_24_cmp_pInit_32, b(30)=>gen_24_cmp_pInit_32, b(29)=>
      gen_24_cmp_pInit_32, b(28)=>gen_24_cmp_pInit_32, b(27)=>
      gen_24_cmp_pInit_32, b(26)=>gen_24_cmp_pInit_32, b(25)=>
      gen_24_cmp_pInit_32, b(24)=>gen_24_cmp_pInit_32, b(23)=>
      gen_24_cmp_pInit_32, b(22)=>gen_24_cmp_pInit_32, b(21)=>
      gen_24_cmp_pInit_32, b(20)=>gen_24_cmp_pInit_32, b(19)=>
      gen_24_cmp_pInit_32, b(18)=>gen_24_cmp_pInit_32, b(17)=>
      gen_24_cmp_pInit_32, b(16)=>gen_24_cmp_pInit_32, b(15)=>
      gen_24_cmp_pInit_32, b(14)=>gen_24_cmp_pInit_32, b(13)=>
      gen_24_cmp_pInit_32, b(12)=>gen_24_cmp_pInit_32, b(11)=>
      gen_24_cmp_pInit_32, b(10)=>gen_24_cmp_pInit_32, b(9)=>
      gen_24_cmp_pInit_32, b(8)=>filter_19_7, b(7)=>filter_19_6, b(6)=>
      filter_19_5, b(5)=>filter_19_4, b(4)=>filter_19_3, b(3)=>filter_19_2, 
      b(2)=>filter_19_1, b(1)=>filter_19_0, b(0)=>gen_24_cmp_pInit_32, sel=>
      nx11898, f(32)=>DANGLING(27), f(31)=>DANGLING(28), f(30)=>
      gen_19_cmp_pMux_30, f(29)=>gen_19_cmp_pMux_29, f(28)=>
      gen_19_cmp_pMux_28, f(27)=>gen_19_cmp_pMux_27, f(26)=>
      gen_19_cmp_pMux_26, f(25)=>gen_19_cmp_pMux_25, f(24)=>
      gen_19_cmp_pMux_24, f(23)=>gen_19_cmp_pMux_23, f(22)=>
      gen_19_cmp_pMux_22, f(21)=>gen_19_cmp_pMux_21, f(20)=>
      gen_19_cmp_pMux_20, f(19)=>gen_19_cmp_pMux_19, f(18)=>
      gen_19_cmp_pMux_18, f(17)=>gen_19_cmp_pMux_17, f(16)=>
      gen_19_cmp_pMux_16, f(15)=>gen_19_cmp_pMux_15, f(14)=>
      gen_19_cmp_pMux_14, f(13)=>gen_19_cmp_pMux_13, f(12)=>
      gen_19_cmp_pMux_12, f(11)=>gen_19_cmp_pMux_11, f(10)=>
      gen_19_cmp_pMux_10, f(9)=>gen_19_cmp_pMux_9, f(8)=>gen_19_cmp_pMux_8, 
      f(7)=>gen_19_cmp_pMux_7, f(6)=>gen_19_cmp_pMux_6, f(5)=>
      gen_19_cmp_pMux_5, f(4)=>gen_19_cmp_pMux_4, f(3)=>gen_19_cmp_pMux_3, 
      f(2)=>gen_19_cmp_pMux_2, f(1)=>gen_19_cmp_pMux_1, f(0)=>
      gen_19_cmp_pMux_0);
   gen_19_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>
      gen_24_cmp_pInit_32, a(22)=>gen_24_cmp_pInit_32, a(21)=>
      gen_19_cmp_pMux_30, a(20)=>gen_19_cmp_pMux_29, a(19)=>
      gen_19_cmp_pMux_28, a(18)=>gen_19_cmp_pMux_27, a(17)=>
      gen_19_cmp_pMux_26, a(16)=>gen_19_cmp_pMux_25, a(15)=>
      gen_19_cmp_pMux_24, a(14)=>gen_19_cmp_pMux_23, a(13)=>
      gen_19_cmp_pMux_22, a(12)=>gen_19_cmp_pMux_21, a(11)=>
      gen_19_cmp_pMux_20, a(10)=>gen_19_cmp_pMux_19, a(9)=>
      gen_19_cmp_pMux_18, a(8)=>gen_19_cmp_pMux_17, a(7)=>gen_19_cmp_pMux_16, 
      a(6)=>gen_19_cmp_pMux_15, a(5)=>gen_19_cmp_pMux_14, a(4)=>
      gen_19_cmp_pMux_13, a(3)=>gen_19_cmp_pMux_12, a(2)=>gen_19_cmp_pMux_11, 
      a(1)=>gen_19_cmp_pMux_10, a(0)=>gen_19_cmp_pMux_9, b(23)=>nx10494, 
      b(22)=>nx10494, b(21)=>nx10492, b(20)=>nx10500, b(19)=>nx10498, b(18)
      =>nx10496, b(17)=>nx10494, b(16)=>nx10492, b(15)=>
      gen_19_cmp_BSCmp_op2_15, b(14)=>gen_19_cmp_BSCmp_op2_14, b(13)=>
      gen_19_cmp_BSCmp_op2_13, b(12)=>gen_19_cmp_BSCmp_op2_12, b(11)=>
      gen_19_cmp_BSCmp_op2_11, b(10)=>gen_19_cmp_BSCmp_op2_10, b(9)=>
      gen_19_cmp_BSCmp_op2_9, b(8)=>gen_19_cmp_BSCmp_op2_8, b(7)=>
      gen_19_cmp_BSCmp_op2_7, b(6)=>gen_19_cmp_BSCmp_op2_6, b(5)=>
      gen_19_cmp_BSCmp_op2_5, b(4)=>gen_19_cmp_BSCmp_op2_4, b(3)=>
      gen_19_cmp_BSCmp_op2_3, b(2)=>gen_19_cmp_BSCmp_op2_2, b(1)=>
      gen_19_cmp_BSCmp_op2_1, b(0)=>gen_19_cmp_BSCmp_op2_0, carryIn=>
      gen_19_cmp_BSCmp_carryIn, sum(23)=>gen_19_cmp_pBs_30, sum(22)=>
      gen_19_cmp_pBs_29, sum(21)=>gen_19_cmp_pBs_28, sum(20)=>
      gen_19_cmp_pBs_27, sum(19)=>gen_19_cmp_pBs_26, sum(18)=>
      gen_19_cmp_pBs_25, sum(17)=>gen_19_cmp_pBs_24, sum(16)=>
      gen_19_cmp_pBs_23, sum(15)=>outputs_19_15, sum(14)=>outputs_19_14, 
      sum(13)=>outputs_19_13, sum(12)=>outputs_19_12, sum(11)=>outputs_19_11, 
      sum(10)=>outputs_19_10, sum(9)=>outputs_19_9, sum(8)=>outputs_19_8, 
      sum(7)=>outputs_19_7, sum(6)=>outputs_19_6, sum(5)=>outputs_19_5, 
      sum(4)=>outputs_19_4, sum(3)=>outputs_19_3, sum(2)=>outputs_19_2, 
      sum(1)=>outputs_19_1, sum(0)=>outputs_19_0, carryOut=>DANGLING(29));
   gen_18_cmp_pRegCmp : Reg_33 port map ( D(32)=>gen_24_cmp_pInit_32, D(31)
      =>gen_24_cmp_pInit_32, D(30)=>gen_18_cmp_pBs_30, D(29)=>
      gen_18_cmp_pBs_29, D(28)=>gen_18_cmp_pBs_28, D(27)=>gen_18_cmp_pBs_27, 
      D(26)=>gen_18_cmp_pBs_26, D(25)=>gen_18_cmp_pBs_25, D(24)=>
      gen_18_cmp_pBs_24, D(23)=>gen_18_cmp_pBs_23, D(22)=>outputs_18_15, 
      D(21)=>outputs_18_14, D(20)=>outputs_18_13, D(19)=>outputs_18_12, 
      D(18)=>outputs_18_11, D(17)=>outputs_18_10, D(16)=>outputs_18_9, D(15)
      =>outputs_18_8, D(14)=>outputs_18_7, D(13)=>outputs_18_6, D(12)=>
      outputs_18_5, D(11)=>outputs_18_4, D(10)=>outputs_18_3, D(9)=>
      outputs_18_2, D(8)=>outputs_18_1, D(7)=>outputs_18_0, D(6)=>
      gen_18_cmp_pMux_8, D(5)=>gen_18_cmp_pMux_7, D(4)=>gen_18_cmp_pMux_6, 
      D(3)=>gen_18_cmp_pMux_5, D(2)=>gen_18_cmp_pMux_4, D(1)=>
      gen_18_cmp_pMux_3, D(0)=>nx10202, en=>nx10880, clk=>nx10122, rst=>rst, 
      Q(32)=>DANGLING(30), Q(31)=>DANGLING(31), Q(30)=>gen_18_cmp_pReg_30, 
      Q(29)=>gen_18_cmp_pReg_29, Q(28)=>gen_18_cmp_pReg_28, Q(27)=>
      gen_18_cmp_pReg_27, Q(26)=>gen_18_cmp_pReg_26, Q(25)=>
      gen_18_cmp_pReg_25, Q(24)=>gen_18_cmp_pReg_24, Q(23)=>
      gen_18_cmp_pReg_23, Q(22)=>gen_18_cmp_pReg_22, Q(21)=>
      gen_18_cmp_pReg_21, Q(20)=>gen_18_cmp_pReg_20, Q(19)=>
      gen_18_cmp_pReg_19, Q(18)=>gen_18_cmp_pReg_18, Q(17)=>
      gen_18_cmp_pReg_17, Q(16)=>gen_18_cmp_pReg_16, Q(15)=>
      gen_18_cmp_pReg_15, Q(14)=>gen_18_cmp_pReg_14, Q(13)=>
      gen_18_cmp_pReg_13, Q(12)=>gen_18_cmp_pReg_12, Q(11)=>
      gen_18_cmp_pReg_11, Q(10)=>gen_18_cmp_pReg_10, Q(9)=>gen_18_cmp_pReg_9, 
      Q(8)=>gen_18_cmp_pReg_8, Q(7)=>gen_18_cmp_pReg_7, Q(6)=>
      gen_18_cmp_pReg_6, Q(5)=>gen_18_cmp_pReg_5, Q(4)=>gen_18_cmp_pReg_4, 
      Q(3)=>gen_18_cmp_pReg_3, Q(2)=>gen_18_cmp_pReg_2, Q(1)=>
      gen_18_cmp_pReg_1, Q(0)=>gen_18_cmp_pReg_0);
   gen_18_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>gen_24_cmp_pInit_32, 
      a(31)=>gen_24_cmp_pInit_32, a(30)=>gen_18_cmp_pReg_30, a(29)=>
      gen_18_cmp_pReg_29, a(28)=>gen_18_cmp_pReg_28, a(27)=>
      gen_18_cmp_pReg_27, a(26)=>gen_18_cmp_pReg_26, a(25)=>
      gen_18_cmp_pReg_25, a(24)=>gen_18_cmp_pReg_24, a(23)=>
      gen_18_cmp_pReg_23, a(22)=>gen_18_cmp_pReg_22, a(21)=>
      gen_18_cmp_pReg_21, a(20)=>gen_18_cmp_pReg_20, a(19)=>
      gen_18_cmp_pReg_19, a(18)=>gen_18_cmp_pReg_18, a(17)=>
      gen_18_cmp_pReg_17, a(16)=>gen_18_cmp_pReg_16, a(15)=>
      gen_18_cmp_pReg_15, a(14)=>gen_18_cmp_pReg_14, a(13)=>
      gen_18_cmp_pReg_13, a(12)=>gen_18_cmp_pReg_12, a(11)=>
      gen_18_cmp_pReg_11, a(10)=>gen_18_cmp_pReg_10, a(9)=>gen_18_cmp_pReg_9, 
      a(8)=>gen_18_cmp_pReg_8, a(7)=>gen_18_cmp_pReg_7, a(6)=>
      gen_18_cmp_pReg_6, a(5)=>gen_18_cmp_pReg_5, a(4)=>gen_18_cmp_pReg_4, 
      a(3)=>gen_18_cmp_pReg_3, a(2)=>gen_18_cmp_pReg_2, a(1)=>
      gen_18_cmp_pReg_1, a(0)=>gen_18_cmp_pReg_0, b(32)=>gen_24_cmp_pInit_32, 
      b(31)=>gen_24_cmp_pInit_32, b(30)=>gen_24_cmp_pInit_32, b(29)=>
      gen_24_cmp_pInit_32, b(28)=>gen_24_cmp_pInit_32, b(27)=>
      gen_24_cmp_pInit_32, b(26)=>gen_24_cmp_pInit_32, b(25)=>
      gen_24_cmp_pInit_32, b(24)=>gen_24_cmp_pInit_32, b(23)=>
      gen_24_cmp_pInit_32, b(22)=>gen_24_cmp_pInit_32, b(21)=>
      gen_24_cmp_pInit_32, b(20)=>gen_24_cmp_pInit_32, b(19)=>
      gen_24_cmp_pInit_32, b(18)=>gen_24_cmp_pInit_32, b(17)=>
      gen_24_cmp_pInit_32, b(16)=>gen_24_cmp_pInit_32, b(15)=>
      gen_24_cmp_pInit_32, b(14)=>gen_24_cmp_pInit_32, b(13)=>
      gen_24_cmp_pInit_32, b(12)=>gen_24_cmp_pInit_32, b(11)=>
      gen_24_cmp_pInit_32, b(10)=>gen_24_cmp_pInit_32, b(9)=>
      gen_24_cmp_pInit_32, b(8)=>filter_18_7, b(7)=>filter_18_6, b(6)=>
      filter_18_5, b(5)=>filter_18_4, b(4)=>filter_18_3, b(3)=>filter_18_2, 
      b(2)=>filter_18_1, b(1)=>filter_18_0, b(0)=>gen_24_cmp_pInit_32, sel=>
      nx11900, f(32)=>DANGLING(32), f(31)=>DANGLING(33), f(30)=>
      gen_18_cmp_pMux_30, f(29)=>gen_18_cmp_pMux_29, f(28)=>
      gen_18_cmp_pMux_28, f(27)=>gen_18_cmp_pMux_27, f(26)=>
      gen_18_cmp_pMux_26, f(25)=>gen_18_cmp_pMux_25, f(24)=>
      gen_18_cmp_pMux_24, f(23)=>gen_18_cmp_pMux_23, f(22)=>
      gen_18_cmp_pMux_22, f(21)=>gen_18_cmp_pMux_21, f(20)=>
      gen_18_cmp_pMux_20, f(19)=>gen_18_cmp_pMux_19, f(18)=>
      gen_18_cmp_pMux_18, f(17)=>gen_18_cmp_pMux_17, f(16)=>
      gen_18_cmp_pMux_16, f(15)=>gen_18_cmp_pMux_15, f(14)=>
      gen_18_cmp_pMux_14, f(13)=>gen_18_cmp_pMux_13, f(12)=>
      gen_18_cmp_pMux_12, f(11)=>gen_18_cmp_pMux_11, f(10)=>
      gen_18_cmp_pMux_10, f(9)=>gen_18_cmp_pMux_9, f(8)=>gen_18_cmp_pMux_8, 
      f(7)=>gen_18_cmp_pMux_7, f(6)=>gen_18_cmp_pMux_6, f(5)=>
      gen_18_cmp_pMux_5, f(4)=>gen_18_cmp_pMux_4, f(3)=>gen_18_cmp_pMux_3, 
      f(2)=>gen_18_cmp_pMux_2, f(1)=>gen_18_cmp_pMux_1, f(0)=>
      gen_18_cmp_pMux_0);
   gen_18_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>
      gen_24_cmp_pInit_32, a(22)=>gen_24_cmp_pInit_32, a(21)=>
      gen_18_cmp_pMux_30, a(20)=>gen_18_cmp_pMux_29, a(19)=>
      gen_18_cmp_pMux_28, a(18)=>gen_18_cmp_pMux_27, a(17)=>
      gen_18_cmp_pMux_26, a(16)=>gen_18_cmp_pMux_25, a(15)=>
      gen_18_cmp_pMux_24, a(14)=>gen_18_cmp_pMux_23, a(13)=>
      gen_18_cmp_pMux_22, a(12)=>gen_18_cmp_pMux_21, a(11)=>
      gen_18_cmp_pMux_20, a(10)=>gen_18_cmp_pMux_19, a(9)=>
      gen_18_cmp_pMux_18, a(8)=>gen_18_cmp_pMux_17, a(7)=>gen_18_cmp_pMux_16, 
      a(6)=>gen_18_cmp_pMux_15, a(5)=>gen_18_cmp_pMux_14, a(4)=>
      gen_18_cmp_pMux_13, a(3)=>gen_18_cmp_pMux_12, a(2)=>gen_18_cmp_pMux_11, 
      a(1)=>gen_18_cmp_pMux_10, a(0)=>gen_18_cmp_pMux_9, b(23)=>nx10506, 
      b(22)=>nx10506, b(21)=>nx10504, b(20)=>nx10512, b(19)=>nx10510, b(18)
      =>nx10508, b(17)=>nx10506, b(16)=>nx10504, b(15)=>
      gen_18_cmp_BSCmp_op2_15, b(14)=>gen_18_cmp_BSCmp_op2_14, b(13)=>
      gen_18_cmp_BSCmp_op2_13, b(12)=>gen_18_cmp_BSCmp_op2_12, b(11)=>
      gen_18_cmp_BSCmp_op2_11, b(10)=>gen_18_cmp_BSCmp_op2_10, b(9)=>
      gen_18_cmp_BSCmp_op2_9, b(8)=>gen_18_cmp_BSCmp_op2_8, b(7)=>
      gen_18_cmp_BSCmp_op2_7, b(6)=>gen_18_cmp_BSCmp_op2_6, b(5)=>
      gen_18_cmp_BSCmp_op2_5, b(4)=>gen_18_cmp_BSCmp_op2_4, b(3)=>
      gen_18_cmp_BSCmp_op2_3, b(2)=>gen_18_cmp_BSCmp_op2_2, b(1)=>
      gen_18_cmp_BSCmp_op2_1, b(0)=>gen_18_cmp_BSCmp_op2_0, carryIn=>
      gen_18_cmp_BSCmp_carryIn, sum(23)=>gen_18_cmp_pBs_30, sum(22)=>
      gen_18_cmp_pBs_29, sum(21)=>gen_18_cmp_pBs_28, sum(20)=>
      gen_18_cmp_pBs_27, sum(19)=>gen_18_cmp_pBs_26, sum(18)=>
      gen_18_cmp_pBs_25, sum(17)=>gen_18_cmp_pBs_24, sum(16)=>
      gen_18_cmp_pBs_23, sum(15)=>outputs_18_15, sum(14)=>outputs_18_14, 
      sum(13)=>outputs_18_13, sum(12)=>outputs_18_12, sum(11)=>outputs_18_11, 
      sum(10)=>outputs_18_10, sum(9)=>outputs_18_9, sum(8)=>outputs_18_8, 
      sum(7)=>outputs_18_7, sum(6)=>outputs_18_6, sum(5)=>outputs_18_5, 
      sum(4)=>outputs_18_4, sum(3)=>outputs_18_3, sum(2)=>outputs_18_2, 
      sum(1)=>outputs_18_1, sum(0)=>outputs_18_0, carryOut=>DANGLING(34));
   gen_17_cmp_pRegCmp : Reg_33 port map ( D(32)=>gen_24_cmp_pInit_32, D(31)
      =>gen_24_cmp_pInit_32, D(30)=>gen_17_cmp_pBs_30, D(29)=>
      gen_17_cmp_pBs_29, D(28)=>gen_17_cmp_pBs_28, D(27)=>gen_17_cmp_pBs_27, 
      D(26)=>gen_17_cmp_pBs_26, D(25)=>gen_17_cmp_pBs_25, D(24)=>
      gen_17_cmp_pBs_24, D(23)=>gen_17_cmp_pBs_23, D(22)=>outputs_17_15, 
      D(21)=>outputs_17_14, D(20)=>outputs_17_13, D(19)=>outputs_17_12, 
      D(18)=>outputs_17_11, D(17)=>outputs_17_10, D(16)=>outputs_17_9, D(15)
      =>outputs_17_8, D(14)=>outputs_17_7, D(13)=>outputs_17_6, D(12)=>
      outputs_17_5, D(11)=>outputs_17_4, D(10)=>outputs_17_3, D(9)=>
      outputs_17_2, D(8)=>outputs_17_1, D(7)=>outputs_17_0, D(6)=>
      gen_17_cmp_pMux_8, D(5)=>gen_17_cmp_pMux_7, D(4)=>gen_17_cmp_pMux_6, 
      D(3)=>gen_17_cmp_pMux_5, D(2)=>gen_17_cmp_pMux_4, D(1)=>
      gen_17_cmp_pMux_3, D(0)=>nx10214, en=>nx11920, clk=>nx10124, rst=>rst, 
      Q(32)=>DANGLING(35), Q(31)=>DANGLING(36), Q(30)=>gen_17_cmp_pReg_30, 
      Q(29)=>gen_17_cmp_pReg_29, Q(28)=>gen_17_cmp_pReg_28, Q(27)=>
      gen_17_cmp_pReg_27, Q(26)=>gen_17_cmp_pReg_26, Q(25)=>
      gen_17_cmp_pReg_25, Q(24)=>gen_17_cmp_pReg_24, Q(23)=>
      gen_17_cmp_pReg_23, Q(22)=>gen_17_cmp_pReg_22, Q(21)=>
      gen_17_cmp_pReg_21, Q(20)=>gen_17_cmp_pReg_20, Q(19)=>
      gen_17_cmp_pReg_19, Q(18)=>gen_17_cmp_pReg_18, Q(17)=>
      gen_17_cmp_pReg_17, Q(16)=>gen_17_cmp_pReg_16, Q(15)=>
      gen_17_cmp_pReg_15, Q(14)=>gen_17_cmp_pReg_14, Q(13)=>
      gen_17_cmp_pReg_13, Q(12)=>gen_17_cmp_pReg_12, Q(11)=>
      gen_17_cmp_pReg_11, Q(10)=>gen_17_cmp_pReg_10, Q(9)=>gen_17_cmp_pReg_9, 
      Q(8)=>gen_17_cmp_pReg_8, Q(7)=>gen_17_cmp_pReg_7, Q(6)=>
      gen_17_cmp_pReg_6, Q(5)=>gen_17_cmp_pReg_5, Q(4)=>gen_17_cmp_pReg_4, 
      Q(3)=>gen_17_cmp_pReg_3, Q(2)=>gen_17_cmp_pReg_2, Q(1)=>
      gen_17_cmp_pReg_1, Q(0)=>gen_17_cmp_pReg_0);
   gen_17_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>gen_24_cmp_pInit_32, 
      a(31)=>gen_24_cmp_pInit_32, a(30)=>gen_17_cmp_pReg_30, a(29)=>
      gen_17_cmp_pReg_29, a(28)=>gen_17_cmp_pReg_28, a(27)=>
      gen_17_cmp_pReg_27, a(26)=>gen_17_cmp_pReg_26, a(25)=>
      gen_17_cmp_pReg_25, a(24)=>gen_17_cmp_pReg_24, a(23)=>
      gen_17_cmp_pReg_23, a(22)=>gen_17_cmp_pReg_22, a(21)=>
      gen_17_cmp_pReg_21, a(20)=>gen_17_cmp_pReg_20, a(19)=>
      gen_17_cmp_pReg_19, a(18)=>gen_17_cmp_pReg_18, a(17)=>
      gen_17_cmp_pReg_17, a(16)=>gen_17_cmp_pReg_16, a(15)=>
      gen_17_cmp_pReg_15, a(14)=>gen_17_cmp_pReg_14, a(13)=>
      gen_17_cmp_pReg_13, a(12)=>gen_17_cmp_pReg_12, a(11)=>
      gen_17_cmp_pReg_11, a(10)=>gen_17_cmp_pReg_10, a(9)=>gen_17_cmp_pReg_9, 
      a(8)=>gen_17_cmp_pReg_8, a(7)=>gen_17_cmp_pReg_7, a(6)=>
      gen_17_cmp_pReg_6, a(5)=>gen_17_cmp_pReg_5, a(4)=>gen_17_cmp_pReg_4, 
      a(3)=>gen_17_cmp_pReg_3, a(2)=>gen_17_cmp_pReg_2, a(1)=>
      gen_17_cmp_pReg_1, a(0)=>gen_17_cmp_pReg_0, b(32)=>gen_24_cmp_pInit_32, 
      b(31)=>gen_24_cmp_pInit_32, b(30)=>gen_24_cmp_pInit_32, b(29)=>
      gen_24_cmp_pInit_32, b(28)=>gen_24_cmp_pInit_32, b(27)=>
      gen_24_cmp_pInit_32, b(26)=>gen_24_cmp_pInit_32, b(25)=>
      gen_24_cmp_pInit_32, b(24)=>gen_24_cmp_pInit_32, b(23)=>
      gen_24_cmp_pInit_32, b(22)=>gen_24_cmp_pInit_32, b(21)=>
      gen_24_cmp_pInit_32, b(20)=>gen_24_cmp_pInit_32, b(19)=>
      gen_24_cmp_pInit_32, b(18)=>gen_24_cmp_pInit_32, b(17)=>
      gen_24_cmp_pInit_32, b(16)=>gen_24_cmp_pInit_32, b(15)=>
      gen_24_cmp_pInit_32, b(14)=>gen_24_cmp_pInit_32, b(13)=>
      gen_24_cmp_pInit_32, b(12)=>gen_24_cmp_pInit_32, b(11)=>
      gen_24_cmp_pInit_32, b(10)=>gen_24_cmp_pInit_32, b(9)=>
      gen_24_cmp_pInit_32, b(8)=>filter_17_7, b(7)=>filter_17_6, b(6)=>
      filter_17_5, b(5)=>filter_17_4, b(4)=>filter_17_3, b(3)=>filter_17_2, 
      b(2)=>filter_17_1, b(1)=>filter_17_0, b(0)=>gen_24_cmp_pInit_32, sel=>
      nx11902, f(32)=>DANGLING(37), f(31)=>DANGLING(38), f(30)=>
      gen_17_cmp_pMux_30, f(29)=>gen_17_cmp_pMux_29, f(28)=>
      gen_17_cmp_pMux_28, f(27)=>gen_17_cmp_pMux_27, f(26)=>
      gen_17_cmp_pMux_26, f(25)=>gen_17_cmp_pMux_25, f(24)=>
      gen_17_cmp_pMux_24, f(23)=>gen_17_cmp_pMux_23, f(22)=>
      gen_17_cmp_pMux_22, f(21)=>gen_17_cmp_pMux_21, f(20)=>
      gen_17_cmp_pMux_20, f(19)=>gen_17_cmp_pMux_19, f(18)=>
      gen_17_cmp_pMux_18, f(17)=>gen_17_cmp_pMux_17, f(16)=>
      gen_17_cmp_pMux_16, f(15)=>gen_17_cmp_pMux_15, f(14)=>
      gen_17_cmp_pMux_14, f(13)=>gen_17_cmp_pMux_13, f(12)=>
      gen_17_cmp_pMux_12, f(11)=>gen_17_cmp_pMux_11, f(10)=>
      gen_17_cmp_pMux_10, f(9)=>gen_17_cmp_pMux_9, f(8)=>gen_17_cmp_pMux_8, 
      f(7)=>gen_17_cmp_pMux_7, f(6)=>gen_17_cmp_pMux_6, f(5)=>
      gen_17_cmp_pMux_5, f(4)=>gen_17_cmp_pMux_4, f(3)=>gen_17_cmp_pMux_3, 
      f(2)=>gen_17_cmp_pMux_2, f(1)=>gen_17_cmp_pMux_1, f(0)=>
      gen_17_cmp_pMux_0);
   gen_17_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>
      gen_24_cmp_pInit_32, a(22)=>gen_24_cmp_pInit_32, a(21)=>
      gen_17_cmp_pMux_30, a(20)=>gen_17_cmp_pMux_29, a(19)=>
      gen_17_cmp_pMux_28, a(18)=>gen_17_cmp_pMux_27, a(17)=>
      gen_17_cmp_pMux_26, a(16)=>gen_17_cmp_pMux_25, a(15)=>
      gen_17_cmp_pMux_24, a(14)=>gen_17_cmp_pMux_23, a(13)=>
      gen_17_cmp_pMux_22, a(12)=>gen_17_cmp_pMux_21, a(11)=>
      gen_17_cmp_pMux_20, a(10)=>gen_17_cmp_pMux_19, a(9)=>
      gen_17_cmp_pMux_18, a(8)=>gen_17_cmp_pMux_17, a(7)=>gen_17_cmp_pMux_16, 
      a(6)=>gen_17_cmp_pMux_15, a(5)=>gen_17_cmp_pMux_14, a(4)=>
      gen_17_cmp_pMux_13, a(3)=>gen_17_cmp_pMux_12, a(2)=>gen_17_cmp_pMux_11, 
      a(1)=>gen_17_cmp_pMux_10, a(0)=>gen_17_cmp_pMux_9, b(23)=>nx10518, 
      b(22)=>nx10518, b(21)=>nx10516, b(20)=>nx10524, b(19)=>nx10522, b(18)
      =>nx10520, b(17)=>nx10518, b(16)=>nx10516, b(15)=>
      gen_17_cmp_BSCmp_op2_15, b(14)=>gen_17_cmp_BSCmp_op2_14, b(13)=>
      gen_17_cmp_BSCmp_op2_13, b(12)=>gen_17_cmp_BSCmp_op2_12, b(11)=>
      gen_17_cmp_BSCmp_op2_11, b(10)=>gen_17_cmp_BSCmp_op2_10, b(9)=>
      gen_17_cmp_BSCmp_op2_9, b(8)=>gen_17_cmp_BSCmp_op2_8, b(7)=>
      gen_17_cmp_BSCmp_op2_7, b(6)=>gen_17_cmp_BSCmp_op2_6, b(5)=>
      gen_17_cmp_BSCmp_op2_5, b(4)=>gen_17_cmp_BSCmp_op2_4, b(3)=>
      gen_17_cmp_BSCmp_op2_3, b(2)=>gen_17_cmp_BSCmp_op2_2, b(1)=>
      gen_17_cmp_BSCmp_op2_1, b(0)=>gen_17_cmp_BSCmp_op2_0, carryIn=>
      gen_17_cmp_BSCmp_carryIn, sum(23)=>gen_17_cmp_pBs_30, sum(22)=>
      gen_17_cmp_pBs_29, sum(21)=>gen_17_cmp_pBs_28, sum(20)=>
      gen_17_cmp_pBs_27, sum(19)=>gen_17_cmp_pBs_26, sum(18)=>
      gen_17_cmp_pBs_25, sum(17)=>gen_17_cmp_pBs_24, sum(16)=>
      gen_17_cmp_pBs_23, sum(15)=>outputs_17_15, sum(14)=>outputs_17_14, 
      sum(13)=>outputs_17_13, sum(12)=>outputs_17_12, sum(11)=>outputs_17_11, 
      sum(10)=>outputs_17_10, sum(9)=>outputs_17_9, sum(8)=>outputs_17_8, 
      sum(7)=>outputs_17_7, sum(6)=>outputs_17_6, sum(5)=>outputs_17_5, 
      sum(4)=>outputs_17_4, sum(3)=>outputs_17_3, sum(2)=>outputs_17_2, 
      sum(1)=>outputs_17_1, sum(0)=>outputs_17_0, carryOut=>DANGLING(39));
   gen_16_cmp_pRegCmp : Reg_33 port map ( D(32)=>gen_24_cmp_pInit_32, D(31)
      =>gen_24_cmp_pInit_32, D(30)=>gen_16_cmp_pBs_30, D(29)=>
      gen_16_cmp_pBs_29, D(28)=>gen_16_cmp_pBs_28, D(27)=>gen_16_cmp_pBs_27, 
      D(26)=>gen_16_cmp_pBs_26, D(25)=>gen_16_cmp_pBs_25, D(24)=>
      gen_16_cmp_pBs_24, D(23)=>gen_16_cmp_pBs_23, D(22)=>outputs_16_15, 
      D(21)=>outputs_16_14, D(20)=>outputs_16_13, D(19)=>outputs_16_12, 
      D(18)=>outputs_16_11, D(17)=>outputs_16_10, D(16)=>outputs_16_9, D(15)
      =>outputs_16_8, D(14)=>outputs_16_7, D(13)=>outputs_16_6, D(12)=>
      outputs_16_5, D(11)=>outputs_16_4, D(10)=>outputs_16_3, D(9)=>
      outputs_16_2, D(8)=>outputs_16_1, D(7)=>outputs_16_0, D(6)=>
      gen_16_cmp_pMux_8, D(5)=>gen_16_cmp_pMux_7, D(4)=>gen_16_cmp_pMux_6, 
      D(3)=>gen_16_cmp_pMux_5, D(2)=>gen_16_cmp_pMux_4, D(1)=>
      gen_16_cmp_pMux_3, D(0)=>nx10226, en=>nx11920, clk=>nx10124, rst=>rst, 
      Q(32)=>DANGLING(40), Q(31)=>DANGLING(41), Q(30)=>gen_16_cmp_pReg_30, 
      Q(29)=>gen_16_cmp_pReg_29, Q(28)=>gen_16_cmp_pReg_28, Q(27)=>
      gen_16_cmp_pReg_27, Q(26)=>gen_16_cmp_pReg_26, Q(25)=>
      gen_16_cmp_pReg_25, Q(24)=>gen_16_cmp_pReg_24, Q(23)=>
      gen_16_cmp_pReg_23, Q(22)=>gen_16_cmp_pReg_22, Q(21)=>
      gen_16_cmp_pReg_21, Q(20)=>gen_16_cmp_pReg_20, Q(19)=>
      gen_16_cmp_pReg_19, Q(18)=>gen_16_cmp_pReg_18, Q(17)=>
      gen_16_cmp_pReg_17, Q(16)=>gen_16_cmp_pReg_16, Q(15)=>
      gen_16_cmp_pReg_15, Q(14)=>gen_16_cmp_pReg_14, Q(13)=>
      gen_16_cmp_pReg_13, Q(12)=>gen_16_cmp_pReg_12, Q(11)=>
      gen_16_cmp_pReg_11, Q(10)=>gen_16_cmp_pReg_10, Q(9)=>gen_16_cmp_pReg_9, 
      Q(8)=>gen_16_cmp_pReg_8, Q(7)=>gen_16_cmp_pReg_7, Q(6)=>
      gen_16_cmp_pReg_6, Q(5)=>gen_16_cmp_pReg_5, Q(4)=>gen_16_cmp_pReg_4, 
      Q(3)=>gen_16_cmp_pReg_3, Q(2)=>gen_16_cmp_pReg_2, Q(1)=>
      gen_16_cmp_pReg_1, Q(0)=>gen_16_cmp_pReg_0);
   gen_16_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>gen_24_cmp_pInit_32, 
      a(31)=>gen_24_cmp_pInit_32, a(30)=>gen_16_cmp_pReg_30, a(29)=>
      gen_16_cmp_pReg_29, a(28)=>gen_16_cmp_pReg_28, a(27)=>
      gen_16_cmp_pReg_27, a(26)=>gen_16_cmp_pReg_26, a(25)=>
      gen_16_cmp_pReg_25, a(24)=>gen_16_cmp_pReg_24, a(23)=>
      gen_16_cmp_pReg_23, a(22)=>gen_16_cmp_pReg_22, a(21)=>
      gen_16_cmp_pReg_21, a(20)=>gen_16_cmp_pReg_20, a(19)=>
      gen_16_cmp_pReg_19, a(18)=>gen_16_cmp_pReg_18, a(17)=>
      gen_16_cmp_pReg_17, a(16)=>gen_16_cmp_pReg_16, a(15)=>
      gen_16_cmp_pReg_15, a(14)=>gen_16_cmp_pReg_14, a(13)=>
      gen_16_cmp_pReg_13, a(12)=>gen_16_cmp_pReg_12, a(11)=>
      gen_16_cmp_pReg_11, a(10)=>gen_16_cmp_pReg_10, a(9)=>gen_16_cmp_pReg_9, 
      a(8)=>gen_16_cmp_pReg_8, a(7)=>gen_16_cmp_pReg_7, a(6)=>
      gen_16_cmp_pReg_6, a(5)=>gen_16_cmp_pReg_5, a(4)=>gen_16_cmp_pReg_4, 
      a(3)=>gen_16_cmp_pReg_3, a(2)=>gen_16_cmp_pReg_2, a(1)=>
      gen_16_cmp_pReg_1, a(0)=>gen_16_cmp_pReg_0, b(32)=>gen_24_cmp_pInit_32, 
      b(31)=>gen_24_cmp_pInit_32, b(30)=>gen_24_cmp_pInit_32, b(29)=>
      gen_24_cmp_pInit_32, b(28)=>gen_24_cmp_pInit_32, b(27)=>
      gen_24_cmp_pInit_32, b(26)=>gen_24_cmp_pInit_32, b(25)=>
      gen_24_cmp_pInit_32, b(24)=>gen_24_cmp_pInit_32, b(23)=>
      gen_24_cmp_pInit_32, b(22)=>gen_24_cmp_pInit_32, b(21)=>
      gen_24_cmp_pInit_32, b(20)=>gen_24_cmp_pInit_32, b(19)=>
      gen_24_cmp_pInit_32, b(18)=>gen_24_cmp_pInit_32, b(17)=>
      gen_24_cmp_pInit_32, b(16)=>gen_24_cmp_pInit_32, b(15)=>
      gen_24_cmp_pInit_32, b(14)=>gen_24_cmp_pInit_32, b(13)=>
      gen_24_cmp_pInit_32, b(12)=>gen_24_cmp_pInit_32, b(11)=>
      gen_24_cmp_pInit_32, b(10)=>gen_24_cmp_pInit_32, b(9)=>
      gen_24_cmp_pInit_32, b(8)=>filter_16_7, b(7)=>filter_16_6, b(6)=>
      filter_16_5, b(5)=>filter_16_4, b(4)=>filter_16_3, b(3)=>filter_16_2, 
      b(2)=>filter_16_1, b(1)=>filter_16_0, b(0)=>gen_24_cmp_pInit_32, sel=>
      nx11902, f(32)=>DANGLING(42), f(31)=>DANGLING(43), f(30)=>
      gen_16_cmp_pMux_30, f(29)=>gen_16_cmp_pMux_29, f(28)=>
      gen_16_cmp_pMux_28, f(27)=>gen_16_cmp_pMux_27, f(26)=>
      gen_16_cmp_pMux_26, f(25)=>gen_16_cmp_pMux_25, f(24)=>
      gen_16_cmp_pMux_24, f(23)=>gen_16_cmp_pMux_23, f(22)=>
      gen_16_cmp_pMux_22, f(21)=>gen_16_cmp_pMux_21, f(20)=>
      gen_16_cmp_pMux_20, f(19)=>gen_16_cmp_pMux_19, f(18)=>
      gen_16_cmp_pMux_18, f(17)=>gen_16_cmp_pMux_17, f(16)=>
      gen_16_cmp_pMux_16, f(15)=>gen_16_cmp_pMux_15, f(14)=>
      gen_16_cmp_pMux_14, f(13)=>gen_16_cmp_pMux_13, f(12)=>
      gen_16_cmp_pMux_12, f(11)=>gen_16_cmp_pMux_11, f(10)=>
      gen_16_cmp_pMux_10, f(9)=>gen_16_cmp_pMux_9, f(8)=>gen_16_cmp_pMux_8, 
      f(7)=>gen_16_cmp_pMux_7, f(6)=>gen_16_cmp_pMux_6, f(5)=>
      gen_16_cmp_pMux_5, f(4)=>gen_16_cmp_pMux_4, f(3)=>gen_16_cmp_pMux_3, 
      f(2)=>gen_16_cmp_pMux_2, f(1)=>gen_16_cmp_pMux_1, f(0)=>
      gen_16_cmp_pMux_0);
   gen_16_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>
      gen_24_cmp_pInit_32, a(22)=>gen_24_cmp_pInit_32, a(21)=>
      gen_16_cmp_pMux_30, a(20)=>gen_16_cmp_pMux_29, a(19)=>
      gen_16_cmp_pMux_28, a(18)=>gen_16_cmp_pMux_27, a(17)=>
      gen_16_cmp_pMux_26, a(16)=>gen_16_cmp_pMux_25, a(15)=>
      gen_16_cmp_pMux_24, a(14)=>gen_16_cmp_pMux_23, a(13)=>
      gen_16_cmp_pMux_22, a(12)=>gen_16_cmp_pMux_21, a(11)=>
      gen_16_cmp_pMux_20, a(10)=>gen_16_cmp_pMux_19, a(9)=>
      gen_16_cmp_pMux_18, a(8)=>gen_16_cmp_pMux_17, a(7)=>gen_16_cmp_pMux_16, 
      a(6)=>gen_16_cmp_pMux_15, a(5)=>gen_16_cmp_pMux_14, a(4)=>
      gen_16_cmp_pMux_13, a(3)=>gen_16_cmp_pMux_12, a(2)=>gen_16_cmp_pMux_11, 
      a(1)=>gen_16_cmp_pMux_10, a(0)=>gen_16_cmp_pMux_9, b(23)=>nx10530, 
      b(22)=>nx10530, b(21)=>nx10528, b(20)=>nx10536, b(19)=>nx10534, b(18)
      =>nx10532, b(17)=>nx10530, b(16)=>nx10528, b(15)=>
      gen_16_cmp_BSCmp_op2_15, b(14)=>gen_16_cmp_BSCmp_op2_14, b(13)=>
      gen_16_cmp_BSCmp_op2_13, b(12)=>gen_16_cmp_BSCmp_op2_12, b(11)=>
      gen_16_cmp_BSCmp_op2_11, b(10)=>gen_16_cmp_BSCmp_op2_10, b(9)=>
      gen_16_cmp_BSCmp_op2_9, b(8)=>gen_16_cmp_BSCmp_op2_8, b(7)=>
      gen_16_cmp_BSCmp_op2_7, b(6)=>gen_16_cmp_BSCmp_op2_6, b(5)=>
      gen_16_cmp_BSCmp_op2_5, b(4)=>gen_16_cmp_BSCmp_op2_4, b(3)=>
      gen_16_cmp_BSCmp_op2_3, b(2)=>gen_16_cmp_BSCmp_op2_2, b(1)=>
      gen_16_cmp_BSCmp_op2_1, b(0)=>gen_16_cmp_BSCmp_op2_0, carryIn=>
      gen_16_cmp_BSCmp_carryIn, sum(23)=>gen_16_cmp_pBs_30, sum(22)=>
      gen_16_cmp_pBs_29, sum(21)=>gen_16_cmp_pBs_28, sum(20)=>
      gen_16_cmp_pBs_27, sum(19)=>gen_16_cmp_pBs_26, sum(18)=>
      gen_16_cmp_pBs_25, sum(17)=>gen_16_cmp_pBs_24, sum(16)=>
      gen_16_cmp_pBs_23, sum(15)=>outputs_16_15, sum(14)=>outputs_16_14, 
      sum(13)=>outputs_16_13, sum(12)=>outputs_16_12, sum(11)=>outputs_16_11, 
      sum(10)=>outputs_16_10, sum(9)=>outputs_16_9, sum(8)=>outputs_16_8, 
      sum(7)=>outputs_16_7, sum(6)=>outputs_16_6, sum(5)=>outputs_16_5, 
      sum(4)=>outputs_16_4, sum(3)=>outputs_16_3, sum(2)=>outputs_16_2, 
      sum(1)=>outputs_16_1, sum(0)=>outputs_16_0, carryOut=>DANGLING(44));
   gen_15_cmp_pRegCmp : Reg_33 port map ( D(32)=>gen_24_cmp_pInit_32, D(31)
      =>gen_24_cmp_pInit_32, D(30)=>gen_15_cmp_pBs_30, D(29)=>
      gen_15_cmp_pBs_29, D(28)=>gen_15_cmp_pBs_28, D(27)=>gen_15_cmp_pBs_27, 
      D(26)=>gen_15_cmp_pBs_26, D(25)=>gen_15_cmp_pBs_25, D(24)=>
      gen_15_cmp_pBs_24, D(23)=>gen_15_cmp_pBs_23, D(22)=>outputs_15_15, 
      D(21)=>outputs_15_14, D(20)=>outputs_15_13, D(19)=>outputs_15_12, 
      D(18)=>outputs_15_11, D(17)=>outputs_15_10, D(16)=>outputs_15_9, D(15)
      =>outputs_15_8, D(14)=>outputs_15_7, D(13)=>outputs_15_6, D(12)=>
      outputs_15_5, D(11)=>outputs_15_4, D(10)=>outputs_15_3, D(9)=>
      outputs_15_2, D(8)=>outputs_15_1, D(7)=>outputs_15_0, D(6)=>
      gen_15_cmp_pMux_8, D(5)=>gen_15_cmp_pMux_7, D(4)=>gen_15_cmp_pMux_6, 
      D(3)=>gen_15_cmp_pMux_5, D(2)=>gen_15_cmp_pMux_4, D(1)=>
      gen_15_cmp_pMux_3, D(0)=>nx10238, en=>nx11920, clk=>nx10124, rst=>rst, 
      Q(32)=>DANGLING(45), Q(31)=>DANGLING(46), Q(30)=>gen_15_cmp_pReg_30, 
      Q(29)=>gen_15_cmp_pReg_29, Q(28)=>gen_15_cmp_pReg_28, Q(27)=>
      gen_15_cmp_pReg_27, Q(26)=>gen_15_cmp_pReg_26, Q(25)=>
      gen_15_cmp_pReg_25, Q(24)=>gen_15_cmp_pReg_24, Q(23)=>
      gen_15_cmp_pReg_23, Q(22)=>gen_15_cmp_pReg_22, Q(21)=>
      gen_15_cmp_pReg_21, Q(20)=>gen_15_cmp_pReg_20, Q(19)=>
      gen_15_cmp_pReg_19, Q(18)=>gen_15_cmp_pReg_18, Q(17)=>
      gen_15_cmp_pReg_17, Q(16)=>gen_15_cmp_pReg_16, Q(15)=>
      gen_15_cmp_pReg_15, Q(14)=>gen_15_cmp_pReg_14, Q(13)=>
      gen_15_cmp_pReg_13, Q(12)=>gen_15_cmp_pReg_12, Q(11)=>
      gen_15_cmp_pReg_11, Q(10)=>gen_15_cmp_pReg_10, Q(9)=>gen_15_cmp_pReg_9, 
      Q(8)=>gen_15_cmp_pReg_8, Q(7)=>gen_15_cmp_pReg_7, Q(6)=>
      gen_15_cmp_pReg_6, Q(5)=>gen_15_cmp_pReg_5, Q(4)=>gen_15_cmp_pReg_4, 
      Q(3)=>gen_15_cmp_pReg_3, Q(2)=>gen_15_cmp_pReg_2, Q(1)=>
      gen_15_cmp_pReg_1, Q(0)=>gen_15_cmp_pReg_0);
   gen_15_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>gen_24_cmp_pInit_32, 
      a(31)=>gen_24_cmp_pInit_32, a(30)=>gen_15_cmp_pReg_30, a(29)=>
      gen_15_cmp_pReg_29, a(28)=>gen_15_cmp_pReg_28, a(27)=>
      gen_15_cmp_pReg_27, a(26)=>gen_15_cmp_pReg_26, a(25)=>
      gen_15_cmp_pReg_25, a(24)=>gen_15_cmp_pReg_24, a(23)=>
      gen_15_cmp_pReg_23, a(22)=>gen_15_cmp_pReg_22, a(21)=>
      gen_15_cmp_pReg_21, a(20)=>gen_15_cmp_pReg_20, a(19)=>
      gen_15_cmp_pReg_19, a(18)=>gen_15_cmp_pReg_18, a(17)=>
      gen_15_cmp_pReg_17, a(16)=>gen_15_cmp_pReg_16, a(15)=>
      gen_15_cmp_pReg_15, a(14)=>gen_15_cmp_pReg_14, a(13)=>
      gen_15_cmp_pReg_13, a(12)=>gen_15_cmp_pReg_12, a(11)=>
      gen_15_cmp_pReg_11, a(10)=>gen_15_cmp_pReg_10, a(9)=>gen_15_cmp_pReg_9, 
      a(8)=>gen_15_cmp_pReg_8, a(7)=>gen_15_cmp_pReg_7, a(6)=>
      gen_15_cmp_pReg_6, a(5)=>gen_15_cmp_pReg_5, a(4)=>gen_15_cmp_pReg_4, 
      a(3)=>gen_15_cmp_pReg_3, a(2)=>gen_15_cmp_pReg_2, a(1)=>
      gen_15_cmp_pReg_1, a(0)=>gen_15_cmp_pReg_0, b(32)=>gen_24_cmp_pInit_32, 
      b(31)=>gen_24_cmp_pInit_32, b(30)=>gen_24_cmp_pInit_32, b(29)=>
      gen_24_cmp_pInit_32, b(28)=>gen_24_cmp_pInit_32, b(27)=>
      gen_24_cmp_pInit_32, b(26)=>gen_24_cmp_pInit_32, b(25)=>
      gen_24_cmp_pInit_32, b(24)=>gen_24_cmp_pInit_32, b(23)=>
      gen_24_cmp_pInit_32, b(22)=>gen_24_cmp_pInit_32, b(21)=>
      gen_24_cmp_pInit_32, b(20)=>gen_24_cmp_pInit_32, b(19)=>
      gen_24_cmp_pInit_32, b(18)=>gen_24_cmp_pInit_32, b(17)=>
      gen_24_cmp_pInit_32, b(16)=>gen_24_cmp_pInit_32, b(15)=>
      gen_24_cmp_pInit_32, b(14)=>gen_24_cmp_pInit_32, b(13)=>
      gen_24_cmp_pInit_32, b(12)=>gen_24_cmp_pInit_32, b(11)=>
      gen_24_cmp_pInit_32, b(10)=>gen_24_cmp_pInit_32, b(9)=>
      gen_24_cmp_pInit_32, b(8)=>filter_15_7, b(7)=>filter_15_6, b(6)=>
      filter_15_5, b(5)=>filter_15_4, b(4)=>filter_15_3, b(3)=>filter_15_2, 
      b(2)=>filter_15_1, b(1)=>filter_15_0, b(0)=>gen_24_cmp_pInit_32, sel=>
      nx11902, f(32)=>DANGLING(47), f(31)=>DANGLING(48), f(30)=>
      gen_15_cmp_pMux_30, f(29)=>gen_15_cmp_pMux_29, f(28)=>
      gen_15_cmp_pMux_28, f(27)=>gen_15_cmp_pMux_27, f(26)=>
      gen_15_cmp_pMux_26, f(25)=>gen_15_cmp_pMux_25, f(24)=>
      gen_15_cmp_pMux_24, f(23)=>gen_15_cmp_pMux_23, f(22)=>
      gen_15_cmp_pMux_22, f(21)=>gen_15_cmp_pMux_21, f(20)=>
      gen_15_cmp_pMux_20, f(19)=>gen_15_cmp_pMux_19, f(18)=>
      gen_15_cmp_pMux_18, f(17)=>gen_15_cmp_pMux_17, f(16)=>
      gen_15_cmp_pMux_16, f(15)=>gen_15_cmp_pMux_15, f(14)=>
      gen_15_cmp_pMux_14, f(13)=>gen_15_cmp_pMux_13, f(12)=>
      gen_15_cmp_pMux_12, f(11)=>gen_15_cmp_pMux_11, f(10)=>
      gen_15_cmp_pMux_10, f(9)=>gen_15_cmp_pMux_9, f(8)=>gen_15_cmp_pMux_8, 
      f(7)=>gen_15_cmp_pMux_7, f(6)=>gen_15_cmp_pMux_6, f(5)=>
      gen_15_cmp_pMux_5, f(4)=>gen_15_cmp_pMux_4, f(3)=>gen_15_cmp_pMux_3, 
      f(2)=>gen_15_cmp_pMux_2, f(1)=>gen_15_cmp_pMux_1, f(0)=>
      gen_15_cmp_pMux_0);
   gen_15_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>
      gen_24_cmp_pInit_32, a(22)=>gen_24_cmp_pInit_32, a(21)=>
      gen_15_cmp_pMux_30, a(20)=>gen_15_cmp_pMux_29, a(19)=>
      gen_15_cmp_pMux_28, a(18)=>gen_15_cmp_pMux_27, a(17)=>
      gen_15_cmp_pMux_26, a(16)=>gen_15_cmp_pMux_25, a(15)=>
      gen_15_cmp_pMux_24, a(14)=>gen_15_cmp_pMux_23, a(13)=>
      gen_15_cmp_pMux_22, a(12)=>gen_15_cmp_pMux_21, a(11)=>
      gen_15_cmp_pMux_20, a(10)=>gen_15_cmp_pMux_19, a(9)=>
      gen_15_cmp_pMux_18, a(8)=>gen_15_cmp_pMux_17, a(7)=>gen_15_cmp_pMux_16, 
      a(6)=>gen_15_cmp_pMux_15, a(5)=>gen_15_cmp_pMux_14, a(4)=>
      gen_15_cmp_pMux_13, a(3)=>gen_15_cmp_pMux_12, a(2)=>gen_15_cmp_pMux_11, 
      a(1)=>gen_15_cmp_pMux_10, a(0)=>gen_15_cmp_pMux_9, b(23)=>nx10542, 
      b(22)=>nx10542, b(21)=>nx10540, b(20)=>nx10548, b(19)=>nx10546, b(18)
      =>nx10544, b(17)=>nx10542, b(16)=>nx10540, b(15)=>
      gen_15_cmp_BSCmp_op2_15, b(14)=>gen_15_cmp_BSCmp_op2_14, b(13)=>
      gen_15_cmp_BSCmp_op2_13, b(12)=>gen_15_cmp_BSCmp_op2_12, b(11)=>
      gen_15_cmp_BSCmp_op2_11, b(10)=>gen_15_cmp_BSCmp_op2_10, b(9)=>
      gen_15_cmp_BSCmp_op2_9, b(8)=>gen_15_cmp_BSCmp_op2_8, b(7)=>
      gen_15_cmp_BSCmp_op2_7, b(6)=>gen_15_cmp_BSCmp_op2_6, b(5)=>
      gen_15_cmp_BSCmp_op2_5, b(4)=>gen_15_cmp_BSCmp_op2_4, b(3)=>
      gen_15_cmp_BSCmp_op2_3, b(2)=>gen_15_cmp_BSCmp_op2_2, b(1)=>
      gen_15_cmp_BSCmp_op2_1, b(0)=>gen_15_cmp_BSCmp_op2_0, carryIn=>
      gen_15_cmp_BSCmp_carryIn, sum(23)=>gen_15_cmp_pBs_30, sum(22)=>
      gen_15_cmp_pBs_29, sum(21)=>gen_15_cmp_pBs_28, sum(20)=>
      gen_15_cmp_pBs_27, sum(19)=>gen_15_cmp_pBs_26, sum(18)=>
      gen_15_cmp_pBs_25, sum(17)=>gen_15_cmp_pBs_24, sum(16)=>
      gen_15_cmp_pBs_23, sum(15)=>outputs_15_15, sum(14)=>outputs_15_14, 
      sum(13)=>outputs_15_13, sum(12)=>outputs_15_12, sum(11)=>outputs_15_11, 
      sum(10)=>outputs_15_10, sum(9)=>outputs_15_9, sum(8)=>outputs_15_8, 
      sum(7)=>outputs_15_7, sum(6)=>outputs_15_6, sum(5)=>outputs_15_5, 
      sum(4)=>outputs_15_4, sum(3)=>outputs_15_3, sum(2)=>outputs_15_2, 
      sum(1)=>outputs_15_1, sum(0)=>outputs_15_0, carryOut=>DANGLING(49));
   gen_14_cmp_pRegCmp : Reg_33 port map ( D(32)=>gen_24_cmp_pInit_32, D(31)
      =>gen_24_cmp_pInit_32, D(30)=>gen_14_cmp_pBs_30, D(29)=>
      gen_14_cmp_pBs_29, D(28)=>gen_14_cmp_pBs_28, D(27)=>gen_14_cmp_pBs_27, 
      D(26)=>gen_14_cmp_pBs_26, D(25)=>gen_14_cmp_pBs_25, D(24)=>
      gen_14_cmp_pBs_24, D(23)=>gen_14_cmp_pBs_23, D(22)=>outputs_14_15, 
      D(21)=>outputs_14_14, D(20)=>outputs_14_13, D(19)=>outputs_14_12, 
      D(18)=>outputs_14_11, D(17)=>outputs_14_10, D(16)=>outputs_14_9, D(15)
      =>outputs_14_8, D(14)=>outputs_14_7, D(13)=>outputs_14_6, D(12)=>
      outputs_14_5, D(11)=>outputs_14_4, D(10)=>outputs_14_3, D(9)=>
      outputs_14_2, D(8)=>outputs_14_1, D(7)=>outputs_14_0, D(6)=>
      gen_14_cmp_pMux_8, D(5)=>gen_14_cmp_pMux_7, D(4)=>gen_14_cmp_pMux_6, 
      D(3)=>gen_14_cmp_pMux_5, D(2)=>gen_14_cmp_pMux_4, D(1)=>
      gen_14_cmp_pMux_3, D(0)=>nx10250, en=>nx11922, clk=>nx10124, rst=>rst, 
      Q(32)=>DANGLING(50), Q(31)=>DANGLING(51), Q(30)=>gen_14_cmp_pReg_30, 
      Q(29)=>gen_14_cmp_pReg_29, Q(28)=>gen_14_cmp_pReg_28, Q(27)=>
      gen_14_cmp_pReg_27, Q(26)=>gen_14_cmp_pReg_26, Q(25)=>
      gen_14_cmp_pReg_25, Q(24)=>gen_14_cmp_pReg_24, Q(23)=>
      gen_14_cmp_pReg_23, Q(22)=>gen_14_cmp_pReg_22, Q(21)=>
      gen_14_cmp_pReg_21, Q(20)=>gen_14_cmp_pReg_20, Q(19)=>
      gen_14_cmp_pReg_19, Q(18)=>gen_14_cmp_pReg_18, Q(17)=>
      gen_14_cmp_pReg_17, Q(16)=>gen_14_cmp_pReg_16, Q(15)=>
      gen_14_cmp_pReg_15, Q(14)=>gen_14_cmp_pReg_14, Q(13)=>
      gen_14_cmp_pReg_13, Q(12)=>gen_14_cmp_pReg_12, Q(11)=>
      gen_14_cmp_pReg_11, Q(10)=>gen_14_cmp_pReg_10, Q(9)=>gen_14_cmp_pReg_9, 
      Q(8)=>gen_14_cmp_pReg_8, Q(7)=>gen_14_cmp_pReg_7, Q(6)=>
      gen_14_cmp_pReg_6, Q(5)=>gen_14_cmp_pReg_5, Q(4)=>gen_14_cmp_pReg_4, 
      Q(3)=>gen_14_cmp_pReg_3, Q(2)=>gen_14_cmp_pReg_2, Q(1)=>
      gen_14_cmp_pReg_1, Q(0)=>gen_14_cmp_pReg_0);
   gen_14_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>gen_24_cmp_pInit_32, 
      a(31)=>gen_24_cmp_pInit_32, a(30)=>gen_14_cmp_pReg_30, a(29)=>
      gen_14_cmp_pReg_29, a(28)=>gen_14_cmp_pReg_28, a(27)=>
      gen_14_cmp_pReg_27, a(26)=>gen_14_cmp_pReg_26, a(25)=>
      gen_14_cmp_pReg_25, a(24)=>gen_14_cmp_pReg_24, a(23)=>
      gen_14_cmp_pReg_23, a(22)=>gen_14_cmp_pReg_22, a(21)=>
      gen_14_cmp_pReg_21, a(20)=>gen_14_cmp_pReg_20, a(19)=>
      gen_14_cmp_pReg_19, a(18)=>gen_14_cmp_pReg_18, a(17)=>
      gen_14_cmp_pReg_17, a(16)=>gen_14_cmp_pReg_16, a(15)=>
      gen_14_cmp_pReg_15, a(14)=>gen_14_cmp_pReg_14, a(13)=>
      gen_14_cmp_pReg_13, a(12)=>gen_14_cmp_pReg_12, a(11)=>
      gen_14_cmp_pReg_11, a(10)=>gen_14_cmp_pReg_10, a(9)=>gen_14_cmp_pReg_9, 
      a(8)=>gen_14_cmp_pReg_8, a(7)=>gen_14_cmp_pReg_7, a(6)=>
      gen_14_cmp_pReg_6, a(5)=>gen_14_cmp_pReg_5, a(4)=>gen_14_cmp_pReg_4, 
      a(3)=>gen_14_cmp_pReg_3, a(2)=>gen_14_cmp_pReg_2, a(1)=>
      gen_14_cmp_pReg_1, a(0)=>gen_14_cmp_pReg_0, b(32)=>gen_24_cmp_pInit_32, 
      b(31)=>gen_24_cmp_pInit_32, b(30)=>gen_24_cmp_pInit_32, b(29)=>
      gen_24_cmp_pInit_32, b(28)=>gen_24_cmp_pInit_32, b(27)=>
      gen_24_cmp_pInit_32, b(26)=>gen_24_cmp_pInit_32, b(25)=>
      gen_24_cmp_pInit_32, b(24)=>gen_24_cmp_pInit_32, b(23)=>
      gen_24_cmp_pInit_32, b(22)=>gen_24_cmp_pInit_32, b(21)=>
      gen_24_cmp_pInit_32, b(20)=>gen_24_cmp_pInit_32, b(19)=>
      gen_24_cmp_pInit_32, b(18)=>gen_24_cmp_pInit_32, b(17)=>
      gen_24_cmp_pInit_32, b(16)=>gen_24_cmp_pInit_32, b(15)=>
      gen_24_cmp_pInit_32, b(14)=>gen_24_cmp_pInit_32, b(13)=>
      gen_24_cmp_pInit_32, b(12)=>gen_24_cmp_pInit_32, b(11)=>
      gen_24_cmp_pInit_32, b(10)=>gen_24_cmp_pInit_32, b(9)=>
      gen_24_cmp_pInit_32, b(8)=>filter_14_7, b(7)=>filter_14_6, b(6)=>
      filter_14_5, b(5)=>filter_14_4, b(4)=>filter_14_3, b(3)=>filter_14_2, 
      b(2)=>filter_14_1, b(1)=>filter_14_0, b(0)=>gen_24_cmp_pInit_32, sel=>
      nx11904, f(32)=>DANGLING(52), f(31)=>DANGLING(53), f(30)=>
      gen_14_cmp_pMux_30, f(29)=>gen_14_cmp_pMux_29, f(28)=>
      gen_14_cmp_pMux_28, f(27)=>gen_14_cmp_pMux_27, f(26)=>
      gen_14_cmp_pMux_26, f(25)=>gen_14_cmp_pMux_25, f(24)=>
      gen_14_cmp_pMux_24, f(23)=>gen_14_cmp_pMux_23, f(22)=>
      gen_14_cmp_pMux_22, f(21)=>gen_14_cmp_pMux_21, f(20)=>
      gen_14_cmp_pMux_20, f(19)=>gen_14_cmp_pMux_19, f(18)=>
      gen_14_cmp_pMux_18, f(17)=>gen_14_cmp_pMux_17, f(16)=>
      gen_14_cmp_pMux_16, f(15)=>gen_14_cmp_pMux_15, f(14)=>
      gen_14_cmp_pMux_14, f(13)=>gen_14_cmp_pMux_13, f(12)=>
      gen_14_cmp_pMux_12, f(11)=>gen_14_cmp_pMux_11, f(10)=>
      gen_14_cmp_pMux_10, f(9)=>gen_14_cmp_pMux_9, f(8)=>gen_14_cmp_pMux_8, 
      f(7)=>gen_14_cmp_pMux_7, f(6)=>gen_14_cmp_pMux_6, f(5)=>
      gen_14_cmp_pMux_5, f(4)=>gen_14_cmp_pMux_4, f(3)=>gen_14_cmp_pMux_3, 
      f(2)=>gen_14_cmp_pMux_2, f(1)=>gen_14_cmp_pMux_1, f(0)=>
      gen_14_cmp_pMux_0);
   gen_14_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>
      gen_24_cmp_pInit_32, a(22)=>gen_24_cmp_pInit_32, a(21)=>
      gen_14_cmp_pMux_30, a(20)=>gen_14_cmp_pMux_29, a(19)=>
      gen_14_cmp_pMux_28, a(18)=>gen_14_cmp_pMux_27, a(17)=>
      gen_14_cmp_pMux_26, a(16)=>gen_14_cmp_pMux_25, a(15)=>
      gen_14_cmp_pMux_24, a(14)=>gen_14_cmp_pMux_23, a(13)=>
      gen_14_cmp_pMux_22, a(12)=>gen_14_cmp_pMux_21, a(11)=>
      gen_14_cmp_pMux_20, a(10)=>gen_14_cmp_pMux_19, a(9)=>
      gen_14_cmp_pMux_18, a(8)=>gen_14_cmp_pMux_17, a(7)=>gen_14_cmp_pMux_16, 
      a(6)=>gen_14_cmp_pMux_15, a(5)=>gen_14_cmp_pMux_14, a(4)=>
      gen_14_cmp_pMux_13, a(3)=>gen_14_cmp_pMux_12, a(2)=>gen_14_cmp_pMux_11, 
      a(1)=>gen_14_cmp_pMux_10, a(0)=>gen_14_cmp_pMux_9, b(23)=>nx10554, 
      b(22)=>nx10554, b(21)=>nx10552, b(20)=>nx10560, b(19)=>nx10558, b(18)
      =>nx10556, b(17)=>nx10554, b(16)=>nx10552, b(15)=>
      gen_14_cmp_BSCmp_op2_15, b(14)=>gen_14_cmp_BSCmp_op2_14, b(13)=>
      gen_14_cmp_BSCmp_op2_13, b(12)=>gen_14_cmp_BSCmp_op2_12, b(11)=>
      gen_14_cmp_BSCmp_op2_11, b(10)=>gen_14_cmp_BSCmp_op2_10, b(9)=>
      gen_14_cmp_BSCmp_op2_9, b(8)=>gen_14_cmp_BSCmp_op2_8, b(7)=>
      gen_14_cmp_BSCmp_op2_7, b(6)=>gen_14_cmp_BSCmp_op2_6, b(5)=>
      gen_14_cmp_BSCmp_op2_5, b(4)=>gen_14_cmp_BSCmp_op2_4, b(3)=>
      gen_14_cmp_BSCmp_op2_3, b(2)=>gen_14_cmp_BSCmp_op2_2, b(1)=>
      gen_14_cmp_BSCmp_op2_1, b(0)=>gen_14_cmp_BSCmp_op2_0, carryIn=>
      gen_14_cmp_BSCmp_carryIn, sum(23)=>gen_14_cmp_pBs_30, sum(22)=>
      gen_14_cmp_pBs_29, sum(21)=>gen_14_cmp_pBs_28, sum(20)=>
      gen_14_cmp_pBs_27, sum(19)=>gen_14_cmp_pBs_26, sum(18)=>
      gen_14_cmp_pBs_25, sum(17)=>gen_14_cmp_pBs_24, sum(16)=>
      gen_14_cmp_pBs_23, sum(15)=>outputs_14_15, sum(14)=>outputs_14_14, 
      sum(13)=>outputs_14_13, sum(12)=>outputs_14_12, sum(11)=>outputs_14_11, 
      sum(10)=>outputs_14_10, sum(9)=>outputs_14_9, sum(8)=>outputs_14_8, 
      sum(7)=>outputs_14_7, sum(6)=>outputs_14_6, sum(5)=>outputs_14_5, 
      sum(4)=>outputs_14_4, sum(3)=>outputs_14_3, sum(2)=>outputs_14_2, 
      sum(1)=>outputs_14_1, sum(0)=>outputs_14_0, carryOut=>DANGLING(54));
   gen_13_cmp_pRegCmp : Reg_33 port map ( D(32)=>gen_24_cmp_pInit_32, D(31)
      =>gen_24_cmp_pInit_32, D(30)=>gen_13_cmp_pBs_30, D(29)=>
      gen_13_cmp_pBs_29, D(28)=>gen_13_cmp_pBs_28, D(27)=>gen_13_cmp_pBs_27, 
      D(26)=>gen_13_cmp_pBs_26, D(25)=>gen_13_cmp_pBs_25, D(24)=>
      gen_13_cmp_pBs_24, D(23)=>gen_13_cmp_pBs_23, D(22)=>outputs_13_15, 
      D(21)=>outputs_13_14, D(20)=>outputs_13_13, D(19)=>outputs_13_12, 
      D(18)=>outputs_13_11, D(17)=>outputs_13_10, D(16)=>outputs_13_9, D(15)
      =>outputs_13_8, D(14)=>outputs_13_7, D(13)=>outputs_13_6, D(12)=>
      outputs_13_5, D(11)=>outputs_13_4, D(10)=>outputs_13_3, D(9)=>
      outputs_13_2, D(8)=>outputs_13_1, D(7)=>outputs_13_0, D(6)=>
      gen_13_cmp_pMux_8, D(5)=>gen_13_cmp_pMux_7, D(4)=>gen_13_cmp_pMux_6, 
      D(3)=>gen_13_cmp_pMux_5, D(2)=>gen_13_cmp_pMux_4, D(1)=>
      gen_13_cmp_pMux_3, D(0)=>nx10262, en=>nx11922, clk=>nx10124, rst=>rst, 
      Q(32)=>DANGLING(55), Q(31)=>DANGLING(56), Q(30)=>gen_13_cmp_pReg_30, 
      Q(29)=>gen_13_cmp_pReg_29, Q(28)=>gen_13_cmp_pReg_28, Q(27)=>
      gen_13_cmp_pReg_27, Q(26)=>gen_13_cmp_pReg_26, Q(25)=>
      gen_13_cmp_pReg_25, Q(24)=>gen_13_cmp_pReg_24, Q(23)=>
      gen_13_cmp_pReg_23, Q(22)=>gen_13_cmp_pReg_22, Q(21)=>
      gen_13_cmp_pReg_21, Q(20)=>gen_13_cmp_pReg_20, Q(19)=>
      gen_13_cmp_pReg_19, Q(18)=>gen_13_cmp_pReg_18, Q(17)=>
      gen_13_cmp_pReg_17, Q(16)=>gen_13_cmp_pReg_16, Q(15)=>
      gen_13_cmp_pReg_15, Q(14)=>gen_13_cmp_pReg_14, Q(13)=>
      gen_13_cmp_pReg_13, Q(12)=>gen_13_cmp_pReg_12, Q(11)=>
      gen_13_cmp_pReg_11, Q(10)=>gen_13_cmp_pReg_10, Q(9)=>gen_13_cmp_pReg_9, 
      Q(8)=>gen_13_cmp_pReg_8, Q(7)=>gen_13_cmp_pReg_7, Q(6)=>
      gen_13_cmp_pReg_6, Q(5)=>gen_13_cmp_pReg_5, Q(4)=>gen_13_cmp_pReg_4, 
      Q(3)=>gen_13_cmp_pReg_3, Q(2)=>gen_13_cmp_pReg_2, Q(1)=>
      gen_13_cmp_pReg_1, Q(0)=>gen_13_cmp_pReg_0);
   gen_13_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>gen_24_cmp_pInit_32, 
      a(31)=>gen_24_cmp_pInit_32, a(30)=>gen_13_cmp_pReg_30, a(29)=>
      gen_13_cmp_pReg_29, a(28)=>gen_13_cmp_pReg_28, a(27)=>
      gen_13_cmp_pReg_27, a(26)=>gen_13_cmp_pReg_26, a(25)=>
      gen_13_cmp_pReg_25, a(24)=>gen_13_cmp_pReg_24, a(23)=>
      gen_13_cmp_pReg_23, a(22)=>gen_13_cmp_pReg_22, a(21)=>
      gen_13_cmp_pReg_21, a(20)=>gen_13_cmp_pReg_20, a(19)=>
      gen_13_cmp_pReg_19, a(18)=>gen_13_cmp_pReg_18, a(17)=>
      gen_13_cmp_pReg_17, a(16)=>gen_13_cmp_pReg_16, a(15)=>
      gen_13_cmp_pReg_15, a(14)=>gen_13_cmp_pReg_14, a(13)=>
      gen_13_cmp_pReg_13, a(12)=>gen_13_cmp_pReg_12, a(11)=>
      gen_13_cmp_pReg_11, a(10)=>gen_13_cmp_pReg_10, a(9)=>gen_13_cmp_pReg_9, 
      a(8)=>gen_13_cmp_pReg_8, a(7)=>gen_13_cmp_pReg_7, a(6)=>
      gen_13_cmp_pReg_6, a(5)=>gen_13_cmp_pReg_5, a(4)=>gen_13_cmp_pReg_4, 
      a(3)=>gen_13_cmp_pReg_3, a(2)=>gen_13_cmp_pReg_2, a(1)=>
      gen_13_cmp_pReg_1, a(0)=>gen_13_cmp_pReg_0, b(32)=>gen_24_cmp_pInit_32, 
      b(31)=>gen_24_cmp_pInit_32, b(30)=>gen_24_cmp_pInit_32, b(29)=>
      gen_24_cmp_pInit_32, b(28)=>gen_24_cmp_pInit_32, b(27)=>
      gen_24_cmp_pInit_32, b(26)=>gen_24_cmp_pInit_32, b(25)=>
      gen_24_cmp_pInit_32, b(24)=>gen_24_cmp_pInit_32, b(23)=>
      gen_24_cmp_pInit_32, b(22)=>gen_24_cmp_pInit_32, b(21)=>
      gen_24_cmp_pInit_32, b(20)=>gen_24_cmp_pInit_32, b(19)=>
      gen_24_cmp_pInit_32, b(18)=>gen_24_cmp_pInit_32, b(17)=>
      gen_24_cmp_pInit_32, b(16)=>gen_24_cmp_pInit_32, b(15)=>
      gen_24_cmp_pInit_32, b(14)=>gen_24_cmp_pInit_32, b(13)=>
      gen_24_cmp_pInit_32, b(12)=>gen_24_cmp_pInit_32, b(11)=>
      gen_24_cmp_pInit_32, b(10)=>gen_24_cmp_pInit_32, b(9)=>
      gen_24_cmp_pInit_32, b(8)=>filter_13_7, b(7)=>filter_13_6, b(6)=>
      filter_13_5, b(5)=>filter_13_4, b(4)=>filter_13_3, b(3)=>filter_13_2, 
      b(2)=>filter_13_1, b(1)=>filter_13_0, b(0)=>gen_24_cmp_pInit_32, sel=>
      nx11904, f(32)=>DANGLING(57), f(31)=>DANGLING(58), f(30)=>
      gen_13_cmp_pMux_30, f(29)=>gen_13_cmp_pMux_29, f(28)=>
      gen_13_cmp_pMux_28, f(27)=>gen_13_cmp_pMux_27, f(26)=>
      gen_13_cmp_pMux_26, f(25)=>gen_13_cmp_pMux_25, f(24)=>
      gen_13_cmp_pMux_24, f(23)=>gen_13_cmp_pMux_23, f(22)=>
      gen_13_cmp_pMux_22, f(21)=>gen_13_cmp_pMux_21, f(20)=>
      gen_13_cmp_pMux_20, f(19)=>gen_13_cmp_pMux_19, f(18)=>
      gen_13_cmp_pMux_18, f(17)=>gen_13_cmp_pMux_17, f(16)=>
      gen_13_cmp_pMux_16, f(15)=>gen_13_cmp_pMux_15, f(14)=>
      gen_13_cmp_pMux_14, f(13)=>gen_13_cmp_pMux_13, f(12)=>
      gen_13_cmp_pMux_12, f(11)=>gen_13_cmp_pMux_11, f(10)=>
      gen_13_cmp_pMux_10, f(9)=>gen_13_cmp_pMux_9, f(8)=>gen_13_cmp_pMux_8, 
      f(7)=>gen_13_cmp_pMux_7, f(6)=>gen_13_cmp_pMux_6, f(5)=>
      gen_13_cmp_pMux_5, f(4)=>gen_13_cmp_pMux_4, f(3)=>gen_13_cmp_pMux_3, 
      f(2)=>gen_13_cmp_pMux_2, f(1)=>gen_13_cmp_pMux_1, f(0)=>
      gen_13_cmp_pMux_0);
   gen_13_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>
      gen_24_cmp_pInit_32, a(22)=>gen_24_cmp_pInit_32, a(21)=>
      gen_13_cmp_pMux_30, a(20)=>gen_13_cmp_pMux_29, a(19)=>
      gen_13_cmp_pMux_28, a(18)=>gen_13_cmp_pMux_27, a(17)=>
      gen_13_cmp_pMux_26, a(16)=>gen_13_cmp_pMux_25, a(15)=>
      gen_13_cmp_pMux_24, a(14)=>gen_13_cmp_pMux_23, a(13)=>
      gen_13_cmp_pMux_22, a(12)=>gen_13_cmp_pMux_21, a(11)=>
      gen_13_cmp_pMux_20, a(10)=>gen_13_cmp_pMux_19, a(9)=>
      gen_13_cmp_pMux_18, a(8)=>gen_13_cmp_pMux_17, a(7)=>gen_13_cmp_pMux_16, 
      a(6)=>gen_13_cmp_pMux_15, a(5)=>gen_13_cmp_pMux_14, a(4)=>
      gen_13_cmp_pMux_13, a(3)=>gen_13_cmp_pMux_12, a(2)=>gen_13_cmp_pMux_11, 
      a(1)=>gen_13_cmp_pMux_10, a(0)=>gen_13_cmp_pMux_9, b(23)=>nx10566, 
      b(22)=>nx10566, b(21)=>nx10564, b(20)=>nx10572, b(19)=>nx10570, b(18)
      =>nx10568, b(17)=>nx10566, b(16)=>nx10564, b(15)=>
      gen_13_cmp_BSCmp_op2_15, b(14)=>gen_13_cmp_BSCmp_op2_14, b(13)=>
      gen_13_cmp_BSCmp_op2_13, b(12)=>gen_13_cmp_BSCmp_op2_12, b(11)=>
      gen_13_cmp_BSCmp_op2_11, b(10)=>gen_13_cmp_BSCmp_op2_10, b(9)=>
      gen_13_cmp_BSCmp_op2_9, b(8)=>gen_13_cmp_BSCmp_op2_8, b(7)=>
      gen_13_cmp_BSCmp_op2_7, b(6)=>gen_13_cmp_BSCmp_op2_6, b(5)=>
      gen_13_cmp_BSCmp_op2_5, b(4)=>gen_13_cmp_BSCmp_op2_4, b(3)=>
      gen_13_cmp_BSCmp_op2_3, b(2)=>gen_13_cmp_BSCmp_op2_2, b(1)=>
      gen_13_cmp_BSCmp_op2_1, b(0)=>gen_13_cmp_BSCmp_op2_0, carryIn=>
      gen_13_cmp_BSCmp_carryIn, sum(23)=>gen_13_cmp_pBs_30, sum(22)=>
      gen_13_cmp_pBs_29, sum(21)=>gen_13_cmp_pBs_28, sum(20)=>
      gen_13_cmp_pBs_27, sum(19)=>gen_13_cmp_pBs_26, sum(18)=>
      gen_13_cmp_pBs_25, sum(17)=>gen_13_cmp_pBs_24, sum(16)=>
      gen_13_cmp_pBs_23, sum(15)=>outputs_13_15, sum(14)=>outputs_13_14, 
      sum(13)=>outputs_13_13, sum(12)=>outputs_13_12, sum(11)=>outputs_13_11, 
      sum(10)=>outputs_13_10, sum(9)=>outputs_13_9, sum(8)=>outputs_13_8, 
      sum(7)=>outputs_13_7, sum(6)=>outputs_13_6, sum(5)=>outputs_13_5, 
      sum(4)=>outputs_13_4, sum(3)=>outputs_13_3, sum(2)=>outputs_13_2, 
      sum(1)=>outputs_13_1, sum(0)=>outputs_13_0, carryOut=>DANGLING(59));
   gen_12_cmp_pRegCmp : Reg_33 port map ( D(32)=>gen_24_cmp_pInit_32, D(31)
      =>gen_24_cmp_pInit_32, D(30)=>gen_12_cmp_pBs_30, D(29)=>
      gen_12_cmp_pBs_29, D(28)=>gen_12_cmp_pBs_28, D(27)=>gen_12_cmp_pBs_27, 
      D(26)=>gen_12_cmp_pBs_26, D(25)=>gen_12_cmp_pBs_25, D(24)=>
      gen_12_cmp_pBs_24, D(23)=>gen_12_cmp_pBs_23, D(22)=>outputs_12_15, 
      D(21)=>outputs_12_14, D(20)=>outputs_12_13, D(19)=>outputs_12_12, 
      D(18)=>outputs_12_11, D(17)=>outputs_12_10, D(16)=>outputs_12_9, D(15)
      =>outputs_12_8, D(14)=>outputs_12_7, D(13)=>outputs_12_6, D(12)=>
      outputs_12_5, D(11)=>outputs_12_4, D(10)=>outputs_12_3, D(9)=>
      outputs_12_2, D(8)=>outputs_12_1, D(7)=>outputs_12_0, D(6)=>
      gen_12_cmp_pMux_8, D(5)=>gen_12_cmp_pMux_7, D(4)=>gen_12_cmp_pMux_6, 
      D(3)=>gen_12_cmp_pMux_5, D(2)=>gen_12_cmp_pMux_4, D(1)=>
      gen_12_cmp_pMux_3, D(0)=>nx10274, en=>nx11922, clk=>nx10124, rst=>rst, 
      Q(32)=>DANGLING(60), Q(31)=>DANGLING(61), Q(30)=>gen_12_cmp_pReg_30, 
      Q(29)=>gen_12_cmp_pReg_29, Q(28)=>gen_12_cmp_pReg_28, Q(27)=>
      gen_12_cmp_pReg_27, Q(26)=>gen_12_cmp_pReg_26, Q(25)=>
      gen_12_cmp_pReg_25, Q(24)=>gen_12_cmp_pReg_24, Q(23)=>
      gen_12_cmp_pReg_23, Q(22)=>gen_12_cmp_pReg_22, Q(21)=>
      gen_12_cmp_pReg_21, Q(20)=>gen_12_cmp_pReg_20, Q(19)=>
      gen_12_cmp_pReg_19, Q(18)=>gen_12_cmp_pReg_18, Q(17)=>
      gen_12_cmp_pReg_17, Q(16)=>gen_12_cmp_pReg_16, Q(15)=>
      gen_12_cmp_pReg_15, Q(14)=>gen_12_cmp_pReg_14, Q(13)=>
      gen_12_cmp_pReg_13, Q(12)=>gen_12_cmp_pReg_12, Q(11)=>
      gen_12_cmp_pReg_11, Q(10)=>gen_12_cmp_pReg_10, Q(9)=>gen_12_cmp_pReg_9, 
      Q(8)=>gen_12_cmp_pReg_8, Q(7)=>gen_12_cmp_pReg_7, Q(6)=>
      gen_12_cmp_pReg_6, Q(5)=>gen_12_cmp_pReg_5, Q(4)=>gen_12_cmp_pReg_4, 
      Q(3)=>gen_12_cmp_pReg_3, Q(2)=>gen_12_cmp_pReg_2, Q(1)=>
      gen_12_cmp_pReg_1, Q(0)=>gen_12_cmp_pReg_0);
   gen_12_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>gen_24_cmp_pInit_32, 
      a(31)=>gen_24_cmp_pInit_32, a(30)=>gen_12_cmp_pReg_30, a(29)=>
      gen_12_cmp_pReg_29, a(28)=>gen_12_cmp_pReg_28, a(27)=>
      gen_12_cmp_pReg_27, a(26)=>gen_12_cmp_pReg_26, a(25)=>
      gen_12_cmp_pReg_25, a(24)=>gen_12_cmp_pReg_24, a(23)=>
      gen_12_cmp_pReg_23, a(22)=>gen_12_cmp_pReg_22, a(21)=>
      gen_12_cmp_pReg_21, a(20)=>gen_12_cmp_pReg_20, a(19)=>
      gen_12_cmp_pReg_19, a(18)=>gen_12_cmp_pReg_18, a(17)=>
      gen_12_cmp_pReg_17, a(16)=>gen_12_cmp_pReg_16, a(15)=>
      gen_12_cmp_pReg_15, a(14)=>gen_12_cmp_pReg_14, a(13)=>
      gen_12_cmp_pReg_13, a(12)=>gen_12_cmp_pReg_12, a(11)=>
      gen_12_cmp_pReg_11, a(10)=>gen_12_cmp_pReg_10, a(9)=>gen_12_cmp_pReg_9, 
      a(8)=>gen_12_cmp_pReg_8, a(7)=>gen_12_cmp_pReg_7, a(6)=>
      gen_12_cmp_pReg_6, a(5)=>gen_12_cmp_pReg_5, a(4)=>gen_12_cmp_pReg_4, 
      a(3)=>gen_12_cmp_pReg_3, a(2)=>gen_12_cmp_pReg_2, a(1)=>
      gen_12_cmp_pReg_1, a(0)=>gen_12_cmp_pReg_0, b(32)=>gen_24_cmp_pInit_32, 
      b(31)=>gen_24_cmp_pInit_32, b(30)=>gen_24_cmp_pInit_32, b(29)=>
      gen_24_cmp_pInit_32, b(28)=>gen_24_cmp_pInit_32, b(27)=>
      gen_24_cmp_pInit_32, b(26)=>gen_24_cmp_pInit_32, b(25)=>
      gen_24_cmp_pInit_32, b(24)=>gen_24_cmp_pInit_32, b(23)=>
      gen_24_cmp_pInit_32, b(22)=>gen_24_cmp_pInit_32, b(21)=>
      gen_24_cmp_pInit_32, b(20)=>gen_24_cmp_pInit_32, b(19)=>
      gen_24_cmp_pInit_32, b(18)=>gen_24_cmp_pInit_32, b(17)=>
      gen_24_cmp_pInit_32, b(16)=>gen_24_cmp_pInit_32, b(15)=>
      gen_24_cmp_pInit_32, b(14)=>gen_24_cmp_pInit_32, b(13)=>
      gen_24_cmp_pInit_32, b(12)=>gen_24_cmp_pInit_32, b(11)=>
      gen_24_cmp_pInit_32, b(10)=>gen_24_cmp_pInit_32, b(9)=>
      gen_24_cmp_pInit_32, b(8)=>filter_12_7, b(7)=>filter_12_6, b(6)=>
      filter_12_5, b(5)=>filter_12_4, b(4)=>filter_12_3, b(3)=>filter_12_2, 
      b(2)=>filter_12_1, b(1)=>filter_12_0, b(0)=>gen_24_cmp_pInit_32, sel=>
      nx11904, f(32)=>DANGLING(62), f(31)=>DANGLING(63), f(30)=>
      gen_12_cmp_pMux_30, f(29)=>gen_12_cmp_pMux_29, f(28)=>
      gen_12_cmp_pMux_28, f(27)=>gen_12_cmp_pMux_27, f(26)=>
      gen_12_cmp_pMux_26, f(25)=>gen_12_cmp_pMux_25, f(24)=>
      gen_12_cmp_pMux_24, f(23)=>gen_12_cmp_pMux_23, f(22)=>
      gen_12_cmp_pMux_22, f(21)=>gen_12_cmp_pMux_21, f(20)=>
      gen_12_cmp_pMux_20, f(19)=>gen_12_cmp_pMux_19, f(18)=>
      gen_12_cmp_pMux_18, f(17)=>gen_12_cmp_pMux_17, f(16)=>
      gen_12_cmp_pMux_16, f(15)=>gen_12_cmp_pMux_15, f(14)=>
      gen_12_cmp_pMux_14, f(13)=>gen_12_cmp_pMux_13, f(12)=>
      gen_12_cmp_pMux_12, f(11)=>gen_12_cmp_pMux_11, f(10)=>
      gen_12_cmp_pMux_10, f(9)=>gen_12_cmp_pMux_9, f(8)=>gen_12_cmp_pMux_8, 
      f(7)=>gen_12_cmp_pMux_7, f(6)=>gen_12_cmp_pMux_6, f(5)=>
      gen_12_cmp_pMux_5, f(4)=>gen_12_cmp_pMux_4, f(3)=>gen_12_cmp_pMux_3, 
      f(2)=>gen_12_cmp_pMux_2, f(1)=>gen_12_cmp_pMux_1, f(0)=>
      gen_12_cmp_pMux_0);
   gen_12_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>
      gen_24_cmp_pInit_32, a(22)=>gen_24_cmp_pInit_32, a(21)=>
      gen_12_cmp_pMux_30, a(20)=>gen_12_cmp_pMux_29, a(19)=>
      gen_12_cmp_pMux_28, a(18)=>gen_12_cmp_pMux_27, a(17)=>
      gen_12_cmp_pMux_26, a(16)=>gen_12_cmp_pMux_25, a(15)=>
      gen_12_cmp_pMux_24, a(14)=>gen_12_cmp_pMux_23, a(13)=>
      gen_12_cmp_pMux_22, a(12)=>gen_12_cmp_pMux_21, a(11)=>
      gen_12_cmp_pMux_20, a(10)=>gen_12_cmp_pMux_19, a(9)=>
      gen_12_cmp_pMux_18, a(8)=>gen_12_cmp_pMux_17, a(7)=>gen_12_cmp_pMux_16, 
      a(6)=>gen_12_cmp_pMux_15, a(5)=>gen_12_cmp_pMux_14, a(4)=>
      gen_12_cmp_pMux_13, a(3)=>gen_12_cmp_pMux_12, a(2)=>gen_12_cmp_pMux_11, 
      a(1)=>gen_12_cmp_pMux_10, a(0)=>gen_12_cmp_pMux_9, b(23)=>nx10578, 
      b(22)=>nx10578, b(21)=>nx10576, b(20)=>nx10584, b(19)=>nx10582, b(18)
      =>nx10580, b(17)=>nx10578, b(16)=>nx10576, b(15)=>
      gen_12_cmp_BSCmp_op2_15, b(14)=>gen_12_cmp_BSCmp_op2_14, b(13)=>
      gen_12_cmp_BSCmp_op2_13, b(12)=>gen_12_cmp_BSCmp_op2_12, b(11)=>
      gen_12_cmp_BSCmp_op2_11, b(10)=>gen_12_cmp_BSCmp_op2_10, b(9)=>
      gen_12_cmp_BSCmp_op2_9, b(8)=>gen_12_cmp_BSCmp_op2_8, b(7)=>
      gen_12_cmp_BSCmp_op2_7, b(6)=>gen_12_cmp_BSCmp_op2_6, b(5)=>
      gen_12_cmp_BSCmp_op2_5, b(4)=>gen_12_cmp_BSCmp_op2_4, b(3)=>
      gen_12_cmp_BSCmp_op2_3, b(2)=>gen_12_cmp_BSCmp_op2_2, b(1)=>
      gen_12_cmp_BSCmp_op2_1, b(0)=>gen_12_cmp_BSCmp_op2_0, carryIn=>
      gen_12_cmp_BSCmp_carryIn, sum(23)=>gen_12_cmp_pBs_30, sum(22)=>
      gen_12_cmp_pBs_29, sum(21)=>gen_12_cmp_pBs_28, sum(20)=>
      gen_12_cmp_pBs_27, sum(19)=>gen_12_cmp_pBs_26, sum(18)=>
      gen_12_cmp_pBs_25, sum(17)=>gen_12_cmp_pBs_24, sum(16)=>
      gen_12_cmp_pBs_23, sum(15)=>outputs_12_15, sum(14)=>outputs_12_14, 
      sum(13)=>outputs_12_13, sum(12)=>outputs_12_12, sum(11)=>outputs_12_11, 
      sum(10)=>outputs_12_10, sum(9)=>outputs_12_9, sum(8)=>outputs_12_8, 
      sum(7)=>outputs_12_7, sum(6)=>outputs_12_6, sum(5)=>outputs_12_5, 
      sum(4)=>outputs_12_4, sum(3)=>outputs_12_3, sum(2)=>outputs_12_2, 
      sum(1)=>outputs_12_1, sum(0)=>outputs_12_0, carryOut=>DANGLING(64));
   gen_11_cmp_pRegCmp : Reg_33 port map ( D(32)=>gen_24_cmp_pInit_32, D(31)
      =>gen_24_cmp_pInit_32, D(30)=>gen_11_cmp_pBs_30, D(29)=>
      gen_11_cmp_pBs_29, D(28)=>gen_11_cmp_pBs_28, D(27)=>gen_11_cmp_pBs_27, 
      D(26)=>gen_11_cmp_pBs_26, D(25)=>gen_11_cmp_pBs_25, D(24)=>
      gen_11_cmp_pBs_24, D(23)=>gen_11_cmp_pBs_23, D(22)=>outputs_11_15, 
      D(21)=>outputs_11_14, D(20)=>outputs_11_13, D(19)=>outputs_11_12, 
      D(18)=>outputs_11_11, D(17)=>outputs_11_10, D(16)=>outputs_11_9, D(15)
      =>outputs_11_8, D(14)=>outputs_11_7, D(13)=>outputs_11_6, D(12)=>
      outputs_11_5, D(11)=>outputs_11_4, D(10)=>outputs_11_3, D(9)=>
      outputs_11_2, D(8)=>outputs_11_1, D(7)=>outputs_11_0, D(6)=>
      gen_11_cmp_pMux_8, D(5)=>gen_11_cmp_pMux_7, D(4)=>gen_11_cmp_pMux_6, 
      D(3)=>gen_11_cmp_pMux_5, D(2)=>gen_11_cmp_pMux_4, D(1)=>
      gen_11_cmp_pMux_3, D(0)=>nx10286, en=>nx10882, clk=>nx10124, rst=>rst, 
      Q(32)=>DANGLING(65), Q(31)=>DANGLING(66), Q(30)=>gen_11_cmp_pReg_30, 
      Q(29)=>gen_11_cmp_pReg_29, Q(28)=>gen_11_cmp_pReg_28, Q(27)=>
      gen_11_cmp_pReg_27, Q(26)=>gen_11_cmp_pReg_26, Q(25)=>
      gen_11_cmp_pReg_25, Q(24)=>gen_11_cmp_pReg_24, Q(23)=>
      gen_11_cmp_pReg_23, Q(22)=>gen_11_cmp_pReg_22, Q(21)=>
      gen_11_cmp_pReg_21, Q(20)=>gen_11_cmp_pReg_20, Q(19)=>
      gen_11_cmp_pReg_19, Q(18)=>gen_11_cmp_pReg_18, Q(17)=>
      gen_11_cmp_pReg_17, Q(16)=>gen_11_cmp_pReg_16, Q(15)=>
      gen_11_cmp_pReg_15, Q(14)=>gen_11_cmp_pReg_14, Q(13)=>
      gen_11_cmp_pReg_13, Q(12)=>gen_11_cmp_pReg_12, Q(11)=>
      gen_11_cmp_pReg_11, Q(10)=>gen_11_cmp_pReg_10, Q(9)=>gen_11_cmp_pReg_9, 
      Q(8)=>gen_11_cmp_pReg_8, Q(7)=>gen_11_cmp_pReg_7, Q(6)=>
      gen_11_cmp_pReg_6, Q(5)=>gen_11_cmp_pReg_5, Q(4)=>gen_11_cmp_pReg_4, 
      Q(3)=>gen_11_cmp_pReg_3, Q(2)=>gen_11_cmp_pReg_2, Q(1)=>
      gen_11_cmp_pReg_1, Q(0)=>gen_11_cmp_pReg_0);
   gen_11_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>gen_24_cmp_pInit_32, 
      a(31)=>gen_24_cmp_pInit_32, a(30)=>gen_11_cmp_pReg_30, a(29)=>
      gen_11_cmp_pReg_29, a(28)=>gen_11_cmp_pReg_28, a(27)=>
      gen_11_cmp_pReg_27, a(26)=>gen_11_cmp_pReg_26, a(25)=>
      gen_11_cmp_pReg_25, a(24)=>gen_11_cmp_pReg_24, a(23)=>
      gen_11_cmp_pReg_23, a(22)=>gen_11_cmp_pReg_22, a(21)=>
      gen_11_cmp_pReg_21, a(20)=>gen_11_cmp_pReg_20, a(19)=>
      gen_11_cmp_pReg_19, a(18)=>gen_11_cmp_pReg_18, a(17)=>
      gen_11_cmp_pReg_17, a(16)=>gen_11_cmp_pReg_16, a(15)=>
      gen_11_cmp_pReg_15, a(14)=>gen_11_cmp_pReg_14, a(13)=>
      gen_11_cmp_pReg_13, a(12)=>gen_11_cmp_pReg_12, a(11)=>
      gen_11_cmp_pReg_11, a(10)=>gen_11_cmp_pReg_10, a(9)=>gen_11_cmp_pReg_9, 
      a(8)=>gen_11_cmp_pReg_8, a(7)=>gen_11_cmp_pReg_7, a(6)=>
      gen_11_cmp_pReg_6, a(5)=>gen_11_cmp_pReg_5, a(4)=>gen_11_cmp_pReg_4, 
      a(3)=>gen_11_cmp_pReg_3, a(2)=>gen_11_cmp_pReg_2, a(1)=>
      gen_11_cmp_pReg_1, a(0)=>gen_11_cmp_pReg_0, b(32)=>gen_24_cmp_pInit_32, 
      b(31)=>gen_24_cmp_pInit_32, b(30)=>gen_24_cmp_pInit_32, b(29)=>
      gen_24_cmp_pInit_32, b(28)=>gen_24_cmp_pInit_32, b(27)=>
      gen_24_cmp_pInit_32, b(26)=>gen_24_cmp_pInit_32, b(25)=>
      gen_24_cmp_pInit_32, b(24)=>gen_24_cmp_pInit_32, b(23)=>
      gen_24_cmp_pInit_32, b(22)=>gen_24_cmp_pInit_32, b(21)=>
      gen_24_cmp_pInit_32, b(20)=>gen_24_cmp_pInit_32, b(19)=>
      gen_24_cmp_pInit_32, b(18)=>gen_24_cmp_pInit_32, b(17)=>
      gen_24_cmp_pInit_32, b(16)=>gen_24_cmp_pInit_32, b(15)=>
      gen_24_cmp_pInit_32, b(14)=>gen_24_cmp_pInit_32, b(13)=>
      gen_24_cmp_pInit_32, b(12)=>gen_24_cmp_pInit_32, b(11)=>
      gen_24_cmp_pInit_32, b(10)=>gen_24_cmp_pInit_32, b(9)=>
      gen_24_cmp_pInit_32, b(8)=>filter_11_7, b(7)=>filter_11_6, b(6)=>
      filter_11_5, b(5)=>filter_11_4, b(4)=>filter_11_3, b(3)=>filter_11_2, 
      b(2)=>filter_11_1, b(1)=>filter_11_0, b(0)=>gen_24_cmp_pInit_32, sel=>
      nx11906, f(32)=>DANGLING(67), f(31)=>DANGLING(68), f(30)=>
      gen_11_cmp_pMux_30, f(29)=>gen_11_cmp_pMux_29, f(28)=>
      gen_11_cmp_pMux_28, f(27)=>gen_11_cmp_pMux_27, f(26)=>
      gen_11_cmp_pMux_26, f(25)=>gen_11_cmp_pMux_25, f(24)=>
      gen_11_cmp_pMux_24, f(23)=>gen_11_cmp_pMux_23, f(22)=>
      gen_11_cmp_pMux_22, f(21)=>gen_11_cmp_pMux_21, f(20)=>
      gen_11_cmp_pMux_20, f(19)=>gen_11_cmp_pMux_19, f(18)=>
      gen_11_cmp_pMux_18, f(17)=>gen_11_cmp_pMux_17, f(16)=>
      gen_11_cmp_pMux_16, f(15)=>gen_11_cmp_pMux_15, f(14)=>
      gen_11_cmp_pMux_14, f(13)=>gen_11_cmp_pMux_13, f(12)=>
      gen_11_cmp_pMux_12, f(11)=>gen_11_cmp_pMux_11, f(10)=>
      gen_11_cmp_pMux_10, f(9)=>gen_11_cmp_pMux_9, f(8)=>gen_11_cmp_pMux_8, 
      f(7)=>gen_11_cmp_pMux_7, f(6)=>gen_11_cmp_pMux_6, f(5)=>
      gen_11_cmp_pMux_5, f(4)=>gen_11_cmp_pMux_4, f(3)=>gen_11_cmp_pMux_3, 
      f(2)=>gen_11_cmp_pMux_2, f(1)=>gen_11_cmp_pMux_1, f(0)=>
      gen_11_cmp_pMux_0);
   gen_11_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>
      gen_24_cmp_pInit_32, a(22)=>gen_24_cmp_pInit_32, a(21)=>
      gen_11_cmp_pMux_30, a(20)=>gen_11_cmp_pMux_29, a(19)=>
      gen_11_cmp_pMux_28, a(18)=>gen_11_cmp_pMux_27, a(17)=>
      gen_11_cmp_pMux_26, a(16)=>gen_11_cmp_pMux_25, a(15)=>
      gen_11_cmp_pMux_24, a(14)=>gen_11_cmp_pMux_23, a(13)=>
      gen_11_cmp_pMux_22, a(12)=>gen_11_cmp_pMux_21, a(11)=>
      gen_11_cmp_pMux_20, a(10)=>gen_11_cmp_pMux_19, a(9)=>
      gen_11_cmp_pMux_18, a(8)=>gen_11_cmp_pMux_17, a(7)=>gen_11_cmp_pMux_16, 
      a(6)=>gen_11_cmp_pMux_15, a(5)=>gen_11_cmp_pMux_14, a(4)=>
      gen_11_cmp_pMux_13, a(3)=>gen_11_cmp_pMux_12, a(2)=>gen_11_cmp_pMux_11, 
      a(1)=>gen_11_cmp_pMux_10, a(0)=>gen_11_cmp_pMux_9, b(23)=>nx10590, 
      b(22)=>nx10590, b(21)=>nx10588, b(20)=>nx10596, b(19)=>nx10594, b(18)
      =>nx10592, b(17)=>nx10590, b(16)=>nx10588, b(15)=>
      gen_11_cmp_BSCmp_op2_15, b(14)=>gen_11_cmp_BSCmp_op2_14, b(13)=>
      gen_11_cmp_BSCmp_op2_13, b(12)=>gen_11_cmp_BSCmp_op2_12, b(11)=>
      gen_11_cmp_BSCmp_op2_11, b(10)=>gen_11_cmp_BSCmp_op2_10, b(9)=>
      gen_11_cmp_BSCmp_op2_9, b(8)=>gen_11_cmp_BSCmp_op2_8, b(7)=>
      gen_11_cmp_BSCmp_op2_7, b(6)=>gen_11_cmp_BSCmp_op2_6, b(5)=>
      gen_11_cmp_BSCmp_op2_5, b(4)=>gen_11_cmp_BSCmp_op2_4, b(3)=>
      gen_11_cmp_BSCmp_op2_3, b(2)=>gen_11_cmp_BSCmp_op2_2, b(1)=>
      gen_11_cmp_BSCmp_op2_1, b(0)=>gen_11_cmp_BSCmp_op2_0, carryIn=>
      gen_11_cmp_BSCmp_carryIn, sum(23)=>gen_11_cmp_pBs_30, sum(22)=>
      gen_11_cmp_pBs_29, sum(21)=>gen_11_cmp_pBs_28, sum(20)=>
      gen_11_cmp_pBs_27, sum(19)=>gen_11_cmp_pBs_26, sum(18)=>
      gen_11_cmp_pBs_25, sum(17)=>gen_11_cmp_pBs_24, sum(16)=>
      gen_11_cmp_pBs_23, sum(15)=>outputs_11_15, sum(14)=>outputs_11_14, 
      sum(13)=>outputs_11_13, sum(12)=>outputs_11_12, sum(11)=>outputs_11_11, 
      sum(10)=>outputs_11_10, sum(9)=>outputs_11_9, sum(8)=>outputs_11_8, 
      sum(7)=>outputs_11_7, sum(6)=>outputs_11_6, sum(5)=>outputs_11_5, 
      sum(4)=>outputs_11_4, sum(3)=>outputs_11_3, sum(2)=>outputs_11_2, 
      sum(1)=>outputs_11_1, sum(0)=>outputs_11_0, carryOut=>DANGLING(69));
   gen_10_cmp_pRegCmp : Reg_33 port map ( D(32)=>gen_24_cmp_pInit_32, D(31)
      =>gen_24_cmp_pInit_32, D(30)=>gen_10_cmp_pBs_30, D(29)=>
      gen_10_cmp_pBs_29, D(28)=>gen_10_cmp_pBs_28, D(27)=>gen_10_cmp_pBs_27, 
      D(26)=>gen_10_cmp_pBs_26, D(25)=>gen_10_cmp_pBs_25, D(24)=>
      gen_10_cmp_pBs_24, D(23)=>gen_10_cmp_pBs_23, D(22)=>outputs_10_15, 
      D(21)=>outputs_10_14, D(20)=>outputs_10_13, D(19)=>outputs_10_12, 
      D(18)=>outputs_10_11, D(17)=>outputs_10_10, D(16)=>outputs_10_9, D(15)
      =>outputs_10_8, D(14)=>outputs_10_7, D(13)=>outputs_10_6, D(12)=>
      outputs_10_5, D(11)=>outputs_10_4, D(10)=>outputs_10_3, D(9)=>
      outputs_10_2, D(8)=>outputs_10_1, D(7)=>outputs_10_0, D(6)=>
      gen_10_cmp_pMux_8, D(5)=>gen_10_cmp_pMux_7, D(4)=>gen_10_cmp_pMux_6, 
      D(3)=>gen_10_cmp_pMux_5, D(2)=>gen_10_cmp_pMux_4, D(1)=>
      gen_10_cmp_pMux_3, D(0)=>nx10298, en=>nx11924, clk=>nx10126, rst=>rst, 
      Q(32)=>DANGLING(70), Q(31)=>DANGLING(71), Q(30)=>gen_10_cmp_pReg_30, 
      Q(29)=>gen_10_cmp_pReg_29, Q(28)=>gen_10_cmp_pReg_28, Q(27)=>
      gen_10_cmp_pReg_27, Q(26)=>gen_10_cmp_pReg_26, Q(25)=>
      gen_10_cmp_pReg_25, Q(24)=>gen_10_cmp_pReg_24, Q(23)=>
      gen_10_cmp_pReg_23, Q(22)=>gen_10_cmp_pReg_22, Q(21)=>
      gen_10_cmp_pReg_21, Q(20)=>gen_10_cmp_pReg_20, Q(19)=>
      gen_10_cmp_pReg_19, Q(18)=>gen_10_cmp_pReg_18, Q(17)=>
      gen_10_cmp_pReg_17, Q(16)=>gen_10_cmp_pReg_16, Q(15)=>
      gen_10_cmp_pReg_15, Q(14)=>gen_10_cmp_pReg_14, Q(13)=>
      gen_10_cmp_pReg_13, Q(12)=>gen_10_cmp_pReg_12, Q(11)=>
      gen_10_cmp_pReg_11, Q(10)=>gen_10_cmp_pReg_10, Q(9)=>gen_10_cmp_pReg_9, 
      Q(8)=>gen_10_cmp_pReg_8, Q(7)=>gen_10_cmp_pReg_7, Q(6)=>
      gen_10_cmp_pReg_6, Q(5)=>gen_10_cmp_pReg_5, Q(4)=>gen_10_cmp_pReg_4, 
      Q(3)=>gen_10_cmp_pReg_3, Q(2)=>gen_10_cmp_pReg_2, Q(1)=>
      gen_10_cmp_pReg_1, Q(0)=>gen_10_cmp_pReg_0);
   gen_10_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>gen_24_cmp_pInit_32, 
      a(31)=>gen_24_cmp_pInit_32, a(30)=>gen_10_cmp_pReg_30, a(29)=>
      gen_10_cmp_pReg_29, a(28)=>gen_10_cmp_pReg_28, a(27)=>
      gen_10_cmp_pReg_27, a(26)=>gen_10_cmp_pReg_26, a(25)=>
      gen_10_cmp_pReg_25, a(24)=>gen_10_cmp_pReg_24, a(23)=>
      gen_10_cmp_pReg_23, a(22)=>gen_10_cmp_pReg_22, a(21)=>
      gen_10_cmp_pReg_21, a(20)=>gen_10_cmp_pReg_20, a(19)=>
      gen_10_cmp_pReg_19, a(18)=>gen_10_cmp_pReg_18, a(17)=>
      gen_10_cmp_pReg_17, a(16)=>gen_10_cmp_pReg_16, a(15)=>
      gen_10_cmp_pReg_15, a(14)=>gen_10_cmp_pReg_14, a(13)=>
      gen_10_cmp_pReg_13, a(12)=>gen_10_cmp_pReg_12, a(11)=>
      gen_10_cmp_pReg_11, a(10)=>gen_10_cmp_pReg_10, a(9)=>gen_10_cmp_pReg_9, 
      a(8)=>gen_10_cmp_pReg_8, a(7)=>gen_10_cmp_pReg_7, a(6)=>
      gen_10_cmp_pReg_6, a(5)=>gen_10_cmp_pReg_5, a(4)=>gen_10_cmp_pReg_4, 
      a(3)=>gen_10_cmp_pReg_3, a(2)=>gen_10_cmp_pReg_2, a(1)=>
      gen_10_cmp_pReg_1, a(0)=>gen_10_cmp_pReg_0, b(32)=>gen_24_cmp_pInit_32, 
      b(31)=>gen_24_cmp_pInit_32, b(30)=>gen_24_cmp_pInit_32, b(29)=>
      gen_24_cmp_pInit_32, b(28)=>gen_24_cmp_pInit_32, b(27)=>
      gen_24_cmp_pInit_32, b(26)=>gen_24_cmp_pInit_32, b(25)=>
      gen_24_cmp_pInit_32, b(24)=>gen_24_cmp_pInit_32, b(23)=>
      gen_24_cmp_pInit_32, b(22)=>gen_24_cmp_pInit_32, b(21)=>
      gen_24_cmp_pInit_32, b(20)=>gen_24_cmp_pInit_32, b(19)=>
      gen_24_cmp_pInit_32, b(18)=>gen_24_cmp_pInit_32, b(17)=>
      gen_24_cmp_pInit_32, b(16)=>gen_24_cmp_pInit_32, b(15)=>
      gen_24_cmp_pInit_32, b(14)=>gen_24_cmp_pInit_32, b(13)=>
      gen_24_cmp_pInit_32, b(12)=>gen_24_cmp_pInit_32, b(11)=>
      gen_24_cmp_pInit_32, b(10)=>gen_24_cmp_pInit_32, b(9)=>
      gen_24_cmp_pInit_32, b(8)=>filter_10_7, b(7)=>filter_10_6, b(6)=>
      filter_10_5, b(5)=>filter_10_4, b(4)=>filter_10_3, b(3)=>filter_10_2, 
      b(2)=>filter_10_1, b(1)=>filter_10_0, b(0)=>gen_24_cmp_pInit_32, sel=>
      nx11908, f(32)=>DANGLING(72), f(31)=>DANGLING(73), f(30)=>
      gen_10_cmp_pMux_30, f(29)=>gen_10_cmp_pMux_29, f(28)=>
      gen_10_cmp_pMux_28, f(27)=>gen_10_cmp_pMux_27, f(26)=>
      gen_10_cmp_pMux_26, f(25)=>gen_10_cmp_pMux_25, f(24)=>
      gen_10_cmp_pMux_24, f(23)=>gen_10_cmp_pMux_23, f(22)=>
      gen_10_cmp_pMux_22, f(21)=>gen_10_cmp_pMux_21, f(20)=>
      gen_10_cmp_pMux_20, f(19)=>gen_10_cmp_pMux_19, f(18)=>
      gen_10_cmp_pMux_18, f(17)=>gen_10_cmp_pMux_17, f(16)=>
      gen_10_cmp_pMux_16, f(15)=>gen_10_cmp_pMux_15, f(14)=>
      gen_10_cmp_pMux_14, f(13)=>gen_10_cmp_pMux_13, f(12)=>
      gen_10_cmp_pMux_12, f(11)=>gen_10_cmp_pMux_11, f(10)=>
      gen_10_cmp_pMux_10, f(9)=>gen_10_cmp_pMux_9, f(8)=>gen_10_cmp_pMux_8, 
      f(7)=>gen_10_cmp_pMux_7, f(6)=>gen_10_cmp_pMux_6, f(5)=>
      gen_10_cmp_pMux_5, f(4)=>gen_10_cmp_pMux_4, f(3)=>gen_10_cmp_pMux_3, 
      f(2)=>gen_10_cmp_pMux_2, f(1)=>gen_10_cmp_pMux_1, f(0)=>
      gen_10_cmp_pMux_0);
   gen_10_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>
      gen_24_cmp_pInit_32, a(22)=>gen_24_cmp_pInit_32, a(21)=>
      gen_10_cmp_pMux_30, a(20)=>gen_10_cmp_pMux_29, a(19)=>
      gen_10_cmp_pMux_28, a(18)=>gen_10_cmp_pMux_27, a(17)=>
      gen_10_cmp_pMux_26, a(16)=>gen_10_cmp_pMux_25, a(15)=>
      gen_10_cmp_pMux_24, a(14)=>gen_10_cmp_pMux_23, a(13)=>
      gen_10_cmp_pMux_22, a(12)=>gen_10_cmp_pMux_21, a(11)=>
      gen_10_cmp_pMux_20, a(10)=>gen_10_cmp_pMux_19, a(9)=>
      gen_10_cmp_pMux_18, a(8)=>gen_10_cmp_pMux_17, a(7)=>gen_10_cmp_pMux_16, 
      a(6)=>gen_10_cmp_pMux_15, a(5)=>gen_10_cmp_pMux_14, a(4)=>
      gen_10_cmp_pMux_13, a(3)=>gen_10_cmp_pMux_12, a(2)=>gen_10_cmp_pMux_11, 
      a(1)=>gen_10_cmp_pMux_10, a(0)=>gen_10_cmp_pMux_9, b(23)=>nx10602, 
      b(22)=>nx10602, b(21)=>nx10600, b(20)=>nx10608, b(19)=>nx10606, b(18)
      =>nx10604, b(17)=>nx10602, b(16)=>nx10600, b(15)=>
      gen_10_cmp_BSCmp_op2_15, b(14)=>gen_10_cmp_BSCmp_op2_14, b(13)=>
      gen_10_cmp_BSCmp_op2_13, b(12)=>gen_10_cmp_BSCmp_op2_12, b(11)=>
      gen_10_cmp_BSCmp_op2_11, b(10)=>gen_10_cmp_BSCmp_op2_10, b(9)=>
      gen_10_cmp_BSCmp_op2_9, b(8)=>gen_10_cmp_BSCmp_op2_8, b(7)=>
      gen_10_cmp_BSCmp_op2_7, b(6)=>gen_10_cmp_BSCmp_op2_6, b(5)=>
      gen_10_cmp_BSCmp_op2_5, b(4)=>gen_10_cmp_BSCmp_op2_4, b(3)=>
      gen_10_cmp_BSCmp_op2_3, b(2)=>gen_10_cmp_BSCmp_op2_2, b(1)=>
      gen_10_cmp_BSCmp_op2_1, b(0)=>gen_10_cmp_BSCmp_op2_0, carryIn=>
      gen_10_cmp_BSCmp_carryIn, sum(23)=>gen_10_cmp_pBs_30, sum(22)=>
      gen_10_cmp_pBs_29, sum(21)=>gen_10_cmp_pBs_28, sum(20)=>
      gen_10_cmp_pBs_27, sum(19)=>gen_10_cmp_pBs_26, sum(18)=>
      gen_10_cmp_pBs_25, sum(17)=>gen_10_cmp_pBs_24, sum(16)=>
      gen_10_cmp_pBs_23, sum(15)=>outputs_10_15, sum(14)=>outputs_10_14, 
      sum(13)=>outputs_10_13, sum(12)=>outputs_10_12, sum(11)=>outputs_10_11, 
      sum(10)=>outputs_10_10, sum(9)=>outputs_10_9, sum(8)=>outputs_10_8, 
      sum(7)=>outputs_10_7, sum(6)=>outputs_10_6, sum(5)=>outputs_10_5, 
      sum(4)=>outputs_10_4, sum(3)=>outputs_10_3, sum(2)=>outputs_10_2, 
      sum(1)=>outputs_10_1, sum(0)=>outputs_10_0, carryOut=>DANGLING(74));
   gen_9_cmp_pRegCmp : Reg_33 port map ( D(32)=>gen_24_cmp_pInit_32, D(31)=>
      gen_24_cmp_pInit_32, D(30)=>gen_9_cmp_pBs_30, D(29)=>gen_9_cmp_pBs_29, 
      D(28)=>gen_9_cmp_pBs_28, D(27)=>gen_9_cmp_pBs_27, D(26)=>
      gen_9_cmp_pBs_26, D(25)=>gen_9_cmp_pBs_25, D(24)=>gen_9_cmp_pBs_24, 
      D(23)=>gen_9_cmp_pBs_23, D(22)=>outputs_9_15, D(21)=>outputs_9_14, 
      D(20)=>outputs_9_13, D(19)=>outputs_9_12, D(18)=>outputs_9_11, D(17)=>
      outputs_9_10, D(16)=>outputs_9_9, D(15)=>outputs_9_8, D(14)=>
      outputs_9_7, D(13)=>outputs_9_6, D(12)=>outputs_9_5, D(11)=>
      outputs_9_4, D(10)=>outputs_9_3, D(9)=>outputs_9_2, D(8)=>outputs_9_1, 
      D(7)=>outputs_9_0, D(6)=>gen_9_cmp_pMux_8, D(5)=>gen_9_cmp_pMux_7, 
      D(4)=>gen_9_cmp_pMux_6, D(3)=>gen_9_cmp_pMux_5, D(2)=>gen_9_cmp_pMux_4, 
      D(1)=>gen_9_cmp_pMux_3, D(0)=>nx10310, en=>nx11924, clk=>nx10126, rst
      =>rst, Q(32)=>DANGLING(75), Q(31)=>DANGLING(76), Q(30)=>
      gen_9_cmp_pReg_30, Q(29)=>gen_9_cmp_pReg_29, Q(28)=>gen_9_cmp_pReg_28, 
      Q(27)=>gen_9_cmp_pReg_27, Q(26)=>gen_9_cmp_pReg_26, Q(25)=>
      gen_9_cmp_pReg_25, Q(24)=>gen_9_cmp_pReg_24, Q(23)=>gen_9_cmp_pReg_23, 
      Q(22)=>gen_9_cmp_pReg_22, Q(21)=>gen_9_cmp_pReg_21, Q(20)=>
      gen_9_cmp_pReg_20, Q(19)=>gen_9_cmp_pReg_19, Q(18)=>gen_9_cmp_pReg_18, 
      Q(17)=>gen_9_cmp_pReg_17, Q(16)=>gen_9_cmp_pReg_16, Q(15)=>
      gen_9_cmp_pReg_15, Q(14)=>gen_9_cmp_pReg_14, Q(13)=>gen_9_cmp_pReg_13, 
      Q(12)=>gen_9_cmp_pReg_12, Q(11)=>gen_9_cmp_pReg_11, Q(10)=>
      gen_9_cmp_pReg_10, Q(9)=>gen_9_cmp_pReg_9, Q(8)=>gen_9_cmp_pReg_8, 
      Q(7)=>gen_9_cmp_pReg_7, Q(6)=>gen_9_cmp_pReg_6, Q(5)=>gen_9_cmp_pReg_5, 
      Q(4)=>gen_9_cmp_pReg_4, Q(3)=>gen_9_cmp_pReg_3, Q(2)=>gen_9_cmp_pReg_2, 
      Q(1)=>gen_9_cmp_pReg_1, Q(0)=>gen_9_cmp_pReg_0);
   gen_9_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>gen_24_cmp_pInit_32, 
      a(31)=>gen_24_cmp_pInit_32, a(30)=>gen_9_cmp_pReg_30, a(29)=>
      gen_9_cmp_pReg_29, a(28)=>gen_9_cmp_pReg_28, a(27)=>gen_9_cmp_pReg_27, 
      a(26)=>gen_9_cmp_pReg_26, a(25)=>gen_9_cmp_pReg_25, a(24)=>
      gen_9_cmp_pReg_24, a(23)=>gen_9_cmp_pReg_23, a(22)=>gen_9_cmp_pReg_22, 
      a(21)=>gen_9_cmp_pReg_21, a(20)=>gen_9_cmp_pReg_20, a(19)=>
      gen_9_cmp_pReg_19, a(18)=>gen_9_cmp_pReg_18, a(17)=>gen_9_cmp_pReg_17, 
      a(16)=>gen_9_cmp_pReg_16, a(15)=>gen_9_cmp_pReg_15, a(14)=>
      gen_9_cmp_pReg_14, a(13)=>gen_9_cmp_pReg_13, a(12)=>gen_9_cmp_pReg_12, 
      a(11)=>gen_9_cmp_pReg_11, a(10)=>gen_9_cmp_pReg_10, a(9)=>
      gen_9_cmp_pReg_9, a(8)=>gen_9_cmp_pReg_8, a(7)=>gen_9_cmp_pReg_7, a(6)
      =>gen_9_cmp_pReg_6, a(5)=>gen_9_cmp_pReg_5, a(4)=>gen_9_cmp_pReg_4, 
      a(3)=>gen_9_cmp_pReg_3, a(2)=>gen_9_cmp_pReg_2, a(1)=>gen_9_cmp_pReg_1, 
      a(0)=>gen_9_cmp_pReg_0, b(32)=>gen_24_cmp_pInit_32, b(31)=>
      gen_24_cmp_pInit_32, b(30)=>gen_24_cmp_pInit_32, b(29)=>
      gen_24_cmp_pInit_32, b(28)=>gen_24_cmp_pInit_32, b(27)=>
      gen_24_cmp_pInit_32, b(26)=>gen_24_cmp_pInit_32, b(25)=>
      gen_24_cmp_pInit_32, b(24)=>gen_24_cmp_pInit_32, b(23)=>
      gen_24_cmp_pInit_32, b(22)=>gen_24_cmp_pInit_32, b(21)=>
      gen_24_cmp_pInit_32, b(20)=>gen_24_cmp_pInit_32, b(19)=>
      gen_24_cmp_pInit_32, b(18)=>gen_24_cmp_pInit_32, b(17)=>
      gen_24_cmp_pInit_32, b(16)=>gen_24_cmp_pInit_32, b(15)=>
      gen_24_cmp_pInit_32, b(14)=>gen_24_cmp_pInit_32, b(13)=>
      gen_24_cmp_pInit_32, b(12)=>gen_24_cmp_pInit_32, b(11)=>
      gen_24_cmp_pInit_32, b(10)=>gen_24_cmp_pInit_32, b(9)=>
      gen_24_cmp_pInit_32, b(8)=>filter_9_7, b(7)=>filter_9_6, b(6)=>
      filter_9_5, b(5)=>filter_9_4, b(4)=>filter_9_3, b(3)=>filter_9_2, b(2)
      =>filter_9_1, b(1)=>filter_9_0, b(0)=>gen_24_cmp_pInit_32, sel=>
      nx11908, f(32)=>DANGLING(77), f(31)=>DANGLING(78), f(30)=>
      gen_9_cmp_pMux_30, f(29)=>gen_9_cmp_pMux_29, f(28)=>gen_9_cmp_pMux_28, 
      f(27)=>gen_9_cmp_pMux_27, f(26)=>gen_9_cmp_pMux_26, f(25)=>
      gen_9_cmp_pMux_25, f(24)=>gen_9_cmp_pMux_24, f(23)=>gen_9_cmp_pMux_23, 
      f(22)=>gen_9_cmp_pMux_22, f(21)=>gen_9_cmp_pMux_21, f(20)=>
      gen_9_cmp_pMux_20, f(19)=>gen_9_cmp_pMux_19, f(18)=>gen_9_cmp_pMux_18, 
      f(17)=>gen_9_cmp_pMux_17, f(16)=>gen_9_cmp_pMux_16, f(15)=>
      gen_9_cmp_pMux_15, f(14)=>gen_9_cmp_pMux_14, f(13)=>gen_9_cmp_pMux_13, 
      f(12)=>gen_9_cmp_pMux_12, f(11)=>gen_9_cmp_pMux_11, f(10)=>
      gen_9_cmp_pMux_10, f(9)=>gen_9_cmp_pMux_9, f(8)=>gen_9_cmp_pMux_8, 
      f(7)=>gen_9_cmp_pMux_7, f(6)=>gen_9_cmp_pMux_6, f(5)=>gen_9_cmp_pMux_5, 
      f(4)=>gen_9_cmp_pMux_4, f(3)=>gen_9_cmp_pMux_3, f(2)=>gen_9_cmp_pMux_2, 
      f(1)=>gen_9_cmp_pMux_1, f(0)=>gen_9_cmp_pMux_0);
   gen_9_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>
      gen_24_cmp_pInit_32, a(22)=>gen_24_cmp_pInit_32, a(21)=>
      gen_9_cmp_pMux_30, a(20)=>gen_9_cmp_pMux_29, a(19)=>gen_9_cmp_pMux_28, 
      a(18)=>gen_9_cmp_pMux_27, a(17)=>gen_9_cmp_pMux_26, a(16)=>
      gen_9_cmp_pMux_25, a(15)=>gen_9_cmp_pMux_24, a(14)=>gen_9_cmp_pMux_23, 
      a(13)=>gen_9_cmp_pMux_22, a(12)=>gen_9_cmp_pMux_21, a(11)=>
      gen_9_cmp_pMux_20, a(10)=>gen_9_cmp_pMux_19, a(9)=>gen_9_cmp_pMux_18, 
      a(8)=>gen_9_cmp_pMux_17, a(7)=>gen_9_cmp_pMux_16, a(6)=>
      gen_9_cmp_pMux_15, a(5)=>gen_9_cmp_pMux_14, a(4)=>gen_9_cmp_pMux_13, 
      a(3)=>gen_9_cmp_pMux_12, a(2)=>gen_9_cmp_pMux_11, a(1)=>
      gen_9_cmp_pMux_10, a(0)=>gen_9_cmp_pMux_9, b(23)=>nx10614, b(22)=>
      nx10614, b(21)=>nx10612, b(20)=>nx10620, b(19)=>nx10618, b(18)=>
      nx10616, b(17)=>nx10614, b(16)=>nx10612, b(15)=>gen_9_cmp_BSCmp_op2_15, 
      b(14)=>gen_9_cmp_BSCmp_op2_14, b(13)=>gen_9_cmp_BSCmp_op2_13, b(12)=>
      gen_9_cmp_BSCmp_op2_12, b(11)=>gen_9_cmp_BSCmp_op2_11, b(10)=>
      gen_9_cmp_BSCmp_op2_10, b(9)=>gen_9_cmp_BSCmp_op2_9, b(8)=>
      gen_9_cmp_BSCmp_op2_8, b(7)=>gen_9_cmp_BSCmp_op2_7, b(6)=>
      gen_9_cmp_BSCmp_op2_6, b(5)=>gen_9_cmp_BSCmp_op2_5, b(4)=>
      gen_9_cmp_BSCmp_op2_4, b(3)=>gen_9_cmp_BSCmp_op2_3, b(2)=>
      gen_9_cmp_BSCmp_op2_2, b(1)=>gen_9_cmp_BSCmp_op2_1, b(0)=>
      gen_9_cmp_BSCmp_op2_0, carryIn=>gen_9_cmp_BSCmp_carryIn, sum(23)=>
      gen_9_cmp_pBs_30, sum(22)=>gen_9_cmp_pBs_29, sum(21)=>gen_9_cmp_pBs_28, 
      sum(20)=>gen_9_cmp_pBs_27, sum(19)=>gen_9_cmp_pBs_26, sum(18)=>
      gen_9_cmp_pBs_25, sum(17)=>gen_9_cmp_pBs_24, sum(16)=>gen_9_cmp_pBs_23, 
      sum(15)=>outputs_9_15, sum(14)=>outputs_9_14, sum(13)=>outputs_9_13, 
      sum(12)=>outputs_9_12, sum(11)=>outputs_9_11, sum(10)=>outputs_9_10, 
      sum(9)=>outputs_9_9, sum(8)=>outputs_9_8, sum(7)=>outputs_9_7, sum(6)
      =>outputs_9_6, sum(5)=>outputs_9_5, sum(4)=>outputs_9_4, sum(3)=>
      outputs_9_3, sum(2)=>outputs_9_2, sum(1)=>outputs_9_1, sum(0)=>
      outputs_9_0, carryOut=>DANGLING(79));
   gen_8_cmp_pRegCmp : Reg_33 port map ( D(32)=>gen_24_cmp_pInit_32, D(31)=>
      gen_24_cmp_pInit_32, D(30)=>gen_8_cmp_pBs_30, D(29)=>gen_8_cmp_pBs_29, 
      D(28)=>gen_8_cmp_pBs_28, D(27)=>gen_8_cmp_pBs_27, D(26)=>
      gen_8_cmp_pBs_26, D(25)=>gen_8_cmp_pBs_25, D(24)=>gen_8_cmp_pBs_24, 
      D(23)=>gen_8_cmp_pBs_23, D(22)=>outputs_8_15, D(21)=>outputs_8_14, 
      D(20)=>outputs_8_13, D(19)=>outputs_8_12, D(18)=>outputs_8_11, D(17)=>
      outputs_8_10, D(16)=>outputs_8_9, D(15)=>outputs_8_8, D(14)=>
      outputs_8_7, D(13)=>outputs_8_6, D(12)=>outputs_8_5, D(11)=>
      outputs_8_4, D(10)=>outputs_8_3, D(9)=>outputs_8_2, D(8)=>outputs_8_1, 
      D(7)=>outputs_8_0, D(6)=>gen_8_cmp_pMux_8, D(5)=>gen_8_cmp_pMux_7, 
      D(4)=>gen_8_cmp_pMux_6, D(3)=>gen_8_cmp_pMux_5, D(2)=>gen_8_cmp_pMux_4, 
      D(1)=>gen_8_cmp_pMux_3, D(0)=>nx10322, en=>nx11924, clk=>nx10126, rst
      =>rst, Q(32)=>DANGLING(80), Q(31)=>DANGLING(81), Q(30)=>
      gen_8_cmp_pReg_30, Q(29)=>gen_8_cmp_pReg_29, Q(28)=>gen_8_cmp_pReg_28, 
      Q(27)=>gen_8_cmp_pReg_27, Q(26)=>gen_8_cmp_pReg_26, Q(25)=>
      gen_8_cmp_pReg_25, Q(24)=>gen_8_cmp_pReg_24, Q(23)=>gen_8_cmp_pReg_23, 
      Q(22)=>gen_8_cmp_pReg_22, Q(21)=>gen_8_cmp_pReg_21, Q(20)=>
      gen_8_cmp_pReg_20, Q(19)=>gen_8_cmp_pReg_19, Q(18)=>gen_8_cmp_pReg_18, 
      Q(17)=>gen_8_cmp_pReg_17, Q(16)=>gen_8_cmp_pReg_16, Q(15)=>
      gen_8_cmp_pReg_15, Q(14)=>gen_8_cmp_pReg_14, Q(13)=>gen_8_cmp_pReg_13, 
      Q(12)=>gen_8_cmp_pReg_12, Q(11)=>gen_8_cmp_pReg_11, Q(10)=>
      gen_8_cmp_pReg_10, Q(9)=>gen_8_cmp_pReg_9, Q(8)=>gen_8_cmp_pReg_8, 
      Q(7)=>gen_8_cmp_pReg_7, Q(6)=>gen_8_cmp_pReg_6, Q(5)=>gen_8_cmp_pReg_5, 
      Q(4)=>gen_8_cmp_pReg_4, Q(3)=>gen_8_cmp_pReg_3, Q(2)=>gen_8_cmp_pReg_2, 
      Q(1)=>gen_8_cmp_pReg_1, Q(0)=>gen_8_cmp_pReg_0);
   gen_8_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>gen_24_cmp_pInit_32, 
      a(31)=>gen_24_cmp_pInit_32, a(30)=>gen_8_cmp_pReg_30, a(29)=>
      gen_8_cmp_pReg_29, a(28)=>gen_8_cmp_pReg_28, a(27)=>gen_8_cmp_pReg_27, 
      a(26)=>gen_8_cmp_pReg_26, a(25)=>gen_8_cmp_pReg_25, a(24)=>
      gen_8_cmp_pReg_24, a(23)=>gen_8_cmp_pReg_23, a(22)=>gen_8_cmp_pReg_22, 
      a(21)=>gen_8_cmp_pReg_21, a(20)=>gen_8_cmp_pReg_20, a(19)=>
      gen_8_cmp_pReg_19, a(18)=>gen_8_cmp_pReg_18, a(17)=>gen_8_cmp_pReg_17, 
      a(16)=>gen_8_cmp_pReg_16, a(15)=>gen_8_cmp_pReg_15, a(14)=>
      gen_8_cmp_pReg_14, a(13)=>gen_8_cmp_pReg_13, a(12)=>gen_8_cmp_pReg_12, 
      a(11)=>gen_8_cmp_pReg_11, a(10)=>gen_8_cmp_pReg_10, a(9)=>
      gen_8_cmp_pReg_9, a(8)=>gen_8_cmp_pReg_8, a(7)=>gen_8_cmp_pReg_7, a(6)
      =>gen_8_cmp_pReg_6, a(5)=>gen_8_cmp_pReg_5, a(4)=>gen_8_cmp_pReg_4, 
      a(3)=>gen_8_cmp_pReg_3, a(2)=>gen_8_cmp_pReg_2, a(1)=>gen_8_cmp_pReg_1, 
      a(0)=>gen_8_cmp_pReg_0, b(32)=>gen_24_cmp_pInit_32, b(31)=>
      gen_24_cmp_pInit_32, b(30)=>gen_24_cmp_pInit_32, b(29)=>
      gen_24_cmp_pInit_32, b(28)=>gen_24_cmp_pInit_32, b(27)=>
      gen_24_cmp_pInit_32, b(26)=>gen_24_cmp_pInit_32, b(25)=>
      gen_24_cmp_pInit_32, b(24)=>gen_24_cmp_pInit_32, b(23)=>
      gen_24_cmp_pInit_32, b(22)=>gen_24_cmp_pInit_32, b(21)=>
      gen_24_cmp_pInit_32, b(20)=>gen_24_cmp_pInit_32, b(19)=>
      gen_24_cmp_pInit_32, b(18)=>gen_24_cmp_pInit_32, b(17)=>
      gen_24_cmp_pInit_32, b(16)=>gen_24_cmp_pInit_32, b(15)=>
      gen_24_cmp_pInit_32, b(14)=>gen_24_cmp_pInit_32, b(13)=>
      gen_24_cmp_pInit_32, b(12)=>gen_24_cmp_pInit_32, b(11)=>
      gen_24_cmp_pInit_32, b(10)=>gen_24_cmp_pInit_32, b(9)=>
      gen_24_cmp_pInit_32, b(8)=>filter_8_7, b(7)=>filter_8_6, b(6)=>
      filter_8_5, b(5)=>filter_8_4, b(4)=>filter_8_3, b(3)=>filter_8_2, b(2)
      =>filter_8_1, b(1)=>filter_8_0, b(0)=>gen_24_cmp_pInit_32, sel=>
      nx11908, f(32)=>DANGLING(82), f(31)=>DANGLING(83), f(30)=>
      gen_8_cmp_pMux_30, f(29)=>gen_8_cmp_pMux_29, f(28)=>gen_8_cmp_pMux_28, 
      f(27)=>gen_8_cmp_pMux_27, f(26)=>gen_8_cmp_pMux_26, f(25)=>
      gen_8_cmp_pMux_25, f(24)=>gen_8_cmp_pMux_24, f(23)=>gen_8_cmp_pMux_23, 
      f(22)=>gen_8_cmp_pMux_22, f(21)=>gen_8_cmp_pMux_21, f(20)=>
      gen_8_cmp_pMux_20, f(19)=>gen_8_cmp_pMux_19, f(18)=>gen_8_cmp_pMux_18, 
      f(17)=>gen_8_cmp_pMux_17, f(16)=>gen_8_cmp_pMux_16, f(15)=>
      gen_8_cmp_pMux_15, f(14)=>gen_8_cmp_pMux_14, f(13)=>gen_8_cmp_pMux_13, 
      f(12)=>gen_8_cmp_pMux_12, f(11)=>gen_8_cmp_pMux_11, f(10)=>
      gen_8_cmp_pMux_10, f(9)=>gen_8_cmp_pMux_9, f(8)=>gen_8_cmp_pMux_8, 
      f(7)=>gen_8_cmp_pMux_7, f(6)=>gen_8_cmp_pMux_6, f(5)=>gen_8_cmp_pMux_5, 
      f(4)=>gen_8_cmp_pMux_4, f(3)=>gen_8_cmp_pMux_3, f(2)=>gen_8_cmp_pMux_2, 
      f(1)=>gen_8_cmp_pMux_1, f(0)=>gen_8_cmp_pMux_0);
   gen_8_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>
      gen_24_cmp_pInit_32, a(22)=>gen_24_cmp_pInit_32, a(21)=>
      gen_8_cmp_pMux_30, a(20)=>gen_8_cmp_pMux_29, a(19)=>gen_8_cmp_pMux_28, 
      a(18)=>gen_8_cmp_pMux_27, a(17)=>gen_8_cmp_pMux_26, a(16)=>
      gen_8_cmp_pMux_25, a(15)=>gen_8_cmp_pMux_24, a(14)=>gen_8_cmp_pMux_23, 
      a(13)=>gen_8_cmp_pMux_22, a(12)=>gen_8_cmp_pMux_21, a(11)=>
      gen_8_cmp_pMux_20, a(10)=>gen_8_cmp_pMux_19, a(9)=>gen_8_cmp_pMux_18, 
      a(8)=>gen_8_cmp_pMux_17, a(7)=>gen_8_cmp_pMux_16, a(6)=>
      gen_8_cmp_pMux_15, a(5)=>gen_8_cmp_pMux_14, a(4)=>gen_8_cmp_pMux_13, 
      a(3)=>gen_8_cmp_pMux_12, a(2)=>gen_8_cmp_pMux_11, a(1)=>
      gen_8_cmp_pMux_10, a(0)=>gen_8_cmp_pMux_9, b(23)=>nx10626, b(22)=>
      nx10626, b(21)=>nx10624, b(20)=>nx10632, b(19)=>nx10630, b(18)=>
      nx10628, b(17)=>nx10626, b(16)=>nx10624, b(15)=>gen_8_cmp_BSCmp_op2_15, 
      b(14)=>gen_8_cmp_BSCmp_op2_14, b(13)=>gen_8_cmp_BSCmp_op2_13, b(12)=>
      gen_8_cmp_BSCmp_op2_12, b(11)=>gen_8_cmp_BSCmp_op2_11, b(10)=>
      gen_8_cmp_BSCmp_op2_10, b(9)=>gen_8_cmp_BSCmp_op2_9, b(8)=>
      gen_8_cmp_BSCmp_op2_8, b(7)=>gen_8_cmp_BSCmp_op2_7, b(6)=>
      gen_8_cmp_BSCmp_op2_6, b(5)=>gen_8_cmp_BSCmp_op2_5, b(4)=>
      gen_8_cmp_BSCmp_op2_4, b(3)=>gen_8_cmp_BSCmp_op2_3, b(2)=>
      gen_8_cmp_BSCmp_op2_2, b(1)=>gen_8_cmp_BSCmp_op2_1, b(0)=>
      gen_8_cmp_BSCmp_op2_0, carryIn=>gen_8_cmp_BSCmp_carryIn, sum(23)=>
      gen_8_cmp_pBs_30, sum(22)=>gen_8_cmp_pBs_29, sum(21)=>gen_8_cmp_pBs_28, 
      sum(20)=>gen_8_cmp_pBs_27, sum(19)=>gen_8_cmp_pBs_26, sum(18)=>
      gen_8_cmp_pBs_25, sum(17)=>gen_8_cmp_pBs_24, sum(16)=>gen_8_cmp_pBs_23, 
      sum(15)=>outputs_8_15, sum(14)=>outputs_8_14, sum(13)=>outputs_8_13, 
      sum(12)=>outputs_8_12, sum(11)=>outputs_8_11, sum(10)=>outputs_8_10, 
      sum(9)=>outputs_8_9, sum(8)=>outputs_8_8, sum(7)=>outputs_8_7, sum(6)
      =>outputs_8_6, sum(5)=>outputs_8_5, sum(4)=>outputs_8_4, sum(3)=>
      outputs_8_3, sum(2)=>outputs_8_2, sum(1)=>outputs_8_1, sum(0)=>
      outputs_8_0, carryOut=>DANGLING(84));
   gen_7_cmp_pRegCmp : Reg_33 port map ( D(32)=>gen_24_cmp_pInit_32, D(31)=>
      gen_24_cmp_pInit_32, D(30)=>gen_7_cmp_pBs_30, D(29)=>gen_7_cmp_pBs_29, 
      D(28)=>gen_7_cmp_pBs_28, D(27)=>gen_7_cmp_pBs_27, D(26)=>
      gen_7_cmp_pBs_26, D(25)=>gen_7_cmp_pBs_25, D(24)=>gen_7_cmp_pBs_24, 
      D(23)=>gen_7_cmp_pBs_23, D(22)=>outputs_7_15, D(21)=>outputs_7_14, 
      D(20)=>outputs_7_13, D(19)=>outputs_7_12, D(18)=>outputs_7_11, D(17)=>
      outputs_7_10, D(16)=>outputs_7_9, D(15)=>outputs_7_8, D(14)=>
      outputs_7_7, D(13)=>outputs_7_6, D(12)=>outputs_7_5, D(11)=>
      outputs_7_4, D(10)=>outputs_7_3, D(9)=>outputs_7_2, D(8)=>outputs_7_1, 
      D(7)=>outputs_7_0, D(6)=>gen_7_cmp_pMux_8, D(5)=>gen_7_cmp_pMux_7, 
      D(4)=>gen_7_cmp_pMux_6, D(3)=>gen_7_cmp_pMux_5, D(2)=>gen_7_cmp_pMux_4, 
      D(1)=>gen_7_cmp_pMux_3, D(0)=>nx10334, en=>nx11926, clk=>nx10126, rst
      =>rst, Q(32)=>DANGLING(85), Q(31)=>DANGLING(86), Q(30)=>
      gen_7_cmp_pReg_30, Q(29)=>gen_7_cmp_pReg_29, Q(28)=>gen_7_cmp_pReg_28, 
      Q(27)=>gen_7_cmp_pReg_27, Q(26)=>gen_7_cmp_pReg_26, Q(25)=>
      gen_7_cmp_pReg_25, Q(24)=>gen_7_cmp_pReg_24, Q(23)=>gen_7_cmp_pReg_23, 
      Q(22)=>gen_7_cmp_pReg_22, Q(21)=>gen_7_cmp_pReg_21, Q(20)=>
      gen_7_cmp_pReg_20, Q(19)=>gen_7_cmp_pReg_19, Q(18)=>gen_7_cmp_pReg_18, 
      Q(17)=>gen_7_cmp_pReg_17, Q(16)=>gen_7_cmp_pReg_16, Q(15)=>
      gen_7_cmp_pReg_15, Q(14)=>gen_7_cmp_pReg_14, Q(13)=>gen_7_cmp_pReg_13, 
      Q(12)=>gen_7_cmp_pReg_12, Q(11)=>gen_7_cmp_pReg_11, Q(10)=>
      gen_7_cmp_pReg_10, Q(9)=>gen_7_cmp_pReg_9, Q(8)=>gen_7_cmp_pReg_8, 
      Q(7)=>gen_7_cmp_pReg_7, Q(6)=>gen_7_cmp_pReg_6, Q(5)=>gen_7_cmp_pReg_5, 
      Q(4)=>gen_7_cmp_pReg_4, Q(3)=>gen_7_cmp_pReg_3, Q(2)=>gen_7_cmp_pReg_2, 
      Q(1)=>gen_7_cmp_pReg_1, Q(0)=>gen_7_cmp_pReg_0);
   gen_7_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>gen_24_cmp_pInit_32, 
      a(31)=>gen_24_cmp_pInit_32, a(30)=>gen_7_cmp_pReg_30, a(29)=>
      gen_7_cmp_pReg_29, a(28)=>gen_7_cmp_pReg_28, a(27)=>gen_7_cmp_pReg_27, 
      a(26)=>gen_7_cmp_pReg_26, a(25)=>gen_7_cmp_pReg_25, a(24)=>
      gen_7_cmp_pReg_24, a(23)=>gen_7_cmp_pReg_23, a(22)=>gen_7_cmp_pReg_22, 
      a(21)=>gen_7_cmp_pReg_21, a(20)=>gen_7_cmp_pReg_20, a(19)=>
      gen_7_cmp_pReg_19, a(18)=>gen_7_cmp_pReg_18, a(17)=>gen_7_cmp_pReg_17, 
      a(16)=>gen_7_cmp_pReg_16, a(15)=>gen_7_cmp_pReg_15, a(14)=>
      gen_7_cmp_pReg_14, a(13)=>gen_7_cmp_pReg_13, a(12)=>gen_7_cmp_pReg_12, 
      a(11)=>gen_7_cmp_pReg_11, a(10)=>gen_7_cmp_pReg_10, a(9)=>
      gen_7_cmp_pReg_9, a(8)=>gen_7_cmp_pReg_8, a(7)=>gen_7_cmp_pReg_7, a(6)
      =>gen_7_cmp_pReg_6, a(5)=>gen_7_cmp_pReg_5, a(4)=>gen_7_cmp_pReg_4, 
      a(3)=>gen_7_cmp_pReg_3, a(2)=>gen_7_cmp_pReg_2, a(1)=>gen_7_cmp_pReg_1, 
      a(0)=>gen_7_cmp_pReg_0, b(32)=>gen_24_cmp_pInit_32, b(31)=>
      gen_24_cmp_pInit_32, b(30)=>gen_24_cmp_pInit_32, b(29)=>
      gen_24_cmp_pInit_32, b(28)=>gen_24_cmp_pInit_32, b(27)=>
      gen_24_cmp_pInit_32, b(26)=>gen_24_cmp_pInit_32, b(25)=>
      gen_24_cmp_pInit_32, b(24)=>gen_24_cmp_pInit_32, b(23)=>
      gen_24_cmp_pInit_32, b(22)=>gen_24_cmp_pInit_32, b(21)=>
      gen_24_cmp_pInit_32, b(20)=>gen_24_cmp_pInit_32, b(19)=>
      gen_24_cmp_pInit_32, b(18)=>gen_24_cmp_pInit_32, b(17)=>
      gen_24_cmp_pInit_32, b(16)=>gen_24_cmp_pInit_32, b(15)=>
      gen_24_cmp_pInit_32, b(14)=>gen_24_cmp_pInit_32, b(13)=>
      gen_24_cmp_pInit_32, b(12)=>gen_24_cmp_pInit_32, b(11)=>
      gen_24_cmp_pInit_32, b(10)=>gen_24_cmp_pInit_32, b(9)=>
      gen_24_cmp_pInit_32, b(8)=>filter_7_7, b(7)=>filter_7_6, b(6)=>
      filter_7_5, b(5)=>filter_7_4, b(4)=>filter_7_3, b(3)=>filter_7_2, b(2)
      =>filter_7_1, b(1)=>filter_7_0, b(0)=>gen_24_cmp_pInit_32, sel=>
      nx11910, f(32)=>DANGLING(87), f(31)=>DANGLING(88), f(30)=>
      gen_7_cmp_pMux_30, f(29)=>gen_7_cmp_pMux_29, f(28)=>gen_7_cmp_pMux_28, 
      f(27)=>gen_7_cmp_pMux_27, f(26)=>gen_7_cmp_pMux_26, f(25)=>
      gen_7_cmp_pMux_25, f(24)=>gen_7_cmp_pMux_24, f(23)=>gen_7_cmp_pMux_23, 
      f(22)=>gen_7_cmp_pMux_22, f(21)=>gen_7_cmp_pMux_21, f(20)=>
      gen_7_cmp_pMux_20, f(19)=>gen_7_cmp_pMux_19, f(18)=>gen_7_cmp_pMux_18, 
      f(17)=>gen_7_cmp_pMux_17, f(16)=>gen_7_cmp_pMux_16, f(15)=>
      gen_7_cmp_pMux_15, f(14)=>gen_7_cmp_pMux_14, f(13)=>gen_7_cmp_pMux_13, 
      f(12)=>gen_7_cmp_pMux_12, f(11)=>gen_7_cmp_pMux_11, f(10)=>
      gen_7_cmp_pMux_10, f(9)=>gen_7_cmp_pMux_9, f(8)=>gen_7_cmp_pMux_8, 
      f(7)=>gen_7_cmp_pMux_7, f(6)=>gen_7_cmp_pMux_6, f(5)=>gen_7_cmp_pMux_5, 
      f(4)=>gen_7_cmp_pMux_4, f(3)=>gen_7_cmp_pMux_3, f(2)=>gen_7_cmp_pMux_2, 
      f(1)=>gen_7_cmp_pMux_1, f(0)=>gen_7_cmp_pMux_0);
   gen_7_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>
      gen_24_cmp_pInit_32, a(22)=>gen_24_cmp_pInit_32, a(21)=>
      gen_7_cmp_pMux_30, a(20)=>gen_7_cmp_pMux_29, a(19)=>gen_7_cmp_pMux_28, 
      a(18)=>gen_7_cmp_pMux_27, a(17)=>gen_7_cmp_pMux_26, a(16)=>
      gen_7_cmp_pMux_25, a(15)=>gen_7_cmp_pMux_24, a(14)=>gen_7_cmp_pMux_23, 
      a(13)=>gen_7_cmp_pMux_22, a(12)=>gen_7_cmp_pMux_21, a(11)=>
      gen_7_cmp_pMux_20, a(10)=>gen_7_cmp_pMux_19, a(9)=>gen_7_cmp_pMux_18, 
      a(8)=>gen_7_cmp_pMux_17, a(7)=>gen_7_cmp_pMux_16, a(6)=>
      gen_7_cmp_pMux_15, a(5)=>gen_7_cmp_pMux_14, a(4)=>gen_7_cmp_pMux_13, 
      a(3)=>gen_7_cmp_pMux_12, a(2)=>gen_7_cmp_pMux_11, a(1)=>
      gen_7_cmp_pMux_10, a(0)=>gen_7_cmp_pMux_9, b(23)=>nx10638, b(22)=>
      nx10638, b(21)=>nx10636, b(20)=>nx10644, b(19)=>nx10642, b(18)=>
      nx10640, b(17)=>nx10638, b(16)=>nx10636, b(15)=>gen_7_cmp_BSCmp_op2_15, 
      b(14)=>gen_7_cmp_BSCmp_op2_14, b(13)=>gen_7_cmp_BSCmp_op2_13, b(12)=>
      gen_7_cmp_BSCmp_op2_12, b(11)=>gen_7_cmp_BSCmp_op2_11, b(10)=>
      gen_7_cmp_BSCmp_op2_10, b(9)=>gen_7_cmp_BSCmp_op2_9, b(8)=>
      gen_7_cmp_BSCmp_op2_8, b(7)=>gen_7_cmp_BSCmp_op2_7, b(6)=>
      gen_7_cmp_BSCmp_op2_6, b(5)=>gen_7_cmp_BSCmp_op2_5, b(4)=>
      gen_7_cmp_BSCmp_op2_4, b(3)=>gen_7_cmp_BSCmp_op2_3, b(2)=>
      gen_7_cmp_BSCmp_op2_2, b(1)=>gen_7_cmp_BSCmp_op2_1, b(0)=>
      gen_7_cmp_BSCmp_op2_0, carryIn=>gen_7_cmp_BSCmp_carryIn, sum(23)=>
      gen_7_cmp_pBs_30, sum(22)=>gen_7_cmp_pBs_29, sum(21)=>gen_7_cmp_pBs_28, 
      sum(20)=>gen_7_cmp_pBs_27, sum(19)=>gen_7_cmp_pBs_26, sum(18)=>
      gen_7_cmp_pBs_25, sum(17)=>gen_7_cmp_pBs_24, sum(16)=>gen_7_cmp_pBs_23, 
      sum(15)=>outputs_7_15, sum(14)=>outputs_7_14, sum(13)=>outputs_7_13, 
      sum(12)=>outputs_7_12, sum(11)=>outputs_7_11, sum(10)=>outputs_7_10, 
      sum(9)=>outputs_7_9, sum(8)=>outputs_7_8, sum(7)=>outputs_7_7, sum(6)
      =>outputs_7_6, sum(5)=>outputs_7_5, sum(4)=>outputs_7_4, sum(3)=>
      outputs_7_3, sum(2)=>outputs_7_2, sum(1)=>outputs_7_1, sum(0)=>
      outputs_7_0, carryOut=>DANGLING(89));
   gen_6_cmp_pRegCmp : Reg_33 port map ( D(32)=>gen_24_cmp_pInit_32, D(31)=>
      gen_24_cmp_pInit_32, D(30)=>gen_6_cmp_pBs_30, D(29)=>gen_6_cmp_pBs_29, 
      D(28)=>gen_6_cmp_pBs_28, D(27)=>gen_6_cmp_pBs_27, D(26)=>
      gen_6_cmp_pBs_26, D(25)=>gen_6_cmp_pBs_25, D(24)=>gen_6_cmp_pBs_24, 
      D(23)=>gen_6_cmp_pBs_23, D(22)=>outputs_6_15, D(21)=>outputs_6_14, 
      D(20)=>outputs_6_13, D(19)=>outputs_6_12, D(18)=>outputs_6_11, D(17)=>
      outputs_6_10, D(16)=>outputs_6_9, D(15)=>outputs_6_8, D(14)=>
      outputs_6_7, D(13)=>outputs_6_6, D(12)=>outputs_6_5, D(11)=>
      outputs_6_4, D(10)=>outputs_6_3, D(9)=>outputs_6_2, D(8)=>outputs_6_1, 
      D(7)=>outputs_6_0, D(6)=>gen_6_cmp_pMux_8, D(5)=>gen_6_cmp_pMux_7, 
      D(4)=>gen_6_cmp_pMux_6, D(3)=>gen_6_cmp_pMux_5, D(2)=>gen_6_cmp_pMux_4, 
      D(1)=>gen_6_cmp_pMux_3, D(0)=>nx10346, en=>nx11926, clk=>nx10126, rst
      =>rst, Q(32)=>DANGLING(90), Q(31)=>DANGLING(91), Q(30)=>
      gen_6_cmp_pReg_30, Q(29)=>gen_6_cmp_pReg_29, Q(28)=>gen_6_cmp_pReg_28, 
      Q(27)=>gen_6_cmp_pReg_27, Q(26)=>gen_6_cmp_pReg_26, Q(25)=>
      gen_6_cmp_pReg_25, Q(24)=>gen_6_cmp_pReg_24, Q(23)=>gen_6_cmp_pReg_23, 
      Q(22)=>gen_6_cmp_pReg_22, Q(21)=>gen_6_cmp_pReg_21, Q(20)=>
      gen_6_cmp_pReg_20, Q(19)=>gen_6_cmp_pReg_19, Q(18)=>gen_6_cmp_pReg_18, 
      Q(17)=>gen_6_cmp_pReg_17, Q(16)=>gen_6_cmp_pReg_16, Q(15)=>
      gen_6_cmp_pReg_15, Q(14)=>gen_6_cmp_pReg_14, Q(13)=>gen_6_cmp_pReg_13, 
      Q(12)=>gen_6_cmp_pReg_12, Q(11)=>gen_6_cmp_pReg_11, Q(10)=>
      gen_6_cmp_pReg_10, Q(9)=>gen_6_cmp_pReg_9, Q(8)=>gen_6_cmp_pReg_8, 
      Q(7)=>gen_6_cmp_pReg_7, Q(6)=>gen_6_cmp_pReg_6, Q(5)=>gen_6_cmp_pReg_5, 
      Q(4)=>gen_6_cmp_pReg_4, Q(3)=>gen_6_cmp_pReg_3, Q(2)=>gen_6_cmp_pReg_2, 
      Q(1)=>gen_6_cmp_pReg_1, Q(0)=>gen_6_cmp_pReg_0);
   gen_6_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>gen_24_cmp_pInit_32, 
      a(31)=>gen_24_cmp_pInit_32, a(30)=>gen_6_cmp_pReg_30, a(29)=>
      gen_6_cmp_pReg_29, a(28)=>gen_6_cmp_pReg_28, a(27)=>gen_6_cmp_pReg_27, 
      a(26)=>gen_6_cmp_pReg_26, a(25)=>gen_6_cmp_pReg_25, a(24)=>
      gen_6_cmp_pReg_24, a(23)=>gen_6_cmp_pReg_23, a(22)=>gen_6_cmp_pReg_22, 
      a(21)=>gen_6_cmp_pReg_21, a(20)=>gen_6_cmp_pReg_20, a(19)=>
      gen_6_cmp_pReg_19, a(18)=>gen_6_cmp_pReg_18, a(17)=>gen_6_cmp_pReg_17, 
      a(16)=>gen_6_cmp_pReg_16, a(15)=>gen_6_cmp_pReg_15, a(14)=>
      gen_6_cmp_pReg_14, a(13)=>gen_6_cmp_pReg_13, a(12)=>gen_6_cmp_pReg_12, 
      a(11)=>gen_6_cmp_pReg_11, a(10)=>gen_6_cmp_pReg_10, a(9)=>
      gen_6_cmp_pReg_9, a(8)=>gen_6_cmp_pReg_8, a(7)=>gen_6_cmp_pReg_7, a(6)
      =>gen_6_cmp_pReg_6, a(5)=>gen_6_cmp_pReg_5, a(4)=>gen_6_cmp_pReg_4, 
      a(3)=>gen_6_cmp_pReg_3, a(2)=>gen_6_cmp_pReg_2, a(1)=>gen_6_cmp_pReg_1, 
      a(0)=>gen_6_cmp_pReg_0, b(32)=>gen_24_cmp_pInit_32, b(31)=>
      gen_24_cmp_pInit_32, b(30)=>gen_24_cmp_pInit_32, b(29)=>
      gen_24_cmp_pInit_32, b(28)=>gen_24_cmp_pInit_32, b(27)=>
      gen_24_cmp_pInit_32, b(26)=>gen_24_cmp_pInit_32, b(25)=>
      gen_24_cmp_pInit_32, b(24)=>gen_24_cmp_pInit_32, b(23)=>
      gen_24_cmp_pInit_32, b(22)=>gen_24_cmp_pInit_32, b(21)=>
      gen_24_cmp_pInit_32, b(20)=>gen_24_cmp_pInit_32, b(19)=>
      gen_24_cmp_pInit_32, b(18)=>gen_24_cmp_pInit_32, b(17)=>
      gen_24_cmp_pInit_32, b(16)=>gen_24_cmp_pInit_32, b(15)=>
      gen_24_cmp_pInit_32, b(14)=>gen_24_cmp_pInit_32, b(13)=>
      gen_24_cmp_pInit_32, b(12)=>gen_24_cmp_pInit_32, b(11)=>
      gen_24_cmp_pInit_32, b(10)=>gen_24_cmp_pInit_32, b(9)=>
      gen_24_cmp_pInit_32, b(8)=>filter_6_7, b(7)=>filter_6_6, b(6)=>
      filter_6_5, b(5)=>filter_6_4, b(4)=>filter_6_3, b(3)=>filter_6_2, b(2)
      =>filter_6_1, b(1)=>filter_6_0, b(0)=>gen_24_cmp_pInit_32, sel=>
      nx11910, f(32)=>DANGLING(92), f(31)=>DANGLING(93), f(30)=>
      gen_6_cmp_pMux_30, f(29)=>gen_6_cmp_pMux_29, f(28)=>gen_6_cmp_pMux_28, 
      f(27)=>gen_6_cmp_pMux_27, f(26)=>gen_6_cmp_pMux_26, f(25)=>
      gen_6_cmp_pMux_25, f(24)=>gen_6_cmp_pMux_24, f(23)=>gen_6_cmp_pMux_23, 
      f(22)=>gen_6_cmp_pMux_22, f(21)=>gen_6_cmp_pMux_21, f(20)=>
      gen_6_cmp_pMux_20, f(19)=>gen_6_cmp_pMux_19, f(18)=>gen_6_cmp_pMux_18, 
      f(17)=>gen_6_cmp_pMux_17, f(16)=>gen_6_cmp_pMux_16, f(15)=>
      gen_6_cmp_pMux_15, f(14)=>gen_6_cmp_pMux_14, f(13)=>gen_6_cmp_pMux_13, 
      f(12)=>gen_6_cmp_pMux_12, f(11)=>gen_6_cmp_pMux_11, f(10)=>
      gen_6_cmp_pMux_10, f(9)=>gen_6_cmp_pMux_9, f(8)=>gen_6_cmp_pMux_8, 
      f(7)=>gen_6_cmp_pMux_7, f(6)=>gen_6_cmp_pMux_6, f(5)=>gen_6_cmp_pMux_5, 
      f(4)=>gen_6_cmp_pMux_4, f(3)=>gen_6_cmp_pMux_3, f(2)=>gen_6_cmp_pMux_2, 
      f(1)=>gen_6_cmp_pMux_1, f(0)=>gen_6_cmp_pMux_0);
   gen_6_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>
      gen_24_cmp_pInit_32, a(22)=>gen_24_cmp_pInit_32, a(21)=>
      gen_6_cmp_pMux_30, a(20)=>gen_6_cmp_pMux_29, a(19)=>gen_6_cmp_pMux_28, 
      a(18)=>gen_6_cmp_pMux_27, a(17)=>gen_6_cmp_pMux_26, a(16)=>
      gen_6_cmp_pMux_25, a(15)=>gen_6_cmp_pMux_24, a(14)=>gen_6_cmp_pMux_23, 
      a(13)=>gen_6_cmp_pMux_22, a(12)=>gen_6_cmp_pMux_21, a(11)=>
      gen_6_cmp_pMux_20, a(10)=>gen_6_cmp_pMux_19, a(9)=>gen_6_cmp_pMux_18, 
      a(8)=>gen_6_cmp_pMux_17, a(7)=>gen_6_cmp_pMux_16, a(6)=>
      gen_6_cmp_pMux_15, a(5)=>gen_6_cmp_pMux_14, a(4)=>gen_6_cmp_pMux_13, 
      a(3)=>gen_6_cmp_pMux_12, a(2)=>gen_6_cmp_pMux_11, a(1)=>
      gen_6_cmp_pMux_10, a(0)=>gen_6_cmp_pMux_9, b(23)=>nx10650, b(22)=>
      nx10650, b(21)=>nx10648, b(20)=>nx10656, b(19)=>nx10654, b(18)=>
      nx10652, b(17)=>nx10650, b(16)=>nx10648, b(15)=>gen_6_cmp_BSCmp_op2_15, 
      b(14)=>gen_6_cmp_BSCmp_op2_14, b(13)=>gen_6_cmp_BSCmp_op2_13, b(12)=>
      gen_6_cmp_BSCmp_op2_12, b(11)=>gen_6_cmp_BSCmp_op2_11, b(10)=>
      gen_6_cmp_BSCmp_op2_10, b(9)=>gen_6_cmp_BSCmp_op2_9, b(8)=>
      gen_6_cmp_BSCmp_op2_8, b(7)=>gen_6_cmp_BSCmp_op2_7, b(6)=>
      gen_6_cmp_BSCmp_op2_6, b(5)=>gen_6_cmp_BSCmp_op2_5, b(4)=>
      gen_6_cmp_BSCmp_op2_4, b(3)=>gen_6_cmp_BSCmp_op2_3, b(2)=>
      gen_6_cmp_BSCmp_op2_2, b(1)=>gen_6_cmp_BSCmp_op2_1, b(0)=>
      gen_6_cmp_BSCmp_op2_0, carryIn=>gen_6_cmp_BSCmp_carryIn, sum(23)=>
      gen_6_cmp_pBs_30, sum(22)=>gen_6_cmp_pBs_29, sum(21)=>gen_6_cmp_pBs_28, 
      sum(20)=>gen_6_cmp_pBs_27, sum(19)=>gen_6_cmp_pBs_26, sum(18)=>
      gen_6_cmp_pBs_25, sum(17)=>gen_6_cmp_pBs_24, sum(16)=>gen_6_cmp_pBs_23, 
      sum(15)=>outputs_6_15, sum(14)=>outputs_6_14, sum(13)=>outputs_6_13, 
      sum(12)=>outputs_6_12, sum(11)=>outputs_6_11, sum(10)=>outputs_6_10, 
      sum(9)=>outputs_6_9, sum(8)=>outputs_6_8, sum(7)=>outputs_6_7, sum(6)
      =>outputs_6_6, sum(5)=>outputs_6_5, sum(4)=>outputs_6_4, sum(3)=>
      outputs_6_3, sum(2)=>outputs_6_2, sum(1)=>outputs_6_1, sum(0)=>
      outputs_6_0, carryOut=>DANGLING(94));
   gen_5_cmp_pRegCmp : Reg_33 port map ( D(32)=>gen_24_cmp_pInit_32, D(31)=>
      gen_24_cmp_pInit_32, D(30)=>gen_5_cmp_pBs_30, D(29)=>gen_5_cmp_pBs_29, 
      D(28)=>gen_5_cmp_pBs_28, D(27)=>gen_5_cmp_pBs_27, D(26)=>
      gen_5_cmp_pBs_26, D(25)=>gen_5_cmp_pBs_25, D(24)=>gen_5_cmp_pBs_24, 
      D(23)=>gen_5_cmp_pBs_23, D(22)=>outputs_5_15, D(21)=>outputs_5_14, 
      D(20)=>outputs_5_13, D(19)=>outputs_5_12, D(18)=>outputs_5_11, D(17)=>
      outputs_5_10, D(16)=>outputs_5_9, D(15)=>outputs_5_8, D(14)=>
      outputs_5_7, D(13)=>outputs_5_6, D(12)=>outputs_5_5, D(11)=>
      outputs_5_4, D(10)=>outputs_5_3, D(9)=>outputs_5_2, D(8)=>outputs_5_1, 
      D(7)=>outputs_5_0, D(6)=>gen_5_cmp_pMux_8, D(5)=>gen_5_cmp_pMux_7, 
      D(4)=>gen_5_cmp_pMux_6, D(3)=>gen_5_cmp_pMux_5, D(2)=>gen_5_cmp_pMux_4, 
      D(1)=>gen_5_cmp_pMux_3, D(0)=>nx10358, en=>nx11926, clk=>nx10126, rst
      =>rst, Q(32)=>DANGLING(95), Q(31)=>DANGLING(96), Q(30)=>
      gen_5_cmp_pReg_30, Q(29)=>gen_5_cmp_pReg_29, Q(28)=>gen_5_cmp_pReg_28, 
      Q(27)=>gen_5_cmp_pReg_27, Q(26)=>gen_5_cmp_pReg_26, Q(25)=>
      gen_5_cmp_pReg_25, Q(24)=>gen_5_cmp_pReg_24, Q(23)=>gen_5_cmp_pReg_23, 
      Q(22)=>gen_5_cmp_pReg_22, Q(21)=>gen_5_cmp_pReg_21, Q(20)=>
      gen_5_cmp_pReg_20, Q(19)=>gen_5_cmp_pReg_19, Q(18)=>gen_5_cmp_pReg_18, 
      Q(17)=>gen_5_cmp_pReg_17, Q(16)=>gen_5_cmp_pReg_16, Q(15)=>
      gen_5_cmp_pReg_15, Q(14)=>gen_5_cmp_pReg_14, Q(13)=>gen_5_cmp_pReg_13, 
      Q(12)=>gen_5_cmp_pReg_12, Q(11)=>gen_5_cmp_pReg_11, Q(10)=>
      gen_5_cmp_pReg_10, Q(9)=>gen_5_cmp_pReg_9, Q(8)=>gen_5_cmp_pReg_8, 
      Q(7)=>gen_5_cmp_pReg_7, Q(6)=>gen_5_cmp_pReg_6, Q(5)=>gen_5_cmp_pReg_5, 
      Q(4)=>gen_5_cmp_pReg_4, Q(3)=>gen_5_cmp_pReg_3, Q(2)=>gen_5_cmp_pReg_2, 
      Q(1)=>gen_5_cmp_pReg_1, Q(0)=>gen_5_cmp_pReg_0);
   gen_5_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>gen_24_cmp_pInit_32, 
      a(31)=>gen_24_cmp_pInit_32, a(30)=>gen_5_cmp_pReg_30, a(29)=>
      gen_5_cmp_pReg_29, a(28)=>gen_5_cmp_pReg_28, a(27)=>gen_5_cmp_pReg_27, 
      a(26)=>gen_5_cmp_pReg_26, a(25)=>gen_5_cmp_pReg_25, a(24)=>
      gen_5_cmp_pReg_24, a(23)=>gen_5_cmp_pReg_23, a(22)=>gen_5_cmp_pReg_22, 
      a(21)=>gen_5_cmp_pReg_21, a(20)=>gen_5_cmp_pReg_20, a(19)=>
      gen_5_cmp_pReg_19, a(18)=>gen_5_cmp_pReg_18, a(17)=>gen_5_cmp_pReg_17, 
      a(16)=>gen_5_cmp_pReg_16, a(15)=>gen_5_cmp_pReg_15, a(14)=>
      gen_5_cmp_pReg_14, a(13)=>gen_5_cmp_pReg_13, a(12)=>gen_5_cmp_pReg_12, 
      a(11)=>gen_5_cmp_pReg_11, a(10)=>gen_5_cmp_pReg_10, a(9)=>
      gen_5_cmp_pReg_9, a(8)=>gen_5_cmp_pReg_8, a(7)=>gen_5_cmp_pReg_7, a(6)
      =>gen_5_cmp_pReg_6, a(5)=>gen_5_cmp_pReg_5, a(4)=>gen_5_cmp_pReg_4, 
      a(3)=>gen_5_cmp_pReg_3, a(2)=>gen_5_cmp_pReg_2, a(1)=>gen_5_cmp_pReg_1, 
      a(0)=>gen_5_cmp_pReg_0, b(32)=>gen_24_cmp_pInit_32, b(31)=>
      gen_24_cmp_pInit_32, b(30)=>gen_24_cmp_pInit_32, b(29)=>
      gen_24_cmp_pInit_32, b(28)=>gen_24_cmp_pInit_32, b(27)=>
      gen_24_cmp_pInit_32, b(26)=>gen_24_cmp_pInit_32, b(25)=>
      gen_24_cmp_pInit_32, b(24)=>gen_24_cmp_pInit_32, b(23)=>
      gen_24_cmp_pInit_32, b(22)=>gen_24_cmp_pInit_32, b(21)=>
      gen_24_cmp_pInit_32, b(20)=>gen_24_cmp_pInit_32, b(19)=>
      gen_24_cmp_pInit_32, b(18)=>gen_24_cmp_pInit_32, b(17)=>
      gen_24_cmp_pInit_32, b(16)=>gen_24_cmp_pInit_32, b(15)=>
      gen_24_cmp_pInit_32, b(14)=>gen_24_cmp_pInit_32, b(13)=>
      gen_24_cmp_pInit_32, b(12)=>gen_24_cmp_pInit_32, b(11)=>
      gen_24_cmp_pInit_32, b(10)=>gen_24_cmp_pInit_32, b(9)=>
      gen_24_cmp_pInit_32, b(8)=>filter_5_7, b(7)=>filter_5_6, b(6)=>
      filter_5_5, b(5)=>filter_5_4, b(4)=>filter_5_3, b(3)=>filter_5_2, b(2)
      =>filter_5_1, b(1)=>filter_5_0, b(0)=>gen_24_cmp_pInit_32, sel=>
      nx11910, f(32)=>DANGLING(97), f(31)=>DANGLING(98), f(30)=>
      gen_5_cmp_pMux_30, f(29)=>gen_5_cmp_pMux_29, f(28)=>gen_5_cmp_pMux_28, 
      f(27)=>gen_5_cmp_pMux_27, f(26)=>gen_5_cmp_pMux_26, f(25)=>
      gen_5_cmp_pMux_25, f(24)=>gen_5_cmp_pMux_24, f(23)=>gen_5_cmp_pMux_23, 
      f(22)=>gen_5_cmp_pMux_22, f(21)=>gen_5_cmp_pMux_21, f(20)=>
      gen_5_cmp_pMux_20, f(19)=>gen_5_cmp_pMux_19, f(18)=>gen_5_cmp_pMux_18, 
      f(17)=>gen_5_cmp_pMux_17, f(16)=>gen_5_cmp_pMux_16, f(15)=>
      gen_5_cmp_pMux_15, f(14)=>gen_5_cmp_pMux_14, f(13)=>gen_5_cmp_pMux_13, 
      f(12)=>gen_5_cmp_pMux_12, f(11)=>gen_5_cmp_pMux_11, f(10)=>
      gen_5_cmp_pMux_10, f(9)=>gen_5_cmp_pMux_9, f(8)=>gen_5_cmp_pMux_8, 
      f(7)=>gen_5_cmp_pMux_7, f(6)=>gen_5_cmp_pMux_6, f(5)=>gen_5_cmp_pMux_5, 
      f(4)=>gen_5_cmp_pMux_4, f(3)=>gen_5_cmp_pMux_3, f(2)=>gen_5_cmp_pMux_2, 
      f(1)=>gen_5_cmp_pMux_1, f(0)=>gen_5_cmp_pMux_0);
   gen_5_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>
      gen_24_cmp_pInit_32, a(22)=>gen_24_cmp_pInit_32, a(21)=>
      gen_5_cmp_pMux_30, a(20)=>gen_5_cmp_pMux_29, a(19)=>gen_5_cmp_pMux_28, 
      a(18)=>gen_5_cmp_pMux_27, a(17)=>gen_5_cmp_pMux_26, a(16)=>
      gen_5_cmp_pMux_25, a(15)=>gen_5_cmp_pMux_24, a(14)=>gen_5_cmp_pMux_23, 
      a(13)=>gen_5_cmp_pMux_22, a(12)=>gen_5_cmp_pMux_21, a(11)=>
      gen_5_cmp_pMux_20, a(10)=>gen_5_cmp_pMux_19, a(9)=>gen_5_cmp_pMux_18, 
      a(8)=>gen_5_cmp_pMux_17, a(7)=>gen_5_cmp_pMux_16, a(6)=>
      gen_5_cmp_pMux_15, a(5)=>gen_5_cmp_pMux_14, a(4)=>gen_5_cmp_pMux_13, 
      a(3)=>gen_5_cmp_pMux_12, a(2)=>gen_5_cmp_pMux_11, a(1)=>
      gen_5_cmp_pMux_10, a(0)=>gen_5_cmp_pMux_9, b(23)=>nx10662, b(22)=>
      nx10662, b(21)=>nx10660, b(20)=>nx10668, b(19)=>nx10666, b(18)=>
      nx10664, b(17)=>nx10662, b(16)=>nx10660, b(15)=>gen_5_cmp_BSCmp_op2_15, 
      b(14)=>gen_5_cmp_BSCmp_op2_14, b(13)=>gen_5_cmp_BSCmp_op2_13, b(12)=>
      gen_5_cmp_BSCmp_op2_12, b(11)=>gen_5_cmp_BSCmp_op2_11, b(10)=>
      gen_5_cmp_BSCmp_op2_10, b(9)=>gen_5_cmp_BSCmp_op2_9, b(8)=>
      gen_5_cmp_BSCmp_op2_8, b(7)=>gen_5_cmp_BSCmp_op2_7, b(6)=>
      gen_5_cmp_BSCmp_op2_6, b(5)=>gen_5_cmp_BSCmp_op2_5, b(4)=>
      gen_5_cmp_BSCmp_op2_4, b(3)=>gen_5_cmp_BSCmp_op2_3, b(2)=>
      gen_5_cmp_BSCmp_op2_2, b(1)=>gen_5_cmp_BSCmp_op2_1, b(0)=>
      gen_5_cmp_BSCmp_op2_0, carryIn=>gen_5_cmp_BSCmp_carryIn, sum(23)=>
      gen_5_cmp_pBs_30, sum(22)=>gen_5_cmp_pBs_29, sum(21)=>gen_5_cmp_pBs_28, 
      sum(20)=>gen_5_cmp_pBs_27, sum(19)=>gen_5_cmp_pBs_26, sum(18)=>
      gen_5_cmp_pBs_25, sum(17)=>gen_5_cmp_pBs_24, sum(16)=>gen_5_cmp_pBs_23, 
      sum(15)=>outputs_5_15, sum(14)=>outputs_5_14, sum(13)=>outputs_5_13, 
      sum(12)=>outputs_5_12, sum(11)=>outputs_5_11, sum(10)=>outputs_5_10, 
      sum(9)=>outputs_5_9, sum(8)=>outputs_5_8, sum(7)=>outputs_5_7, sum(6)
      =>outputs_5_6, sum(5)=>outputs_5_5, sum(4)=>outputs_5_4, sum(3)=>
      outputs_5_3, sum(2)=>outputs_5_2, sum(1)=>outputs_5_1, sum(0)=>
      outputs_5_0, carryOut=>DANGLING(99));
   gen_4_cmp_pRegCmp : Reg_33 port map ( D(32)=>gen_24_cmp_pInit_32, D(31)=>
      gen_24_cmp_pInit_32, D(30)=>gen_4_cmp_pBs_30, D(29)=>gen_4_cmp_pBs_29, 
      D(28)=>gen_4_cmp_pBs_28, D(27)=>gen_4_cmp_pBs_27, D(26)=>
      gen_4_cmp_pBs_26, D(25)=>gen_4_cmp_pBs_25, D(24)=>gen_4_cmp_pBs_24, 
      D(23)=>gen_4_cmp_pBs_23, D(22)=>outputs_4_15, D(21)=>outputs_4_14, 
      D(20)=>outputs_4_13, D(19)=>outputs_4_12, D(18)=>outputs_4_11, D(17)=>
      outputs_4_10, D(16)=>outputs_4_9, D(15)=>outputs_4_8, D(14)=>
      outputs_4_7, D(13)=>outputs_4_6, D(12)=>outputs_4_5, D(11)=>
      outputs_4_4, D(10)=>outputs_4_3, D(9)=>outputs_4_2, D(8)=>outputs_4_1, 
      D(7)=>outputs_4_0, D(6)=>gen_4_cmp_pMux_8, D(5)=>gen_4_cmp_pMux_7, 
      D(4)=>gen_4_cmp_pMux_6, D(3)=>gen_4_cmp_pMux_5, D(2)=>gen_4_cmp_pMux_4, 
      D(1)=>gen_4_cmp_pMux_3, D(0)=>nx10370, en=>nx10884, clk=>nx10126, rst
      =>rst, Q(32)=>DANGLING(100), Q(31)=>DANGLING(101), Q(30)=>
      gen_4_cmp_pReg_30, Q(29)=>gen_4_cmp_pReg_29, Q(28)=>gen_4_cmp_pReg_28, 
      Q(27)=>gen_4_cmp_pReg_27, Q(26)=>gen_4_cmp_pReg_26, Q(25)=>
      gen_4_cmp_pReg_25, Q(24)=>gen_4_cmp_pReg_24, Q(23)=>gen_4_cmp_pReg_23, 
      Q(22)=>gen_4_cmp_pReg_22, Q(21)=>gen_4_cmp_pReg_21, Q(20)=>
      gen_4_cmp_pReg_20, Q(19)=>gen_4_cmp_pReg_19, Q(18)=>gen_4_cmp_pReg_18, 
      Q(17)=>gen_4_cmp_pReg_17, Q(16)=>gen_4_cmp_pReg_16, Q(15)=>
      gen_4_cmp_pReg_15, Q(14)=>gen_4_cmp_pReg_14, Q(13)=>gen_4_cmp_pReg_13, 
      Q(12)=>gen_4_cmp_pReg_12, Q(11)=>gen_4_cmp_pReg_11, Q(10)=>
      gen_4_cmp_pReg_10, Q(9)=>gen_4_cmp_pReg_9, Q(8)=>gen_4_cmp_pReg_8, 
      Q(7)=>gen_4_cmp_pReg_7, Q(6)=>gen_4_cmp_pReg_6, Q(5)=>gen_4_cmp_pReg_5, 
      Q(4)=>gen_4_cmp_pReg_4, Q(3)=>gen_4_cmp_pReg_3, Q(2)=>gen_4_cmp_pReg_2, 
      Q(1)=>gen_4_cmp_pReg_1, Q(0)=>gen_4_cmp_pReg_0);
   gen_4_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>gen_24_cmp_pInit_32, 
      a(31)=>gen_24_cmp_pInit_32, a(30)=>gen_4_cmp_pReg_30, a(29)=>
      gen_4_cmp_pReg_29, a(28)=>gen_4_cmp_pReg_28, a(27)=>gen_4_cmp_pReg_27, 
      a(26)=>gen_4_cmp_pReg_26, a(25)=>gen_4_cmp_pReg_25, a(24)=>
      gen_4_cmp_pReg_24, a(23)=>gen_4_cmp_pReg_23, a(22)=>gen_4_cmp_pReg_22, 
      a(21)=>gen_4_cmp_pReg_21, a(20)=>gen_4_cmp_pReg_20, a(19)=>
      gen_4_cmp_pReg_19, a(18)=>gen_4_cmp_pReg_18, a(17)=>gen_4_cmp_pReg_17, 
      a(16)=>gen_4_cmp_pReg_16, a(15)=>gen_4_cmp_pReg_15, a(14)=>
      gen_4_cmp_pReg_14, a(13)=>gen_4_cmp_pReg_13, a(12)=>gen_4_cmp_pReg_12, 
      a(11)=>gen_4_cmp_pReg_11, a(10)=>gen_4_cmp_pReg_10, a(9)=>
      gen_4_cmp_pReg_9, a(8)=>gen_4_cmp_pReg_8, a(7)=>gen_4_cmp_pReg_7, a(6)
      =>gen_4_cmp_pReg_6, a(5)=>gen_4_cmp_pReg_5, a(4)=>gen_4_cmp_pReg_4, 
      a(3)=>gen_4_cmp_pReg_3, a(2)=>gen_4_cmp_pReg_2, a(1)=>gen_4_cmp_pReg_1, 
      a(0)=>gen_4_cmp_pReg_0, b(32)=>gen_24_cmp_pInit_32, b(31)=>
      gen_24_cmp_pInit_32, b(30)=>gen_24_cmp_pInit_32, b(29)=>
      gen_24_cmp_pInit_32, b(28)=>gen_24_cmp_pInit_32, b(27)=>
      gen_24_cmp_pInit_32, b(26)=>gen_24_cmp_pInit_32, b(25)=>
      gen_24_cmp_pInit_32, b(24)=>gen_24_cmp_pInit_32, b(23)=>
      gen_24_cmp_pInit_32, b(22)=>gen_24_cmp_pInit_32, b(21)=>
      gen_24_cmp_pInit_32, b(20)=>gen_24_cmp_pInit_32, b(19)=>
      gen_24_cmp_pInit_32, b(18)=>gen_24_cmp_pInit_32, b(17)=>
      gen_24_cmp_pInit_32, b(16)=>gen_24_cmp_pInit_32, b(15)=>
      gen_24_cmp_pInit_32, b(14)=>gen_24_cmp_pInit_32, b(13)=>
      gen_24_cmp_pInit_32, b(12)=>gen_24_cmp_pInit_32, b(11)=>
      gen_24_cmp_pInit_32, b(10)=>gen_24_cmp_pInit_32, b(9)=>
      gen_24_cmp_pInit_32, b(8)=>filter_4_7, b(7)=>filter_4_6, b(6)=>
      filter_4_5, b(5)=>filter_4_4, b(4)=>filter_4_3, b(3)=>filter_4_2, b(2)
      =>filter_4_1, b(1)=>filter_4_0, b(0)=>gen_24_cmp_pInit_32, sel=>
      nx11912, f(32)=>DANGLING(102), f(31)=>DANGLING(103), f(30)=>
      gen_4_cmp_pMux_30, f(29)=>gen_4_cmp_pMux_29, f(28)=>gen_4_cmp_pMux_28, 
      f(27)=>gen_4_cmp_pMux_27, f(26)=>gen_4_cmp_pMux_26, f(25)=>
      gen_4_cmp_pMux_25, f(24)=>gen_4_cmp_pMux_24, f(23)=>gen_4_cmp_pMux_23, 
      f(22)=>gen_4_cmp_pMux_22, f(21)=>gen_4_cmp_pMux_21, f(20)=>
      gen_4_cmp_pMux_20, f(19)=>gen_4_cmp_pMux_19, f(18)=>gen_4_cmp_pMux_18, 
      f(17)=>gen_4_cmp_pMux_17, f(16)=>gen_4_cmp_pMux_16, f(15)=>
      gen_4_cmp_pMux_15, f(14)=>gen_4_cmp_pMux_14, f(13)=>gen_4_cmp_pMux_13, 
      f(12)=>gen_4_cmp_pMux_12, f(11)=>gen_4_cmp_pMux_11, f(10)=>
      gen_4_cmp_pMux_10, f(9)=>gen_4_cmp_pMux_9, f(8)=>gen_4_cmp_pMux_8, 
      f(7)=>gen_4_cmp_pMux_7, f(6)=>gen_4_cmp_pMux_6, f(5)=>gen_4_cmp_pMux_5, 
      f(4)=>gen_4_cmp_pMux_4, f(3)=>gen_4_cmp_pMux_3, f(2)=>gen_4_cmp_pMux_2, 
      f(1)=>gen_4_cmp_pMux_1, f(0)=>gen_4_cmp_pMux_0);
   gen_4_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>
      gen_24_cmp_pInit_32, a(22)=>gen_24_cmp_pInit_32, a(21)=>
      gen_4_cmp_pMux_30, a(20)=>gen_4_cmp_pMux_29, a(19)=>gen_4_cmp_pMux_28, 
      a(18)=>gen_4_cmp_pMux_27, a(17)=>gen_4_cmp_pMux_26, a(16)=>
      gen_4_cmp_pMux_25, a(15)=>gen_4_cmp_pMux_24, a(14)=>gen_4_cmp_pMux_23, 
      a(13)=>gen_4_cmp_pMux_22, a(12)=>gen_4_cmp_pMux_21, a(11)=>
      gen_4_cmp_pMux_20, a(10)=>gen_4_cmp_pMux_19, a(9)=>gen_4_cmp_pMux_18, 
      a(8)=>gen_4_cmp_pMux_17, a(7)=>gen_4_cmp_pMux_16, a(6)=>
      gen_4_cmp_pMux_15, a(5)=>gen_4_cmp_pMux_14, a(4)=>gen_4_cmp_pMux_13, 
      a(3)=>gen_4_cmp_pMux_12, a(2)=>gen_4_cmp_pMux_11, a(1)=>
      gen_4_cmp_pMux_10, a(0)=>gen_4_cmp_pMux_9, b(23)=>nx10674, b(22)=>
      nx10674, b(21)=>nx10672, b(20)=>nx10680, b(19)=>nx10678, b(18)=>
      nx10676, b(17)=>nx10674, b(16)=>nx10672, b(15)=>gen_4_cmp_BSCmp_op2_15, 
      b(14)=>gen_4_cmp_BSCmp_op2_14, b(13)=>gen_4_cmp_BSCmp_op2_13, b(12)=>
      gen_4_cmp_BSCmp_op2_12, b(11)=>gen_4_cmp_BSCmp_op2_11, b(10)=>
      gen_4_cmp_BSCmp_op2_10, b(9)=>gen_4_cmp_BSCmp_op2_9, b(8)=>
      gen_4_cmp_BSCmp_op2_8, b(7)=>gen_4_cmp_BSCmp_op2_7, b(6)=>
      gen_4_cmp_BSCmp_op2_6, b(5)=>gen_4_cmp_BSCmp_op2_5, b(4)=>
      gen_4_cmp_BSCmp_op2_4, b(3)=>gen_4_cmp_BSCmp_op2_3, b(2)=>
      gen_4_cmp_BSCmp_op2_2, b(1)=>gen_4_cmp_BSCmp_op2_1, b(0)=>
      gen_4_cmp_BSCmp_op2_0, carryIn=>gen_4_cmp_BSCmp_carryIn, sum(23)=>
      gen_4_cmp_pBs_30, sum(22)=>gen_4_cmp_pBs_29, sum(21)=>gen_4_cmp_pBs_28, 
      sum(20)=>gen_4_cmp_pBs_27, sum(19)=>gen_4_cmp_pBs_26, sum(18)=>
      gen_4_cmp_pBs_25, sum(17)=>gen_4_cmp_pBs_24, sum(16)=>gen_4_cmp_pBs_23, 
      sum(15)=>outputs_4_15, sum(14)=>outputs_4_14, sum(13)=>outputs_4_13, 
      sum(12)=>outputs_4_12, sum(11)=>outputs_4_11, sum(10)=>outputs_4_10, 
      sum(9)=>outputs_4_9, sum(8)=>outputs_4_8, sum(7)=>outputs_4_7, sum(6)
      =>outputs_4_6, sum(5)=>outputs_4_5, sum(4)=>outputs_4_4, sum(3)=>
      outputs_4_3, sum(2)=>outputs_4_2, sum(1)=>outputs_4_1, sum(0)=>
      outputs_4_0, carryOut=>DANGLING(104));
   gen_3_cmp_pRegCmp : Reg_33 port map ( D(32)=>gen_24_cmp_pInit_32, D(31)=>
      gen_24_cmp_pInit_32, D(30)=>gen_3_cmp_pBs_30, D(29)=>gen_3_cmp_pBs_29, 
      D(28)=>gen_3_cmp_pBs_28, D(27)=>gen_3_cmp_pBs_27, D(26)=>
      gen_3_cmp_pBs_26, D(25)=>gen_3_cmp_pBs_25, D(24)=>gen_3_cmp_pBs_24, 
      D(23)=>gen_3_cmp_pBs_23, D(22)=>outputs_3_15, D(21)=>outputs_3_14, 
      D(20)=>outputs_3_13, D(19)=>outputs_3_12, D(18)=>outputs_3_11, D(17)=>
      outputs_3_10, D(16)=>outputs_3_9, D(15)=>outputs_3_8, D(14)=>
      outputs_3_7, D(13)=>outputs_3_6, D(12)=>outputs_3_5, D(11)=>
      outputs_3_4, D(10)=>outputs_3_3, D(9)=>outputs_3_2, D(8)=>outputs_3_1, 
      D(7)=>outputs_3_0, D(6)=>gen_3_cmp_pMux_8, D(5)=>gen_3_cmp_pMux_7, 
      D(4)=>gen_3_cmp_pMux_6, D(3)=>gen_3_cmp_pMux_5, D(2)=>gen_3_cmp_pMux_4, 
      D(1)=>gen_3_cmp_pMux_3, D(0)=>nx10382, en=>nx11928, clk=>nx10128, rst
      =>rst, Q(32)=>DANGLING(105), Q(31)=>DANGLING(106), Q(30)=>
      gen_3_cmp_pReg_30, Q(29)=>gen_3_cmp_pReg_29, Q(28)=>gen_3_cmp_pReg_28, 
      Q(27)=>gen_3_cmp_pReg_27, Q(26)=>gen_3_cmp_pReg_26, Q(25)=>
      gen_3_cmp_pReg_25, Q(24)=>gen_3_cmp_pReg_24, Q(23)=>gen_3_cmp_pReg_23, 
      Q(22)=>gen_3_cmp_pReg_22, Q(21)=>gen_3_cmp_pReg_21, Q(20)=>
      gen_3_cmp_pReg_20, Q(19)=>gen_3_cmp_pReg_19, Q(18)=>gen_3_cmp_pReg_18, 
      Q(17)=>gen_3_cmp_pReg_17, Q(16)=>gen_3_cmp_pReg_16, Q(15)=>
      gen_3_cmp_pReg_15, Q(14)=>gen_3_cmp_pReg_14, Q(13)=>gen_3_cmp_pReg_13, 
      Q(12)=>gen_3_cmp_pReg_12, Q(11)=>gen_3_cmp_pReg_11, Q(10)=>
      gen_3_cmp_pReg_10, Q(9)=>gen_3_cmp_pReg_9, Q(8)=>gen_3_cmp_pReg_8, 
      Q(7)=>gen_3_cmp_pReg_7, Q(6)=>gen_3_cmp_pReg_6, Q(5)=>gen_3_cmp_pReg_5, 
      Q(4)=>gen_3_cmp_pReg_4, Q(3)=>gen_3_cmp_pReg_3, Q(2)=>gen_3_cmp_pReg_2, 
      Q(1)=>gen_3_cmp_pReg_1, Q(0)=>gen_3_cmp_pReg_0);
   gen_3_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>gen_24_cmp_pInit_32, 
      a(31)=>gen_24_cmp_pInit_32, a(30)=>gen_3_cmp_pReg_30, a(29)=>
      gen_3_cmp_pReg_29, a(28)=>gen_3_cmp_pReg_28, a(27)=>gen_3_cmp_pReg_27, 
      a(26)=>gen_3_cmp_pReg_26, a(25)=>gen_3_cmp_pReg_25, a(24)=>
      gen_3_cmp_pReg_24, a(23)=>gen_3_cmp_pReg_23, a(22)=>gen_3_cmp_pReg_22, 
      a(21)=>gen_3_cmp_pReg_21, a(20)=>gen_3_cmp_pReg_20, a(19)=>
      gen_3_cmp_pReg_19, a(18)=>gen_3_cmp_pReg_18, a(17)=>gen_3_cmp_pReg_17, 
      a(16)=>gen_3_cmp_pReg_16, a(15)=>gen_3_cmp_pReg_15, a(14)=>
      gen_3_cmp_pReg_14, a(13)=>gen_3_cmp_pReg_13, a(12)=>gen_3_cmp_pReg_12, 
      a(11)=>gen_3_cmp_pReg_11, a(10)=>gen_3_cmp_pReg_10, a(9)=>
      gen_3_cmp_pReg_9, a(8)=>gen_3_cmp_pReg_8, a(7)=>gen_3_cmp_pReg_7, a(6)
      =>gen_3_cmp_pReg_6, a(5)=>gen_3_cmp_pReg_5, a(4)=>gen_3_cmp_pReg_4, 
      a(3)=>gen_3_cmp_pReg_3, a(2)=>gen_3_cmp_pReg_2, a(1)=>gen_3_cmp_pReg_1, 
      a(0)=>gen_3_cmp_pReg_0, b(32)=>gen_24_cmp_pInit_32, b(31)=>
      gen_24_cmp_pInit_32, b(30)=>gen_24_cmp_pInit_32, b(29)=>
      gen_24_cmp_pInit_32, b(28)=>gen_24_cmp_pInit_32, b(27)=>
      gen_24_cmp_pInit_32, b(26)=>gen_24_cmp_pInit_32, b(25)=>
      gen_24_cmp_pInit_32, b(24)=>gen_24_cmp_pInit_32, b(23)=>
      gen_24_cmp_pInit_32, b(22)=>gen_24_cmp_pInit_32, b(21)=>
      gen_24_cmp_pInit_32, b(20)=>gen_24_cmp_pInit_32, b(19)=>
      gen_24_cmp_pInit_32, b(18)=>gen_24_cmp_pInit_32, b(17)=>
      gen_24_cmp_pInit_32, b(16)=>gen_24_cmp_pInit_32, b(15)=>
      gen_24_cmp_pInit_32, b(14)=>gen_24_cmp_pInit_32, b(13)=>
      gen_24_cmp_pInit_32, b(12)=>gen_24_cmp_pInit_32, b(11)=>
      gen_24_cmp_pInit_32, b(10)=>gen_24_cmp_pInit_32, b(9)=>
      gen_24_cmp_pInit_32, b(8)=>filter_3_7, b(7)=>filter_3_6, b(6)=>
      filter_3_5, b(5)=>filter_3_4, b(4)=>filter_3_3, b(3)=>filter_3_2, b(2)
      =>filter_3_1, b(1)=>filter_3_0, b(0)=>gen_24_cmp_pInit_32, sel=>
      nx11914, f(32)=>DANGLING(107), f(31)=>DANGLING(108), f(30)=>
      gen_3_cmp_pMux_30, f(29)=>gen_3_cmp_pMux_29, f(28)=>gen_3_cmp_pMux_28, 
      f(27)=>gen_3_cmp_pMux_27, f(26)=>gen_3_cmp_pMux_26, f(25)=>
      gen_3_cmp_pMux_25, f(24)=>gen_3_cmp_pMux_24, f(23)=>gen_3_cmp_pMux_23, 
      f(22)=>gen_3_cmp_pMux_22, f(21)=>gen_3_cmp_pMux_21, f(20)=>
      gen_3_cmp_pMux_20, f(19)=>gen_3_cmp_pMux_19, f(18)=>gen_3_cmp_pMux_18, 
      f(17)=>gen_3_cmp_pMux_17, f(16)=>gen_3_cmp_pMux_16, f(15)=>
      gen_3_cmp_pMux_15, f(14)=>gen_3_cmp_pMux_14, f(13)=>gen_3_cmp_pMux_13, 
      f(12)=>gen_3_cmp_pMux_12, f(11)=>gen_3_cmp_pMux_11, f(10)=>
      gen_3_cmp_pMux_10, f(9)=>gen_3_cmp_pMux_9, f(8)=>gen_3_cmp_pMux_8, 
      f(7)=>gen_3_cmp_pMux_7, f(6)=>gen_3_cmp_pMux_6, f(5)=>gen_3_cmp_pMux_5, 
      f(4)=>gen_3_cmp_pMux_4, f(3)=>gen_3_cmp_pMux_3, f(2)=>gen_3_cmp_pMux_2, 
      f(1)=>gen_3_cmp_pMux_1, f(0)=>gen_3_cmp_pMux_0);
   gen_3_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>
      gen_24_cmp_pInit_32, a(22)=>gen_24_cmp_pInit_32, a(21)=>
      gen_3_cmp_pMux_30, a(20)=>gen_3_cmp_pMux_29, a(19)=>gen_3_cmp_pMux_28, 
      a(18)=>gen_3_cmp_pMux_27, a(17)=>gen_3_cmp_pMux_26, a(16)=>
      gen_3_cmp_pMux_25, a(15)=>gen_3_cmp_pMux_24, a(14)=>gen_3_cmp_pMux_23, 
      a(13)=>gen_3_cmp_pMux_22, a(12)=>gen_3_cmp_pMux_21, a(11)=>
      gen_3_cmp_pMux_20, a(10)=>gen_3_cmp_pMux_19, a(9)=>gen_3_cmp_pMux_18, 
      a(8)=>gen_3_cmp_pMux_17, a(7)=>gen_3_cmp_pMux_16, a(6)=>
      gen_3_cmp_pMux_15, a(5)=>gen_3_cmp_pMux_14, a(4)=>gen_3_cmp_pMux_13, 
      a(3)=>gen_3_cmp_pMux_12, a(2)=>gen_3_cmp_pMux_11, a(1)=>
      gen_3_cmp_pMux_10, a(0)=>gen_3_cmp_pMux_9, b(23)=>nx10686, b(22)=>
      nx10686, b(21)=>nx10684, b(20)=>nx10692, b(19)=>nx10690, b(18)=>
      nx10688, b(17)=>nx10686, b(16)=>nx10684, b(15)=>gen_3_cmp_BSCmp_op2_15, 
      b(14)=>gen_3_cmp_BSCmp_op2_14, b(13)=>gen_3_cmp_BSCmp_op2_13, b(12)=>
      gen_3_cmp_BSCmp_op2_12, b(11)=>gen_3_cmp_BSCmp_op2_11, b(10)=>
      gen_3_cmp_BSCmp_op2_10, b(9)=>gen_3_cmp_BSCmp_op2_9, b(8)=>
      gen_3_cmp_BSCmp_op2_8, b(7)=>gen_3_cmp_BSCmp_op2_7, b(6)=>
      gen_3_cmp_BSCmp_op2_6, b(5)=>gen_3_cmp_BSCmp_op2_5, b(4)=>
      gen_3_cmp_BSCmp_op2_4, b(3)=>gen_3_cmp_BSCmp_op2_3, b(2)=>
      gen_3_cmp_BSCmp_op2_2, b(1)=>gen_3_cmp_BSCmp_op2_1, b(0)=>
      gen_3_cmp_BSCmp_op2_0, carryIn=>gen_3_cmp_BSCmp_carryIn, sum(23)=>
      gen_3_cmp_pBs_30, sum(22)=>gen_3_cmp_pBs_29, sum(21)=>gen_3_cmp_pBs_28, 
      sum(20)=>gen_3_cmp_pBs_27, sum(19)=>gen_3_cmp_pBs_26, sum(18)=>
      gen_3_cmp_pBs_25, sum(17)=>gen_3_cmp_pBs_24, sum(16)=>gen_3_cmp_pBs_23, 
      sum(15)=>outputs_3_15, sum(14)=>outputs_3_14, sum(13)=>outputs_3_13, 
      sum(12)=>outputs_3_12, sum(11)=>outputs_3_11, sum(10)=>outputs_3_10, 
      sum(9)=>outputs_3_9, sum(8)=>outputs_3_8, sum(7)=>outputs_3_7, sum(6)
      =>outputs_3_6, sum(5)=>outputs_3_5, sum(4)=>outputs_3_4, sum(3)=>
      outputs_3_3, sum(2)=>outputs_3_2, sum(1)=>outputs_3_1, sum(0)=>
      outputs_3_0, carryOut=>DANGLING(109));
   gen_2_cmp_pRegCmp : Reg_33 port map ( D(32)=>gen_24_cmp_pInit_32, D(31)=>
      gen_24_cmp_pInit_32, D(30)=>gen_2_cmp_pBs_30, D(29)=>gen_2_cmp_pBs_29, 
      D(28)=>gen_2_cmp_pBs_28, D(27)=>gen_2_cmp_pBs_27, D(26)=>
      gen_2_cmp_pBs_26, D(25)=>gen_2_cmp_pBs_25, D(24)=>gen_2_cmp_pBs_24, 
      D(23)=>gen_2_cmp_pBs_23, D(22)=>outputs_2_15, D(21)=>outputs_2_14, 
      D(20)=>outputs_2_13, D(19)=>outputs_2_12, D(18)=>outputs_2_11, D(17)=>
      outputs_2_10, D(16)=>outputs_2_9, D(15)=>outputs_2_8, D(14)=>
      outputs_2_7, D(13)=>outputs_2_6, D(12)=>outputs_2_5, D(11)=>
      outputs_2_4, D(10)=>outputs_2_3, D(9)=>outputs_2_2, D(8)=>outputs_2_1, 
      D(7)=>outputs_2_0, D(6)=>gen_2_cmp_pMux_8, D(5)=>gen_2_cmp_pMux_7, 
      D(4)=>gen_2_cmp_pMux_6, D(3)=>gen_2_cmp_pMux_5, D(2)=>gen_2_cmp_pMux_4, 
      D(1)=>gen_2_cmp_pMux_3, D(0)=>nx10394, en=>nx11928, clk=>nx10128, rst
      =>rst, Q(32)=>DANGLING(110), Q(31)=>DANGLING(111), Q(30)=>
      gen_2_cmp_pReg_30, Q(29)=>gen_2_cmp_pReg_29, Q(28)=>gen_2_cmp_pReg_28, 
      Q(27)=>gen_2_cmp_pReg_27, Q(26)=>gen_2_cmp_pReg_26, Q(25)=>
      gen_2_cmp_pReg_25, Q(24)=>gen_2_cmp_pReg_24, Q(23)=>gen_2_cmp_pReg_23, 
      Q(22)=>gen_2_cmp_pReg_22, Q(21)=>gen_2_cmp_pReg_21, Q(20)=>
      gen_2_cmp_pReg_20, Q(19)=>gen_2_cmp_pReg_19, Q(18)=>gen_2_cmp_pReg_18, 
      Q(17)=>gen_2_cmp_pReg_17, Q(16)=>gen_2_cmp_pReg_16, Q(15)=>
      gen_2_cmp_pReg_15, Q(14)=>gen_2_cmp_pReg_14, Q(13)=>gen_2_cmp_pReg_13, 
      Q(12)=>gen_2_cmp_pReg_12, Q(11)=>gen_2_cmp_pReg_11, Q(10)=>
      gen_2_cmp_pReg_10, Q(9)=>gen_2_cmp_pReg_9, Q(8)=>gen_2_cmp_pReg_8, 
      Q(7)=>gen_2_cmp_pReg_7, Q(6)=>gen_2_cmp_pReg_6, Q(5)=>gen_2_cmp_pReg_5, 
      Q(4)=>gen_2_cmp_pReg_4, Q(3)=>gen_2_cmp_pReg_3, Q(2)=>gen_2_cmp_pReg_2, 
      Q(1)=>gen_2_cmp_pReg_1, Q(0)=>gen_2_cmp_pReg_0);
   gen_2_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>gen_24_cmp_pInit_32, 
      a(31)=>gen_24_cmp_pInit_32, a(30)=>gen_2_cmp_pReg_30, a(29)=>
      gen_2_cmp_pReg_29, a(28)=>gen_2_cmp_pReg_28, a(27)=>gen_2_cmp_pReg_27, 
      a(26)=>gen_2_cmp_pReg_26, a(25)=>gen_2_cmp_pReg_25, a(24)=>
      gen_2_cmp_pReg_24, a(23)=>gen_2_cmp_pReg_23, a(22)=>gen_2_cmp_pReg_22, 
      a(21)=>gen_2_cmp_pReg_21, a(20)=>gen_2_cmp_pReg_20, a(19)=>
      gen_2_cmp_pReg_19, a(18)=>gen_2_cmp_pReg_18, a(17)=>gen_2_cmp_pReg_17, 
      a(16)=>gen_2_cmp_pReg_16, a(15)=>gen_2_cmp_pReg_15, a(14)=>
      gen_2_cmp_pReg_14, a(13)=>gen_2_cmp_pReg_13, a(12)=>gen_2_cmp_pReg_12, 
      a(11)=>gen_2_cmp_pReg_11, a(10)=>gen_2_cmp_pReg_10, a(9)=>
      gen_2_cmp_pReg_9, a(8)=>gen_2_cmp_pReg_8, a(7)=>gen_2_cmp_pReg_7, a(6)
      =>gen_2_cmp_pReg_6, a(5)=>gen_2_cmp_pReg_5, a(4)=>gen_2_cmp_pReg_4, 
      a(3)=>gen_2_cmp_pReg_3, a(2)=>gen_2_cmp_pReg_2, a(1)=>gen_2_cmp_pReg_1, 
      a(0)=>gen_2_cmp_pReg_0, b(32)=>gen_24_cmp_pInit_32, b(31)=>
      gen_24_cmp_pInit_32, b(30)=>gen_24_cmp_pInit_32, b(29)=>
      gen_24_cmp_pInit_32, b(28)=>gen_24_cmp_pInit_32, b(27)=>
      gen_24_cmp_pInit_32, b(26)=>gen_24_cmp_pInit_32, b(25)=>
      gen_24_cmp_pInit_32, b(24)=>gen_24_cmp_pInit_32, b(23)=>
      gen_24_cmp_pInit_32, b(22)=>gen_24_cmp_pInit_32, b(21)=>
      gen_24_cmp_pInit_32, b(20)=>gen_24_cmp_pInit_32, b(19)=>
      gen_24_cmp_pInit_32, b(18)=>gen_24_cmp_pInit_32, b(17)=>
      gen_24_cmp_pInit_32, b(16)=>gen_24_cmp_pInit_32, b(15)=>
      gen_24_cmp_pInit_32, b(14)=>gen_24_cmp_pInit_32, b(13)=>
      gen_24_cmp_pInit_32, b(12)=>gen_24_cmp_pInit_32, b(11)=>
      gen_24_cmp_pInit_32, b(10)=>gen_24_cmp_pInit_32, b(9)=>
      gen_24_cmp_pInit_32, b(8)=>filter_2_7, b(7)=>filter_2_6, b(6)=>
      filter_2_5, b(5)=>filter_2_4, b(4)=>filter_2_3, b(3)=>filter_2_2, b(2)
      =>filter_2_1, b(1)=>filter_2_0, b(0)=>gen_24_cmp_pInit_32, sel=>
      nx11914, f(32)=>DANGLING(112), f(31)=>DANGLING(113), f(30)=>
      gen_2_cmp_pMux_30, f(29)=>gen_2_cmp_pMux_29, f(28)=>gen_2_cmp_pMux_28, 
      f(27)=>gen_2_cmp_pMux_27, f(26)=>gen_2_cmp_pMux_26, f(25)=>
      gen_2_cmp_pMux_25, f(24)=>gen_2_cmp_pMux_24, f(23)=>gen_2_cmp_pMux_23, 
      f(22)=>gen_2_cmp_pMux_22, f(21)=>gen_2_cmp_pMux_21, f(20)=>
      gen_2_cmp_pMux_20, f(19)=>gen_2_cmp_pMux_19, f(18)=>gen_2_cmp_pMux_18, 
      f(17)=>gen_2_cmp_pMux_17, f(16)=>gen_2_cmp_pMux_16, f(15)=>
      gen_2_cmp_pMux_15, f(14)=>gen_2_cmp_pMux_14, f(13)=>gen_2_cmp_pMux_13, 
      f(12)=>gen_2_cmp_pMux_12, f(11)=>gen_2_cmp_pMux_11, f(10)=>
      gen_2_cmp_pMux_10, f(9)=>gen_2_cmp_pMux_9, f(8)=>gen_2_cmp_pMux_8, 
      f(7)=>gen_2_cmp_pMux_7, f(6)=>gen_2_cmp_pMux_6, f(5)=>gen_2_cmp_pMux_5, 
      f(4)=>gen_2_cmp_pMux_4, f(3)=>gen_2_cmp_pMux_3, f(2)=>gen_2_cmp_pMux_2, 
      f(1)=>gen_2_cmp_pMux_1, f(0)=>gen_2_cmp_pMux_0);
   gen_2_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>
      gen_24_cmp_pInit_32, a(22)=>gen_24_cmp_pInit_32, a(21)=>
      gen_2_cmp_pMux_30, a(20)=>gen_2_cmp_pMux_29, a(19)=>gen_2_cmp_pMux_28, 
      a(18)=>gen_2_cmp_pMux_27, a(17)=>gen_2_cmp_pMux_26, a(16)=>
      gen_2_cmp_pMux_25, a(15)=>gen_2_cmp_pMux_24, a(14)=>gen_2_cmp_pMux_23, 
      a(13)=>gen_2_cmp_pMux_22, a(12)=>gen_2_cmp_pMux_21, a(11)=>
      gen_2_cmp_pMux_20, a(10)=>gen_2_cmp_pMux_19, a(9)=>gen_2_cmp_pMux_18, 
      a(8)=>gen_2_cmp_pMux_17, a(7)=>gen_2_cmp_pMux_16, a(6)=>
      gen_2_cmp_pMux_15, a(5)=>gen_2_cmp_pMux_14, a(4)=>gen_2_cmp_pMux_13, 
      a(3)=>gen_2_cmp_pMux_12, a(2)=>gen_2_cmp_pMux_11, a(1)=>
      gen_2_cmp_pMux_10, a(0)=>gen_2_cmp_pMux_9, b(23)=>nx10698, b(22)=>
      nx10698, b(21)=>nx10696, b(20)=>nx10704, b(19)=>nx10702, b(18)=>
      nx10700, b(17)=>nx10698, b(16)=>nx10696, b(15)=>gen_2_cmp_BSCmp_op2_15, 
      b(14)=>gen_2_cmp_BSCmp_op2_14, b(13)=>gen_2_cmp_BSCmp_op2_13, b(12)=>
      gen_2_cmp_BSCmp_op2_12, b(11)=>gen_2_cmp_BSCmp_op2_11, b(10)=>
      gen_2_cmp_BSCmp_op2_10, b(9)=>gen_2_cmp_BSCmp_op2_9, b(8)=>
      gen_2_cmp_BSCmp_op2_8, b(7)=>gen_2_cmp_BSCmp_op2_7, b(6)=>
      gen_2_cmp_BSCmp_op2_6, b(5)=>gen_2_cmp_BSCmp_op2_5, b(4)=>
      gen_2_cmp_BSCmp_op2_4, b(3)=>gen_2_cmp_BSCmp_op2_3, b(2)=>
      gen_2_cmp_BSCmp_op2_2, b(1)=>gen_2_cmp_BSCmp_op2_1, b(0)=>
      gen_2_cmp_BSCmp_op2_0, carryIn=>gen_2_cmp_BSCmp_carryIn, sum(23)=>
      gen_2_cmp_pBs_30, sum(22)=>gen_2_cmp_pBs_29, sum(21)=>gen_2_cmp_pBs_28, 
      sum(20)=>gen_2_cmp_pBs_27, sum(19)=>gen_2_cmp_pBs_26, sum(18)=>
      gen_2_cmp_pBs_25, sum(17)=>gen_2_cmp_pBs_24, sum(16)=>gen_2_cmp_pBs_23, 
      sum(15)=>outputs_2_15, sum(14)=>outputs_2_14, sum(13)=>outputs_2_13, 
      sum(12)=>outputs_2_12, sum(11)=>outputs_2_11, sum(10)=>outputs_2_10, 
      sum(9)=>outputs_2_9, sum(8)=>outputs_2_8, sum(7)=>outputs_2_7, sum(6)
      =>outputs_2_6, sum(5)=>outputs_2_5, sum(4)=>outputs_2_4, sum(3)=>
      outputs_2_3, sum(2)=>outputs_2_2, sum(1)=>outputs_2_1, sum(0)=>
      outputs_2_0, carryOut=>DANGLING(114));
   gen_1_cmp_pRegCmp : Reg_33 port map ( D(32)=>gen_24_cmp_pInit_32, D(31)=>
      gen_24_cmp_pInit_32, D(30)=>gen_1_cmp_pBs_30, D(29)=>gen_1_cmp_pBs_29, 
      D(28)=>gen_1_cmp_pBs_28, D(27)=>gen_1_cmp_pBs_27, D(26)=>
      gen_1_cmp_pBs_26, D(25)=>gen_1_cmp_pBs_25, D(24)=>gen_1_cmp_pBs_24, 
      D(23)=>gen_1_cmp_pBs_23, D(22)=>outputs_1_15, D(21)=>outputs_1_14, 
      D(20)=>outputs_1_13, D(19)=>outputs_1_12, D(18)=>outputs_1_11, D(17)=>
      outputs_1_10, D(16)=>outputs_1_9, D(15)=>outputs_1_8, D(14)=>
      outputs_1_7, D(13)=>outputs_1_6, D(12)=>outputs_1_5, D(11)=>
      outputs_1_4, D(10)=>outputs_1_3, D(9)=>outputs_1_2, D(8)=>outputs_1_1, 
      D(7)=>outputs_1_0, D(6)=>gen_1_cmp_pMux_8, D(5)=>gen_1_cmp_pMux_7, 
      D(4)=>gen_1_cmp_pMux_6, D(3)=>gen_1_cmp_pMux_5, D(2)=>gen_1_cmp_pMux_4, 
      D(1)=>gen_1_cmp_pMux_3, D(0)=>nx10406, en=>nx11928, clk=>nx10128, rst
      =>rst, Q(32)=>DANGLING(115), Q(31)=>DANGLING(116), Q(30)=>
      gen_1_cmp_pReg_30, Q(29)=>gen_1_cmp_pReg_29, Q(28)=>gen_1_cmp_pReg_28, 
      Q(27)=>gen_1_cmp_pReg_27, Q(26)=>gen_1_cmp_pReg_26, Q(25)=>
      gen_1_cmp_pReg_25, Q(24)=>gen_1_cmp_pReg_24, Q(23)=>gen_1_cmp_pReg_23, 
      Q(22)=>gen_1_cmp_pReg_22, Q(21)=>gen_1_cmp_pReg_21, Q(20)=>
      gen_1_cmp_pReg_20, Q(19)=>gen_1_cmp_pReg_19, Q(18)=>gen_1_cmp_pReg_18, 
      Q(17)=>gen_1_cmp_pReg_17, Q(16)=>gen_1_cmp_pReg_16, Q(15)=>
      gen_1_cmp_pReg_15, Q(14)=>gen_1_cmp_pReg_14, Q(13)=>gen_1_cmp_pReg_13, 
      Q(12)=>gen_1_cmp_pReg_12, Q(11)=>gen_1_cmp_pReg_11, Q(10)=>
      gen_1_cmp_pReg_10, Q(9)=>gen_1_cmp_pReg_9, Q(8)=>gen_1_cmp_pReg_8, 
      Q(7)=>gen_1_cmp_pReg_7, Q(6)=>gen_1_cmp_pReg_6, Q(5)=>gen_1_cmp_pReg_5, 
      Q(4)=>gen_1_cmp_pReg_4, Q(3)=>gen_1_cmp_pReg_3, Q(2)=>gen_1_cmp_pReg_2, 
      Q(1)=>gen_1_cmp_pReg_1, Q(0)=>gen_1_cmp_pReg_0);
   gen_1_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>gen_24_cmp_pInit_32, 
      a(31)=>gen_24_cmp_pInit_32, a(30)=>gen_1_cmp_pReg_30, a(29)=>
      gen_1_cmp_pReg_29, a(28)=>gen_1_cmp_pReg_28, a(27)=>gen_1_cmp_pReg_27, 
      a(26)=>gen_1_cmp_pReg_26, a(25)=>gen_1_cmp_pReg_25, a(24)=>
      gen_1_cmp_pReg_24, a(23)=>gen_1_cmp_pReg_23, a(22)=>gen_1_cmp_pReg_22, 
      a(21)=>gen_1_cmp_pReg_21, a(20)=>gen_1_cmp_pReg_20, a(19)=>
      gen_1_cmp_pReg_19, a(18)=>gen_1_cmp_pReg_18, a(17)=>gen_1_cmp_pReg_17, 
      a(16)=>gen_1_cmp_pReg_16, a(15)=>gen_1_cmp_pReg_15, a(14)=>
      gen_1_cmp_pReg_14, a(13)=>gen_1_cmp_pReg_13, a(12)=>gen_1_cmp_pReg_12, 
      a(11)=>gen_1_cmp_pReg_11, a(10)=>gen_1_cmp_pReg_10, a(9)=>
      gen_1_cmp_pReg_9, a(8)=>gen_1_cmp_pReg_8, a(7)=>gen_1_cmp_pReg_7, a(6)
      =>gen_1_cmp_pReg_6, a(5)=>gen_1_cmp_pReg_5, a(4)=>gen_1_cmp_pReg_4, 
      a(3)=>gen_1_cmp_pReg_3, a(2)=>gen_1_cmp_pReg_2, a(1)=>gen_1_cmp_pReg_1, 
      a(0)=>gen_1_cmp_pReg_0, b(32)=>gen_24_cmp_pInit_32, b(31)=>
      gen_24_cmp_pInit_32, b(30)=>gen_24_cmp_pInit_32, b(29)=>
      gen_24_cmp_pInit_32, b(28)=>gen_24_cmp_pInit_32, b(27)=>
      gen_24_cmp_pInit_32, b(26)=>gen_24_cmp_pInit_32, b(25)=>
      gen_24_cmp_pInit_32, b(24)=>gen_24_cmp_pInit_32, b(23)=>
      gen_24_cmp_pInit_32, b(22)=>gen_24_cmp_pInit_32, b(21)=>
      gen_24_cmp_pInit_32, b(20)=>gen_24_cmp_pInit_32, b(19)=>
      gen_24_cmp_pInit_32, b(18)=>gen_24_cmp_pInit_32, b(17)=>
      gen_24_cmp_pInit_32, b(16)=>gen_24_cmp_pInit_32, b(15)=>
      gen_24_cmp_pInit_32, b(14)=>gen_24_cmp_pInit_32, b(13)=>
      gen_24_cmp_pInit_32, b(12)=>gen_24_cmp_pInit_32, b(11)=>
      gen_24_cmp_pInit_32, b(10)=>gen_24_cmp_pInit_32, b(9)=>
      gen_24_cmp_pInit_32, b(8)=>filter_1_7, b(7)=>filter_1_6, b(6)=>
      filter_1_5, b(5)=>filter_1_4, b(4)=>filter_1_3, b(3)=>filter_1_2, b(2)
      =>filter_1_1, b(1)=>filter_1_0, b(0)=>gen_24_cmp_pInit_32, sel=>
      nx10120, f(32)=>DANGLING(117), f(31)=>DANGLING(118), f(30)=>
      gen_1_cmp_pMux_30, f(29)=>gen_1_cmp_pMux_29, f(28)=>gen_1_cmp_pMux_28, 
      f(27)=>gen_1_cmp_pMux_27, f(26)=>gen_1_cmp_pMux_26, f(25)=>
      gen_1_cmp_pMux_25, f(24)=>gen_1_cmp_pMux_24, f(23)=>gen_1_cmp_pMux_23, 
      f(22)=>gen_1_cmp_pMux_22, f(21)=>gen_1_cmp_pMux_21, f(20)=>
      gen_1_cmp_pMux_20, f(19)=>gen_1_cmp_pMux_19, f(18)=>gen_1_cmp_pMux_18, 
      f(17)=>gen_1_cmp_pMux_17, f(16)=>gen_1_cmp_pMux_16, f(15)=>
      gen_1_cmp_pMux_15, f(14)=>gen_1_cmp_pMux_14, f(13)=>gen_1_cmp_pMux_13, 
      f(12)=>gen_1_cmp_pMux_12, f(11)=>gen_1_cmp_pMux_11, f(10)=>
      gen_1_cmp_pMux_10, f(9)=>gen_1_cmp_pMux_9, f(8)=>gen_1_cmp_pMux_8, 
      f(7)=>gen_1_cmp_pMux_7, f(6)=>gen_1_cmp_pMux_6, f(5)=>gen_1_cmp_pMux_5, 
      f(4)=>gen_1_cmp_pMux_4, f(3)=>gen_1_cmp_pMux_3, f(2)=>gen_1_cmp_pMux_2, 
      f(1)=>gen_1_cmp_pMux_1, f(0)=>gen_1_cmp_pMux_0);
   gen_1_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>
      gen_24_cmp_pInit_32, a(22)=>gen_24_cmp_pInit_32, a(21)=>
      gen_1_cmp_pMux_30, a(20)=>gen_1_cmp_pMux_29, a(19)=>gen_1_cmp_pMux_28, 
      a(18)=>gen_1_cmp_pMux_27, a(17)=>gen_1_cmp_pMux_26, a(16)=>
      gen_1_cmp_pMux_25, a(15)=>gen_1_cmp_pMux_24, a(14)=>gen_1_cmp_pMux_23, 
      a(13)=>gen_1_cmp_pMux_22, a(12)=>gen_1_cmp_pMux_21, a(11)=>
      gen_1_cmp_pMux_20, a(10)=>gen_1_cmp_pMux_19, a(9)=>gen_1_cmp_pMux_18, 
      a(8)=>gen_1_cmp_pMux_17, a(7)=>gen_1_cmp_pMux_16, a(6)=>
      gen_1_cmp_pMux_15, a(5)=>gen_1_cmp_pMux_14, a(4)=>gen_1_cmp_pMux_13, 
      a(3)=>gen_1_cmp_pMux_12, a(2)=>gen_1_cmp_pMux_11, a(1)=>
      gen_1_cmp_pMux_10, a(0)=>gen_1_cmp_pMux_9, b(23)=>nx10710, b(22)=>
      nx10710, b(21)=>nx10708, b(20)=>nx10716, b(19)=>nx10714, b(18)=>
      nx10712, b(17)=>nx10710, b(16)=>nx10708, b(15)=>gen_1_cmp_BSCmp_op2_15, 
      b(14)=>gen_1_cmp_BSCmp_op2_14, b(13)=>gen_1_cmp_BSCmp_op2_13, b(12)=>
      gen_1_cmp_BSCmp_op2_12, b(11)=>gen_1_cmp_BSCmp_op2_11, b(10)=>
      gen_1_cmp_BSCmp_op2_10, b(9)=>gen_1_cmp_BSCmp_op2_9, b(8)=>
      gen_1_cmp_BSCmp_op2_8, b(7)=>gen_1_cmp_BSCmp_op2_7, b(6)=>
      gen_1_cmp_BSCmp_op2_6, b(5)=>gen_1_cmp_BSCmp_op2_5, b(4)=>
      gen_1_cmp_BSCmp_op2_4, b(3)=>gen_1_cmp_BSCmp_op2_3, b(2)=>
      gen_1_cmp_BSCmp_op2_2, b(1)=>gen_1_cmp_BSCmp_op2_1, b(0)=>
      gen_1_cmp_BSCmp_op2_0, carryIn=>gen_1_cmp_BSCmp_carryIn, sum(23)=>
      gen_1_cmp_pBs_30, sum(22)=>gen_1_cmp_pBs_29, sum(21)=>gen_1_cmp_pBs_28, 
      sum(20)=>gen_1_cmp_pBs_27, sum(19)=>gen_1_cmp_pBs_26, sum(18)=>
      gen_1_cmp_pBs_25, sum(17)=>gen_1_cmp_pBs_24, sum(16)=>gen_1_cmp_pBs_23, 
      sum(15)=>outputs_1_15, sum(14)=>outputs_1_14, sum(13)=>outputs_1_13, 
      sum(12)=>outputs_1_12, sum(11)=>outputs_1_11, sum(10)=>outputs_1_10, 
      sum(9)=>outputs_1_9, sum(8)=>outputs_1_8, sum(7)=>outputs_1_7, sum(6)
      =>outputs_1_6, sum(5)=>outputs_1_5, sum(4)=>outputs_1_4, sum(3)=>
      outputs_1_3, sum(2)=>outputs_1_2, sum(1)=>outputs_1_1, sum(0)=>
      outputs_1_0, carryOut=>DANGLING(119));
   gen_0_cmp_pRegCmp : Reg_33 port map ( D(32)=>gen_24_cmp_pInit_32, D(31)=>
      gen_24_cmp_pInit_32, D(30)=>gen_0_cmp_pBs_30, D(29)=>gen_0_cmp_pBs_29, 
      D(28)=>gen_0_cmp_pBs_28, D(27)=>gen_0_cmp_pBs_27, D(26)=>
      gen_0_cmp_pBs_26, D(25)=>gen_0_cmp_pBs_25, D(24)=>gen_0_cmp_pBs_24, 
      D(23)=>gen_0_cmp_pBs_23, D(22)=>outputs_0_15, D(21)=>outputs_0_14, 
      D(20)=>outputs_0_13, D(19)=>outputs_0_12, D(18)=>outputs_0_11, D(17)=>
      outputs_0_10, D(16)=>outputs_0_9, D(15)=>outputs_0_8, D(14)=>
      outputs_0_7, D(13)=>outputs_0_6, D(12)=>outputs_0_5, D(11)=>
      outputs_0_4, D(10)=>outputs_0_3, D(9)=>outputs_0_2, D(8)=>outputs_0_1, 
      D(7)=>outputs_0_0, D(6)=>gen_0_cmp_pMux_8, D(5)=>gen_0_cmp_pMux_7, 
      D(4)=>gen_0_cmp_pMux_6, D(3)=>gen_0_cmp_pMux_5, D(2)=>gen_0_cmp_pMux_4, 
      D(1)=>gen_0_cmp_pMux_3, D(0)=>nx10418, en=>nx10886, clk=>nx10128, rst
      =>rst, Q(32)=>DANGLING(120), Q(31)=>DANGLING(121), Q(30)=>
      gen_0_cmp_pReg_30, Q(29)=>gen_0_cmp_pReg_29, Q(28)=>gen_0_cmp_pReg_28, 
      Q(27)=>gen_0_cmp_pReg_27, Q(26)=>gen_0_cmp_pReg_26, Q(25)=>
      gen_0_cmp_pReg_25, Q(24)=>gen_0_cmp_pReg_24, Q(23)=>gen_0_cmp_pReg_23, 
      Q(22)=>gen_0_cmp_pReg_22, Q(21)=>gen_0_cmp_pReg_21, Q(20)=>
      gen_0_cmp_pReg_20, Q(19)=>gen_0_cmp_pReg_19, Q(18)=>gen_0_cmp_pReg_18, 
      Q(17)=>gen_0_cmp_pReg_17, Q(16)=>gen_0_cmp_pReg_16, Q(15)=>
      gen_0_cmp_pReg_15, Q(14)=>gen_0_cmp_pReg_14, Q(13)=>gen_0_cmp_pReg_13, 
      Q(12)=>gen_0_cmp_pReg_12, Q(11)=>gen_0_cmp_pReg_11, Q(10)=>
      gen_0_cmp_pReg_10, Q(9)=>gen_0_cmp_pReg_9, Q(8)=>gen_0_cmp_pReg_8, 
      Q(7)=>gen_0_cmp_pReg_7, Q(6)=>gen_0_cmp_pReg_6, Q(5)=>gen_0_cmp_pReg_5, 
      Q(4)=>gen_0_cmp_pReg_4, Q(3)=>gen_0_cmp_pReg_3, Q(2)=>gen_0_cmp_pReg_2, 
      Q(1)=>gen_0_cmp_pReg_1, Q(0)=>gen_0_cmp_pReg_0);
   gen_0_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>gen_24_cmp_pInit_32, 
      a(31)=>gen_24_cmp_pInit_32, a(30)=>gen_0_cmp_pReg_30, a(29)=>
      gen_0_cmp_pReg_29, a(28)=>gen_0_cmp_pReg_28, a(27)=>gen_0_cmp_pReg_27, 
      a(26)=>gen_0_cmp_pReg_26, a(25)=>gen_0_cmp_pReg_25, a(24)=>
      gen_0_cmp_pReg_24, a(23)=>gen_0_cmp_pReg_23, a(22)=>gen_0_cmp_pReg_22, 
      a(21)=>gen_0_cmp_pReg_21, a(20)=>gen_0_cmp_pReg_20, a(19)=>
      gen_0_cmp_pReg_19, a(18)=>gen_0_cmp_pReg_18, a(17)=>gen_0_cmp_pReg_17, 
      a(16)=>gen_0_cmp_pReg_16, a(15)=>gen_0_cmp_pReg_15, a(14)=>
      gen_0_cmp_pReg_14, a(13)=>gen_0_cmp_pReg_13, a(12)=>gen_0_cmp_pReg_12, 
      a(11)=>gen_0_cmp_pReg_11, a(10)=>gen_0_cmp_pReg_10, a(9)=>
      gen_0_cmp_pReg_9, a(8)=>gen_0_cmp_pReg_8, a(7)=>gen_0_cmp_pReg_7, a(6)
      =>gen_0_cmp_pReg_6, a(5)=>gen_0_cmp_pReg_5, a(4)=>gen_0_cmp_pReg_4, 
      a(3)=>gen_0_cmp_pReg_3, a(2)=>gen_0_cmp_pReg_2, a(1)=>gen_0_cmp_pReg_1, 
      a(0)=>gen_0_cmp_pReg_0, b(32)=>gen_24_cmp_pInit_32, b(31)=>
      gen_24_cmp_pInit_32, b(30)=>gen_24_cmp_pInit_32, b(29)=>
      gen_24_cmp_pInit_32, b(28)=>gen_24_cmp_pInit_32, b(27)=>
      gen_24_cmp_pInit_32, b(26)=>gen_24_cmp_pInit_32, b(25)=>
      gen_24_cmp_pInit_32, b(24)=>gen_24_cmp_pInit_32, b(23)=>
      gen_24_cmp_pInit_32, b(22)=>gen_24_cmp_pInit_32, b(21)=>
      gen_24_cmp_pInit_32, b(20)=>gen_24_cmp_pInit_32, b(19)=>
      gen_24_cmp_pInit_32, b(18)=>gen_24_cmp_pInit_32, b(17)=>
      gen_24_cmp_pInit_32, b(16)=>gen_24_cmp_pInit_32, b(15)=>
      gen_24_cmp_pInit_32, b(14)=>gen_24_cmp_pInit_32, b(13)=>
      gen_24_cmp_pInit_32, b(12)=>gen_24_cmp_pInit_32, b(11)=>
      gen_24_cmp_pInit_32, b(10)=>gen_24_cmp_pInit_32, b(9)=>
      gen_24_cmp_pInit_32, b(8)=>filter_0_7, b(7)=>filter_0_6, b(6)=>
      filter_0_5, b(5)=>filter_0_4, b(4)=>filter_0_3, b(3)=>filter_0_2, b(2)
      =>filter_0_1, b(1)=>filter_0_0, b(0)=>gen_24_cmp_pInit_32, sel=>
      nx10120, f(32)=>DANGLING(122), f(31)=>DANGLING(123), f(30)=>
      gen_0_cmp_pMux_30, f(29)=>gen_0_cmp_pMux_29, f(28)=>gen_0_cmp_pMux_28, 
      f(27)=>gen_0_cmp_pMux_27, f(26)=>gen_0_cmp_pMux_26, f(25)=>
      gen_0_cmp_pMux_25, f(24)=>gen_0_cmp_pMux_24, f(23)=>gen_0_cmp_pMux_23, 
      f(22)=>gen_0_cmp_pMux_22, f(21)=>gen_0_cmp_pMux_21, f(20)=>
      gen_0_cmp_pMux_20, f(19)=>gen_0_cmp_pMux_19, f(18)=>gen_0_cmp_pMux_18, 
      f(17)=>gen_0_cmp_pMux_17, f(16)=>gen_0_cmp_pMux_16, f(15)=>
      gen_0_cmp_pMux_15, f(14)=>gen_0_cmp_pMux_14, f(13)=>gen_0_cmp_pMux_13, 
      f(12)=>gen_0_cmp_pMux_12, f(11)=>gen_0_cmp_pMux_11, f(10)=>
      gen_0_cmp_pMux_10, f(9)=>gen_0_cmp_pMux_9, f(8)=>gen_0_cmp_pMux_8, 
      f(7)=>gen_0_cmp_pMux_7, f(6)=>gen_0_cmp_pMux_6, f(5)=>gen_0_cmp_pMux_5, 
      f(4)=>gen_0_cmp_pMux_4, f(3)=>gen_0_cmp_pMux_3, f(2)=>gen_0_cmp_pMux_2, 
      f(1)=>gen_0_cmp_pMux_1, f(0)=>gen_0_cmp_pMux_0);
   gen_0_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>
      gen_24_cmp_pInit_32, a(22)=>gen_24_cmp_pInit_32, a(21)=>
      gen_0_cmp_pMux_30, a(20)=>gen_0_cmp_pMux_29, a(19)=>gen_0_cmp_pMux_28, 
      a(18)=>gen_0_cmp_pMux_27, a(17)=>gen_0_cmp_pMux_26, a(16)=>
      gen_0_cmp_pMux_25, a(15)=>gen_0_cmp_pMux_24, a(14)=>gen_0_cmp_pMux_23, 
      a(13)=>gen_0_cmp_pMux_22, a(12)=>gen_0_cmp_pMux_21, a(11)=>
      gen_0_cmp_pMux_20, a(10)=>gen_0_cmp_pMux_19, a(9)=>gen_0_cmp_pMux_18, 
      a(8)=>gen_0_cmp_pMux_17, a(7)=>gen_0_cmp_pMux_16, a(6)=>
      gen_0_cmp_pMux_15, a(5)=>gen_0_cmp_pMux_14, a(4)=>gen_0_cmp_pMux_13, 
      a(3)=>gen_0_cmp_pMux_12, a(2)=>gen_0_cmp_pMux_11, a(1)=>
      gen_0_cmp_pMux_10, a(0)=>gen_0_cmp_pMux_9, b(23)=>nx10722, b(22)=>
      nx10722, b(21)=>nx10720, b(20)=>nx10728, b(19)=>nx10726, b(18)=>
      nx10724, b(17)=>nx10722, b(16)=>nx10720, b(15)=>gen_0_cmp_BSCmp_op2_15, 
      b(14)=>gen_0_cmp_BSCmp_op2_14, b(13)=>gen_0_cmp_BSCmp_op2_13, b(12)=>
      gen_0_cmp_BSCmp_op2_12, b(11)=>gen_0_cmp_BSCmp_op2_11, b(10)=>
      gen_0_cmp_BSCmp_op2_10, b(9)=>gen_0_cmp_BSCmp_op2_9, b(8)=>
      gen_0_cmp_BSCmp_op2_8, b(7)=>gen_0_cmp_BSCmp_op2_7, b(6)=>
      gen_0_cmp_BSCmp_op2_6, b(5)=>gen_0_cmp_BSCmp_op2_5, b(4)=>
      gen_0_cmp_BSCmp_op2_4, b(3)=>gen_0_cmp_BSCmp_op2_3, b(2)=>
      gen_0_cmp_BSCmp_op2_2, b(1)=>gen_0_cmp_BSCmp_op2_1, b(0)=>
      gen_0_cmp_BSCmp_op2_0, carryIn=>gen_0_cmp_BSCmp_carryIn, sum(23)=>
      gen_0_cmp_pBs_30, sum(22)=>gen_0_cmp_pBs_29, sum(21)=>gen_0_cmp_pBs_28, 
      sum(20)=>gen_0_cmp_pBs_27, sum(19)=>gen_0_cmp_pBs_26, sum(18)=>
      gen_0_cmp_pBs_25, sum(17)=>gen_0_cmp_pBs_24, sum(16)=>gen_0_cmp_pBs_23, 
      sum(15)=>outputs_0_15, sum(14)=>outputs_0_14, sum(13)=>outputs_0_13, 
      sum(12)=>outputs_0_12, sum(11)=>outputs_0_11, sum(10)=>outputs_0_10, 
      sum(9)=>outputs_0_9, sum(8)=>outputs_0_8, sum(7)=>outputs_0_7, sum(6)
      =>outputs_0_6, sum(5)=>outputs_0_5, sum(4)=>outputs_0_4, sum(3)=>
      outputs_0_3, sum(2)=>outputs_0_2, sum(1)=>outputs_0_1, sum(0)=>
      outputs_0_0, carryOut=>DANGLING(124));
   ix3692 : nand02 port map ( Y=>nx3691, A0=>nx11928, A1=>nx3729);
   CounterCmp_reg_outp_3 : dffr port map ( Q=>done, QB=>OPEN, D=>nx3691, CLK
      =>clk, R=>nx9666);
   ix9667 : inv01 port map ( Y=>nx9666, A=>nx3713);
   ix3714 : nor02_2x port map ( Y=>nx3713, A0=>restartDetection, A1=>rst);
   StartCaptuerCmp_reg_f : dffr port map ( Q=>restartDetection, QB=>OPEN, D
      =>nx9650, CLK=>start, R=>nx9660);
   ix9651 : fake_vcc port map ( Y=>nx9650);
   ix9661 : inv01 port map ( Y=>nx9660, A=>nx3720);
   ix3721 : nor02_2x port map ( Y=>nx3720, A0=>StartCaptuerCmp_d, A1=>rst);
   StartCaptuerCmp_reg_d : dff port map ( Q=>StartCaptuerCmp_d, QB=>OPEN, D
      =>restartDetection, CLK=>nx10128);
   CounterCmp_reg_outp_2 : dffr port map ( Q=>OPEN, QB=>nx3729, D=>nx3681, 
      CLK=>clk, R=>nx9666);
   ix3682 : mux21 port map ( Y=>nx3681, A0=>nx3733, A1=>nx3729, S0=>nx11934
   );
   ix3672 : nand02 port map ( Y=>nx3671, A0=>nx3737, A1=>nx3741);
   ix3738 : nand02 port map ( Y=>nx3737, A0=>CounterCmp_outp_1, A1=>nx11934
   );
   CounterCmp_reg_outp_1 : dffr port map ( Q=>CounterCmp_outp_1, QB=>nx3733, 
      D=>nx3671, CLK=>clk, R=>nx9666);
   ix3742 : nand02 port map ( Y=>nx3741, A0=>nx11914, A1=>nx10886);
   ix3698 : nor02_2x port map ( Y=>nx3697, A0=>nx11938, A1=>nx10886);
   CounterCmp_reg_outp_0 : dffs_ni port map ( Q=>OPEN, QB=>nx3745, D=>nx3697, 
      CLK=>clk, S=>nx9666);
   ix3184 : fake_gnd port map ( Y=>gen_24_cmp_pInit_32);
   ix67 : nand02 port map ( Y=>gen_0_cmp_BSCmp_op2_1, A0=>nx3751, A1=>nx3771
   );
   ix3752 : nor02_2x port map ( Y=>nx3751, A0=>nx62, A1=>nx58);
   ix63 : nor03_2x port map ( Y=>nx62, A0=>gen_0_cmp_mReg_0, A1=>nx10424, A2
      =>nx10890);
   gen_0_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_0_cmp_mReg_0, QB=>
      nx3757, D=>window_0_0, CLK=>start, R=>rst);
   ix3762 : inv01 port map ( Y=>nx3761, A=>gen_0_cmp_pMux_0);
   ix59 : nor03_2x port map ( Y=>nx58, A0=>nx3757, A1=>nx10896, A2=>nx10906
   );
   ix3770 : inv02 port map ( Y=>nx3769, A=>gen_0_cmp_pMux_2);
   ix3772 : nor02_2x port map ( Y=>nx3771, A0=>nx48, A1=>nx46);
   ix49 : nor03_2x port map ( Y=>nx48, A0=>nx3775, A1=>nx10418, A2=>nx10914
   );
   gen_0_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_0_cmp_mReg_1, QB=>
      nx3775, D=>window_0_1, CLK=>start, R=>rst);
   ix47 : nor03_2x port map ( Y=>nx46, A0=>gen_0_cmp_mReg_1, A1=>nx10730, A2
      =>nx10922);
   ix7 : nor03_2x port map ( Y=>nx6, A0=>nx10424, A1=>nx3769, A2=>
      gen_0_cmp_pMux_0);
   ix89 : nand02 port map ( Y=>gen_0_cmp_BSCmp_op2_2, A0=>nx3786, A1=>nx3791
   );
   ix3787 : nor02_2x port map ( Y=>nx3786, A0=>nx84, A1=>nx80);
   ix85 : nor03_2x port map ( Y=>nx84, A0=>gen_0_cmp_mReg_1, A1=>nx10424, A2
      =>nx10890);
   ix81 : nor03_2x port map ( Y=>nx80, A0=>nx3775, A1=>nx10896, A2=>nx10906
   );
   ix3792 : nor02_2x port map ( Y=>nx3791, A0=>nx76, A1=>nx74);
   ix77 : nor03_2x port map ( Y=>nx76, A0=>nx3795, A1=>nx10418, A2=>nx10914
   );
   gen_0_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_0_cmp_mReg_2, QB=>
      nx3795, D=>window_0_2, CLK=>start, R=>rst);
   ix75 : nor03_2x port map ( Y=>nx74, A0=>gen_0_cmp_mReg_2, A1=>nx10730, A2
      =>nx10922);
   ix111 : nand02 port map ( Y=>gen_0_cmp_BSCmp_op2_3, A0=>nx3801, A1=>
      nx3807);
   ix3802 : nor02_2x port map ( Y=>nx3801, A0=>nx106, A1=>nx102);
   ix107 : nor03_2x port map ( Y=>nx106, A0=>gen_0_cmp_mReg_2, A1=>nx10424, 
      A2=>nx10890);
   ix103 : nor03_2x port map ( Y=>nx102, A0=>nx3795, A1=>nx10896, A2=>
      nx10906);
   ix3808 : nor02_2x port map ( Y=>nx3807, A0=>nx98, A1=>nx96);
   ix99 : nor03_2x port map ( Y=>nx98, A0=>nx3810, A1=>nx10418, A2=>nx10914
   );
   gen_0_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_0_cmp_mReg_3, QB=>
      nx3810, D=>window_0_3, CLK=>start, R=>rst);
   ix97 : nor03_2x port map ( Y=>nx96, A0=>gen_0_cmp_mReg_3, A1=>nx10730, A2
      =>nx10922);
   ix133 : nand02 port map ( Y=>gen_0_cmp_BSCmp_op2_4, A0=>nx3817, A1=>
      nx3823);
   ix3818 : nor02_2x port map ( Y=>nx3817, A0=>nx128, A1=>nx124);
   ix129 : nor03_2x port map ( Y=>nx128, A0=>gen_0_cmp_mReg_3, A1=>nx10424, 
      A2=>nx10890);
   ix125 : nor03_2x port map ( Y=>nx124, A0=>nx3810, A1=>nx10896, A2=>
      nx10906);
   ix3824 : nor02_2x port map ( Y=>nx3823, A0=>nx120, A1=>nx118);
   ix121 : nor03_2x port map ( Y=>nx120, A0=>nx3827, A1=>nx10418, A2=>
      nx10914);
   gen_0_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_0_cmp_mReg_4, QB=>
      nx3827, D=>window_0_4, CLK=>start, R=>rst);
   ix119 : nor03_2x port map ( Y=>nx118, A0=>gen_0_cmp_mReg_4, A1=>nx10730, 
      A2=>nx10922);
   ix155 : nand02 port map ( Y=>gen_0_cmp_BSCmp_op2_5, A0=>nx3831, A1=>
      nx3837);
   ix3832 : nor02_2x port map ( Y=>nx3831, A0=>nx150, A1=>nx146);
   ix151 : nor03_2x port map ( Y=>nx150, A0=>gen_0_cmp_mReg_4, A1=>nx10424, 
      A2=>nx10890);
   ix147 : nor03_2x port map ( Y=>nx146, A0=>nx3827, A1=>nx10896, A2=>
      nx10906);
   ix3838 : nor02_2x port map ( Y=>nx3837, A0=>nx142, A1=>nx140);
   ix143 : nor03_2x port map ( Y=>nx142, A0=>nx3841, A1=>nx10420, A2=>
      nx10914);
   gen_0_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_0_cmp_mReg_5, QB=>
      nx3841, D=>window_0_5, CLK=>start, R=>rst);
   ix141 : nor03_2x port map ( Y=>nx140, A0=>gen_0_cmp_mReg_5, A1=>nx10730, 
      A2=>nx10922);
   ix177 : nand02 port map ( Y=>gen_0_cmp_BSCmp_op2_6, A0=>nx3845, A1=>
      nx3851);
   ix3846 : nor02_2x port map ( Y=>nx3845, A0=>nx172, A1=>nx168);
   ix173 : nor03_2x port map ( Y=>nx172, A0=>gen_0_cmp_mReg_5, A1=>nx10426, 
      A2=>nx10890);
   ix169 : nor03_2x port map ( Y=>nx168, A0=>nx3841, A1=>nx10896, A2=>
      nx10906);
   ix3852 : nor02_2x port map ( Y=>nx3851, A0=>nx164, A1=>nx162);
   ix165 : nor03_2x port map ( Y=>nx164, A0=>nx3855, A1=>nx10420, A2=>
      nx10914);
   gen_0_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_0_cmp_mReg_6, QB=>
      nx3855, D=>window_0_6, CLK=>start, R=>rst);
   ix163 : nor03_2x port map ( Y=>nx162, A0=>gen_0_cmp_mReg_6, A1=>nx10730, 
      A2=>nx10922);
   ix199 : nand02 port map ( Y=>gen_0_cmp_BSCmp_op2_7, A0=>nx3861, A1=>
      nx3867);
   ix3862 : nor02_2x port map ( Y=>nx3861, A0=>nx194, A1=>nx190);
   ix195 : nor03_2x port map ( Y=>nx194, A0=>gen_0_cmp_mReg_6, A1=>nx10426, 
      A2=>nx10892);
   ix191 : nor03_2x port map ( Y=>nx190, A0=>nx3855, A1=>nx10898, A2=>
      nx10908);
   ix3868 : nor02_2x port map ( Y=>nx3867, A0=>nx186, A1=>nx184);
   ix187 : nor03_2x port map ( Y=>nx186, A0=>nx3870, A1=>nx10420, A2=>
      nx10916);
   gen_0_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_0_cmp_mReg_7, QB=>
      nx3870, D=>window_0_7, CLK=>start, R=>rst);
   ix185 : nor03_2x port map ( Y=>nx184, A0=>gen_0_cmp_mReg_7, A1=>nx10730, 
      A2=>nx10924);
   ix221 : nand02 port map ( Y=>gen_0_cmp_BSCmp_op2_8, A0=>nx3874, A1=>
      nx3879);
   ix3875 : nor02_2x port map ( Y=>nx3874, A0=>nx216, A1=>nx212);
   ix217 : nor03_2x port map ( Y=>nx216, A0=>gen_0_cmp_mReg_7, A1=>nx10426, 
      A2=>nx10892);
   ix213 : nor03_2x port map ( Y=>nx212, A0=>nx3870, A1=>nx10898, A2=>
      nx10908);
   ix3880 : nor02_2x port map ( Y=>nx3879, A0=>nx208, A1=>nx206);
   ix209 : nor03_2x port map ( Y=>nx208, A0=>nx3883, A1=>nx10420, A2=>
      nx10916);
   gen_0_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_0_cmp_mReg_8, QB=>
      nx3883, D=>window_0_8, CLK=>start, R=>rst);
   ix207 : nor03_2x port map ( Y=>nx206, A0=>gen_0_cmp_mReg_8, A1=>nx10732, 
      A2=>nx10924);
   ix243 : nand02 port map ( Y=>gen_0_cmp_BSCmp_op2_9, A0=>nx3889, A1=>
      nx3895);
   ix3890 : nor02_2x port map ( Y=>nx3889, A0=>nx238, A1=>nx234);
   ix239 : nor03_2x port map ( Y=>nx238, A0=>gen_0_cmp_mReg_8, A1=>nx10426, 
      A2=>nx10892);
   ix235 : nor03_2x port map ( Y=>nx234, A0=>nx3883, A1=>nx10898, A2=>
      nx10908);
   ix3896 : nor02_2x port map ( Y=>nx3895, A0=>nx230, A1=>nx228);
   ix231 : nor03_2x port map ( Y=>nx230, A0=>nx3899, A1=>nx10420, A2=>
      nx10916);
   gen_0_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_0_cmp_mReg_9, QB=>
      nx3899, D=>window_0_9, CLK=>start, R=>rst);
   ix229 : nor03_2x port map ( Y=>nx228, A0=>gen_0_cmp_mReg_9, A1=>nx10732, 
      A2=>nx10924);
   ix265 : nand02 port map ( Y=>gen_0_cmp_BSCmp_op2_10, A0=>nx3903, A1=>
      nx3909);
   ix3904 : nor02_2x port map ( Y=>nx3903, A0=>nx260, A1=>nx256);
   ix261 : nor03_2x port map ( Y=>nx260, A0=>gen_0_cmp_mReg_9, A1=>nx10426, 
      A2=>nx10892);
   ix257 : nor03_2x port map ( Y=>nx256, A0=>nx3899, A1=>nx10898, A2=>
      nx10908);
   ix3910 : nor02_2x port map ( Y=>nx3909, A0=>nx252, A1=>nx250);
   ix253 : nor03_2x port map ( Y=>nx252, A0=>nx3913, A1=>nx10420, A2=>
      nx10916);
   gen_0_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_0_cmp_mReg_10, QB=>
      nx3913, D=>window_0_10, CLK=>start, R=>rst);
   ix251 : nor03_2x port map ( Y=>nx250, A0=>gen_0_cmp_mReg_10, A1=>nx10732, 
      A2=>nx10924);
   ix287 : nand02 port map ( Y=>gen_0_cmp_BSCmp_op2_11, A0=>nx3919, A1=>
      nx3923);
   ix3920 : nor02_2x port map ( Y=>nx3919, A0=>nx282, A1=>nx278);
   ix283 : nor03_2x port map ( Y=>nx282, A0=>gen_0_cmp_mReg_10, A1=>nx10426, 
      A2=>nx10892);
   ix279 : nor03_2x port map ( Y=>nx278, A0=>nx3913, A1=>nx10898, A2=>
      nx10908);
   ix3924 : nor02_2x port map ( Y=>nx3923, A0=>nx274, A1=>nx272);
   ix275 : nor03_2x port map ( Y=>nx274, A0=>nx3927, A1=>nx10420, A2=>
      nx10916);
   gen_0_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_0_cmp_mReg_11, QB=>
      nx3927, D=>window_0_11, CLK=>start, R=>rst);
   ix273 : nor03_2x port map ( Y=>nx272, A0=>gen_0_cmp_mReg_11, A1=>nx10732, 
      A2=>nx10924);
   ix309 : nand02 port map ( Y=>gen_0_cmp_BSCmp_op2_12, A0=>nx3931, A1=>
      nx3937);
   ix3932 : nor02_2x port map ( Y=>nx3931, A0=>nx304, A1=>nx300);
   ix305 : nor03_2x port map ( Y=>nx304, A0=>gen_0_cmp_mReg_11, A1=>nx10426, 
      A2=>nx10892);
   ix301 : nor03_2x port map ( Y=>nx300, A0=>nx3927, A1=>nx10898, A2=>
      nx10908);
   ix3938 : nor02_2x port map ( Y=>nx3937, A0=>nx296, A1=>nx294);
   ix297 : nor03_2x port map ( Y=>nx296, A0=>nx3941, A1=>nx10422, A2=>
      nx10916);
   gen_0_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_0_cmp_mReg_12, QB=>
      nx3941, D=>window_0_12, CLK=>start, R=>rst);
   ix295 : nor03_2x port map ( Y=>nx294, A0=>gen_0_cmp_mReg_12, A1=>nx10732, 
      A2=>nx10924);
   ix331 : nand02 port map ( Y=>gen_0_cmp_BSCmp_op2_13, A0=>nx3945, A1=>
      nx3951);
   ix3946 : nor02_2x port map ( Y=>nx3945, A0=>nx326, A1=>nx322);
   ix327 : nor03_2x port map ( Y=>nx326, A0=>gen_0_cmp_mReg_12, A1=>nx10428, 
      A2=>nx10894);
   ix323 : nor03_2x port map ( Y=>nx322, A0=>nx3941, A1=>nx10898, A2=>
      nx10910);
   ix3952 : nor02_2x port map ( Y=>nx3951, A0=>nx318, A1=>nx316);
   ix319 : nor03_2x port map ( Y=>nx318, A0=>nx3954, A1=>nx10422, A2=>
      nx10918);
   gen_0_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_0_cmp_mReg_13, QB=>
      nx3954, D=>window_0_13, CLK=>start, R=>rst);
   ix317 : nor03_2x port map ( Y=>nx316, A0=>gen_0_cmp_mReg_13, A1=>nx10732, 
      A2=>nx10926);
   ix353 : nand02 port map ( Y=>gen_0_cmp_BSCmp_op2_14, A0=>nx3961, A1=>
      nx3967);
   ix3962 : nor02_2x port map ( Y=>nx3961, A0=>nx348, A1=>nx344);
   ix349 : nor03_2x port map ( Y=>nx348, A0=>gen_0_cmp_mReg_13, A1=>nx10428, 
      A2=>nx10894);
   ix345 : nor03_2x port map ( Y=>nx344, A0=>nx3954, A1=>nx10900, A2=>
      nx10910);
   ix3968 : nor02_2x port map ( Y=>nx3967, A0=>nx340, A1=>nx338);
   ix341 : nor03_2x port map ( Y=>nx340, A0=>nx3971, A1=>nx10422, A2=>
      nx10918);
   gen_0_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_0_cmp_mReg_14, QB=>
      nx3971, D=>window_0_14, CLK=>start, R=>rst);
   ix339 : nor03_2x port map ( Y=>nx338, A0=>gen_0_cmp_mReg_14, A1=>nx10732, 
      A2=>nx10926);
   ix375 : nand02 port map ( Y=>gen_0_cmp_BSCmp_op2_15, A0=>nx3975, A1=>
      nx3981);
   ix3976 : nor02_2x port map ( Y=>nx3975, A0=>nx370, A1=>nx366);
   ix371 : nor03_2x port map ( Y=>nx370, A0=>gen_0_cmp_mReg_14, A1=>nx10428, 
      A2=>nx10894);
   ix367 : nor03_2x port map ( Y=>nx366, A0=>nx3971, A1=>nx10900, A2=>
      nx10910);
   ix3982 : nor02_2x port map ( Y=>nx3981, A0=>nx362, A1=>nx360);
   ix363 : nor03_2x port map ( Y=>nx362, A0=>nx3985, A1=>nx10422, A2=>
      nx10918);
   gen_0_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_0_cmp_mReg_15, QB=>
      nx3985, D=>window_0_15, CLK=>start, R=>rst);
   ix361 : nor03_2x port map ( Y=>nx360, A0=>gen_0_cmp_mReg_15, A1=>nx10734, 
      A2=>nx10926);
   ix385 : nand02 port map ( Y=>gen_0_cmp_BSCmp_op2_16, A0=>nx3989, A1=>
      nx3981);
   ix3990 : nor02_2x port map ( Y=>nx3989, A0=>nx380, A1=>nx376);
   ix381 : nor03_2x port map ( Y=>nx380, A0=>gen_0_cmp_mReg_15, A1=>nx10428, 
      A2=>nx10894);
   ix377 : nor03_2x port map ( Y=>nx376, A0=>nx3985, A1=>nx10900, A2=>
      nx10910);
   ix453 : nand02 port map ( Y=>gen_1_cmp_BSCmp_op2_1, A0=>nx3996, A1=>
      nx4015);
   ix3997 : nor02_2x port map ( Y=>nx3996, A0=>nx448, A1=>nx444);
   ix449 : nor03_2x port map ( Y=>nx448, A0=>gen_1_cmp_mReg_0, A1=>nx10412, 
      A2=>nx10930);
   gen_1_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_1_cmp_mReg_0, QB=>
      nx4001, D=>window_1_0, CLK=>start, R=>rst);
   ix4006 : inv01 port map ( Y=>nx4005, A=>gen_1_cmp_pMux_0);
   ix445 : nor03_2x port map ( Y=>nx444, A0=>nx4001, A1=>nx10936, A2=>
      nx10946);
   ix4014 : inv02 port map ( Y=>nx4013, A=>gen_1_cmp_pMux_2);
   ix4016 : nor02_2x port map ( Y=>nx4015, A0=>nx434, A1=>nx432);
   ix435 : nor03_2x port map ( Y=>nx434, A0=>nx4018, A1=>nx10406, A2=>
      nx10954);
   gen_1_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_1_cmp_mReg_1, QB=>
      nx4018, D=>window_1_1, CLK=>start, R=>rst);
   ix433 : nor03_2x port map ( Y=>nx432, A0=>gen_1_cmp_mReg_1, A1=>nx10736, 
      A2=>nx10962);
   ix393 : nor03_2x port map ( Y=>nx392, A0=>nx10412, A1=>nx4013, A2=>
      gen_1_cmp_pMux_0);
   ix475 : nand02 port map ( Y=>gen_1_cmp_BSCmp_op2_2, A0=>nx4031, A1=>
      nx4037);
   ix4032 : nor02_2x port map ( Y=>nx4031, A0=>nx470, A1=>nx466);
   ix471 : nor03_2x port map ( Y=>nx470, A0=>gen_1_cmp_mReg_1, A1=>nx10412, 
      A2=>nx10930);
   ix467 : nor03_2x port map ( Y=>nx466, A0=>nx4018, A1=>nx10936, A2=>
      nx10946);
   ix4038 : nor02_2x port map ( Y=>nx4037, A0=>nx462, A1=>nx460);
   ix463 : nor03_2x port map ( Y=>nx462, A0=>nx4040, A1=>nx10406, A2=>
      nx10954);
   gen_1_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_1_cmp_mReg_2, QB=>
      nx4040, D=>window_1_2, CLK=>start, R=>rst);
   ix461 : nor03_2x port map ( Y=>nx460, A0=>gen_1_cmp_mReg_2, A1=>nx10736, 
      A2=>nx10962);
   ix497 : nand02 port map ( Y=>gen_1_cmp_BSCmp_op2_3, A0=>nx4045, A1=>
      nx4051);
   ix4046 : nor02_2x port map ( Y=>nx4045, A0=>nx492, A1=>nx488);
   ix493 : nor03_2x port map ( Y=>nx492, A0=>gen_1_cmp_mReg_2, A1=>nx10412, 
      A2=>nx10930);
   ix489 : nor03_2x port map ( Y=>nx488, A0=>nx4040, A1=>nx10936, A2=>
      nx10946);
   ix4052 : nor02_2x port map ( Y=>nx4051, A0=>nx484, A1=>nx482);
   ix485 : nor03_2x port map ( Y=>nx484, A0=>nx4055, A1=>nx10406, A2=>
      nx10954);
   gen_1_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_1_cmp_mReg_3, QB=>
      nx4055, D=>window_1_3, CLK=>start, R=>rst);
   ix483 : nor03_2x port map ( Y=>nx482, A0=>gen_1_cmp_mReg_3, A1=>nx10736, 
      A2=>nx10962);
   ix519 : nand02 port map ( Y=>gen_1_cmp_BSCmp_op2_4, A0=>nx4061, A1=>
      nx4065);
   ix4062 : nor02_2x port map ( Y=>nx4061, A0=>nx514, A1=>nx510);
   ix515 : nor03_2x port map ( Y=>nx514, A0=>gen_1_cmp_mReg_3, A1=>nx10412, 
      A2=>nx10930);
   ix511 : nor03_2x port map ( Y=>nx510, A0=>nx4055, A1=>nx10936, A2=>
      nx10946);
   ix4066 : nor02_2x port map ( Y=>nx4065, A0=>nx506, A1=>nx504);
   ix507 : nor03_2x port map ( Y=>nx506, A0=>nx4069, A1=>nx10406, A2=>
      nx10954);
   gen_1_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_1_cmp_mReg_4, QB=>
      nx4069, D=>window_1_4, CLK=>start, R=>rst);
   ix505 : nor03_2x port map ( Y=>nx504, A0=>gen_1_cmp_mReg_4, A1=>nx10736, 
      A2=>nx10962);
   ix541 : nand02 port map ( Y=>gen_1_cmp_BSCmp_op2_5, A0=>nx4075, A1=>
      nx4081);
   ix4076 : nor02_2x port map ( Y=>nx4075, A0=>nx536, A1=>nx532);
   ix537 : nor03_2x port map ( Y=>nx536, A0=>gen_1_cmp_mReg_4, A1=>nx10412, 
      A2=>nx10930);
   ix533 : nor03_2x port map ( Y=>nx532, A0=>nx4069, A1=>nx10936, A2=>
      nx10946);
   ix4082 : nor02_2x port map ( Y=>nx4081, A0=>nx528, A1=>nx526);
   ix529 : nor03_2x port map ( Y=>nx528, A0=>nx4084, A1=>nx10408, A2=>
      nx10954);
   gen_1_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_1_cmp_mReg_5, QB=>
      nx4084, D=>window_1_5, CLK=>start, R=>rst);
   ix527 : nor03_2x port map ( Y=>nx526, A0=>gen_1_cmp_mReg_5, A1=>nx10736, 
      A2=>nx10962);
   ix563 : nand02 port map ( Y=>gen_1_cmp_BSCmp_op2_6, A0=>nx4089, A1=>
      nx4095);
   ix4090 : nor02_2x port map ( Y=>nx4089, A0=>nx558, A1=>nx554);
   ix559 : nor03_2x port map ( Y=>nx558, A0=>gen_1_cmp_mReg_5, A1=>nx10414, 
      A2=>nx10930);
   ix555 : nor03_2x port map ( Y=>nx554, A0=>nx4084, A1=>nx10936, A2=>
      nx10946);
   ix4096 : nor02_2x port map ( Y=>nx4095, A0=>nx550, A1=>nx548);
   ix551 : nor03_2x port map ( Y=>nx550, A0=>nx4099, A1=>nx10408, A2=>
      nx10954);
   gen_1_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_1_cmp_mReg_6, QB=>
      nx4099, D=>window_1_6, CLK=>start, R=>rst);
   ix549 : nor03_2x port map ( Y=>nx548, A0=>gen_1_cmp_mReg_6, A1=>nx10736, 
      A2=>nx10962);
   ix585 : nand02 port map ( Y=>gen_1_cmp_BSCmp_op2_7, A0=>nx4105, A1=>
      nx4109);
   ix4106 : nor02_2x port map ( Y=>nx4105, A0=>nx580, A1=>nx576);
   ix581 : nor03_2x port map ( Y=>nx580, A0=>gen_1_cmp_mReg_6, A1=>nx10414, 
      A2=>nx10932);
   ix577 : nor03_2x port map ( Y=>nx576, A0=>nx4099, A1=>nx10938, A2=>
      nx10948);
   ix4110 : nor02_2x port map ( Y=>nx4109, A0=>nx572, A1=>nx570);
   ix573 : nor03_2x port map ( Y=>nx572, A0=>nx4113, A1=>nx10408, A2=>
      nx10956);
   gen_1_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_1_cmp_mReg_7, QB=>
      nx4113, D=>window_1_7, CLK=>start, R=>rst);
   ix571 : nor03_2x port map ( Y=>nx570, A0=>gen_1_cmp_mReg_7, A1=>nx10736, 
      A2=>nx10964);
   ix607 : nand02 port map ( Y=>gen_1_cmp_BSCmp_op2_8, A0=>nx4119, A1=>
      nx4125);
   ix4120 : nor02_2x port map ( Y=>nx4119, A0=>nx602, A1=>nx598);
   ix603 : nor03_2x port map ( Y=>nx602, A0=>gen_1_cmp_mReg_7, A1=>nx10414, 
      A2=>nx10932);
   ix599 : nor03_2x port map ( Y=>nx598, A0=>nx4113, A1=>nx10938, A2=>
      nx10948);
   ix4126 : nor02_2x port map ( Y=>nx4125, A0=>nx594, A1=>nx592);
   ix595 : nor03_2x port map ( Y=>nx594, A0=>nx4128, A1=>nx10408, A2=>
      nx10956);
   gen_1_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_1_cmp_mReg_8, QB=>
      nx4128, D=>window_1_8, CLK=>start, R=>rst);
   ix593 : nor03_2x port map ( Y=>nx592, A0=>gen_1_cmp_mReg_8, A1=>nx10738, 
      A2=>nx10964);
   ix629 : nand02 port map ( Y=>gen_1_cmp_BSCmp_op2_9, A0=>nx4133, A1=>
      nx4139);
   ix4134 : nor02_2x port map ( Y=>nx4133, A0=>nx624, A1=>nx620);
   ix625 : nor03_2x port map ( Y=>nx624, A0=>gen_1_cmp_mReg_8, A1=>nx10414, 
      A2=>nx10932);
   ix621 : nor03_2x port map ( Y=>nx620, A0=>nx4128, A1=>nx10938, A2=>
      nx10948);
   ix4140 : nor02_2x port map ( Y=>nx4139, A0=>nx616, A1=>nx614);
   ix617 : nor03_2x port map ( Y=>nx616, A0=>nx4143, A1=>nx10408, A2=>
      nx10956);
   gen_1_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_1_cmp_mReg_9, QB=>
      nx4143, D=>window_1_9, CLK=>start, R=>rst);
   ix615 : nor03_2x port map ( Y=>nx614, A0=>gen_1_cmp_mReg_9, A1=>nx10738, 
      A2=>nx10964);
   ix651 : nand02 port map ( Y=>gen_1_cmp_BSCmp_op2_10, A0=>nx4149, A1=>
      nx4153);
   ix4150 : nor02_2x port map ( Y=>nx4149, A0=>nx646, A1=>nx642);
   ix647 : nor03_2x port map ( Y=>nx646, A0=>gen_1_cmp_mReg_9, A1=>nx10414, 
      A2=>nx10932);
   ix643 : nor03_2x port map ( Y=>nx642, A0=>nx4143, A1=>nx10938, A2=>
      nx10948);
   ix4154 : nor02_2x port map ( Y=>nx4153, A0=>nx638, A1=>nx636);
   ix639 : nor03_2x port map ( Y=>nx638, A0=>nx4157, A1=>nx10408, A2=>
      nx10956);
   gen_1_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_1_cmp_mReg_10, QB=>
      nx4157, D=>window_1_10, CLK=>start, R=>rst);
   ix637 : nor03_2x port map ( Y=>nx636, A0=>gen_1_cmp_mReg_10, A1=>nx10738, 
      A2=>nx10964);
   ix673 : nand02 port map ( Y=>gen_1_cmp_BSCmp_op2_11, A0=>nx4163, A1=>
      nx4169);
   ix4164 : nor02_2x port map ( Y=>nx4163, A0=>nx668, A1=>nx664);
   ix669 : nor03_2x port map ( Y=>nx668, A0=>gen_1_cmp_mReg_10, A1=>nx10414, 
      A2=>nx10932);
   ix665 : nor03_2x port map ( Y=>nx664, A0=>nx4157, A1=>nx10938, A2=>
      nx10948);
   ix4170 : nor02_2x port map ( Y=>nx4169, A0=>nx660, A1=>nx658);
   ix661 : nor03_2x port map ( Y=>nx660, A0=>nx4172, A1=>nx10408, A2=>
      nx10956);
   gen_1_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_1_cmp_mReg_11, QB=>
      nx4172, D=>window_1_11, CLK=>start, R=>rst);
   ix659 : nor03_2x port map ( Y=>nx658, A0=>gen_1_cmp_mReg_11, A1=>nx10738, 
      A2=>nx10964);
   ix695 : nand02 port map ( Y=>gen_1_cmp_BSCmp_op2_12, A0=>nx4177, A1=>
      nx4183);
   ix4178 : nor02_2x port map ( Y=>nx4177, A0=>nx690, A1=>nx686);
   ix691 : nor03_2x port map ( Y=>nx690, A0=>gen_1_cmp_mReg_11, A1=>nx10414, 
      A2=>nx10932);
   ix687 : nor03_2x port map ( Y=>nx686, A0=>nx4172, A1=>nx10938, A2=>
      nx10948);
   ix4184 : nor02_2x port map ( Y=>nx4183, A0=>nx682, A1=>nx680);
   ix683 : nor03_2x port map ( Y=>nx682, A0=>nx4187, A1=>nx10410, A2=>
      nx10956);
   gen_1_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_1_cmp_mReg_12, QB=>
      nx4187, D=>window_1_12, CLK=>start, R=>rst);
   ix681 : nor03_2x port map ( Y=>nx680, A0=>gen_1_cmp_mReg_12, A1=>nx10738, 
      A2=>nx10964);
   ix717 : nand02 port map ( Y=>gen_1_cmp_BSCmp_op2_13, A0=>nx4193, A1=>
      nx4197);
   ix4194 : nor02_2x port map ( Y=>nx4193, A0=>nx712, A1=>nx708);
   ix713 : nor03_2x port map ( Y=>nx712, A0=>gen_1_cmp_mReg_12, A1=>nx10416, 
      A2=>nx10934);
   ix709 : nor03_2x port map ( Y=>nx708, A0=>nx4187, A1=>nx10938, A2=>
      nx10950);
   ix4198 : nor02_2x port map ( Y=>nx4197, A0=>nx704, A1=>nx702);
   ix705 : nor03_2x port map ( Y=>nx704, A0=>nx4201, A1=>nx10410, A2=>
      nx10958);
   gen_1_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_1_cmp_mReg_13, QB=>
      nx4201, D=>window_1_13, CLK=>start, R=>rst);
   ix703 : nor03_2x port map ( Y=>nx702, A0=>gen_1_cmp_mReg_13, A1=>nx10738, 
      A2=>nx10966);
   ix739 : nand02 port map ( Y=>gen_1_cmp_BSCmp_op2_14, A0=>nx4207, A1=>
      nx4213);
   ix4208 : nor02_2x port map ( Y=>nx4207, A0=>nx734, A1=>nx730);
   ix735 : nor03_2x port map ( Y=>nx734, A0=>gen_1_cmp_mReg_13, A1=>nx10416, 
      A2=>nx10934);
   ix731 : nor03_2x port map ( Y=>nx730, A0=>nx4201, A1=>nx10940, A2=>
      nx10950);
   ix4214 : nor02_2x port map ( Y=>nx4213, A0=>nx726, A1=>nx724);
   ix727 : nor03_2x port map ( Y=>nx726, A0=>nx4216, A1=>nx10410, A2=>
      nx10958);
   gen_1_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_1_cmp_mReg_14, QB=>
      nx4216, D=>window_1_14, CLK=>start, R=>rst);
   ix725 : nor03_2x port map ( Y=>nx724, A0=>gen_1_cmp_mReg_14, A1=>nx10738, 
      A2=>nx10966);
   ix761 : nand02 port map ( Y=>gen_1_cmp_BSCmp_op2_15, A0=>nx4221, A1=>
      nx4227);
   ix4222 : nor02_2x port map ( Y=>nx4221, A0=>nx756, A1=>nx752);
   ix757 : nor03_2x port map ( Y=>nx756, A0=>gen_1_cmp_mReg_14, A1=>nx10416, 
      A2=>nx10934);
   ix753 : nor03_2x port map ( Y=>nx752, A0=>nx4216, A1=>nx10940, A2=>
      nx10950);
   ix4228 : nor02_2x port map ( Y=>nx4227, A0=>nx748, A1=>nx746);
   ix749 : nor03_2x port map ( Y=>nx748, A0=>nx4231, A1=>nx10410, A2=>
      nx10958);
   gen_1_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_1_cmp_mReg_15, QB=>
      nx4231, D=>window_1_15, CLK=>start, R=>rst);
   ix747 : nor03_2x port map ( Y=>nx746, A0=>gen_1_cmp_mReg_15, A1=>nx10740, 
      A2=>nx10966);
   ix771 : nand02 port map ( Y=>gen_1_cmp_BSCmp_op2_16, A0=>nx4237, A1=>
      nx4227);
   ix4238 : nor02_2x port map ( Y=>nx4237, A0=>nx766, A1=>nx762);
   ix767 : nor03_2x port map ( Y=>nx766, A0=>gen_1_cmp_mReg_15, A1=>nx10416, 
      A2=>nx10934);
   ix763 : nor03_2x port map ( Y=>nx762, A0=>nx4231, A1=>nx10940, A2=>
      nx10950);
   ix839 : nand02 port map ( Y=>gen_2_cmp_BSCmp_op2_1, A0=>nx4243, A1=>
      nx4263);
   ix4244 : nor02_2x port map ( Y=>nx4243, A0=>nx834, A1=>nx830);
   ix835 : nor03_2x port map ( Y=>nx834, A0=>gen_2_cmp_mReg_0, A1=>nx10400, 
      A2=>nx10970);
   gen_2_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_2_cmp_mReg_0, QB=>
      nx4249, D=>window_2_0, CLK=>start, R=>rst);
   ix4254 : inv01 port map ( Y=>nx4253, A=>gen_2_cmp_pMux_0);
   ix831 : nor03_2x port map ( Y=>nx830, A0=>nx4249, A1=>nx10976, A2=>
      nx10986);
   ix4261 : inv02 port map ( Y=>nx4260, A=>gen_2_cmp_pMux_2);
   ix4264 : nor02_2x port map ( Y=>nx4263, A0=>nx820, A1=>nx818);
   ix821 : nor03_2x port map ( Y=>nx820, A0=>nx4267, A1=>nx10394, A2=>
      nx10994);
   gen_2_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_2_cmp_mReg_1, QB=>
      nx4267, D=>window_2_1, CLK=>start, R=>rst);
   ix819 : nor03_2x port map ( Y=>nx818, A0=>gen_2_cmp_mReg_1, A1=>nx10742, 
      A2=>nx11002);
   ix779 : nor03_2x port map ( Y=>nx778, A0=>nx10400, A1=>nx4260, A2=>
      gen_2_cmp_pMux_0);
   ix861 : nand02 port map ( Y=>gen_2_cmp_BSCmp_op2_2, A0=>nx4279, A1=>
      nx4285);
   ix4280 : nor02_2x port map ( Y=>nx4279, A0=>nx856, A1=>nx852);
   ix857 : nor03_2x port map ( Y=>nx856, A0=>gen_2_cmp_mReg_1, A1=>nx10400, 
      A2=>nx10970);
   ix853 : nor03_2x port map ( Y=>nx852, A0=>nx4267, A1=>nx10976, A2=>
      nx10986);
   ix4286 : nor02_2x port map ( Y=>nx4285, A0=>nx848, A1=>nx846);
   ix849 : nor03_2x port map ( Y=>nx848, A0=>nx4288, A1=>nx10394, A2=>
      nx10994);
   gen_2_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_2_cmp_mReg_2, QB=>
      nx4288, D=>window_2_2, CLK=>start, R=>rst);
   ix847 : nor03_2x port map ( Y=>nx846, A0=>gen_2_cmp_mReg_2, A1=>nx10742, 
      A2=>nx11002);
   ix883 : nand02 port map ( Y=>gen_2_cmp_BSCmp_op2_3, A0=>nx4293, A1=>
      nx4299);
   ix4294 : nor02_2x port map ( Y=>nx4293, A0=>nx878, A1=>nx874);
   ix879 : nor03_2x port map ( Y=>nx878, A0=>gen_2_cmp_mReg_2, A1=>nx10400, 
      A2=>nx10970);
   ix875 : nor03_2x port map ( Y=>nx874, A0=>nx4288, A1=>nx10976, A2=>
      nx10986);
   ix4300 : nor02_2x port map ( Y=>nx4299, A0=>nx870, A1=>nx868);
   ix871 : nor03_2x port map ( Y=>nx870, A0=>nx4303, A1=>nx10394, A2=>
      nx10994);
   gen_2_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_2_cmp_mReg_3, QB=>
      nx4303, D=>window_2_3, CLK=>start, R=>rst);
   ix869 : nor03_2x port map ( Y=>nx868, A0=>gen_2_cmp_mReg_3, A1=>nx10742, 
      A2=>nx11002);
   ix905 : nand02 port map ( Y=>gen_2_cmp_BSCmp_op2_4, A0=>nx4309, A1=>
      nx4315);
   ix4310 : nor02_2x port map ( Y=>nx4309, A0=>nx900, A1=>nx896);
   ix901 : nor03_2x port map ( Y=>nx900, A0=>gen_2_cmp_mReg_3, A1=>nx10400, 
      A2=>nx10970);
   ix897 : nor03_2x port map ( Y=>nx896, A0=>nx4303, A1=>nx10976, A2=>
      nx10986);
   ix4316 : nor02_2x port map ( Y=>nx4315, A0=>nx892, A1=>nx890);
   ix893 : nor03_2x port map ( Y=>nx892, A0=>nx4318, A1=>nx10394, A2=>
      nx10994);
   gen_2_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_2_cmp_mReg_4, QB=>
      nx4318, D=>window_2_4, CLK=>start, R=>rst);
   ix891 : nor03_2x port map ( Y=>nx890, A0=>gen_2_cmp_mReg_4, A1=>nx10742, 
      A2=>nx11002);
   ix927 : nand02 port map ( Y=>gen_2_cmp_BSCmp_op2_5, A0=>nx4325, A1=>
      nx4331);
   ix4326 : nor02_2x port map ( Y=>nx4325, A0=>nx922, A1=>nx918);
   ix923 : nor03_2x port map ( Y=>nx922, A0=>gen_2_cmp_mReg_4, A1=>nx10400, 
      A2=>nx10970);
   ix919 : nor03_2x port map ( Y=>nx918, A0=>nx4318, A1=>nx10976, A2=>
      nx10986);
   ix4332 : nor02_2x port map ( Y=>nx4331, A0=>nx914, A1=>nx912);
   ix915 : nor03_2x port map ( Y=>nx914, A0=>nx4335, A1=>nx10396, A2=>
      nx10994);
   gen_2_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_2_cmp_mReg_5, QB=>
      nx4335, D=>window_2_5, CLK=>start, R=>rst);
   ix913 : nor03_2x port map ( Y=>nx912, A0=>gen_2_cmp_mReg_5, A1=>nx10742, 
      A2=>nx11002);
   ix949 : nand02 port map ( Y=>gen_2_cmp_BSCmp_op2_6, A0=>nx4339, A1=>
      nx4345);
   ix4340 : nor02_2x port map ( Y=>nx4339, A0=>nx944, A1=>nx940);
   ix945 : nor03_2x port map ( Y=>nx944, A0=>gen_2_cmp_mReg_5, A1=>nx10402, 
      A2=>nx10970);
   ix941 : nor03_2x port map ( Y=>nx940, A0=>nx4335, A1=>nx10976, A2=>
      nx10986);
   ix4346 : nor02_2x port map ( Y=>nx4345, A0=>nx936, A1=>nx934);
   ix937 : nor03_2x port map ( Y=>nx936, A0=>nx4349, A1=>nx10396, A2=>
      nx10994);
   gen_2_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_2_cmp_mReg_6, QB=>
      nx4349, D=>window_2_6, CLK=>start, R=>rst);
   ix935 : nor03_2x port map ( Y=>nx934, A0=>gen_2_cmp_mReg_6, A1=>nx10742, 
      A2=>nx11002);
   ix971 : nand02 port map ( Y=>gen_2_cmp_BSCmp_op2_7, A0=>nx4353, A1=>
      nx4359);
   ix4354 : nor02_2x port map ( Y=>nx4353, A0=>nx966, A1=>nx962);
   ix967 : nor03_2x port map ( Y=>nx966, A0=>gen_2_cmp_mReg_6, A1=>nx10402, 
      A2=>nx10972);
   ix963 : nor03_2x port map ( Y=>nx962, A0=>nx4349, A1=>nx10978, A2=>
      nx10988);
   ix4360 : nor02_2x port map ( Y=>nx4359, A0=>nx958, A1=>nx956);
   ix959 : nor03_2x port map ( Y=>nx958, A0=>nx4362, A1=>nx10396, A2=>
      nx10996);
   gen_2_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_2_cmp_mReg_7, QB=>
      nx4362, D=>window_2_7, CLK=>start, R=>rst);
   ix957 : nor03_2x port map ( Y=>nx956, A0=>gen_2_cmp_mReg_7, A1=>nx10742, 
      A2=>nx11004);
   ix993 : nand02 port map ( Y=>gen_2_cmp_BSCmp_op2_8, A0=>nx4369, A1=>
      nx4375);
   ix4370 : nor02_2x port map ( Y=>nx4369, A0=>nx988, A1=>nx984);
   ix989 : nor03_2x port map ( Y=>nx988, A0=>gen_2_cmp_mReg_7, A1=>nx10402, 
      A2=>nx10972);
   ix985 : nor03_2x port map ( Y=>nx984, A0=>nx4362, A1=>nx10978, A2=>
      nx10988);
   ix4376 : nor02_2x port map ( Y=>nx4375, A0=>nx980, A1=>nx978);
   ix981 : nor03_2x port map ( Y=>nx980, A0=>nx4379, A1=>nx10396, A2=>
      nx10996);
   gen_2_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_2_cmp_mReg_8, QB=>
      nx4379, D=>window_2_8, CLK=>start, R=>rst);
   ix979 : nor03_2x port map ( Y=>nx978, A0=>gen_2_cmp_mReg_8, A1=>nx10744, 
      A2=>nx11004);
   ix1015 : nand02 port map ( Y=>gen_2_cmp_BSCmp_op2_9, A0=>nx4383, A1=>
      nx4389);
   ix4384 : nor02_2x port map ( Y=>nx4383, A0=>nx1010, A1=>nx1006);
   ix1011 : nor03_2x port map ( Y=>nx1010, A0=>gen_2_cmp_mReg_8, A1=>nx10402, 
      A2=>nx10972);
   ix1007 : nor03_2x port map ( Y=>nx1006, A0=>nx4379, A1=>nx10978, A2=>
      nx10988);
   ix4390 : nor02_2x port map ( Y=>nx4389, A0=>nx1002, A1=>nx1000);
   ix1003 : nor03_2x port map ( Y=>nx1002, A0=>nx4393, A1=>nx10396, A2=>
      nx10996);
   gen_2_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_2_cmp_mReg_9, QB=>
      nx4393, D=>window_2_9, CLK=>start, R=>rst);
   ix1001 : nor03_2x port map ( Y=>nx1000, A0=>gen_2_cmp_mReg_9, A1=>nx10744, 
      A2=>nx11004);
   ix1037 : nand02 port map ( Y=>gen_2_cmp_BSCmp_op2_10, A0=>nx4397, A1=>
      nx4403);
   ix4398 : nor02_2x port map ( Y=>nx4397, A0=>nx1032, A1=>nx1028);
   ix1033 : nor03_2x port map ( Y=>nx1032, A0=>gen_2_cmp_mReg_9, A1=>nx10402, 
      A2=>nx10972);
   ix1029 : nor03_2x port map ( Y=>nx1028, A0=>nx4393, A1=>nx10978, A2=>
      nx10988);
   ix4404 : nor02_2x port map ( Y=>nx4403, A0=>nx1024, A1=>nx1022);
   ix1025 : nor03_2x port map ( Y=>nx1024, A0=>nx4406, A1=>nx10396, A2=>
      nx10996);
   gen_2_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_2_cmp_mReg_10, QB=>
      nx4406, D=>window_2_10, CLK=>start, R=>rst);
   ix1023 : nor03_2x port map ( Y=>nx1022, A0=>gen_2_cmp_mReg_10, A1=>
      nx10744, A2=>nx11004);
   ix1059 : nand02 port map ( Y=>gen_2_cmp_BSCmp_op2_11, A0=>nx4413, A1=>
      nx4419);
   ix4414 : nor02_2x port map ( Y=>nx4413, A0=>nx1054, A1=>nx1050);
   ix1055 : nor03_2x port map ( Y=>nx1054, A0=>gen_2_cmp_mReg_10, A1=>
      nx10402, A2=>nx10972);
   ix1051 : nor03_2x port map ( Y=>nx1050, A0=>nx4406, A1=>nx10978, A2=>
      nx10988);
   ix4420 : nor02_2x port map ( Y=>nx4419, A0=>nx1046, A1=>nx1044);
   ix1047 : nor03_2x port map ( Y=>nx1046, A0=>nx4423, A1=>nx10396, A2=>
      nx10996);
   gen_2_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_2_cmp_mReg_11, QB=>
      nx4423, D=>window_2_11, CLK=>start, R=>rst);
   ix1045 : nor03_2x port map ( Y=>nx1044, A0=>gen_2_cmp_mReg_11, A1=>
      nx10744, A2=>nx11004);
   ix1081 : nand02 port map ( Y=>gen_2_cmp_BSCmp_op2_12, A0=>nx4427, A1=>
      nx4433);
   ix4428 : nor02_2x port map ( Y=>nx4427, A0=>nx1076, A1=>nx1072);
   ix1077 : nor03_2x port map ( Y=>nx1076, A0=>gen_2_cmp_mReg_11, A1=>
      nx10402, A2=>nx10972);
   ix1073 : nor03_2x port map ( Y=>nx1072, A0=>nx4423, A1=>nx10978, A2=>
      nx10988);
   ix4434 : nor02_2x port map ( Y=>nx4433, A0=>nx1068, A1=>nx1066);
   ix1069 : nor03_2x port map ( Y=>nx1068, A0=>nx4437, A1=>nx10398, A2=>
      nx10996);
   gen_2_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_2_cmp_mReg_12, QB=>
      nx4437, D=>window_2_12, CLK=>start, R=>rst);
   ix1067 : nor03_2x port map ( Y=>nx1066, A0=>gen_2_cmp_mReg_12, A1=>
      nx10744, A2=>nx11004);
   ix1103 : nand02 port map ( Y=>gen_2_cmp_BSCmp_op2_13, A0=>nx4441, A1=>
      nx4447);
   ix4442 : nor02_2x port map ( Y=>nx4441, A0=>nx1098, A1=>nx1094);
   ix1099 : nor03_2x port map ( Y=>nx1098, A0=>gen_2_cmp_mReg_12, A1=>
      nx10404, A2=>nx10974);
   ix1095 : nor03_2x port map ( Y=>nx1094, A0=>nx4437, A1=>nx10978, A2=>
      nx10990);
   ix4448 : nor02_2x port map ( Y=>nx4447, A0=>nx1090, A1=>nx1088);
   ix1091 : nor03_2x port map ( Y=>nx1090, A0=>nx4450, A1=>nx10398, A2=>
      nx10998);
   gen_2_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_2_cmp_mReg_13, QB=>
      nx4450, D=>window_2_13, CLK=>start, R=>rst);
   ix1089 : nor03_2x port map ( Y=>nx1088, A0=>gen_2_cmp_mReg_13, A1=>
      nx10744, A2=>nx11006);
   ix1125 : nand02 port map ( Y=>gen_2_cmp_BSCmp_op2_14, A0=>nx4457, A1=>
      nx4463);
   ix4458 : nor02_2x port map ( Y=>nx4457, A0=>nx1120, A1=>nx1116);
   ix1121 : nor03_2x port map ( Y=>nx1120, A0=>gen_2_cmp_mReg_13, A1=>
      nx10404, A2=>nx10974);
   ix1117 : nor03_2x port map ( Y=>nx1116, A0=>nx4450, A1=>nx10980, A2=>
      nx10990);
   ix4464 : nor02_2x port map ( Y=>nx4463, A0=>nx1112, A1=>nx1110);
   ix1113 : nor03_2x port map ( Y=>nx1112, A0=>nx4467, A1=>nx10398, A2=>
      nx10998);
   gen_2_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_2_cmp_mReg_14, QB=>
      nx4467, D=>window_2_14, CLK=>start, R=>rst);
   ix1111 : nor03_2x port map ( Y=>nx1110, A0=>gen_2_cmp_mReg_14, A1=>
      nx10744, A2=>nx11006);
   ix1147 : nand02 port map ( Y=>gen_2_cmp_BSCmp_op2_15, A0=>nx4471, A1=>
      nx4477);
   ix4472 : nor02_2x port map ( Y=>nx4471, A0=>nx1142, A1=>nx1138);
   ix1143 : nor03_2x port map ( Y=>nx1142, A0=>gen_2_cmp_mReg_14, A1=>
      nx10404, A2=>nx10974);
   ix1139 : nor03_2x port map ( Y=>nx1138, A0=>nx4467, A1=>nx10980, A2=>
      nx10990);
   ix4478 : nor02_2x port map ( Y=>nx4477, A0=>nx1134, A1=>nx1132);
   ix1135 : nor03_2x port map ( Y=>nx1134, A0=>nx4481, A1=>nx10398, A2=>
      nx10998);
   gen_2_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_2_cmp_mReg_15, QB=>
      nx4481, D=>window_2_15, CLK=>start, R=>rst);
   ix1133 : nor03_2x port map ( Y=>nx1132, A0=>gen_2_cmp_mReg_15, A1=>
      nx10746, A2=>nx11006);
   ix1157 : nand02 port map ( Y=>gen_2_cmp_BSCmp_op2_16, A0=>nx4485, A1=>
      nx4477);
   ix4486 : nor02_2x port map ( Y=>nx4485, A0=>nx1152, A1=>nx1148);
   ix1153 : nor03_2x port map ( Y=>nx1152, A0=>gen_2_cmp_mReg_15, A1=>
      nx10404, A2=>nx10974);
   ix1149 : nor03_2x port map ( Y=>nx1148, A0=>nx4481, A1=>nx10980, A2=>
      nx10990);
   ix1225 : nand02 port map ( Y=>gen_3_cmp_BSCmp_op2_1, A0=>nx4492, A1=>
      nx4511);
   ix4493 : nor02_2x port map ( Y=>nx4492, A0=>nx1220, A1=>nx1216);
   ix1221 : nor03_2x port map ( Y=>nx1220, A0=>gen_3_cmp_mReg_0, A1=>nx10388, 
      A2=>nx11010);
   gen_3_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_3_cmp_mReg_0, QB=>
      nx4497, D=>window_3_0, CLK=>start, R=>rst);
   ix4502 : inv01 port map ( Y=>nx4501, A=>gen_3_cmp_pMux_0);
   ix1217 : nor03_2x port map ( Y=>nx1216, A0=>nx4497, A1=>nx11016, A2=>
      nx11026);
   ix4510 : inv02 port map ( Y=>nx4509, A=>gen_3_cmp_pMux_2);
   ix4512 : nor02_2x port map ( Y=>nx4511, A0=>nx1206, A1=>nx1204);
   ix1207 : nor03_2x port map ( Y=>nx1206, A0=>nx4514, A1=>nx10382, A2=>
      nx11034);
   gen_3_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_3_cmp_mReg_1, QB=>
      nx4514, D=>window_3_1, CLK=>start, R=>rst);
   ix1205 : nor03_2x port map ( Y=>nx1204, A0=>gen_3_cmp_mReg_1, A1=>nx10748, 
      A2=>nx11042);
   ix1165 : nor03_2x port map ( Y=>nx1164, A0=>nx10388, A1=>nx4509, A2=>
      gen_3_cmp_pMux_0);
   ix1247 : nand02 port map ( Y=>gen_3_cmp_BSCmp_op2_2, A0=>nx4527, A1=>
      nx4533);
   ix4528 : nor02_2x port map ( Y=>nx4527, A0=>nx1242, A1=>nx1238);
   ix1243 : nor03_2x port map ( Y=>nx1242, A0=>gen_3_cmp_mReg_1, A1=>nx10388, 
      A2=>nx11010);
   ix1239 : nor03_2x port map ( Y=>nx1238, A0=>nx4514, A1=>nx11016, A2=>
      nx11026);
   ix4534 : nor02_2x port map ( Y=>nx4533, A0=>nx1234, A1=>nx1232);
   ix1235 : nor03_2x port map ( Y=>nx1234, A0=>nx4536, A1=>nx10382, A2=>
      nx11034);
   gen_3_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_3_cmp_mReg_2, QB=>
      nx4536, D=>window_3_2, CLK=>start, R=>rst);
   ix1233 : nor03_2x port map ( Y=>nx1232, A0=>gen_3_cmp_mReg_2, A1=>nx10748, 
      A2=>nx11042);
   ix1269 : nand02 port map ( Y=>gen_3_cmp_BSCmp_op2_3, A0=>nx4541, A1=>
      nx4547);
   ix4542 : nor02_2x port map ( Y=>nx4541, A0=>nx1264, A1=>nx1260);
   ix1265 : nor03_2x port map ( Y=>nx1264, A0=>gen_3_cmp_mReg_2, A1=>nx10388, 
      A2=>nx11010);
   ix1261 : nor03_2x port map ( Y=>nx1260, A0=>nx4536, A1=>nx11016, A2=>
      nx11026);
   ix4548 : nor02_2x port map ( Y=>nx4547, A0=>nx1256, A1=>nx1254);
   ix1257 : nor03_2x port map ( Y=>nx1256, A0=>nx4551, A1=>nx10382, A2=>
      nx11034);
   gen_3_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_3_cmp_mReg_3, QB=>
      nx4551, D=>window_3_3, CLK=>start, R=>rst);
   ix1255 : nor03_2x port map ( Y=>nx1254, A0=>gen_3_cmp_mReg_3, A1=>nx10748, 
      A2=>nx11042);
   ix1291 : nand02 port map ( Y=>gen_3_cmp_BSCmp_op2_4, A0=>nx4557, A1=>
      nx4561);
   ix4558 : nor02_2x port map ( Y=>nx4557, A0=>nx1286, A1=>nx1282);
   ix1287 : nor03_2x port map ( Y=>nx1286, A0=>gen_3_cmp_mReg_3, A1=>nx10388, 
      A2=>nx11010);
   ix1283 : nor03_2x port map ( Y=>nx1282, A0=>nx4551, A1=>nx11016, A2=>
      nx11026);
   ix4562 : nor02_2x port map ( Y=>nx4561, A0=>nx1278, A1=>nx1276);
   ix1279 : nor03_2x port map ( Y=>nx1278, A0=>nx4565, A1=>nx10382, A2=>
      nx11034);
   gen_3_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_3_cmp_mReg_4, QB=>
      nx4565, D=>window_3_4, CLK=>start, R=>rst);
   ix1277 : nor03_2x port map ( Y=>nx1276, A0=>gen_3_cmp_mReg_4, A1=>nx10748, 
      A2=>nx11042);
   ix1313 : nand02 port map ( Y=>gen_3_cmp_BSCmp_op2_5, A0=>nx4571, A1=>
      nx4577);
   ix4572 : nor02_2x port map ( Y=>nx4571, A0=>nx1308, A1=>nx1304);
   ix1309 : nor03_2x port map ( Y=>nx1308, A0=>gen_3_cmp_mReg_4, A1=>nx10388, 
      A2=>nx11010);
   ix1305 : nor03_2x port map ( Y=>nx1304, A0=>nx4565, A1=>nx11016, A2=>
      nx11026);
   ix4578 : nor02_2x port map ( Y=>nx4577, A0=>nx1300, A1=>nx1298);
   ix1301 : nor03_2x port map ( Y=>nx1300, A0=>nx4580, A1=>nx10384, A2=>
      nx11034);
   gen_3_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_3_cmp_mReg_5, QB=>
      nx4580, D=>window_3_5, CLK=>start, R=>rst);
   ix1299 : nor03_2x port map ( Y=>nx1298, A0=>gen_3_cmp_mReg_5, A1=>nx10748, 
      A2=>nx11042);
   ix1335 : nand02 port map ( Y=>gen_3_cmp_BSCmp_op2_6, A0=>nx4585, A1=>
      nx4591);
   ix4586 : nor02_2x port map ( Y=>nx4585, A0=>nx1330, A1=>nx1326);
   ix1331 : nor03_2x port map ( Y=>nx1330, A0=>gen_3_cmp_mReg_5, A1=>nx10390, 
      A2=>nx11010);
   ix1327 : nor03_2x port map ( Y=>nx1326, A0=>nx4580, A1=>nx11016, A2=>
      nx11026);
   ix4592 : nor02_2x port map ( Y=>nx4591, A0=>nx1322, A1=>nx1320);
   ix1323 : nor03_2x port map ( Y=>nx1322, A0=>nx4595, A1=>nx10384, A2=>
      nx11034);
   gen_3_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_3_cmp_mReg_6, QB=>
      nx4595, D=>window_3_6, CLK=>start, R=>rst);
   ix1321 : nor03_2x port map ( Y=>nx1320, A0=>gen_3_cmp_mReg_6, A1=>nx10748, 
      A2=>nx11042);
   ix1357 : nand02 port map ( Y=>gen_3_cmp_BSCmp_op2_7, A0=>nx4601, A1=>
      nx4605);
   ix4602 : nor02_2x port map ( Y=>nx4601, A0=>nx1352, A1=>nx1348);
   ix1353 : nor03_2x port map ( Y=>nx1352, A0=>gen_3_cmp_mReg_6, A1=>nx10390, 
      A2=>nx11012);
   ix1349 : nor03_2x port map ( Y=>nx1348, A0=>nx4595, A1=>nx11018, A2=>
      nx11028);
   ix4606 : nor02_2x port map ( Y=>nx4605, A0=>nx1344, A1=>nx1342);
   ix1345 : nor03_2x port map ( Y=>nx1344, A0=>nx4609, A1=>nx10384, A2=>
      nx11036);
   gen_3_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_3_cmp_mReg_7, QB=>
      nx4609, D=>window_3_7, CLK=>start, R=>rst);
   ix1343 : nor03_2x port map ( Y=>nx1342, A0=>gen_3_cmp_mReg_7, A1=>nx10748, 
      A2=>nx11044);
   ix1379 : nand02 port map ( Y=>gen_3_cmp_BSCmp_op2_8, A0=>nx4615, A1=>
      nx4621);
   ix4616 : nor02_2x port map ( Y=>nx4615, A0=>nx1374, A1=>nx1370);
   ix1375 : nor03_2x port map ( Y=>nx1374, A0=>gen_3_cmp_mReg_7, A1=>nx10390, 
      A2=>nx11012);
   ix1371 : nor03_2x port map ( Y=>nx1370, A0=>nx4609, A1=>nx11018, A2=>
      nx11028);
   ix4622 : nor02_2x port map ( Y=>nx4621, A0=>nx1366, A1=>nx1364);
   ix1367 : nor03_2x port map ( Y=>nx1366, A0=>nx4625, A1=>nx10384, A2=>
      nx11036);
   gen_3_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_3_cmp_mReg_8, QB=>
      nx4625, D=>window_3_8, CLK=>start, R=>rst);
   ix1365 : nor03_2x port map ( Y=>nx1364, A0=>gen_3_cmp_mReg_8, A1=>nx10750, 
      A2=>nx11044);
   ix1401 : nand02 port map ( Y=>gen_3_cmp_BSCmp_op2_9, A0=>nx4631, A1=>
      nx4637);
   ix4632 : nor02_2x port map ( Y=>nx4631, A0=>nx1396, A1=>nx1392);
   ix1397 : nor03_2x port map ( Y=>nx1396, A0=>gen_3_cmp_mReg_8, A1=>nx10390, 
      A2=>nx11012);
   ix1393 : nor03_2x port map ( Y=>nx1392, A0=>nx4625, A1=>nx11018, A2=>
      nx11028);
   ix4638 : nor02_2x port map ( Y=>nx4637, A0=>nx1388, A1=>nx1386);
   ix1389 : nor03_2x port map ( Y=>nx1388, A0=>nx4641, A1=>nx10384, A2=>
      nx11036);
   gen_3_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_3_cmp_mReg_9, QB=>
      nx4641, D=>window_3_9, CLK=>start, R=>rst);
   ix1387 : nor03_2x port map ( Y=>nx1386, A0=>gen_3_cmp_mReg_9, A1=>nx10750, 
      A2=>nx11044);
   ix1423 : nand02 port map ( Y=>gen_3_cmp_BSCmp_op2_10, A0=>nx4645, A1=>
      nx4649);
   ix4646 : nor02_2x port map ( Y=>nx4645, A0=>nx1418, A1=>nx1414);
   ix1419 : nor03_2x port map ( Y=>nx1418, A0=>gen_3_cmp_mReg_9, A1=>nx10390, 
      A2=>nx11012);
   ix1415 : nor03_2x port map ( Y=>nx1414, A0=>nx4641, A1=>nx11018, A2=>
      nx11028);
   ix4650 : nor02_2x port map ( Y=>nx4649, A0=>nx1410, A1=>nx1408);
   ix1411 : nor03_2x port map ( Y=>nx1410, A0=>nx4653, A1=>nx10384, A2=>
      nx11036);
   gen_3_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_3_cmp_mReg_10, QB=>
      nx4653, D=>window_3_10, CLK=>start, R=>rst);
   ix1409 : nor03_2x port map ( Y=>nx1408, A0=>gen_3_cmp_mReg_10, A1=>
      nx10750, A2=>nx11044);
   ix1445 : nand02 port map ( Y=>gen_3_cmp_BSCmp_op2_11, A0=>nx4659, A1=>
      nx4665);
   ix4660 : nor02_2x port map ( Y=>nx4659, A0=>nx1440, A1=>nx1436);
   ix1441 : nor03_2x port map ( Y=>nx1440, A0=>gen_3_cmp_mReg_10, A1=>
      nx10390, A2=>nx11012);
   ix1437 : nor03_2x port map ( Y=>nx1436, A0=>nx4653, A1=>nx11018, A2=>
      nx11028);
   ix4666 : nor02_2x port map ( Y=>nx4665, A0=>nx1432, A1=>nx1430);
   ix1433 : nor03_2x port map ( Y=>nx1432, A0=>nx4669, A1=>nx10384, A2=>
      nx11036);
   gen_3_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_3_cmp_mReg_11, QB=>
      nx4669, D=>window_3_11, CLK=>start, R=>rst);
   ix1431 : nor03_2x port map ( Y=>nx1430, A0=>gen_3_cmp_mReg_11, A1=>
      nx10750, A2=>nx11044);
   ix1467 : nand02 port map ( Y=>gen_3_cmp_BSCmp_op2_12, A0=>nx4674, A1=>
      nx4679);
   ix4675 : nor02_2x port map ( Y=>nx4674, A0=>nx1462, A1=>nx1458);
   ix1463 : nor03_2x port map ( Y=>nx1462, A0=>gen_3_cmp_mReg_11, A1=>
      nx10390, A2=>nx11012);
   ix1459 : nor03_2x port map ( Y=>nx1458, A0=>nx4669, A1=>nx11018, A2=>
      nx11028);
   ix4680 : nor02_2x port map ( Y=>nx4679, A0=>nx1454, A1=>nx1452);
   ix1455 : nor03_2x port map ( Y=>nx1454, A0=>nx4683, A1=>nx10386, A2=>
      nx11036);
   gen_3_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_3_cmp_mReg_12, QB=>
      nx4683, D=>window_3_12, CLK=>start, R=>rst);
   ix1453 : nor03_2x port map ( Y=>nx1452, A0=>gen_3_cmp_mReg_12, A1=>
      nx10750, A2=>nx11044);
   ix1489 : nand02 port map ( Y=>gen_3_cmp_BSCmp_op2_13, A0=>nx4687, A1=>
      nx4693);
   ix4688 : nor02_2x port map ( Y=>nx4687, A0=>nx1484, A1=>nx1480);
   ix1485 : nor03_2x port map ( Y=>nx1484, A0=>gen_3_cmp_mReg_12, A1=>
      nx10392, A2=>nx11014);
   ix1481 : nor03_2x port map ( Y=>nx1480, A0=>nx4683, A1=>nx11018, A2=>
      nx11030);
   ix4694 : nor02_2x port map ( Y=>nx4693, A0=>nx1476, A1=>nx1474);
   ix1477 : nor03_2x port map ( Y=>nx1476, A0=>nx4697, A1=>nx10386, A2=>
      nx11038);
   gen_3_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_3_cmp_mReg_13, QB=>
      nx4697, D=>window_3_13, CLK=>start, R=>rst);
   ix1475 : nor03_2x port map ( Y=>nx1474, A0=>gen_3_cmp_mReg_13, A1=>
      nx10750, A2=>nx11046);
   ix1511 : nand02 port map ( Y=>gen_3_cmp_BSCmp_op2_14, A0=>nx4702, A1=>
      nx4707);
   ix4703 : nor02_2x port map ( Y=>nx4702, A0=>nx1506, A1=>nx1502);
   ix1507 : nor03_2x port map ( Y=>nx1506, A0=>gen_3_cmp_mReg_13, A1=>
      nx10392, A2=>nx11014);
   ix1503 : nor03_2x port map ( Y=>nx1502, A0=>nx4697, A1=>nx11020, A2=>
      nx11030);
   ix4708 : nor02_2x port map ( Y=>nx4707, A0=>nx1498, A1=>nx1496);
   ix1499 : nor03_2x port map ( Y=>nx1498, A0=>nx4711, A1=>nx10386, A2=>
      nx11038);
   gen_3_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_3_cmp_mReg_14, QB=>
      nx4711, D=>window_3_14, CLK=>start, R=>rst);
   ix1497 : nor03_2x port map ( Y=>nx1496, A0=>gen_3_cmp_mReg_14, A1=>
      nx10750, A2=>nx11046);
   ix1533 : nand02 port map ( Y=>gen_3_cmp_BSCmp_op2_15, A0=>nx4717, A1=>
      nx4723);
   ix4718 : nor02_2x port map ( Y=>nx4717, A0=>nx1528, A1=>nx1524);
   ix1529 : nor03_2x port map ( Y=>nx1528, A0=>gen_3_cmp_mReg_14, A1=>
      nx10392, A2=>nx11014);
   ix1525 : nor03_2x port map ( Y=>nx1524, A0=>nx4711, A1=>nx11020, A2=>
      nx11030);
   ix4724 : nor02_2x port map ( Y=>nx4723, A0=>nx1520, A1=>nx1518);
   ix1521 : nor03_2x port map ( Y=>nx1520, A0=>nx4726, A1=>nx10386, A2=>
      nx11038);
   gen_3_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_3_cmp_mReg_15, QB=>
      nx4726, D=>window_3_15, CLK=>start, R=>rst);
   ix1519 : nor03_2x port map ( Y=>nx1518, A0=>gen_3_cmp_mReg_15, A1=>
      nx10752, A2=>nx11046);
   ix1543 : nand02 port map ( Y=>gen_3_cmp_BSCmp_op2_16, A0=>nx4733, A1=>
      nx4723);
   ix4734 : nor02_2x port map ( Y=>nx4733, A0=>nx1538, A1=>nx1534);
   ix1539 : nor03_2x port map ( Y=>nx1538, A0=>gen_3_cmp_mReg_15, A1=>
      nx10392, A2=>nx11014);
   ix1535 : nor03_2x port map ( Y=>nx1534, A0=>nx4726, A1=>nx11020, A2=>
      nx11030);
   ix1611 : nand02 port map ( Y=>gen_4_cmp_BSCmp_op2_1, A0=>nx4739, A1=>
      nx4759);
   ix4740 : nor02_2x port map ( Y=>nx4739, A0=>nx1606, A1=>nx1602);
   ix1607 : nor03_2x port map ( Y=>nx1606, A0=>gen_4_cmp_mReg_0, A1=>nx10376, 
      A2=>nx11050);
   gen_4_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_4_cmp_mReg_0, QB=>
      nx4745, D=>window_4_0, CLK=>start, R=>rst);
   ix4750 : inv01 port map ( Y=>nx4748, A=>gen_4_cmp_pMux_0);
   ix1603 : nor03_2x port map ( Y=>nx1602, A0=>nx4745, A1=>nx11056, A2=>
      nx11066);
   ix4758 : inv02 port map ( Y=>nx4757, A=>gen_4_cmp_pMux_2);
   ix4760 : nor02_2x port map ( Y=>nx4759, A0=>nx1592, A1=>nx1590);
   ix1593 : nor03_2x port map ( Y=>nx1592, A0=>nx4763, A1=>nx10370, A2=>
      nx11074);
   gen_4_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_4_cmp_mReg_1, QB=>
      nx4763, D=>window_4_1, CLK=>start, R=>rst);
   ix1591 : nor03_2x port map ( Y=>nx1590, A0=>gen_4_cmp_mReg_1, A1=>nx10754, 
      A2=>nx11082);
   ix1551 : nor03_2x port map ( Y=>nx1550, A0=>nx10376, A1=>nx4757, A2=>
      gen_4_cmp_pMux_0);
   ix1633 : nand02 port map ( Y=>gen_4_cmp_BSCmp_op2_2, A0=>nx4773, A1=>
      nx4779);
   ix4774 : nor02_2x port map ( Y=>nx4773, A0=>nx1628, A1=>nx1624);
   ix1629 : nor03_2x port map ( Y=>nx1628, A0=>gen_4_cmp_mReg_1, A1=>nx10376, 
      A2=>nx11050);
   ix1625 : nor03_2x port map ( Y=>nx1624, A0=>nx4763, A1=>nx11056, A2=>
      nx11066);
   ix4780 : nor02_2x port map ( Y=>nx4779, A0=>nx1620, A1=>nx1618);
   ix1621 : nor03_2x port map ( Y=>nx1620, A0=>nx4783, A1=>nx10370, A2=>
      nx11074);
   gen_4_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_4_cmp_mReg_2, QB=>
      nx4783, D=>window_4_2, CLK=>start, R=>rst);
   ix1619 : nor03_2x port map ( Y=>nx1618, A0=>gen_4_cmp_mReg_2, A1=>nx10754, 
      A2=>nx11082);
   ix1655 : nand02 port map ( Y=>gen_4_cmp_BSCmp_op2_3, A0=>nx4789, A1=>
      nx4793);
   ix4790 : nor02_2x port map ( Y=>nx4789, A0=>nx1650, A1=>nx1646);
   ix1651 : nor03_2x port map ( Y=>nx1650, A0=>gen_4_cmp_mReg_2, A1=>nx10376, 
      A2=>nx11050);
   ix1647 : nor03_2x port map ( Y=>nx1646, A0=>nx4783, A1=>nx11056, A2=>
      nx11066);
   ix4794 : nor02_2x port map ( Y=>nx4793, A0=>nx1642, A1=>nx1640);
   ix1643 : nor03_2x port map ( Y=>nx1642, A0=>nx4797, A1=>nx10370, A2=>
      nx11074);
   gen_4_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_4_cmp_mReg_3, QB=>
      nx4797, D=>window_4_3, CLK=>start, R=>rst);
   ix1641 : nor03_2x port map ( Y=>nx1640, A0=>gen_4_cmp_mReg_3, A1=>nx10754, 
      A2=>nx11082);
   ix1677 : nand02 port map ( Y=>gen_4_cmp_BSCmp_op2_4, A0=>nx4803, A1=>
      nx4809);
   ix4804 : nor02_2x port map ( Y=>nx4803, A0=>nx1672, A1=>nx1668);
   ix1673 : nor03_2x port map ( Y=>nx1672, A0=>gen_4_cmp_mReg_3, A1=>nx10376, 
      A2=>nx11050);
   ix1669 : nor03_2x port map ( Y=>nx1668, A0=>nx4797, A1=>nx11056, A2=>
      nx11066);
   ix4810 : nor02_2x port map ( Y=>nx4809, A0=>nx1664, A1=>nx1662);
   ix1665 : nor03_2x port map ( Y=>nx1664, A0=>nx4812, A1=>nx10370, A2=>
      nx11074);
   gen_4_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_4_cmp_mReg_4, QB=>
      nx4812, D=>window_4_4, CLK=>start, R=>rst);
   ix1663 : nor03_2x port map ( Y=>nx1662, A0=>gen_4_cmp_mReg_4, A1=>nx10754, 
      A2=>nx11082);
   ix1699 : nand02 port map ( Y=>gen_4_cmp_BSCmp_op2_5, A0=>nx4817, A1=>
      nx4823);
   ix4818 : nor02_2x port map ( Y=>nx4817, A0=>nx1694, A1=>nx1690);
   ix1695 : nor03_2x port map ( Y=>nx1694, A0=>gen_4_cmp_mReg_4, A1=>nx10376, 
      A2=>nx11050);
   ix1691 : nor03_2x port map ( Y=>nx1690, A0=>nx4812, A1=>nx11056, A2=>
      nx11066);
   ix4824 : nor02_2x port map ( Y=>nx4823, A0=>nx1686, A1=>nx1684);
   ix1687 : nor03_2x port map ( Y=>nx1686, A0=>nx4827, A1=>nx10372, A2=>
      nx11074);
   gen_4_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_4_cmp_mReg_5, QB=>
      nx4827, D=>window_4_5, CLK=>start, R=>rst);
   ix1685 : nor03_2x port map ( Y=>nx1684, A0=>gen_4_cmp_mReg_5, A1=>nx10754, 
      A2=>nx11082);
   ix1721 : nand02 port map ( Y=>gen_4_cmp_BSCmp_op2_6, A0=>nx4833, A1=>
      nx4837);
   ix4834 : nor02_2x port map ( Y=>nx4833, A0=>nx1716, A1=>nx1712);
   ix1717 : nor03_2x port map ( Y=>nx1716, A0=>gen_4_cmp_mReg_5, A1=>nx10378, 
      A2=>nx11050);
   ix1713 : nor03_2x port map ( Y=>nx1712, A0=>nx4827, A1=>nx11056, A2=>
      nx11066);
   ix4838 : nor02_2x port map ( Y=>nx4837, A0=>nx1708, A1=>nx1706);
   ix1709 : nor03_2x port map ( Y=>nx1708, A0=>nx4841, A1=>nx10372, A2=>
      nx11074);
   gen_4_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_4_cmp_mReg_6, QB=>
      nx4841, D=>window_4_6, CLK=>start, R=>rst);
   ix1707 : nor03_2x port map ( Y=>nx1706, A0=>gen_4_cmp_mReg_6, A1=>nx10754, 
      A2=>nx11082);
   ix1743 : nand02 port map ( Y=>gen_4_cmp_BSCmp_op2_7, A0=>nx4847, A1=>
      nx4853);
   ix4848 : nor02_2x port map ( Y=>nx4847, A0=>nx1738, A1=>nx1734);
   ix1739 : nor03_2x port map ( Y=>nx1738, A0=>gen_4_cmp_mReg_6, A1=>nx10378, 
      A2=>nx11052);
   ix1735 : nor03_2x port map ( Y=>nx1734, A0=>nx4841, A1=>nx11058, A2=>
      nx11068);
   ix4854 : nor02_2x port map ( Y=>nx4853, A0=>nx1730, A1=>nx1728);
   ix1731 : nor03_2x port map ( Y=>nx1730, A0=>nx4856, A1=>nx10372, A2=>
      nx11076);
   gen_4_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_4_cmp_mReg_7, QB=>
      nx4856, D=>window_4_7, CLK=>start, R=>rst);
   ix1729 : nor03_2x port map ( Y=>nx1728, A0=>gen_4_cmp_mReg_7, A1=>nx10754, 
      A2=>nx11084);
   ix1765 : nand02 port map ( Y=>gen_4_cmp_BSCmp_op2_8, A0=>nx4861, A1=>
      nx4867);
   ix4862 : nor02_2x port map ( Y=>nx4861, A0=>nx1760, A1=>nx1756);
   ix1761 : nor03_2x port map ( Y=>nx1760, A0=>gen_4_cmp_mReg_7, A1=>nx10378, 
      A2=>nx11052);
   ix1757 : nor03_2x port map ( Y=>nx1756, A0=>nx4856, A1=>nx11058, A2=>
      nx11068);
   ix4868 : nor02_2x port map ( Y=>nx4867, A0=>nx1752, A1=>nx1750);
   ix1753 : nor03_2x port map ( Y=>nx1752, A0=>nx4871, A1=>nx10372, A2=>
      nx11076);
   gen_4_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_4_cmp_mReg_8, QB=>
      nx4871, D=>window_4_8, CLK=>start, R=>rst);
   ix1751 : nor03_2x port map ( Y=>nx1750, A0=>gen_4_cmp_mReg_8, A1=>nx10756, 
      A2=>nx11084);
   ix1787 : nand02 port map ( Y=>gen_4_cmp_BSCmp_op2_9, A0=>nx4877, A1=>
      nx4881);
   ix4878 : nor02_2x port map ( Y=>nx4877, A0=>nx1782, A1=>nx1778);
   ix1783 : nor03_2x port map ( Y=>nx1782, A0=>gen_4_cmp_mReg_8, A1=>nx10378, 
      A2=>nx11052);
   ix1779 : nor03_2x port map ( Y=>nx1778, A0=>nx4871, A1=>nx11058, A2=>
      nx11068);
   ix4882 : nor02_2x port map ( Y=>nx4881, A0=>nx1774, A1=>nx1772);
   ix1775 : nor03_2x port map ( Y=>nx1774, A0=>nx4885, A1=>nx10372, A2=>
      nx11076);
   gen_4_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_4_cmp_mReg_9, QB=>
      nx4885, D=>window_4_9, CLK=>start, R=>rst);
   ix1773 : nor03_2x port map ( Y=>nx1772, A0=>gen_4_cmp_mReg_9, A1=>nx10756, 
      A2=>nx11084);
   ix1809 : nand02 port map ( Y=>gen_4_cmp_BSCmp_op2_10, A0=>nx4891, A1=>
      nx4897);
   ix4892 : nor02_2x port map ( Y=>nx4891, A0=>nx1804, A1=>nx1800);
   ix1805 : nor03_2x port map ( Y=>nx1804, A0=>gen_4_cmp_mReg_9, A1=>nx10378, 
      A2=>nx11052);
   ix1801 : nor03_2x port map ( Y=>nx1800, A0=>nx4885, A1=>nx11058, A2=>
      nx11068);
   ix4898 : nor02_2x port map ( Y=>nx4897, A0=>nx1796, A1=>nx1794);
   ix1797 : nor03_2x port map ( Y=>nx1796, A0=>nx4900, A1=>nx10372, A2=>
      nx11076);
   gen_4_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_4_cmp_mReg_10, QB=>
      nx4900, D=>window_4_10, CLK=>start, R=>rst);
   ix1795 : nor03_2x port map ( Y=>nx1794, A0=>gen_4_cmp_mReg_10, A1=>
      nx10756, A2=>nx11084);
   ix1831 : nand02 port map ( Y=>gen_4_cmp_BSCmp_op2_11, A0=>nx4905, A1=>
      nx4911);
   ix4906 : nor02_2x port map ( Y=>nx4905, A0=>nx1826, A1=>nx1822);
   ix1827 : nor03_2x port map ( Y=>nx1826, A0=>gen_4_cmp_mReg_10, A1=>
      nx10378, A2=>nx11052);
   ix1823 : nor03_2x port map ( Y=>nx1822, A0=>nx4900, A1=>nx11058, A2=>
      nx11068);
   ix4912 : nor02_2x port map ( Y=>nx4911, A0=>nx1818, A1=>nx1816);
   ix1819 : nor03_2x port map ( Y=>nx1818, A0=>nx4915, A1=>nx10372, A2=>
      nx11076);
   gen_4_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_4_cmp_mReg_11, QB=>
      nx4915, D=>window_4_11, CLK=>start, R=>rst);
   ix1817 : nor03_2x port map ( Y=>nx1816, A0=>gen_4_cmp_mReg_11, A1=>
      nx10756, A2=>nx11084);
   ix1853 : nand02 port map ( Y=>gen_4_cmp_BSCmp_op2_12, A0=>nx4921, A1=>
      nx4925);
   ix4922 : nor02_2x port map ( Y=>nx4921, A0=>nx1848, A1=>nx1844);
   ix1849 : nor03_2x port map ( Y=>nx1848, A0=>gen_4_cmp_mReg_11, A1=>
      nx10378, A2=>nx11052);
   ix1845 : nor03_2x port map ( Y=>nx1844, A0=>nx4915, A1=>nx11058, A2=>
      nx11068);
   ix4926 : nor02_2x port map ( Y=>nx4925, A0=>nx1840, A1=>nx1838);
   ix1841 : nor03_2x port map ( Y=>nx1840, A0=>nx4929, A1=>nx10374, A2=>
      nx11076);
   gen_4_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_4_cmp_mReg_12, QB=>
      nx4929, D=>window_4_12, CLK=>start, R=>rst);
   ix1839 : nor03_2x port map ( Y=>nx1838, A0=>gen_4_cmp_mReg_12, A1=>
      nx10756, A2=>nx11084);
   ix1875 : nand02 port map ( Y=>gen_4_cmp_BSCmp_op2_13, A0=>nx4935, A1=>
      nx4941);
   ix4936 : nor02_2x port map ( Y=>nx4935, A0=>nx1870, A1=>nx1866);
   ix1871 : nor03_2x port map ( Y=>nx1870, A0=>gen_4_cmp_mReg_12, A1=>
      nx10380, A2=>nx11054);
   ix1867 : nor03_2x port map ( Y=>nx1866, A0=>nx4929, A1=>nx11058, A2=>
      nx11070);
   ix4942 : nor02_2x port map ( Y=>nx4941, A0=>nx1862, A1=>nx1860);
   ix1863 : nor03_2x port map ( Y=>nx1862, A0=>nx4944, A1=>nx10374, A2=>
      nx11078);
   gen_4_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_4_cmp_mReg_13, QB=>
      nx4944, D=>window_4_13, CLK=>start, R=>rst);
   ix1861 : nor03_2x port map ( Y=>nx1860, A0=>gen_4_cmp_mReg_13, A1=>
      nx10756, A2=>nx11086);
   ix1897 : nand02 port map ( Y=>gen_4_cmp_BSCmp_op2_14, A0=>nx4949, A1=>
      nx4955);
   ix4950 : nor02_2x port map ( Y=>nx4949, A0=>nx1892, A1=>nx1888);
   ix1893 : nor03_2x port map ( Y=>nx1892, A0=>gen_4_cmp_mReg_13, A1=>
      nx10380, A2=>nx11054);
   ix1889 : nor03_2x port map ( Y=>nx1888, A0=>nx4944, A1=>nx11060, A2=>
      nx11070);
   ix4956 : nor02_2x port map ( Y=>nx4955, A0=>nx1884, A1=>nx1882);
   ix1885 : nor03_2x port map ( Y=>nx1884, A0=>nx4959, A1=>nx10374, A2=>
      nx11078);
   gen_4_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_4_cmp_mReg_14, QB=>
      nx4959, D=>window_4_14, CLK=>start, R=>rst);
   ix1883 : nor03_2x port map ( Y=>nx1882, A0=>gen_4_cmp_mReg_14, A1=>
      nx10756, A2=>nx11086);
   ix1919 : nand02 port map ( Y=>gen_4_cmp_BSCmp_op2_15, A0=>nx4965, A1=>
      nx4969);
   ix4966 : nor02_2x port map ( Y=>nx4965, A0=>nx1914, A1=>nx1910);
   ix1915 : nor03_2x port map ( Y=>nx1914, A0=>gen_4_cmp_mReg_14, A1=>
      nx10380, A2=>nx11054);
   ix1911 : nor03_2x port map ( Y=>nx1910, A0=>nx4959, A1=>nx11060, A2=>
      nx11070);
   ix4970 : nor02_2x port map ( Y=>nx4969, A0=>nx1906, A1=>nx1904);
   ix1907 : nor03_2x port map ( Y=>nx1906, A0=>nx4973, A1=>nx10374, A2=>
      nx11078);
   gen_4_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_4_cmp_mReg_15, QB=>
      nx4973, D=>window_4_15, CLK=>start, R=>rst);
   ix1905 : nor03_2x port map ( Y=>nx1904, A0=>gen_4_cmp_mReg_15, A1=>
      nx10758, A2=>nx11086);
   ix1929 : nand02 port map ( Y=>gen_4_cmp_BSCmp_op2_16, A0=>nx4979, A1=>
      nx4969);
   ix4980 : nor02_2x port map ( Y=>nx4979, A0=>nx1924, A1=>nx1920);
   ix1925 : nor03_2x port map ( Y=>nx1924, A0=>gen_4_cmp_mReg_15, A1=>
      nx10380, A2=>nx11054);
   ix1921 : nor03_2x port map ( Y=>nx1920, A0=>nx4973, A1=>nx11060, A2=>
      nx11070);
   ix1997 : nand02 port map ( Y=>gen_5_cmp_BSCmp_op2_1, A0=>nx4987, A1=>
      nx5005);
   ix4988 : nor02_2x port map ( Y=>nx4987, A0=>nx1992, A1=>nx1988);
   ix1993 : nor03_2x port map ( Y=>nx1992, A0=>gen_5_cmp_mReg_0, A1=>nx10364, 
      A2=>nx11090);
   gen_5_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_5_cmp_mReg_0, QB=>
      nx4991, D=>window_5_0, CLK=>start, R=>rst);
   ix4996 : inv01 port map ( Y=>nx4995, A=>gen_5_cmp_pMux_0);
   ix1989 : nor03_2x port map ( Y=>nx1988, A0=>nx4991, A1=>nx11096, A2=>
      nx11106);
   ix5004 : inv02 port map ( Y=>nx5003, A=>gen_5_cmp_pMux_2);
   ix5006 : nor02_2x port map ( Y=>nx5005, A0=>nx1978, A1=>nx1976);
   ix1979 : nor03_2x port map ( Y=>nx1978, A0=>nx5009, A1=>nx10358, A2=>
      nx11114);
   gen_5_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_5_cmp_mReg_1, QB=>
      nx5009, D=>window_5_1, CLK=>start, R=>rst);
   ix1977 : nor03_2x port map ( Y=>nx1976, A0=>gen_5_cmp_mReg_1, A1=>nx10760, 
      A2=>nx11122);
   ix1937 : nor03_2x port map ( Y=>nx1936, A0=>nx10364, A1=>nx5003, A2=>
      gen_5_cmp_pMux_0);
   ix2019 : nand02 port map ( Y=>gen_5_cmp_BSCmp_op2_2, A0=>nx5021, A1=>
      nx5027);
   ix5022 : nor02_2x port map ( Y=>nx5021, A0=>nx2014, A1=>nx2010);
   ix2015 : nor03_2x port map ( Y=>nx2014, A0=>gen_5_cmp_mReg_1, A1=>nx10364, 
      A2=>nx11090);
   ix2011 : nor03_2x port map ( Y=>nx2010, A0=>nx5009, A1=>nx11096, A2=>
      nx11106);
   ix5028 : nor02_2x port map ( Y=>nx5027, A0=>nx2006, A1=>nx2004);
   ix2007 : nor03_2x port map ( Y=>nx2006, A0=>nx5030, A1=>nx10358, A2=>
      nx11114);
   gen_5_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_5_cmp_mReg_2, QB=>
      nx5030, D=>window_5_2, CLK=>start, R=>rst);
   ix2005 : nor03_2x port map ( Y=>nx2004, A0=>gen_5_cmp_mReg_2, A1=>nx10760, 
      A2=>nx11122);
   ix2041 : nand02 port map ( Y=>gen_5_cmp_BSCmp_op2_3, A0=>nx5035, A1=>
      nx5041);
   ix5036 : nor02_2x port map ( Y=>nx5035, A0=>nx2036, A1=>nx2032);
   ix2037 : nor03_2x port map ( Y=>nx2036, A0=>gen_5_cmp_mReg_2, A1=>nx10364, 
      A2=>nx11090);
   ix2033 : nor03_2x port map ( Y=>nx2032, A0=>nx5030, A1=>nx11096, A2=>
      nx11106);
   ix5042 : nor02_2x port map ( Y=>nx5041, A0=>nx2028, A1=>nx2026);
   ix2029 : nor03_2x port map ( Y=>nx2028, A0=>nx5045, A1=>nx10358, A2=>
      nx11114);
   gen_5_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_5_cmp_mReg_3, QB=>
      nx5045, D=>window_5_3, CLK=>start, R=>rst);
   ix2027 : nor03_2x port map ( Y=>nx2026, A0=>gen_5_cmp_mReg_3, A1=>nx10760, 
      A2=>nx11122);
   ix2063 : nand02 port map ( Y=>gen_5_cmp_BSCmp_op2_4, A0=>nx5051, A1=>
      nx5057);
   ix5052 : nor02_2x port map ( Y=>nx5051, A0=>nx2058, A1=>nx2054);
   ix2059 : nor03_2x port map ( Y=>nx2058, A0=>gen_5_cmp_mReg_3, A1=>nx10364, 
      A2=>nx11090);
   ix2055 : nor03_2x port map ( Y=>nx2054, A0=>nx5045, A1=>nx11096, A2=>
      nx11106);
   ix5058 : nor02_2x port map ( Y=>nx5057, A0=>nx2050, A1=>nx2048);
   ix2051 : nor03_2x port map ( Y=>nx2050, A0=>nx5060, A1=>nx10358, A2=>
      nx11114);
   gen_5_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_5_cmp_mReg_4, QB=>
      nx5060, D=>window_5_4, CLK=>start, R=>rst);
   ix2049 : nor03_2x port map ( Y=>nx2048, A0=>gen_5_cmp_mReg_4, A1=>nx10760, 
      A2=>nx11122);
   ix2085 : nand02 port map ( Y=>gen_5_cmp_BSCmp_op2_5, A0=>nx5065, A1=>
      nx5071);
   ix5066 : nor02_2x port map ( Y=>nx5065, A0=>nx2080, A1=>nx2076);
   ix2081 : nor03_2x port map ( Y=>nx2080, A0=>gen_5_cmp_mReg_4, A1=>nx10364, 
      A2=>nx11090);
   ix2077 : nor03_2x port map ( Y=>nx2076, A0=>nx5060, A1=>nx11096, A2=>
      nx11106);
   ix5072 : nor02_2x port map ( Y=>nx5071, A0=>nx2072, A1=>nx2070);
   ix2073 : nor03_2x port map ( Y=>nx2072, A0=>nx5075, A1=>nx10360, A2=>
      nx11114);
   gen_5_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_5_cmp_mReg_5, QB=>
      nx5075, D=>window_5_5, CLK=>start, R=>rst);
   ix2071 : nor03_2x port map ( Y=>nx2070, A0=>gen_5_cmp_mReg_5, A1=>nx10760, 
      A2=>nx11122);
   ix2107 : nand02 port map ( Y=>gen_5_cmp_BSCmp_op2_6, A0=>nx5081, A1=>
      nx5087);
   ix5082 : nor02_2x port map ( Y=>nx5081, A0=>nx2102, A1=>nx2098);
   ix2103 : nor03_2x port map ( Y=>nx2102, A0=>gen_5_cmp_mReg_5, A1=>nx10366, 
      A2=>nx11090);
   ix2099 : nor03_2x port map ( Y=>nx2098, A0=>nx5075, A1=>nx11096, A2=>
      nx11106);
   ix5088 : nor02_2x port map ( Y=>nx5087, A0=>nx2094, A1=>nx2092);
   ix2095 : nor03_2x port map ( Y=>nx2094, A0=>nx5090, A1=>nx10360, A2=>
      nx11114);
   gen_5_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_5_cmp_mReg_6, QB=>
      nx5090, D=>window_5_6, CLK=>start, R=>rst);
   ix2093 : nor03_2x port map ( Y=>nx2092, A0=>gen_5_cmp_mReg_6, A1=>nx10760, 
      A2=>nx11122);
   ix2129 : nand02 port map ( Y=>gen_5_cmp_BSCmp_op2_7, A0=>nx5097, A1=>
      nx5103);
   ix5098 : nor02_2x port map ( Y=>nx5097, A0=>nx2124, A1=>nx2120);
   ix2125 : nor03_2x port map ( Y=>nx2124, A0=>gen_5_cmp_mReg_6, A1=>nx10366, 
      A2=>nx11092);
   ix2121 : nor03_2x port map ( Y=>nx2120, A0=>nx5090, A1=>nx11098, A2=>
      nx11108);
   ix5104 : nor02_2x port map ( Y=>nx5103, A0=>nx2116, A1=>nx2114);
   ix2117 : nor03_2x port map ( Y=>nx2116, A0=>nx5107, A1=>nx10360, A2=>
      nx11116);
   gen_5_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_5_cmp_mReg_7, QB=>
      nx5107, D=>window_5_7, CLK=>start, R=>rst);
   ix2115 : nor03_2x port map ( Y=>nx2114, A0=>gen_5_cmp_mReg_7, A1=>nx10760, 
      A2=>nx11124);
   ix2151 : nand02 port map ( Y=>gen_5_cmp_BSCmp_op2_8, A0=>nx5111, A1=>
      nx5117);
   ix5112 : nor02_2x port map ( Y=>nx5111, A0=>nx2146, A1=>nx2142);
   ix2147 : nor03_2x port map ( Y=>nx2146, A0=>gen_5_cmp_mReg_7, A1=>nx10366, 
      A2=>nx11092);
   ix2143 : nor03_2x port map ( Y=>nx2142, A0=>nx5107, A1=>nx11098, A2=>
      nx11108);
   ix5118 : nor02_2x port map ( Y=>nx5117, A0=>nx2138, A1=>nx2136);
   ix2139 : nor03_2x port map ( Y=>nx2138, A0=>nx5121, A1=>nx10360, A2=>
      nx11116);
   gen_5_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_5_cmp_mReg_8, QB=>
      nx5121, D=>window_5_8, CLK=>start, R=>rst);
   ix2137 : nor03_2x port map ( Y=>nx2136, A0=>gen_5_cmp_mReg_8, A1=>nx10762, 
      A2=>nx11124);
   ix2173 : nand02 port map ( Y=>gen_5_cmp_BSCmp_op2_9, A0=>nx5125, A1=>
      nx5131);
   ix5126 : nor02_2x port map ( Y=>nx5125, A0=>nx2168, A1=>nx2164);
   ix2169 : nor03_2x port map ( Y=>nx2168, A0=>gen_5_cmp_mReg_8, A1=>nx10366, 
      A2=>nx11092);
   ix2165 : nor03_2x port map ( Y=>nx2164, A0=>nx5121, A1=>nx11098, A2=>
      nx11108);
   ix5132 : nor02_2x port map ( Y=>nx5131, A0=>nx2160, A1=>nx2158);
   ix2161 : nor03_2x port map ( Y=>nx2160, A0=>nx5134, A1=>nx10360, A2=>
      nx11116);
   gen_5_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_5_cmp_mReg_9, QB=>
      nx5134, D=>window_5_9, CLK=>start, R=>rst);
   ix2159 : nor03_2x port map ( Y=>nx2158, A0=>gen_5_cmp_mReg_9, A1=>nx10762, 
      A2=>nx11124);
   ix2195 : nand02 port map ( Y=>gen_5_cmp_BSCmp_op2_10, A0=>nx5141, A1=>
      nx5147);
   ix5142 : nor02_2x port map ( Y=>nx5141, A0=>nx2190, A1=>nx2186);
   ix2191 : nor03_2x port map ( Y=>nx2190, A0=>gen_5_cmp_mReg_9, A1=>nx10366, 
      A2=>nx11092);
   ix2187 : nor03_2x port map ( Y=>nx2186, A0=>nx5134, A1=>nx11098, A2=>
      nx11108);
   ix5148 : nor02_2x port map ( Y=>nx5147, A0=>nx2182, A1=>nx2180);
   ix2183 : nor03_2x port map ( Y=>nx2182, A0=>nx5151, A1=>nx10360, A2=>
      nx11116);
   gen_5_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_5_cmp_mReg_10, QB=>
      nx5151, D=>window_5_10, CLK=>start, R=>rst);
   ix2181 : nor03_2x port map ( Y=>nx2180, A0=>gen_5_cmp_mReg_10, A1=>
      nx10762, A2=>nx11124);
   ix2217 : nand02 port map ( Y=>gen_5_cmp_BSCmp_op2_11, A0=>nx5155, A1=>
      nx5161);
   ix5156 : nor02_2x port map ( Y=>nx5155, A0=>nx2212, A1=>nx2208);
   ix2213 : nor03_2x port map ( Y=>nx2212, A0=>gen_5_cmp_mReg_10, A1=>
      nx10366, A2=>nx11092);
   ix2209 : nor03_2x port map ( Y=>nx2208, A0=>nx5151, A1=>nx11098, A2=>
      nx11108);
   ix5162 : nor02_2x port map ( Y=>nx5161, A0=>nx2204, A1=>nx2202);
   ix2205 : nor03_2x port map ( Y=>nx2204, A0=>nx5165, A1=>nx10360, A2=>
      nx11116);
   gen_5_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_5_cmp_mReg_11, QB=>
      nx5165, D=>window_5_11, CLK=>start, R=>rst);
   ix2203 : nor03_2x port map ( Y=>nx2202, A0=>gen_5_cmp_mReg_11, A1=>
      nx10762, A2=>nx11124);
   ix2239 : nand02 port map ( Y=>gen_5_cmp_BSCmp_op2_12, A0=>nx5169, A1=>
      nx5175);
   ix5170 : nor02_2x port map ( Y=>nx5169, A0=>nx2234, A1=>nx2230);
   ix2235 : nor03_2x port map ( Y=>nx2234, A0=>gen_5_cmp_mReg_11, A1=>
      nx10366, A2=>nx11092);
   ix2231 : nor03_2x port map ( Y=>nx2230, A0=>nx5165, A1=>nx11098, A2=>
      nx11108);
   ix5176 : nor02_2x port map ( Y=>nx5175, A0=>nx2226, A1=>nx2224);
   ix2227 : nor03_2x port map ( Y=>nx2226, A0=>nx5178, A1=>nx10362, A2=>
      nx11116);
   gen_5_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_5_cmp_mReg_12, QB=>
      nx5178, D=>window_5_12, CLK=>start, R=>rst);
   ix2225 : nor03_2x port map ( Y=>nx2224, A0=>gen_5_cmp_mReg_12, A1=>
      nx10762, A2=>nx11124);
   ix2261 : nand02 port map ( Y=>gen_5_cmp_BSCmp_op2_13, A0=>nx5185, A1=>
      nx5191);
   ix5186 : nor02_2x port map ( Y=>nx5185, A0=>nx2256, A1=>nx2252);
   ix2257 : nor03_2x port map ( Y=>nx2256, A0=>gen_5_cmp_mReg_12, A1=>
      nx10368, A2=>nx11094);
   ix2253 : nor03_2x port map ( Y=>nx2252, A0=>nx5178, A1=>nx11098, A2=>
      nx11110);
   ix5192 : nor02_2x port map ( Y=>nx5191, A0=>nx2248, A1=>nx2246);
   ix2249 : nor03_2x port map ( Y=>nx2248, A0=>nx5195, A1=>nx10362, A2=>
      nx11118);
   gen_5_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_5_cmp_mReg_13, QB=>
      nx5195, D=>window_5_13, CLK=>start, R=>rst);
   ix2247 : nor03_2x port map ( Y=>nx2246, A0=>gen_5_cmp_mReg_13, A1=>
      nx10762, A2=>nx11126);
   ix2283 : nand02 port map ( Y=>gen_5_cmp_BSCmp_op2_14, A0=>nx5199, A1=>
      nx5205);
   ix5200 : nor02_2x port map ( Y=>nx5199, A0=>nx2278, A1=>nx2274);
   ix2279 : nor03_2x port map ( Y=>nx2278, A0=>gen_5_cmp_mReg_13, A1=>
      nx10368, A2=>nx11094);
   ix2275 : nor03_2x port map ( Y=>nx2274, A0=>nx5195, A1=>nx11100, A2=>
      nx11110);
   ix5206 : nor02_2x port map ( Y=>nx5205, A0=>nx2270, A1=>nx2268);
   ix2271 : nor03_2x port map ( Y=>nx2270, A0=>nx5209, A1=>nx10362, A2=>
      nx11118);
   gen_5_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_5_cmp_mReg_14, QB=>
      nx5209, D=>window_5_14, CLK=>start, R=>rst);
   ix2269 : nor03_2x port map ( Y=>nx2268, A0=>gen_5_cmp_mReg_14, A1=>
      nx10762, A2=>nx11126);
   ix2305 : nand02 port map ( Y=>gen_5_cmp_BSCmp_op2_15, A0=>nx5213, A1=>
      nx5219);
   ix5214 : nor02_2x port map ( Y=>nx5213, A0=>nx2300, A1=>nx2296);
   ix2301 : nor03_2x port map ( Y=>nx2300, A0=>gen_5_cmp_mReg_14, A1=>
      nx10368, A2=>nx11094);
   ix2297 : nor03_2x port map ( Y=>nx2296, A0=>nx5209, A1=>nx11100, A2=>
      nx11110);
   ix5220 : nor02_2x port map ( Y=>nx5219, A0=>nx2292, A1=>nx2290);
   ix2293 : nor03_2x port map ( Y=>nx2292, A0=>nx5222, A1=>nx10362, A2=>
      nx11118);
   gen_5_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_5_cmp_mReg_15, QB=>
      nx5222, D=>window_5_15, CLK=>start, R=>rst);
   ix2291 : nor03_2x port map ( Y=>nx2290, A0=>gen_5_cmp_mReg_15, A1=>
      nx10764, A2=>nx11126);
   ix2315 : nand02 port map ( Y=>gen_5_cmp_BSCmp_op2_16, A0=>nx5229, A1=>
      nx5219);
   ix5230 : nor02_2x port map ( Y=>nx5229, A0=>nx2310, A1=>nx2306);
   ix2311 : nor03_2x port map ( Y=>nx2310, A0=>gen_5_cmp_mReg_15, A1=>
      nx10368, A2=>nx11094);
   ix2307 : nor03_2x port map ( Y=>nx2306, A0=>nx5222, A1=>nx11100, A2=>
      nx11110);
   ix2383 : nand02 port map ( Y=>gen_6_cmp_BSCmp_op2_1, A0=>nx5235, A1=>
      nx5255);
   ix5236 : nor02_2x port map ( Y=>nx5235, A0=>nx2378, A1=>nx2374);
   ix2379 : nor03_2x port map ( Y=>nx2378, A0=>gen_6_cmp_mReg_0, A1=>nx10352, 
      A2=>nx11130);
   gen_6_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_6_cmp_mReg_0, QB=>
      nx5241, D=>window_6_0, CLK=>start, R=>rst);
   ix5246 : inv01 port map ( Y=>nx5244, A=>gen_6_cmp_pMux_0);
   ix2375 : nor03_2x port map ( Y=>nx2374, A0=>nx5241, A1=>nx11136, A2=>
      nx11146);
   ix5254 : inv02 port map ( Y=>nx5253, A=>gen_6_cmp_pMux_2);
   ix5256 : nor02_2x port map ( Y=>nx5255, A0=>nx2364, A1=>nx2362);
   ix2365 : nor03_2x port map ( Y=>nx2364, A0=>nx5259, A1=>nx10346, A2=>
      nx11154);
   gen_6_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_6_cmp_mReg_1, QB=>
      nx5259, D=>window_6_1, CLK=>start, R=>rst);
   ix2363 : nor03_2x port map ( Y=>nx2362, A0=>gen_6_cmp_mReg_1, A1=>nx10766, 
      A2=>nx11162);
   ix2323 : nor03_2x port map ( Y=>nx2322, A0=>nx10352, A1=>nx5253, A2=>
      gen_6_cmp_pMux_0);
   ix2405 : nand02 port map ( Y=>gen_6_cmp_BSCmp_op2_2, A0=>nx5269, A1=>
      nx5275);
   ix5270 : nor02_2x port map ( Y=>nx5269, A0=>nx2400, A1=>nx2396);
   ix2401 : nor03_2x port map ( Y=>nx2400, A0=>gen_6_cmp_mReg_1, A1=>nx10352, 
      A2=>nx11130);
   ix2397 : nor03_2x port map ( Y=>nx2396, A0=>nx5259, A1=>nx11136, A2=>
      nx11146);
   ix5276 : nor02_2x port map ( Y=>nx5275, A0=>nx2392, A1=>nx2390);
   ix2393 : nor03_2x port map ( Y=>nx2392, A0=>nx5279, A1=>nx10346, A2=>
      nx11154);
   gen_6_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_6_cmp_mReg_2, QB=>
      nx5279, D=>window_6_2, CLK=>start, R=>rst);
   ix2391 : nor03_2x port map ( Y=>nx2390, A0=>gen_6_cmp_mReg_2, A1=>nx10766, 
      A2=>nx11162);
   ix2427 : nand02 port map ( Y=>gen_6_cmp_BSCmp_op2_3, A0=>nx5285, A1=>
      nx5289);
   ix5286 : nor02_2x port map ( Y=>nx5285, A0=>nx2422, A1=>nx2418);
   ix2423 : nor03_2x port map ( Y=>nx2422, A0=>gen_6_cmp_mReg_2, A1=>nx10352, 
      A2=>nx11130);
   ix2419 : nor03_2x port map ( Y=>nx2418, A0=>nx5279, A1=>nx11136, A2=>
      nx11146);
   ix5290 : nor02_2x port map ( Y=>nx5289, A0=>nx2414, A1=>nx2412);
   ix2415 : nor03_2x port map ( Y=>nx2414, A0=>nx5293, A1=>nx10346, A2=>
      nx11154);
   gen_6_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_6_cmp_mReg_3, QB=>
      nx5293, D=>window_6_3, CLK=>start, R=>rst);
   ix2413 : nor03_2x port map ( Y=>nx2412, A0=>gen_6_cmp_mReg_3, A1=>nx10766, 
      A2=>nx11162);
   ix2449 : nand02 port map ( Y=>gen_6_cmp_BSCmp_op2_4, A0=>nx5299, A1=>
      nx5305);
   ix5300 : nor02_2x port map ( Y=>nx5299, A0=>nx2444, A1=>nx2440);
   ix2445 : nor03_2x port map ( Y=>nx2444, A0=>gen_6_cmp_mReg_3, A1=>nx10352, 
      A2=>nx11130);
   ix2441 : nor03_2x port map ( Y=>nx2440, A0=>nx5293, A1=>nx11136, A2=>
      nx11146);
   ix5306 : nor02_2x port map ( Y=>nx5305, A0=>nx2436, A1=>nx2434);
   ix2437 : nor03_2x port map ( Y=>nx2436, A0=>nx5308, A1=>nx10346, A2=>
      nx11154);
   gen_6_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_6_cmp_mReg_4, QB=>
      nx5308, D=>window_6_4, CLK=>start, R=>rst);
   ix2435 : nor03_2x port map ( Y=>nx2434, A0=>gen_6_cmp_mReg_4, A1=>nx10766, 
      A2=>nx11162);
   ix2471 : nand02 port map ( Y=>gen_6_cmp_BSCmp_op2_5, A0=>nx5313, A1=>
      nx5319);
   ix5314 : nor02_2x port map ( Y=>nx5313, A0=>nx2466, A1=>nx2462);
   ix2467 : nor03_2x port map ( Y=>nx2466, A0=>gen_6_cmp_mReg_4, A1=>nx10352, 
      A2=>nx11130);
   ix2463 : nor03_2x port map ( Y=>nx2462, A0=>nx5308, A1=>nx11136, A2=>
      nx11146);
   ix5320 : nor02_2x port map ( Y=>nx5319, A0=>nx2458, A1=>nx2456);
   ix2459 : nor03_2x port map ( Y=>nx2458, A0=>nx5323, A1=>nx10348, A2=>
      nx11154);
   gen_6_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_6_cmp_mReg_5, QB=>
      nx5323, D=>window_6_5, CLK=>start, R=>rst);
   ix2457 : nor03_2x port map ( Y=>nx2456, A0=>gen_6_cmp_mReg_5, A1=>nx10766, 
      A2=>nx11162);
   ix2493 : nand02 port map ( Y=>gen_6_cmp_BSCmp_op2_6, A0=>nx5329, A1=>
      nx5333);
   ix5330 : nor02_2x port map ( Y=>nx5329, A0=>nx2488, A1=>nx2484);
   ix2489 : nor03_2x port map ( Y=>nx2488, A0=>gen_6_cmp_mReg_5, A1=>nx10354, 
      A2=>nx11130);
   ix2485 : nor03_2x port map ( Y=>nx2484, A0=>nx5323, A1=>nx11136, A2=>
      nx11146);
   ix5334 : nor02_2x port map ( Y=>nx5333, A0=>nx2480, A1=>nx2478);
   ix2481 : nor03_2x port map ( Y=>nx2480, A0=>nx5337, A1=>nx10348, A2=>
      nx11154);
   gen_6_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_6_cmp_mReg_6, QB=>
      nx5337, D=>window_6_6, CLK=>start, R=>rst);
   ix2479 : nor03_2x port map ( Y=>nx2478, A0=>gen_6_cmp_mReg_6, A1=>nx10766, 
      A2=>nx11162);
   ix2515 : nand02 port map ( Y=>gen_6_cmp_BSCmp_op2_7, A0=>nx5343, A1=>
      nx5349);
   ix5344 : nor02_2x port map ( Y=>nx5343, A0=>nx2510, A1=>nx2506);
   ix2511 : nor03_2x port map ( Y=>nx2510, A0=>gen_6_cmp_mReg_6, A1=>nx10354, 
      A2=>nx11132);
   ix2507 : nor03_2x port map ( Y=>nx2506, A0=>nx5337, A1=>nx11138, A2=>
      nx11148);
   ix5350 : nor02_2x port map ( Y=>nx5349, A0=>nx2502, A1=>nx2500);
   ix2503 : nor03_2x port map ( Y=>nx2502, A0=>nx5352, A1=>nx10348, A2=>
      nx11156);
   gen_6_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_6_cmp_mReg_7, QB=>
      nx5352, D=>window_6_7, CLK=>start, R=>rst);
   ix2501 : nor03_2x port map ( Y=>nx2500, A0=>gen_6_cmp_mReg_7, A1=>nx10766, 
      A2=>nx11164);
   ix2537 : nand02 port map ( Y=>gen_6_cmp_BSCmp_op2_8, A0=>nx5357, A1=>
      nx5363);
   ix5358 : nor02_2x port map ( Y=>nx5357, A0=>nx2532, A1=>nx2528);
   ix2533 : nor03_2x port map ( Y=>nx2532, A0=>gen_6_cmp_mReg_7, A1=>nx10354, 
      A2=>nx11132);
   ix2529 : nor03_2x port map ( Y=>nx2528, A0=>nx5352, A1=>nx11138, A2=>
      nx11148);
   ix5364 : nor02_2x port map ( Y=>nx5363, A0=>nx2524, A1=>nx2522);
   ix2525 : nor03_2x port map ( Y=>nx2524, A0=>nx5367, A1=>nx10348, A2=>
      nx11156);
   gen_6_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_6_cmp_mReg_8, QB=>
      nx5367, D=>window_6_8, CLK=>start, R=>rst);
   ix2523 : nor03_2x port map ( Y=>nx2522, A0=>gen_6_cmp_mReg_8, A1=>nx10768, 
      A2=>nx11164);
   ix2559 : nand02 port map ( Y=>gen_6_cmp_BSCmp_op2_9, A0=>nx5373, A1=>
      nx5377);
   ix5374 : nor02_2x port map ( Y=>nx5373, A0=>nx2554, A1=>nx2550);
   ix2555 : nor03_2x port map ( Y=>nx2554, A0=>gen_6_cmp_mReg_8, A1=>nx10354, 
      A2=>nx11132);
   ix2551 : nor03_2x port map ( Y=>nx2550, A0=>nx5367, A1=>nx11138, A2=>
      nx11148);
   ix5378 : nor02_2x port map ( Y=>nx5377, A0=>nx2546, A1=>nx2544);
   ix2547 : nor03_2x port map ( Y=>nx2546, A0=>nx5381, A1=>nx10348, A2=>
      nx11156);
   gen_6_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_6_cmp_mReg_9, QB=>
      nx5381, D=>window_6_9, CLK=>start, R=>rst);
   ix2545 : nor03_2x port map ( Y=>nx2544, A0=>gen_6_cmp_mReg_9, A1=>nx10768, 
      A2=>nx11164);
   ix2581 : nand02 port map ( Y=>gen_6_cmp_BSCmp_op2_10, A0=>nx5387, A1=>
      nx5393);
   ix5388 : nor02_2x port map ( Y=>nx5387, A0=>nx2576, A1=>nx2572);
   ix2577 : nor03_2x port map ( Y=>nx2576, A0=>gen_6_cmp_mReg_9, A1=>nx10354, 
      A2=>nx11132);
   ix2573 : nor03_2x port map ( Y=>nx2572, A0=>nx5381, A1=>nx11138, A2=>
      nx11148);
   ix5394 : nor02_2x port map ( Y=>nx5393, A0=>nx2568, A1=>nx2566);
   ix2569 : nor03_2x port map ( Y=>nx2568, A0=>nx5397, A1=>nx10348, A2=>
      nx11156);
   gen_6_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_6_cmp_mReg_10, QB=>
      nx5397, D=>window_6_10, CLK=>start, R=>rst);
   ix2567 : nor03_2x port map ( Y=>nx2566, A0=>gen_6_cmp_mReg_10, A1=>
      nx10768, A2=>nx11164);
   ix2603 : nand02 port map ( Y=>gen_6_cmp_BSCmp_op2_11, A0=>nx5403, A1=>
      nx5409);
   ix5404 : nor02_2x port map ( Y=>nx5403, A0=>nx2598, A1=>nx2594);
   ix2599 : nor03_2x port map ( Y=>nx2598, A0=>gen_6_cmp_mReg_10, A1=>
      nx10354, A2=>nx11132);
   ix2595 : nor03_2x port map ( Y=>nx2594, A0=>nx5397, A1=>nx11138, A2=>
      nx11148);
   ix5410 : nor02_2x port map ( Y=>nx5409, A0=>nx2590, A1=>nx2588);
   ix2591 : nor03_2x port map ( Y=>nx2590, A0=>nx5413, A1=>nx10348, A2=>
      nx11156);
   gen_6_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_6_cmp_mReg_11, QB=>
      nx5413, D=>window_6_11, CLK=>start, R=>rst);
   ix2589 : nor03_2x port map ( Y=>nx2588, A0=>gen_6_cmp_mReg_11, A1=>
      nx10768, A2=>nx11164);
   ix2625 : nand02 port map ( Y=>gen_6_cmp_BSCmp_op2_12, A0=>nx5417, A1=>
      nx5421);
   ix5418 : nor02_2x port map ( Y=>nx5417, A0=>nx2620, A1=>nx2616);
   ix2621 : nor03_2x port map ( Y=>nx2620, A0=>gen_6_cmp_mReg_11, A1=>
      nx10354, A2=>nx11132);
   ix2617 : nor03_2x port map ( Y=>nx2616, A0=>nx5413, A1=>nx11138, A2=>
      nx11148);
   ix5422 : nor02_2x port map ( Y=>nx5421, A0=>nx2612, A1=>nx2610);
   ix2613 : nor03_2x port map ( Y=>nx2612, A0=>nx5425, A1=>nx10350, A2=>
      nx11156);
   gen_6_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_6_cmp_mReg_12, QB=>
      nx5425, D=>window_6_12, CLK=>start, R=>rst);
   ix2611 : nor03_2x port map ( Y=>nx2610, A0=>gen_6_cmp_mReg_12, A1=>
      nx10768, A2=>nx11164);
   ix2647 : nand02 port map ( Y=>gen_6_cmp_BSCmp_op2_13, A0=>nx5431, A1=>
      nx5437);
   ix5432 : nor02_2x port map ( Y=>nx5431, A0=>nx2642, A1=>nx2638);
   ix2643 : nor03_2x port map ( Y=>nx2642, A0=>gen_6_cmp_mReg_12, A1=>
      nx10356, A2=>nx11134);
   ix2639 : nor03_2x port map ( Y=>nx2638, A0=>nx5425, A1=>nx11138, A2=>
      nx11150);
   ix5438 : nor02_2x port map ( Y=>nx5437, A0=>nx2634, A1=>nx2632);
   ix2635 : nor03_2x port map ( Y=>nx2634, A0=>nx5441, A1=>nx10350, A2=>
      nx11158);
   gen_6_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_6_cmp_mReg_13, QB=>
      nx5441, D=>window_6_13, CLK=>start, R=>rst);
   ix2633 : nor03_2x port map ( Y=>nx2632, A0=>gen_6_cmp_mReg_13, A1=>
      nx10768, A2=>nx11166);
   ix2669 : nand02 port map ( Y=>gen_6_cmp_BSCmp_op2_14, A0=>nx5446, A1=>
      nx5451);
   ix5447 : nor02_2x port map ( Y=>nx5446, A0=>nx2664, A1=>nx2660);
   ix2665 : nor03_2x port map ( Y=>nx2664, A0=>gen_6_cmp_mReg_13, A1=>
      nx10356, A2=>nx11134);
   ix2661 : nor03_2x port map ( Y=>nx2660, A0=>nx5441, A1=>nx11140, A2=>
      nx11150);
   ix5452 : nor02_2x port map ( Y=>nx5451, A0=>nx2656, A1=>nx2654);
   ix2657 : nor03_2x port map ( Y=>nx2656, A0=>nx5455, A1=>nx10350, A2=>
      nx11158);
   gen_6_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_6_cmp_mReg_14, QB=>
      nx5455, D=>window_6_14, CLK=>start, R=>rst);
   ix2655 : nor03_2x port map ( Y=>nx2654, A0=>gen_6_cmp_mReg_14, A1=>
      nx10768, A2=>nx11166);
   ix2691 : nand02 port map ( Y=>gen_6_cmp_BSCmp_op2_15, A0=>nx5459, A1=>
      nx5465);
   ix5460 : nor02_2x port map ( Y=>nx5459, A0=>nx2686, A1=>nx2682);
   ix2687 : nor03_2x port map ( Y=>nx2686, A0=>gen_6_cmp_mReg_14, A1=>
      nx10356, A2=>nx11134);
   ix2683 : nor03_2x port map ( Y=>nx2682, A0=>nx5455, A1=>nx11140, A2=>
      nx11150);
   ix5466 : nor02_2x port map ( Y=>nx5465, A0=>nx2678, A1=>nx2676);
   ix2679 : nor03_2x port map ( Y=>nx2678, A0=>nx5469, A1=>nx10350, A2=>
      nx11158);
   gen_6_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_6_cmp_mReg_15, QB=>
      nx5469, D=>window_6_15, CLK=>start, R=>rst);
   ix2677 : nor03_2x port map ( Y=>nx2676, A0=>gen_6_cmp_mReg_15, A1=>
      nx10770, A2=>nx11166);
   ix2701 : nand02 port map ( Y=>gen_6_cmp_BSCmp_op2_16, A0=>nx5474, A1=>
      nx5465);
   ix5475 : nor02_2x port map ( Y=>nx5474, A0=>nx2696, A1=>nx2692);
   ix2697 : nor03_2x port map ( Y=>nx2696, A0=>gen_6_cmp_mReg_15, A1=>
      nx10356, A2=>nx11134);
   ix2693 : nor03_2x port map ( Y=>nx2692, A0=>nx5469, A1=>nx11140, A2=>
      nx11150);
   ix2769 : nand02 port map ( Y=>gen_7_cmp_BSCmp_op2_1, A0=>nx5481, A1=>
      nx5501);
   ix5482 : nor02_2x port map ( Y=>nx5481, A0=>nx2764, A1=>nx2760);
   ix2765 : nor03_2x port map ( Y=>nx2764, A0=>gen_7_cmp_mReg_0, A1=>nx10340, 
      A2=>nx11170);
   gen_7_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_7_cmp_mReg_0, QB=>
      nx5487, D=>window_7_0, CLK=>start, R=>rst);
   ix5492 : inv01 port map ( Y=>nx5491, A=>gen_7_cmp_pMux_0);
   ix2761 : nor03_2x port map ( Y=>nx2760, A0=>nx5487, A1=>nx11176, A2=>
      nx11186);
   ix5500 : inv02 port map ( Y=>nx5499, A=>gen_7_cmp_pMux_2);
   ix5502 : nor02_2x port map ( Y=>nx5501, A0=>nx2750, A1=>nx2748);
   ix2751 : nor03_2x port map ( Y=>nx2750, A0=>nx5505, A1=>nx10334, A2=>
      nx11194);
   gen_7_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_7_cmp_mReg_1, QB=>
      nx5505, D=>window_7_1, CLK=>start, R=>rst);
   ix2749 : nor03_2x port map ( Y=>nx2748, A0=>gen_7_cmp_mReg_1, A1=>nx10772, 
      A2=>nx11202);
   ix2709 : nor03_2x port map ( Y=>nx2708, A0=>nx10340, A1=>nx5499, A2=>
      gen_7_cmp_pMux_0);
   ix2791 : nand02 port map ( Y=>gen_7_cmp_BSCmp_op2_2, A0=>nx5515, A1=>
      nx5519);
   ix5516 : nor02_2x port map ( Y=>nx5515, A0=>nx2786, A1=>nx2782);
   ix2787 : nor03_2x port map ( Y=>nx2786, A0=>gen_7_cmp_mReg_1, A1=>nx10340, 
      A2=>nx11170);
   ix2783 : nor03_2x port map ( Y=>nx2782, A0=>nx5505, A1=>nx11176, A2=>
      nx11186);
   ix5520 : nor02_2x port map ( Y=>nx5519, A0=>nx2778, A1=>nx2776);
   ix2779 : nor03_2x port map ( Y=>nx2778, A0=>nx5523, A1=>nx10334, A2=>
      nx11194);
   gen_7_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_7_cmp_mReg_2, QB=>
      nx5523, D=>window_7_2, CLK=>start, R=>rst);
   ix2777 : nor03_2x port map ( Y=>nx2776, A0=>gen_7_cmp_mReg_2, A1=>nx10772, 
      A2=>nx11202);
   ix2813 : nand02 port map ( Y=>gen_7_cmp_BSCmp_op2_3, A0=>nx5529, A1=>
      nx5533);
   ix5530 : nor02_2x port map ( Y=>nx5529, A0=>nx2808, A1=>nx2804);
   ix2809 : nor03_2x port map ( Y=>nx2808, A0=>gen_7_cmp_mReg_2, A1=>nx10340, 
      A2=>nx11170);
   ix2805 : nor03_2x port map ( Y=>nx2804, A0=>nx5523, A1=>nx11176, A2=>
      nx11186);
   ix5534 : nor02_2x port map ( Y=>nx5533, A0=>nx2800, A1=>nx2798);
   ix2801 : nor03_2x port map ( Y=>nx2800, A0=>nx5537, A1=>nx10334, A2=>
      nx11194);
   gen_7_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_7_cmp_mReg_3, QB=>
      nx5537, D=>window_7_3, CLK=>start, R=>rst);
   ix2799 : nor03_2x port map ( Y=>nx2798, A0=>gen_7_cmp_mReg_3, A1=>nx10772, 
      A2=>nx11202);
   ix2835 : nand02 port map ( Y=>gen_7_cmp_BSCmp_op2_4, A0=>nx5541, A1=>
      nx5547);
   ix5542 : nor02_2x port map ( Y=>nx5541, A0=>nx2830, A1=>nx2826);
   ix2831 : nor03_2x port map ( Y=>nx2830, A0=>gen_7_cmp_mReg_3, A1=>nx10340, 
      A2=>nx11170);
   ix2827 : nor03_2x port map ( Y=>nx2826, A0=>nx5537, A1=>nx11176, A2=>
      nx11186);
   ix5548 : nor02_2x port map ( Y=>nx5547, A0=>nx2822, A1=>nx2820);
   ix2823 : nor03_2x port map ( Y=>nx2822, A0=>nx5551, A1=>nx10334, A2=>
      nx11194);
   gen_7_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_7_cmp_mReg_4, QB=>
      nx5551, D=>window_7_4, CLK=>start, R=>rst);
   ix2821 : nor03_2x port map ( Y=>nx2820, A0=>gen_7_cmp_mReg_4, A1=>nx10772, 
      A2=>nx11202);
   ix2857 : nand02 port map ( Y=>gen_7_cmp_BSCmp_op2_5, A0=>nx5555, A1=>
      nx5561);
   ix5556 : nor02_2x port map ( Y=>nx5555, A0=>nx2852, A1=>nx2848);
   ix2853 : nor03_2x port map ( Y=>nx2852, A0=>gen_7_cmp_mReg_4, A1=>nx10340, 
      A2=>nx11170);
   ix2849 : nor03_2x port map ( Y=>nx2848, A0=>nx5551, A1=>nx11176, A2=>
      nx11186);
   ix5562 : nor02_2x port map ( Y=>nx5561, A0=>nx2844, A1=>nx2842);
   ix2845 : nor03_2x port map ( Y=>nx2844, A0=>nx5564, A1=>nx10336, A2=>
      nx11194);
   gen_7_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_7_cmp_mReg_5, QB=>
      nx5564, D=>window_7_5, CLK=>start, R=>rst);
   ix2843 : nor03_2x port map ( Y=>nx2842, A0=>gen_7_cmp_mReg_5, A1=>nx10772, 
      A2=>nx11202);
   ix2879 : nand02 port map ( Y=>gen_7_cmp_BSCmp_op2_6, A0=>nx5571, A1=>
      nx5577);
   ix5572 : nor02_2x port map ( Y=>nx5571, A0=>nx2874, A1=>nx2870);
   ix2875 : nor03_2x port map ( Y=>nx2874, A0=>gen_7_cmp_mReg_5, A1=>nx10342, 
      A2=>nx11170);
   ix2871 : nor03_2x port map ( Y=>nx2870, A0=>nx5564, A1=>nx11176, A2=>
      nx11186);
   ix5578 : nor02_2x port map ( Y=>nx5577, A0=>nx2866, A1=>nx2864);
   ix2867 : nor03_2x port map ( Y=>nx2866, A0=>nx5581, A1=>nx10336, A2=>
      nx11194);
   gen_7_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_7_cmp_mReg_6, QB=>
      nx5581, D=>window_7_6, CLK=>start, R=>rst);
   ix2865 : nor03_2x port map ( Y=>nx2864, A0=>gen_7_cmp_mReg_6, A1=>nx10772, 
      A2=>nx11202);
   ix2901 : nand02 port map ( Y=>gen_7_cmp_BSCmp_op2_7, A0=>nx5585, A1=>
      nx5591);
   ix5586 : nor02_2x port map ( Y=>nx5585, A0=>nx2896, A1=>nx2892);
   ix2897 : nor03_2x port map ( Y=>nx2896, A0=>gen_7_cmp_mReg_6, A1=>nx10342, 
      A2=>nx11172);
   ix2893 : nor03_2x port map ( Y=>nx2892, A0=>nx5581, A1=>nx11178, A2=>
      nx11188);
   ix5592 : nor02_2x port map ( Y=>nx5591, A0=>nx2888, A1=>nx2886);
   ix2889 : nor03_2x port map ( Y=>nx2888, A0=>nx5595, A1=>nx10336, A2=>
      nx11196);
   gen_7_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_7_cmp_mReg_7, QB=>
      nx5595, D=>window_7_7, CLK=>start, R=>rst);
   ix2887 : nor03_2x port map ( Y=>nx2886, A0=>gen_7_cmp_mReg_7, A1=>nx10772, 
      A2=>nx11204);
   ix2923 : nand02 port map ( Y=>gen_7_cmp_BSCmp_op2_8, A0=>nx5599, A1=>
      nx5605);
   ix5600 : nor02_2x port map ( Y=>nx5599, A0=>nx2918, A1=>nx2914);
   ix2919 : nor03_2x port map ( Y=>nx2918, A0=>gen_7_cmp_mReg_7, A1=>nx10342, 
      A2=>nx11172);
   ix2915 : nor03_2x port map ( Y=>nx2914, A0=>nx5595, A1=>nx11178, A2=>
      nx11188);
   ix5606 : nor02_2x port map ( Y=>nx5605, A0=>nx2910, A1=>nx2908);
   ix2911 : nor03_2x port map ( Y=>nx2910, A0=>nx5608, A1=>nx10336, A2=>
      nx11196);
   gen_7_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_7_cmp_mReg_8, QB=>
      nx5608, D=>window_7_8, CLK=>start, R=>rst);
   ix2909 : nor03_2x port map ( Y=>nx2908, A0=>gen_7_cmp_mReg_8, A1=>nx10774, 
      A2=>nx11204);
   ix2945 : nand02 port map ( Y=>gen_7_cmp_BSCmp_op2_9, A0=>nx5615, A1=>
      nx5621);
   ix5616 : nor02_2x port map ( Y=>nx5615, A0=>nx2940, A1=>nx2936);
   ix2941 : nor03_2x port map ( Y=>nx2940, A0=>gen_7_cmp_mReg_8, A1=>nx10342, 
      A2=>nx11172);
   ix2937 : nor03_2x port map ( Y=>nx2936, A0=>nx5608, A1=>nx11178, A2=>
      nx11188);
   ix5622 : nor02_2x port map ( Y=>nx5621, A0=>nx2932, A1=>nx2930);
   ix2933 : nor03_2x port map ( Y=>nx2932, A0=>nx5625, A1=>nx10336, A2=>
      nx11196);
   gen_7_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_7_cmp_mReg_9, QB=>
      nx5625, D=>window_7_9, CLK=>start, R=>rst);
   ix2931 : nor03_2x port map ( Y=>nx2930, A0=>gen_7_cmp_mReg_9, A1=>nx10774, 
      A2=>nx11204);
   ix2967 : nand02 port map ( Y=>gen_7_cmp_BSCmp_op2_10, A0=>nx5629, A1=>
      nx5635);
   ix5630 : nor02_2x port map ( Y=>nx5629, A0=>nx2962, A1=>nx2958);
   ix2963 : nor03_2x port map ( Y=>nx2962, A0=>gen_7_cmp_mReg_9, A1=>nx10342, 
      A2=>nx11172);
   ix2959 : nor03_2x port map ( Y=>nx2958, A0=>nx5625, A1=>nx11178, A2=>
      nx11188);
   ix5636 : nor02_2x port map ( Y=>nx5635, A0=>nx2954, A1=>nx2952);
   ix2955 : nor03_2x port map ( Y=>nx2954, A0=>nx5639, A1=>nx10336, A2=>
      nx11196);
   gen_7_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_7_cmp_mReg_10, QB=>
      nx5639, D=>window_7_10, CLK=>start, R=>rst);
   ix2953 : nor03_2x port map ( Y=>nx2952, A0=>gen_7_cmp_mReg_10, A1=>
      nx10774, A2=>nx11204);
   ix2989 : nand02 port map ( Y=>gen_7_cmp_BSCmp_op2_11, A0=>nx5643, A1=>
      nx5649);
   ix5644 : nor02_2x port map ( Y=>nx5643, A0=>nx2984, A1=>nx2980);
   ix2985 : nor03_2x port map ( Y=>nx2984, A0=>gen_7_cmp_mReg_10, A1=>
      nx10342, A2=>nx11172);
   ix2981 : nor03_2x port map ( Y=>nx2980, A0=>nx5639, A1=>nx11178, A2=>
      nx11188);
   ix5650 : nor02_2x port map ( Y=>nx5649, A0=>nx2976, A1=>nx2974);
   ix2977 : nor03_2x port map ( Y=>nx2976, A0=>nx5652, A1=>nx10336, A2=>
      nx11196);
   gen_7_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_7_cmp_mReg_11, QB=>
      nx5652, D=>window_7_11, CLK=>start, R=>rst);
   ix2975 : nor03_2x port map ( Y=>nx2974, A0=>gen_7_cmp_mReg_11, A1=>
      nx10774, A2=>nx11204);
   ix3011 : nand02 port map ( Y=>gen_7_cmp_BSCmp_op2_12, A0=>nx5659, A1=>
      nx5665);
   ix5660 : nor02_2x port map ( Y=>nx5659, A0=>nx3006, A1=>nx3002);
   ix3007 : nor03_2x port map ( Y=>nx3006, A0=>gen_7_cmp_mReg_11, A1=>
      nx10342, A2=>nx11172);
   ix3003 : nor03_2x port map ( Y=>nx3002, A0=>nx5652, A1=>nx11178, A2=>
      nx11188);
   ix5666 : nor02_2x port map ( Y=>nx5665, A0=>nx2998, A1=>nx2996);
   ix2999 : nor03_2x port map ( Y=>nx2998, A0=>nx5669, A1=>nx10338, A2=>
      nx11196);
   gen_7_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_7_cmp_mReg_12, QB=>
      nx5669, D=>window_7_12, CLK=>start, R=>rst);
   ix2997 : nor03_2x port map ( Y=>nx2996, A0=>gen_7_cmp_mReg_12, A1=>
      nx10774, A2=>nx11204);
   ix3033 : nand02 port map ( Y=>gen_7_cmp_BSCmp_op2_13, A0=>nx5673, A1=>
      nx5679);
   ix5674 : nor02_2x port map ( Y=>nx5673, A0=>nx3028, A1=>nx3024);
   ix3029 : nor03_2x port map ( Y=>nx3028, A0=>gen_7_cmp_mReg_12, A1=>
      nx10344, A2=>nx11174);
   ix3025 : nor03_2x port map ( Y=>nx3024, A0=>nx5669, A1=>nx11178, A2=>
      nx11190);
   ix5680 : nor02_2x port map ( Y=>nx5679, A0=>nx3020, A1=>nx3018);
   ix3021 : nor03_2x port map ( Y=>nx3020, A0=>nx5683, A1=>nx10338, A2=>
      nx11198);
   gen_7_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_7_cmp_mReg_13, QB=>
      nx5683, D=>window_7_13, CLK=>start, R=>rst);
   ix3019 : nor03_2x port map ( Y=>nx3018, A0=>gen_7_cmp_mReg_13, A1=>
      nx10774, A2=>nx11206);
   ix3055 : nand02 port map ( Y=>gen_7_cmp_BSCmp_op2_14, A0=>nx5687, A1=>
      nx5693);
   ix5688 : nor02_2x port map ( Y=>nx5687, A0=>nx3050, A1=>nx3046);
   ix3051 : nor03_2x port map ( Y=>nx3050, A0=>gen_7_cmp_mReg_13, A1=>
      nx10344, A2=>nx11174);
   ix3047 : nor03_2x port map ( Y=>nx3046, A0=>nx5683, A1=>nx11180, A2=>
      nx11190);
   ix5694 : nor02_2x port map ( Y=>nx5693, A0=>nx3042, A1=>nx3040);
   ix3043 : nor03_2x port map ( Y=>nx3042, A0=>nx5696, A1=>nx10338, A2=>
      nx11198);
   gen_7_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_7_cmp_mReg_14, QB=>
      nx5696, D=>window_7_14, CLK=>start, R=>rst);
   ix3041 : nor03_2x port map ( Y=>nx3040, A0=>gen_7_cmp_mReg_14, A1=>
      nx10774, A2=>nx11206);
   ix3077 : nand02 port map ( Y=>gen_7_cmp_BSCmp_op2_15, A0=>nx5703, A1=>
      nx5709);
   ix5704 : nor02_2x port map ( Y=>nx5703, A0=>nx3072, A1=>nx3068);
   ix3073 : nor03_2x port map ( Y=>nx3072, A0=>gen_7_cmp_mReg_14, A1=>
      nx10344, A2=>nx11174);
   ix3069 : nor03_2x port map ( Y=>nx3068, A0=>nx5696, A1=>nx11180, A2=>
      nx11190);
   ix5710 : nor02_2x port map ( Y=>nx5709, A0=>nx3064, A1=>nx3062);
   ix3065 : nor03_2x port map ( Y=>nx3064, A0=>nx5713, A1=>nx10338, A2=>
      nx11198);
   gen_7_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_7_cmp_mReg_15, QB=>
      nx5713, D=>window_7_15, CLK=>start, R=>rst);
   ix3063 : nor03_2x port map ( Y=>nx3062, A0=>gen_7_cmp_mReg_15, A1=>
      nx10776, A2=>nx11206);
   ix3087 : nand02 port map ( Y=>gen_7_cmp_BSCmp_op2_16, A0=>nx5717, A1=>
      nx5709);
   ix5718 : nor02_2x port map ( Y=>nx5717, A0=>nx3082, A1=>nx3078);
   ix3083 : nor03_2x port map ( Y=>nx3082, A0=>gen_7_cmp_mReg_15, A1=>
      nx10344, A2=>nx11174);
   ix3079 : nor03_2x port map ( Y=>nx3078, A0=>nx5713, A1=>nx11180, A2=>
      nx11190);
   ix3155 : nand02 port map ( Y=>gen_8_cmp_BSCmp_op2_1, A0=>nx5725, A1=>
      nx5745);
   ix5726 : nor02_2x port map ( Y=>nx5725, A0=>nx3150, A1=>nx3146);
   ix3151 : nor03_2x port map ( Y=>nx3150, A0=>gen_8_cmp_mReg_0, A1=>nx10328, 
      A2=>nx11210);
   gen_8_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_8_cmp_mReg_0, QB=>
      nx5731, D=>window_8_0, CLK=>start, R=>rst);
   ix5736 : inv01 port map ( Y=>nx5735, A=>gen_8_cmp_pMux_0);
   ix3147 : nor03_2x port map ( Y=>nx3146, A0=>nx5731, A1=>nx11216, A2=>
      nx11226);
   ix5744 : inv02 port map ( Y=>nx5743, A=>gen_8_cmp_pMux_2);
   ix5746 : nor02_2x port map ( Y=>nx5745, A0=>nx3136, A1=>nx3134);
   ix3137 : nor03_2x port map ( Y=>nx3136, A0=>nx5749, A1=>nx10322, A2=>
      nx11234);
   gen_8_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_8_cmp_mReg_1, QB=>
      nx5749, D=>window_8_1, CLK=>start, R=>rst);
   ix3135 : nor03_2x port map ( Y=>nx3134, A0=>gen_8_cmp_mReg_1, A1=>nx10778, 
      A2=>nx11242);
   ix3095 : nor03_2x port map ( Y=>nx3094, A0=>nx10328, A1=>nx5743, A2=>
      gen_8_cmp_pMux_0);
   ix3177 : nand02 port map ( Y=>gen_8_cmp_BSCmp_op2_2, A0=>nx5760, A1=>
      nx5765);
   ix5761 : nor02_2x port map ( Y=>nx5760, A0=>nx3172, A1=>nx3168);
   ix3173 : nor03_2x port map ( Y=>nx3172, A0=>gen_8_cmp_mReg_1, A1=>nx10328, 
      A2=>nx11210);
   ix3169 : nor03_2x port map ( Y=>nx3168, A0=>nx5749, A1=>nx11216, A2=>
      nx11226);
   ix5766 : nor02_2x port map ( Y=>nx5765, A0=>nx3164, A1=>nx3162);
   ix3165 : nor03_2x port map ( Y=>nx3164, A0=>nx5769, A1=>nx10322, A2=>
      nx11234);
   gen_8_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_8_cmp_mReg_2, QB=>
      nx5769, D=>window_8_2, CLK=>start, R=>rst);
   ix3163 : nor03_2x port map ( Y=>nx3162, A0=>gen_8_cmp_mReg_2, A1=>nx10778, 
      A2=>nx11242);
   ix3199 : nand02 port map ( Y=>gen_8_cmp_BSCmp_op2_3, A0=>nx5775, A1=>
      nx5781);
   ix5776 : nor02_2x port map ( Y=>nx5775, A0=>nx3194, A1=>nx3190);
   ix3195 : nor03_2x port map ( Y=>nx3194, A0=>gen_8_cmp_mReg_2, A1=>nx10328, 
      A2=>nx11210);
   ix3191 : nor03_2x port map ( Y=>nx3190, A0=>nx5769, A1=>nx11216, A2=>
      nx11226);
   ix5782 : nor02_2x port map ( Y=>nx5781, A0=>nx3186, A1=>nx3184);
   ix3187 : nor03_2x port map ( Y=>nx3186, A0=>nx5785, A1=>nx10322, A2=>
      nx11234);
   gen_8_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_8_cmp_mReg_3, QB=>
      nx5785, D=>window_8_3, CLK=>start, R=>rst);
   ix3185 : nor03_2x port map ( Y=>nx3184, A0=>gen_8_cmp_mReg_3, A1=>nx10778, 
      A2=>nx11242);
   ix3221 : nand02 port map ( Y=>gen_8_cmp_BSCmp_op2_4, A0=>nx5791, A1=>
      nx5797);
   ix5792 : nor02_2x port map ( Y=>nx5791, A0=>nx3216, A1=>nx3212);
   ix3217 : nor03_2x port map ( Y=>nx3216, A0=>gen_8_cmp_mReg_3, A1=>nx10328, 
      A2=>nx11210);
   ix3213 : nor03_2x port map ( Y=>nx3212, A0=>nx5785, A1=>nx11216, A2=>
      nx11226);
   ix5798 : nor02_2x port map ( Y=>nx5797, A0=>nx3208, A1=>nx3206);
   ix3209 : nor03_2x port map ( Y=>nx3208, A0=>nx5800, A1=>nx10322, A2=>
      nx11234);
   gen_8_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_8_cmp_mReg_4, QB=>
      nx5800, D=>window_8_4, CLK=>start, R=>rst);
   ix3207 : nor03_2x port map ( Y=>nx3206, A0=>gen_8_cmp_mReg_4, A1=>nx10778, 
      A2=>nx11242);
   ix3243 : nand02 port map ( Y=>gen_8_cmp_BSCmp_op2_5, A0=>nx5804, A1=>
      nx5809);
   ix5805 : nor02_2x port map ( Y=>nx5804, A0=>nx3238, A1=>nx3234);
   ix3239 : nor03_2x port map ( Y=>nx3238, A0=>gen_8_cmp_mReg_4, A1=>nx10328, 
      A2=>nx11210);
   ix3235 : nor03_2x port map ( Y=>nx3234, A0=>nx5800, A1=>nx11216, A2=>
      nx11226);
   ix5810 : nor02_2x port map ( Y=>nx5809, A0=>nx3230, A1=>nx3228);
   ix3231 : nor03_2x port map ( Y=>nx3230, A0=>nx5813, A1=>nx10324, A2=>
      nx11234);
   gen_8_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_8_cmp_mReg_5, QB=>
      nx5813, D=>window_8_5, CLK=>start, R=>rst);
   ix3229 : nor03_2x port map ( Y=>nx3228, A0=>gen_8_cmp_mReg_5, A1=>nx10778, 
      A2=>nx11242);
   ix3265 : nand02 port map ( Y=>gen_8_cmp_BSCmp_op2_6, A0=>nx5819, A1=>
      nx5825);
   ix5820 : nor02_2x port map ( Y=>nx5819, A0=>nx3260, A1=>nx3256);
   ix3261 : nor03_2x port map ( Y=>nx3260, A0=>gen_8_cmp_mReg_5, A1=>nx10330, 
      A2=>nx11210);
   ix3257 : nor03_2x port map ( Y=>nx3256, A0=>nx5813, A1=>nx11216, A2=>
      nx11226);
   ix5826 : nor02_2x port map ( Y=>nx5825, A0=>nx3252, A1=>nx3250);
   ix3253 : nor03_2x port map ( Y=>nx3252, A0=>nx5829, A1=>nx10324, A2=>
      nx11234);
   gen_8_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_8_cmp_mReg_6, QB=>
      nx5829, D=>window_8_6, CLK=>start, R=>rst);
   ix3251 : nor03_2x port map ( Y=>nx3250, A0=>gen_8_cmp_mReg_6, A1=>nx10778, 
      A2=>nx11242);
   ix3287 : nand02 port map ( Y=>gen_8_cmp_BSCmp_op2_7, A0=>nx5833, A1=>
      nx5839);
   ix5834 : nor02_2x port map ( Y=>nx5833, A0=>nx3282, A1=>nx3278);
   ix3283 : nor03_2x port map ( Y=>nx3282, A0=>gen_8_cmp_mReg_6, A1=>nx10330, 
      A2=>nx11212);
   ix3279 : nor03_2x port map ( Y=>nx3278, A0=>nx5829, A1=>nx11218, A2=>
      nx11228);
   ix5840 : nor02_2x port map ( Y=>nx5839, A0=>nx3274, A1=>nx3272);
   ix3275 : nor03_2x port map ( Y=>nx3274, A0=>nx5843, A1=>nx10324, A2=>
      nx11236);
   gen_8_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_8_cmp_mReg_7, QB=>
      nx5843, D=>window_8_7, CLK=>start, R=>rst);
   ix3273 : nor03_2x port map ( Y=>nx3272, A0=>gen_8_cmp_mReg_7, A1=>nx10778, 
      A2=>nx11244);
   ix3309 : nand02 port map ( Y=>gen_8_cmp_BSCmp_op2_8, A0=>nx5849, A1=>
      nx5853);
   ix5850 : nor02_2x port map ( Y=>nx5849, A0=>nx3304, A1=>nx3300);
   ix3305 : nor03_2x port map ( Y=>nx3304, A0=>gen_8_cmp_mReg_7, A1=>nx10330, 
      A2=>nx11212);
   ix3301 : nor03_2x port map ( Y=>nx3300, A0=>nx5843, A1=>nx11218, A2=>
      nx11228);
   ix5854 : nor02_2x port map ( Y=>nx5853, A0=>nx3296, A1=>nx3294);
   ix3297 : nor03_2x port map ( Y=>nx3296, A0=>nx5857, A1=>nx10324, A2=>
      nx11236);
   gen_8_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_8_cmp_mReg_8, QB=>
      nx5857, D=>window_8_8, CLK=>start, R=>rst);
   ix3295 : nor03_2x port map ( Y=>nx3294, A0=>gen_8_cmp_mReg_8, A1=>nx10780, 
      A2=>nx11244);
   ix3331 : nand02 port map ( Y=>gen_8_cmp_BSCmp_op2_9, A0=>nx5861, A1=>
      nx5867);
   ix5862 : nor02_2x port map ( Y=>nx5861, A0=>nx3326, A1=>nx3322);
   ix3327 : nor03_2x port map ( Y=>nx3326, A0=>gen_8_cmp_mReg_8, A1=>nx10330, 
      A2=>nx11212);
   ix3323 : nor03_2x port map ( Y=>nx3322, A0=>nx5857, A1=>nx11218, A2=>
      nx11228);
   ix5868 : nor02_2x port map ( Y=>nx5867, A0=>nx3318, A1=>nx3316);
   ix3319 : nor03_2x port map ( Y=>nx3318, A0=>nx5871, A1=>nx10324, A2=>
      nx11236);
   gen_8_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_8_cmp_mReg_9, QB=>
      nx5871, D=>window_8_9, CLK=>start, R=>rst);
   ix3317 : nor03_2x port map ( Y=>nx3316, A0=>gen_8_cmp_mReg_9, A1=>nx10780, 
      A2=>nx11244);
   ix3353 : nand02 port map ( Y=>gen_8_cmp_BSCmp_op2_10, A0=>nx5875, A1=>
      nx5881);
   ix5876 : nor02_2x port map ( Y=>nx5875, A0=>nx3348, A1=>nx3344);
   ix3349 : nor03_2x port map ( Y=>nx3348, A0=>gen_8_cmp_mReg_9, A1=>nx10330, 
      A2=>nx11212);
   ix3345 : nor03_2x port map ( Y=>nx3344, A0=>nx5871, A1=>nx11218, A2=>
      nx11228);
   ix5882 : nor02_2x port map ( Y=>nx5881, A0=>nx3340, A1=>nx3338);
   ix3341 : nor03_2x port map ( Y=>nx3340, A0=>nx5884, A1=>nx10324, A2=>
      nx11236);
   gen_8_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_8_cmp_mReg_10, QB=>
      nx5884, D=>window_8_10, CLK=>start, R=>rst);
   ix3339 : nor03_2x port map ( Y=>nx3338, A0=>gen_8_cmp_mReg_10, A1=>
      nx10780, A2=>nx11244);
   ix3375 : nand02 port map ( Y=>gen_8_cmp_BSCmp_op2_11, A0=>nx5891, A1=>
      nx5897);
   ix5892 : nor02_2x port map ( Y=>nx5891, A0=>nx3370, A1=>nx3366);
   ix3371 : nor03_2x port map ( Y=>nx3370, A0=>gen_8_cmp_mReg_10, A1=>
      nx10330, A2=>nx11212);
   ix3367 : nor03_2x port map ( Y=>nx3366, A0=>nx5884, A1=>nx11218, A2=>
      nx11228);
   ix5898 : nor02_2x port map ( Y=>nx5897, A0=>nx3362, A1=>nx3360);
   ix3363 : nor03_2x port map ( Y=>nx3362, A0=>nx5901, A1=>nx10324, A2=>
      nx11236);
   gen_8_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_8_cmp_mReg_11, QB=>
      nx5901, D=>window_8_11, CLK=>start, R=>rst);
   ix3361 : nor03_2x port map ( Y=>nx3360, A0=>gen_8_cmp_mReg_11, A1=>
      nx10780, A2=>nx11244);
   ix3397 : nand02 port map ( Y=>gen_8_cmp_BSCmp_op2_12, A0=>nx5905, A1=>
      nx5911);
   ix5906 : nor02_2x port map ( Y=>nx5905, A0=>nx3392, A1=>nx3388);
   ix3393 : nor03_2x port map ( Y=>nx3392, A0=>gen_8_cmp_mReg_11, A1=>
      nx10330, A2=>nx11212);
   ix3389 : nor03_2x port map ( Y=>nx3388, A0=>nx5901, A1=>nx11218, A2=>
      nx11228);
   ix5912 : nor02_2x port map ( Y=>nx5911, A0=>nx3384, A1=>nx3382);
   ix3385 : nor03_2x port map ( Y=>nx3384, A0=>nx5915, A1=>nx10326, A2=>
      nx11236);
   gen_8_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_8_cmp_mReg_12, QB=>
      nx5915, D=>window_8_12, CLK=>start, R=>rst);
   ix3383 : nor03_2x port map ( Y=>nx3382, A0=>gen_8_cmp_mReg_12, A1=>
      nx10780, A2=>nx11244);
   ix3419 : nand02 port map ( Y=>gen_8_cmp_BSCmp_op2_13, A0=>nx5919, A1=>
      nx5925);
   ix5920 : nor02_2x port map ( Y=>nx5919, A0=>nx3414, A1=>nx3410);
   ix3415 : nor03_2x port map ( Y=>nx3414, A0=>gen_8_cmp_mReg_12, A1=>
      nx10332, A2=>nx11214);
   ix3411 : nor03_2x port map ( Y=>nx3410, A0=>nx5915, A1=>nx11218, A2=>
      nx11230);
   ix5926 : nor02_2x port map ( Y=>nx5925, A0=>nx3406, A1=>nx3404);
   ix3407 : nor03_2x port map ( Y=>nx3406, A0=>nx5928, A1=>nx10326, A2=>
      nx11238);
   gen_8_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_8_cmp_mReg_13, QB=>
      nx5928, D=>window_8_13, CLK=>start, R=>rst);
   ix3405 : nor03_2x port map ( Y=>nx3404, A0=>gen_8_cmp_mReg_13, A1=>
      nx10780, A2=>nx11246);
   ix3441 : nand02 port map ( Y=>gen_8_cmp_BSCmp_op2_14, A0=>nx5935, A1=>
      nx5941);
   ix5936 : nor02_2x port map ( Y=>nx5935, A0=>nx3436, A1=>nx3432);
   ix3437 : nor03_2x port map ( Y=>nx3436, A0=>gen_8_cmp_mReg_13, A1=>
      nx10332, A2=>nx11214);
   ix3433 : nor03_2x port map ( Y=>nx3432, A0=>nx5928, A1=>nx11220, A2=>
      nx11230);
   ix5942 : nor02_2x port map ( Y=>nx5941, A0=>nx3428, A1=>nx3426);
   ix3429 : nor03_2x port map ( Y=>nx3428, A0=>nx5945, A1=>nx10326, A2=>
      nx11238);
   gen_8_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_8_cmp_mReg_14, QB=>
      nx5945, D=>window_8_14, CLK=>start, R=>rst);
   ix3427 : nor03_2x port map ( Y=>nx3426, A0=>gen_8_cmp_mReg_14, A1=>
      nx10780, A2=>nx11246);
   ix3463 : nand02 port map ( Y=>gen_8_cmp_BSCmp_op2_15, A0=>nx5949, A1=>
      nx5955);
   ix5950 : nor02_2x port map ( Y=>nx5949, A0=>nx3458, A1=>nx3454);
   ix3459 : nor03_2x port map ( Y=>nx3458, A0=>gen_8_cmp_mReg_14, A1=>
      nx10332, A2=>nx11214);
   ix3455 : nor03_2x port map ( Y=>nx3454, A0=>nx5945, A1=>nx11220, A2=>
      nx11230);
   ix5956 : nor02_2x port map ( Y=>nx5955, A0=>nx3450, A1=>nx3448);
   ix3451 : nor03_2x port map ( Y=>nx3450, A0=>nx5959, A1=>nx10326, A2=>
      nx11238);
   gen_8_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_8_cmp_mReg_15, QB=>
      nx5959, D=>window_8_15, CLK=>start, R=>rst);
   ix3449 : nor03_2x port map ( Y=>nx3448, A0=>gen_8_cmp_mReg_15, A1=>
      nx10782, A2=>nx11246);
   ix3473 : nand02 port map ( Y=>gen_8_cmp_BSCmp_op2_16, A0=>nx5963, A1=>
      nx5955);
   ix5964 : nor02_2x port map ( Y=>nx5963, A0=>nx3468, A1=>nx3464);
   ix3469 : nor03_2x port map ( Y=>nx3468, A0=>gen_8_cmp_mReg_15, A1=>
      nx10332, A2=>nx11214);
   ix3465 : nor03_2x port map ( Y=>nx3464, A0=>nx5959, A1=>nx11220, A2=>
      nx11230);
   ix3541 : nand02 port map ( Y=>gen_9_cmp_BSCmp_op2_1, A0=>nx5970, A1=>
      nx5989);
   ix5971 : nor02_2x port map ( Y=>nx5970, A0=>nx3536, A1=>nx3532);
   ix3537 : nor03_2x port map ( Y=>nx3536, A0=>gen_9_cmp_mReg_0, A1=>nx10316, 
      A2=>nx11250);
   gen_9_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_9_cmp_mReg_0, QB=>
      nx5975, D=>window_9_0, CLK=>start, R=>rst);
   ix5980 : inv01 port map ( Y=>nx5979, A=>gen_9_cmp_pMux_0);
   ix3533 : nor03_2x port map ( Y=>nx3532, A0=>nx5975, A1=>nx11256, A2=>
      nx11266);
   ix5988 : inv02 port map ( Y=>nx5987, A=>gen_9_cmp_pMux_2);
   ix5990 : nor02_2x port map ( Y=>nx5989, A0=>nx3522, A1=>nx3520);
   ix3523 : nor03_2x port map ( Y=>nx3522, A0=>nx5992, A1=>nx10310, A2=>
      nx11274);
   gen_9_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_9_cmp_mReg_1, QB=>
      nx5992, D=>window_9_1, CLK=>start, R=>rst);
   ix3521 : nor03_2x port map ( Y=>nx3520, A0=>gen_9_cmp_mReg_1, A1=>nx10784, 
      A2=>nx11282);
   ix3481 : nor03_2x port map ( Y=>nx3480, A0=>nx10316, A1=>nx5987, A2=>
      gen_9_cmp_pMux_0);
   ix3563 : nand02 port map ( Y=>gen_9_cmp_BSCmp_op2_2, A0=>nx6005, A1=>
      nx6011);
   ix6006 : nor02_2x port map ( Y=>nx6005, A0=>nx3558, A1=>nx3554);
   ix3559 : nor03_2x port map ( Y=>nx3558, A0=>gen_9_cmp_mReg_1, A1=>nx10316, 
      A2=>nx11250);
   ix3555 : nor03_2x port map ( Y=>nx3554, A0=>nx5992, A1=>nx11256, A2=>
      nx11266);
   ix6012 : nor02_2x port map ( Y=>nx6011, A0=>nx3550, A1=>nx3548);
   ix3551 : nor03_2x port map ( Y=>nx3550, A0=>nx6014, A1=>nx10310, A2=>
      nx11274);
   gen_9_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_9_cmp_mReg_2, QB=>
      nx6014, D=>window_9_2, CLK=>start, R=>rst);
   ix3549 : nor03_2x port map ( Y=>nx3548, A0=>gen_9_cmp_mReg_2, A1=>nx10784, 
      A2=>nx11282);
   ix3585 : nand02 port map ( Y=>gen_9_cmp_BSCmp_op2_3, A0=>nx6019, A1=>
      nx6025);
   ix6020 : nor02_2x port map ( Y=>nx6019, A0=>nx3580, A1=>nx3576);
   ix3581 : nor03_2x port map ( Y=>nx3580, A0=>gen_9_cmp_mReg_2, A1=>nx10316, 
      A2=>nx11250);
   ix3577 : nor03_2x port map ( Y=>nx3576, A0=>nx6014, A1=>nx11256, A2=>
      nx11266);
   ix6026 : nor02_2x port map ( Y=>nx6025, A0=>nx3572, A1=>nx3570);
   ix3573 : nor03_2x port map ( Y=>nx3572, A0=>nx6029, A1=>nx10310, A2=>
      nx11274);
   gen_9_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_9_cmp_mReg_3, QB=>
      nx6029, D=>window_9_3, CLK=>start, R=>rst);
   ix3571 : nor03_2x port map ( Y=>nx3570, A0=>gen_9_cmp_mReg_3, A1=>nx10784, 
      A2=>nx11282);
   ix3607 : nand02 port map ( Y=>gen_9_cmp_BSCmp_op2_4, A0=>nx6035, A1=>
      nx6039);
   ix6036 : nor02_2x port map ( Y=>nx6035, A0=>nx3602, A1=>nx3598);
   ix3603 : nor03_2x port map ( Y=>nx3602, A0=>gen_9_cmp_mReg_3, A1=>nx10316, 
      A2=>nx11250);
   ix3599 : nor03_2x port map ( Y=>nx3598, A0=>nx6029, A1=>nx11256, A2=>
      nx11266);
   ix6040 : nor02_2x port map ( Y=>nx6039, A0=>nx3594, A1=>nx3592);
   ix3595 : nor03_2x port map ( Y=>nx3594, A0=>nx6043, A1=>nx10310, A2=>
      nx11274);
   gen_9_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_9_cmp_mReg_4, QB=>
      nx6043, D=>window_9_4, CLK=>start, R=>rst);
   ix3593 : nor03_2x port map ( Y=>nx3592, A0=>gen_9_cmp_mReg_4, A1=>nx10784, 
      A2=>nx11282);
   ix3629 : nand02 port map ( Y=>gen_9_cmp_BSCmp_op2_5, A0=>nx6049, A1=>
      nx6055);
   ix6050 : nor02_2x port map ( Y=>nx6049, A0=>nx3624, A1=>nx3620);
   ix3625 : nor03_2x port map ( Y=>nx3624, A0=>gen_9_cmp_mReg_4, A1=>nx10316, 
      A2=>nx11250);
   ix3621 : nor03_2x port map ( Y=>nx3620, A0=>nx6043, A1=>nx11256, A2=>
      nx11266);
   ix6056 : nor02_2x port map ( Y=>nx6055, A0=>nx3616, A1=>nx3614);
   ix3617 : nor03_2x port map ( Y=>nx3616, A0=>nx6058, A1=>nx10312, A2=>
      nx11274);
   gen_9_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_9_cmp_mReg_5, QB=>
      nx6058, D=>window_9_5, CLK=>start, R=>rst);
   ix3615 : nor03_2x port map ( Y=>nx3614, A0=>gen_9_cmp_mReg_5, A1=>nx10784, 
      A2=>nx11282);
   ix3651 : nand02 port map ( Y=>gen_9_cmp_BSCmp_op2_6, A0=>nx6063, A1=>
      nx6069);
   ix6064 : nor02_2x port map ( Y=>nx6063, A0=>nx3646, A1=>nx3642);
   ix3647 : nor03_2x port map ( Y=>nx3646, A0=>gen_9_cmp_mReg_5, A1=>nx10318, 
      A2=>nx11250);
   ix3643 : nor03_2x port map ( Y=>nx3642, A0=>nx6058, A1=>nx11256, A2=>
      nx11266);
   ix6070 : nor02_2x port map ( Y=>nx6069, A0=>nx3638, A1=>nx3636);
   ix3639 : nor03_2x port map ( Y=>nx3638, A0=>nx6073, A1=>nx10312, A2=>
      nx11274);
   gen_9_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_9_cmp_mReg_6, QB=>
      nx6073, D=>window_9_6, CLK=>start, R=>rst);
   ix3637 : nor03_2x port map ( Y=>nx3636, A0=>gen_9_cmp_mReg_6, A1=>nx10784, 
      A2=>nx11282);
   ix3673 : nand02 port map ( Y=>gen_9_cmp_BSCmp_op2_7, A0=>nx6079, A1=>
      nx6083);
   ix6080 : nor02_2x port map ( Y=>nx6079, A0=>nx3668, A1=>nx3664);
   ix3669 : nor03_2x port map ( Y=>nx3668, A0=>gen_9_cmp_mReg_6, A1=>nx10318, 
      A2=>nx11252);
   ix3665 : nor03_2x port map ( Y=>nx3664, A0=>nx6073, A1=>nx11258, A2=>
      nx11268);
   ix6084 : nor02_2x port map ( Y=>nx6083, A0=>nx3660, A1=>nx3658);
   ix3661 : nor03_2x port map ( Y=>nx3660, A0=>nx6087, A1=>nx10312, A2=>
      nx11276);
   gen_9_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_9_cmp_mReg_7, QB=>
      nx6087, D=>window_9_7, CLK=>start, R=>rst);
   ix3659 : nor03_2x port map ( Y=>nx3658, A0=>gen_9_cmp_mReg_7, A1=>nx10784, 
      A2=>nx11284);
   ix3695 : nand02 port map ( Y=>gen_9_cmp_BSCmp_op2_8, A0=>nx6093, A1=>
      nx6099);
   ix6094 : nor02_2x port map ( Y=>nx6093, A0=>nx3690, A1=>nx3686);
   ix3691 : nor03_2x port map ( Y=>nx3690, A0=>gen_9_cmp_mReg_7, A1=>nx10318, 
      A2=>nx11252);
   ix3687 : nor03_2x port map ( Y=>nx3686, A0=>nx6087, A1=>nx11258, A2=>
      nx11268);
   ix6100 : nor02_2x port map ( Y=>nx6099, A0=>nx3682, A1=>nx3680);
   ix3683 : nor03_2x port map ( Y=>nx3682, A0=>nx6102, A1=>nx10312, A2=>
      nx11276);
   gen_9_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_9_cmp_mReg_8, QB=>
      nx6102, D=>window_9_8, CLK=>start, R=>rst);
   ix3681 : nor03_2x port map ( Y=>nx3680, A0=>gen_9_cmp_mReg_8, A1=>nx10786, 
      A2=>nx11284);
   ix3717 : nand02 port map ( Y=>gen_9_cmp_BSCmp_op2_9, A0=>nx6107, A1=>
      nx6113);
   ix6108 : nor02_2x port map ( Y=>nx6107, A0=>nx3712, A1=>nx3708);
   ix3713 : nor03_2x port map ( Y=>nx3712, A0=>gen_9_cmp_mReg_8, A1=>nx10318, 
      A2=>nx11252);
   ix3709 : nor03_2x port map ( Y=>nx3708, A0=>nx6102, A1=>nx11258, A2=>
      nx11268);
   ix6114 : nor02_2x port map ( Y=>nx6113, A0=>nx3704, A1=>nx3702);
   ix3705 : nor03_2x port map ( Y=>nx3704, A0=>nx6117, A1=>nx10312, A2=>
      nx11276);
   gen_9_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_9_cmp_mReg_9, QB=>
      nx6117, D=>window_9_9, CLK=>start, R=>rst);
   ix3703 : nor03_2x port map ( Y=>nx3702, A0=>gen_9_cmp_mReg_9, A1=>nx10786, 
      A2=>nx11284);
   ix3739 : nand02 port map ( Y=>gen_9_cmp_BSCmp_op2_10, A0=>nx6123, A1=>
      nx6127);
   ix6124 : nor02_2x port map ( Y=>nx6123, A0=>nx3734, A1=>nx3730);
   ix3735 : nor03_2x port map ( Y=>nx3734, A0=>gen_9_cmp_mReg_9, A1=>nx10318, 
      A2=>nx11252);
   ix3731 : nor03_2x port map ( Y=>nx3730, A0=>nx6117, A1=>nx11258, A2=>
      nx11268);
   ix6128 : nor02_2x port map ( Y=>nx6127, A0=>nx3726, A1=>nx3724);
   ix3727 : nor03_2x port map ( Y=>nx3726, A0=>nx6131, A1=>nx10312, A2=>
      nx11276);
   gen_9_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_9_cmp_mReg_10, QB=>
      nx6131, D=>window_9_10, CLK=>start, R=>rst);
   ix3725 : nor03_2x port map ( Y=>nx3724, A0=>gen_9_cmp_mReg_10, A1=>
      nx10786, A2=>nx11284);
   ix3761 : nand02 port map ( Y=>gen_9_cmp_BSCmp_op2_11, A0=>nx6137, A1=>
      nx6143);
   ix6138 : nor02_2x port map ( Y=>nx6137, A0=>nx3756, A1=>nx3752);
   ix3757 : nor03_2x port map ( Y=>nx3756, A0=>gen_9_cmp_mReg_10, A1=>
      nx10318, A2=>nx11252);
   ix3753 : nor03_2x port map ( Y=>nx3752, A0=>nx6131, A1=>nx11258, A2=>
      nx11268);
   ix6144 : nor02_2x port map ( Y=>nx6143, A0=>nx3748, A1=>nx3746);
   ix3749 : nor03_2x port map ( Y=>nx3748, A0=>nx6146, A1=>nx10312, A2=>
      nx11276);
   gen_9_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_9_cmp_mReg_11, QB=>
      nx6146, D=>window_9_11, CLK=>start, R=>rst);
   ix3747 : nor03_2x port map ( Y=>nx3746, A0=>gen_9_cmp_mReg_11, A1=>
      nx10786, A2=>nx11284);
   ix3783 : nand02 port map ( Y=>gen_9_cmp_BSCmp_op2_12, A0=>nx6151, A1=>
      nx6157);
   ix6152 : nor02_2x port map ( Y=>nx6151, A0=>nx3778, A1=>nx3774);
   ix3779 : nor03_2x port map ( Y=>nx3778, A0=>gen_9_cmp_mReg_11, A1=>
      nx10318, A2=>nx11252);
   ix3775 : nor03_2x port map ( Y=>nx3774, A0=>nx6146, A1=>nx11258, A2=>
      nx11268);
   ix6158 : nor02_2x port map ( Y=>nx6157, A0=>nx3770, A1=>nx3768);
   ix3771 : nor03_2x port map ( Y=>nx3770, A0=>nx6161, A1=>nx10314, A2=>
      nx11276);
   gen_9_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_9_cmp_mReg_12, QB=>
      nx6161, D=>window_9_12, CLK=>start, R=>rst);
   ix3769 : nor03_2x port map ( Y=>nx3768, A0=>gen_9_cmp_mReg_12, A1=>
      nx10786, A2=>nx11284);
   ix3805 : nand02 port map ( Y=>gen_9_cmp_BSCmp_op2_13, A0=>nx6167, A1=>
      nx6171);
   ix6168 : nor02_2x port map ( Y=>nx6167, A0=>nx3800, A1=>nx3796);
   ix3801 : nor03_2x port map ( Y=>nx3800, A0=>gen_9_cmp_mReg_12, A1=>
      nx10320, A2=>nx11254);
   ix3797 : nor03_2x port map ( Y=>nx3796, A0=>nx6161, A1=>nx11258, A2=>
      nx11270);
   ix6172 : nor02_2x port map ( Y=>nx6171, A0=>nx3792, A1=>nx3790);
   ix3793 : nor03_2x port map ( Y=>nx3792, A0=>nx6175, A1=>nx10314, A2=>
      nx11278);
   gen_9_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_9_cmp_mReg_13, QB=>
      nx6175, D=>window_9_13, CLK=>start, R=>rst);
   ix3791 : nor03_2x port map ( Y=>nx3790, A0=>gen_9_cmp_mReg_13, A1=>
      nx10786, A2=>nx11286);
   ix3827 : nand02 port map ( Y=>gen_9_cmp_BSCmp_op2_14, A0=>nx6181, A1=>
      nx6186);
   ix6182 : nor02_2x port map ( Y=>nx6181, A0=>nx3822, A1=>nx3818);
   ix3823 : nor03_2x port map ( Y=>nx3822, A0=>gen_9_cmp_mReg_13, A1=>
      nx10320, A2=>nx11254);
   ix3819 : nor03_2x port map ( Y=>nx3818, A0=>nx6175, A1=>nx11260, A2=>
      nx11270);
   ix6187 : nor02_2x port map ( Y=>nx6186, A0=>nx3814, A1=>nx3812);
   ix3815 : nor03_2x port map ( Y=>nx3814, A0=>nx6189, A1=>nx10314, A2=>
      nx11278);
   gen_9_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_9_cmp_mReg_14, QB=>
      nx6189, D=>window_9_14, CLK=>start, R=>rst);
   ix3813 : nor03_2x port map ( Y=>nx3812, A0=>gen_9_cmp_mReg_14, A1=>
      nx10786, A2=>nx11286);
   ix3849 : nand02 port map ( Y=>gen_9_cmp_BSCmp_op2_15, A0=>nx6193, A1=>
      nx6199);
   ix6194 : nor02_2x port map ( Y=>nx6193, A0=>nx3844, A1=>nx3840);
   ix3845 : nor03_2x port map ( Y=>nx3844, A0=>gen_9_cmp_mReg_14, A1=>
      nx10320, A2=>nx11254);
   ix3841 : nor03_2x port map ( Y=>nx3840, A0=>nx6189, A1=>nx11260, A2=>
      nx11270);
   ix6200 : nor02_2x port map ( Y=>nx6199, A0=>nx3836, A1=>nx3834);
   ix3837 : nor03_2x port map ( Y=>nx3836, A0=>nx6203, A1=>nx10314, A2=>
      nx11278);
   gen_9_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_9_cmp_mReg_15, QB=>
      nx6203, D=>window_9_15, CLK=>start, R=>rst);
   ix3835 : nor03_2x port map ( Y=>nx3834, A0=>gen_9_cmp_mReg_15, A1=>
      nx10788, A2=>nx11286);
   ix3859 : nand02 port map ( Y=>gen_9_cmp_BSCmp_op2_16, A0=>nx6209, A1=>
      nx6199);
   ix6210 : nor02_2x port map ( Y=>nx6209, A0=>nx3854, A1=>nx3850);
   ix3855 : nor03_2x port map ( Y=>nx3854, A0=>gen_9_cmp_mReg_15, A1=>
      nx10320, A2=>nx11254);
   ix3851 : nor03_2x port map ( Y=>nx3850, A0=>nx6203, A1=>nx11260, A2=>
      nx11270);
   ix3927 : nand02 port map ( Y=>gen_10_cmp_BSCmp_op2_1, A0=>nx6217, A1=>
      nx6235);
   ix6218 : nor02_2x port map ( Y=>nx6217, A0=>nx3922, A1=>nx3918);
   ix3923 : nor03_2x port map ( Y=>nx3922, A0=>gen_10_cmp_mReg_0, A1=>
      nx10304, A2=>nx11290);
   gen_10_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_10_cmp_mReg_0, QB=>
      nx6221, D=>window_10_0, CLK=>start, R=>rst);
   ix6226 : inv01 port map ( Y=>nx6225, A=>gen_10_cmp_pMux_0);
   ix3919 : nor03_2x port map ( Y=>nx3918, A0=>nx6221, A1=>nx11296, A2=>
      nx11306);
   ix6234 : inv02 port map ( Y=>nx6233, A=>gen_10_cmp_pMux_2);
   ix6236 : nor02_2x port map ( Y=>nx6235, A0=>nx3908, A1=>nx3906);
   ix3909 : nor03_2x port map ( Y=>nx3908, A0=>nx6239, A1=>nx10298, A2=>
      nx11314);
   gen_10_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_10_cmp_mReg_1, QB=>
      nx6239, D=>window_10_1, CLK=>start, R=>rst);
   ix3907 : nor03_2x port map ( Y=>nx3906, A0=>gen_10_cmp_mReg_1, A1=>
      nx10790, A2=>nx11322);
   ix3867 : nor03_2x port map ( Y=>nx3866, A0=>nx10304, A1=>nx6233, A2=>
      gen_10_cmp_pMux_0);
   ix3949 : nand02 port map ( Y=>gen_10_cmp_BSCmp_op2_2, A0=>nx6249, A1=>
      nx6255);
   ix6250 : nor02_2x port map ( Y=>nx6249, A0=>nx3944, A1=>nx3940);
   ix3945 : nor03_2x port map ( Y=>nx3944, A0=>gen_10_cmp_mReg_1, A1=>
      nx10304, A2=>nx11290);
   ix3941 : nor03_2x port map ( Y=>nx3940, A0=>nx6239, A1=>nx11296, A2=>
      nx11306);
   ix6256 : nor02_2x port map ( Y=>nx6255, A0=>nx3936, A1=>nx3934);
   ix3937 : nor03_2x port map ( Y=>nx3936, A0=>nx6259, A1=>nx10298, A2=>
      nx11314);
   gen_10_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_10_cmp_mReg_2, QB=>
      nx6259, D=>window_10_2, CLK=>start, R=>rst);
   ix3935 : nor03_2x port map ( Y=>nx3934, A0=>gen_10_cmp_mReg_2, A1=>
      nx10790, A2=>nx11322);
   ix3971 : nand02 port map ( Y=>gen_10_cmp_BSCmp_op2_3, A0=>nx6265, A1=>
      nx6269);
   ix6266 : nor02_2x port map ( Y=>nx6265, A0=>nx3966, A1=>nx3962);
   ix3967 : nor03_2x port map ( Y=>nx3966, A0=>gen_10_cmp_mReg_2, A1=>
      nx10304, A2=>nx11290);
   ix3963 : nor03_2x port map ( Y=>nx3962, A0=>nx6259, A1=>nx11296, A2=>
      nx11306);
   ix6270 : nor02_2x port map ( Y=>nx6269, A0=>nx3958, A1=>nx3956);
   ix3959 : nor03_2x port map ( Y=>nx3958, A0=>nx6273, A1=>nx10298, A2=>
      nx11314);
   gen_10_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_10_cmp_mReg_3, QB=>
      nx6273, D=>window_10_3, CLK=>start, R=>rst);
   ix3957 : nor03_2x port map ( Y=>nx3956, A0=>gen_10_cmp_mReg_3, A1=>
      nx10790, A2=>nx11322);
   ix3993 : nand02 port map ( Y=>gen_10_cmp_BSCmp_op2_4, A0=>nx6279, A1=>
      nx6283);
   ix6280 : nor02_2x port map ( Y=>nx6279, A0=>nx3988, A1=>nx3984);
   ix3989 : nor03_2x port map ( Y=>nx3988, A0=>gen_10_cmp_mReg_3, A1=>
      nx10304, A2=>nx11290);
   ix3985 : nor03_2x port map ( Y=>nx3984, A0=>nx6273, A1=>nx11296, A2=>
      nx11306);
   ix6284 : nor02_2x port map ( Y=>nx6283, A0=>nx3980, A1=>nx3978);
   ix3981 : nor03_2x port map ( Y=>nx3980, A0=>nx6287, A1=>nx10298, A2=>
      nx11314);
   gen_10_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_10_cmp_mReg_4, QB=>
      nx6287, D=>window_10_4, CLK=>start, R=>rst);
   ix3979 : nor03_2x port map ( Y=>nx3978, A0=>gen_10_cmp_mReg_4, A1=>
      nx10790, A2=>nx11322);
   ix4015 : nand02 port map ( Y=>gen_10_cmp_BSCmp_op2_5, A0=>nx6291, A1=>
      nx6297);
   ix6292 : nor02_2x port map ( Y=>nx6291, A0=>nx4010, A1=>nx4006);
   ix4011 : nor03_2x port map ( Y=>nx4010, A0=>gen_10_cmp_mReg_4, A1=>
      nx10304, A2=>nx11290);
   ix4007 : nor03_2x port map ( Y=>nx4006, A0=>nx6287, A1=>nx11296, A2=>
      nx11306);
   ix6298 : nor02_2x port map ( Y=>nx6297, A0=>nx4002, A1=>nx4000);
   ix4003 : nor03_2x port map ( Y=>nx4002, A0=>nx6301, A1=>nx10300, A2=>
      nx11314);
   gen_10_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_10_cmp_mReg_5, QB=>
      nx6301, D=>window_10_5, CLK=>start, R=>rst);
   ix4001 : nor03_2x port map ( Y=>nx4000, A0=>gen_10_cmp_mReg_5, A1=>
      nx10790, A2=>nx11322);
   ix4037 : nand02 port map ( Y=>gen_10_cmp_BSCmp_op2_6, A0=>nx6305, A1=>
      nx6311);
   ix6306 : nor02_2x port map ( Y=>nx6305, A0=>nx4032, A1=>nx4028);
   ix4033 : nor03_2x port map ( Y=>nx4032, A0=>gen_10_cmp_mReg_5, A1=>
      nx10306, A2=>nx11290);
   ix4029 : nor03_2x port map ( Y=>nx4028, A0=>nx6301, A1=>nx11296, A2=>
      nx11306);
   ix6312 : nor02_2x port map ( Y=>nx6311, A0=>nx4024, A1=>nx4022);
   ix4025 : nor03_2x port map ( Y=>nx4024, A0=>nx6314, A1=>nx10300, A2=>
      nx11314);
   gen_10_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_10_cmp_mReg_6, QB=>
      nx6314, D=>window_10_6, CLK=>start, R=>rst);
   ix4023 : nor03_2x port map ( Y=>nx4022, A0=>gen_10_cmp_mReg_6, A1=>
      nx10790, A2=>nx11322);
   ix4059 : nand02 port map ( Y=>gen_10_cmp_BSCmp_op2_7, A0=>nx6321, A1=>
      nx6327);
   ix6322 : nor02_2x port map ( Y=>nx6321, A0=>nx4054, A1=>nx4050);
   ix4055 : nor03_2x port map ( Y=>nx4054, A0=>gen_10_cmp_mReg_6, A1=>
      nx10306, A2=>nx11292);
   ix4051 : nor03_2x port map ( Y=>nx4050, A0=>nx6314, A1=>nx11298, A2=>
      nx11308);
   ix6328 : nor02_2x port map ( Y=>nx6327, A0=>nx4046, A1=>nx4044);
   ix4047 : nor03_2x port map ( Y=>nx4046, A0=>nx6331, A1=>nx10300, A2=>
      nx11316);
   gen_10_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_10_cmp_mReg_7, QB=>
      nx6331, D=>window_10_7, CLK=>start, R=>rst);
   ix4045 : nor03_2x port map ( Y=>nx4044, A0=>gen_10_cmp_mReg_7, A1=>
      nx10790, A2=>nx11324);
   ix4081 : nand02 port map ( Y=>gen_10_cmp_BSCmp_op2_8, A0=>nx6335, A1=>
      nx6341);
   ix6336 : nor02_2x port map ( Y=>nx6335, A0=>nx4076, A1=>nx4072);
   ix4077 : nor03_2x port map ( Y=>nx4076, A0=>gen_10_cmp_mReg_7, A1=>
      nx10306, A2=>nx11292);
   ix4073 : nor03_2x port map ( Y=>nx4072, A0=>nx6331, A1=>nx11298, A2=>
      nx11308);
   ix6342 : nor02_2x port map ( Y=>nx6341, A0=>nx4068, A1=>nx4066);
   ix4069 : nor03_2x port map ( Y=>nx4068, A0=>nx6345, A1=>nx10300, A2=>
      nx11316);
   gen_10_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_10_cmp_mReg_8, QB=>
      nx6345, D=>window_10_8, CLK=>start, R=>rst);
   ix4067 : nor03_2x port map ( Y=>nx4066, A0=>gen_10_cmp_mReg_8, A1=>
      nx10792, A2=>nx11324);
   ix4103 : nand02 port map ( Y=>gen_10_cmp_BSCmp_op2_9, A0=>nx6349, A1=>
      nx6355);
   ix6350 : nor02_2x port map ( Y=>nx6349, A0=>nx4098, A1=>nx4094);
   ix4099 : nor03_2x port map ( Y=>nx4098, A0=>gen_10_cmp_mReg_8, A1=>
      nx10306, A2=>nx11292);
   ix4095 : nor03_2x port map ( Y=>nx4094, A0=>nx6345, A1=>nx11298, A2=>
      nx11308);
   ix6356 : nor02_2x port map ( Y=>nx6355, A0=>nx4090, A1=>nx4088);
   ix4091 : nor03_2x port map ( Y=>nx4090, A0=>nx6358, A1=>nx10300, A2=>
      nx11316);
   gen_10_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_10_cmp_mReg_9, QB=>
      nx6358, D=>window_10_9, CLK=>start, R=>rst);
   ix4089 : nor03_2x port map ( Y=>nx4088, A0=>gen_10_cmp_mReg_9, A1=>
      nx10792, A2=>nx11324);
   ix4125 : nand02 port map ( Y=>gen_10_cmp_BSCmp_op2_10, A0=>nx6365, A1=>
      nx6371);
   ix6366 : nor02_2x port map ( Y=>nx6365, A0=>nx4120, A1=>nx4116);
   ix4121 : nor03_2x port map ( Y=>nx4120, A0=>gen_10_cmp_mReg_9, A1=>
      nx10306, A2=>nx11292);
   ix4117 : nor03_2x port map ( Y=>nx4116, A0=>nx6358, A1=>nx11298, A2=>
      nx11308);
   ix6372 : nor02_2x port map ( Y=>nx6371, A0=>nx4112, A1=>nx4110);
   ix4113 : nor03_2x port map ( Y=>nx4112, A0=>nx6375, A1=>nx10300, A2=>
      nx11316);
   gen_10_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_10_cmp_mReg_10, QB=>
      nx6375, D=>window_10_10, CLK=>start, R=>rst);
   ix4111 : nor03_2x port map ( Y=>nx4110, A0=>gen_10_cmp_mReg_10, A1=>
      nx10792, A2=>nx11324);
   ix4147 : nand02 port map ( Y=>gen_10_cmp_BSCmp_op2_11, A0=>nx6379, A1=>
      nx6385);
   ix6380 : nor02_2x port map ( Y=>nx6379, A0=>nx4142, A1=>nx4138);
   ix4143 : nor03_2x port map ( Y=>nx4142, A0=>gen_10_cmp_mReg_10, A1=>
      nx10306, A2=>nx11292);
   ix4139 : nor03_2x port map ( Y=>nx4138, A0=>nx6375, A1=>nx11298, A2=>
      nx11308);
   ix6386 : nor02_2x port map ( Y=>nx6385, A0=>nx4134, A1=>nx4132);
   ix4135 : nor03_2x port map ( Y=>nx4134, A0=>nx6389, A1=>nx10300, A2=>
      nx11316);
   gen_10_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_10_cmp_mReg_11, QB=>
      nx6389, D=>window_10_11, CLK=>start, R=>rst);
   ix4133 : nor03_2x port map ( Y=>nx4132, A0=>gen_10_cmp_mReg_11, A1=>
      nx10792, A2=>nx11324);
   ix4169 : nand02 port map ( Y=>gen_10_cmp_BSCmp_op2_12, A0=>nx6393, A1=>
      nx6399);
   ix6394 : nor02_2x port map ( Y=>nx6393, A0=>nx4164, A1=>nx4160);
   ix4165 : nor03_2x port map ( Y=>nx4164, A0=>gen_10_cmp_mReg_11, A1=>
      nx10306, A2=>nx11292);
   ix4161 : nor03_2x port map ( Y=>nx4160, A0=>nx6389, A1=>nx11298, A2=>
      nx11308);
   ix6400 : nor02_2x port map ( Y=>nx6399, A0=>nx4156, A1=>nx4154);
   ix4157 : nor03_2x port map ( Y=>nx4156, A0=>nx6402, A1=>nx10302, A2=>
      nx11316);
   gen_10_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_10_cmp_mReg_12, QB=>
      nx6402, D=>window_10_12, CLK=>start, R=>rst);
   ix4155 : nor03_2x port map ( Y=>nx4154, A0=>gen_10_cmp_mReg_12, A1=>
      nx10792, A2=>nx11324);
   ix4191 : nand02 port map ( Y=>gen_10_cmp_BSCmp_op2_13, A0=>nx6409, A1=>
      nx6415);
   ix6410 : nor02_2x port map ( Y=>nx6409, A0=>nx4186, A1=>nx4182);
   ix4187 : nor03_2x port map ( Y=>nx4186, A0=>gen_10_cmp_mReg_12, A1=>
      nx10308, A2=>nx11294);
   ix4183 : nor03_2x port map ( Y=>nx4182, A0=>nx6402, A1=>nx11298, A2=>
      nx11310);
   ix6416 : nor02_2x port map ( Y=>nx6415, A0=>nx4178, A1=>nx4176);
   ix4179 : nor03_2x port map ( Y=>nx4178, A0=>nx6419, A1=>nx10302, A2=>
      nx11318);
   gen_10_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_10_cmp_mReg_13, QB=>
      nx6419, D=>window_10_13, CLK=>start, R=>rst);
   ix4177 : nor03_2x port map ( Y=>nx4176, A0=>gen_10_cmp_mReg_13, A1=>
      nx10792, A2=>nx11326);
   ix4213 : nand02 port map ( Y=>gen_10_cmp_BSCmp_op2_14, A0=>nx6423, A1=>
      nx6429);
   ix6424 : nor02_2x port map ( Y=>nx6423, A0=>nx4208, A1=>nx4204);
   ix4209 : nor03_2x port map ( Y=>nx4208, A0=>gen_10_cmp_mReg_13, A1=>
      nx10308, A2=>nx11294);
   ix4205 : nor03_2x port map ( Y=>nx4204, A0=>nx6419, A1=>nx11300, A2=>
      nx11310);
   ix6430 : nor02_2x port map ( Y=>nx6429, A0=>nx4200, A1=>nx4198);
   ix4201 : nor03_2x port map ( Y=>nx4200, A0=>nx6433, A1=>nx10302, A2=>
      nx11318);
   gen_10_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_10_cmp_mReg_14, QB=>
      nx6433, D=>window_10_14, CLK=>start, R=>rst);
   ix4199 : nor03_2x port map ( Y=>nx4198, A0=>gen_10_cmp_mReg_14, A1=>
      nx10792, A2=>nx11326);
   ix4235 : nand02 port map ( Y=>gen_10_cmp_BSCmp_op2_15, A0=>nx6437, A1=>
      nx6443);
   ix6438 : nor02_2x port map ( Y=>nx6437, A0=>nx4230, A1=>nx4226);
   ix4231 : nor03_2x port map ( Y=>nx4230, A0=>gen_10_cmp_mReg_14, A1=>
      nx10308, A2=>nx11294);
   ix4227 : nor03_2x port map ( Y=>nx4226, A0=>nx6433, A1=>nx11300, A2=>
      nx11310);
   ix6444 : nor02_2x port map ( Y=>nx6443, A0=>nx4222, A1=>nx4220);
   ix4223 : nor03_2x port map ( Y=>nx4222, A0=>nx6446, A1=>nx10302, A2=>
      nx11318);
   gen_10_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_10_cmp_mReg_15, QB=>
      nx6446, D=>window_10_15, CLK=>start, R=>rst);
   ix4221 : nor03_2x port map ( Y=>nx4220, A0=>gen_10_cmp_mReg_15, A1=>
      nx10794, A2=>nx11326);
   ix4245 : nand02 port map ( Y=>gen_10_cmp_BSCmp_op2_16, A0=>nx6453, A1=>
      nx6443);
   ix6454 : nor02_2x port map ( Y=>nx6453, A0=>nx4240, A1=>nx4236);
   ix4241 : nor03_2x port map ( Y=>nx4240, A0=>gen_10_cmp_mReg_15, A1=>
      nx10308, A2=>nx11294);
   ix4237 : nor03_2x port map ( Y=>nx4236, A0=>nx6446, A1=>nx11300, A2=>
      nx11310);
   ix4313 : nand02 port map ( Y=>gen_11_cmp_BSCmp_op2_1, A0=>nx6459, A1=>
      nx6479);
   ix6460 : nor02_2x port map ( Y=>nx6459, A0=>nx4308, A1=>nx4304);
   ix4309 : nor03_2x port map ( Y=>nx4308, A0=>gen_11_cmp_mReg_0, A1=>
      nx10292, A2=>nx11330);
   gen_11_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_11_cmp_mReg_0, QB=>
      nx6465, D=>window_11_0, CLK=>start, R=>rst);
   ix6470 : inv01 port map ( Y=>nx6468, A=>gen_11_cmp_pMux_0);
   ix4305 : nor03_2x port map ( Y=>nx4304, A0=>nx6465, A1=>nx11336, A2=>
      nx11346);
   ix6478 : inv02 port map ( Y=>nx6477, A=>gen_11_cmp_pMux_2);
   ix6480 : nor02_2x port map ( Y=>nx6479, A0=>nx4294, A1=>nx4292);
   ix4295 : nor03_2x port map ( Y=>nx4294, A0=>nx6483, A1=>nx10286, A2=>
      nx11354);
   gen_11_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_11_cmp_mReg_1, QB=>
      nx6483, D=>window_11_1, CLK=>start, R=>rst);
   ix4293 : nor03_2x port map ( Y=>nx4292, A0=>gen_11_cmp_mReg_1, A1=>
      nx10796, A2=>nx11362);
   ix4253 : nor03_2x port map ( Y=>nx4252, A0=>nx10292, A1=>nx6477, A2=>
      gen_11_cmp_pMux_0);
   ix4335 : nand02 port map ( Y=>gen_11_cmp_BSCmp_op2_2, A0=>nx6493, A1=>
      nx6499);
   ix6494 : nor02_2x port map ( Y=>nx6493, A0=>nx4330, A1=>nx4326);
   ix4331 : nor03_2x port map ( Y=>nx4330, A0=>gen_11_cmp_mReg_1, A1=>
      nx10292, A2=>nx11330);
   ix4327 : nor03_2x port map ( Y=>nx4326, A0=>nx6483, A1=>nx11336, A2=>
      nx11346);
   ix6500 : nor02_2x port map ( Y=>nx6499, A0=>nx4322, A1=>nx4320);
   ix4323 : nor03_2x port map ( Y=>nx4322, A0=>nx6503, A1=>nx10286, A2=>
      nx11354);
   gen_11_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_11_cmp_mReg_2, QB=>
      nx6503, D=>window_11_2, CLK=>start, R=>rst);
   ix4321 : nor03_2x port map ( Y=>nx4320, A0=>gen_11_cmp_mReg_2, A1=>
      nx10796, A2=>nx11362);
   ix4357 : nand02 port map ( Y=>gen_11_cmp_BSCmp_op2_3, A0=>nx6509, A1=>
      nx6513);
   ix6510 : nor02_2x port map ( Y=>nx6509, A0=>nx4352, A1=>nx4348);
   ix4353 : nor03_2x port map ( Y=>nx4352, A0=>gen_11_cmp_mReg_2, A1=>
      nx10292, A2=>nx11330);
   ix4349 : nor03_2x port map ( Y=>nx4348, A0=>nx6503, A1=>nx11336, A2=>
      nx11346);
   ix6514 : nor02_2x port map ( Y=>nx6513, A0=>nx4344, A1=>nx4342);
   ix4345 : nor03_2x port map ( Y=>nx4344, A0=>nx6517, A1=>nx10286, A2=>
      nx11354);
   gen_11_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_11_cmp_mReg_3, QB=>
      nx6517, D=>window_11_3, CLK=>start, R=>rst);
   ix4343 : nor03_2x port map ( Y=>nx4342, A0=>gen_11_cmp_mReg_3, A1=>
      nx10796, A2=>nx11362);
   ix4379 : nand02 port map ( Y=>gen_11_cmp_BSCmp_op2_4, A0=>nx6523, A1=>
      nx6529);
   ix6524 : nor02_2x port map ( Y=>nx6523, A0=>nx4374, A1=>nx4370);
   ix4375 : nor03_2x port map ( Y=>nx4374, A0=>gen_11_cmp_mReg_3, A1=>
      nx10292, A2=>nx11330);
   ix4371 : nor03_2x port map ( Y=>nx4370, A0=>nx6517, A1=>nx11336, A2=>
      nx11346);
   ix6530 : nor02_2x port map ( Y=>nx6529, A0=>nx4366, A1=>nx4364);
   ix4367 : nor03_2x port map ( Y=>nx4366, A0=>nx6532, A1=>nx10286, A2=>
      nx11354);
   gen_11_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_11_cmp_mReg_4, QB=>
      nx6532, D=>window_11_4, CLK=>start, R=>rst);
   ix4365 : nor03_2x port map ( Y=>nx4364, A0=>gen_11_cmp_mReg_4, A1=>
      nx10796, A2=>nx11362);
   ix4401 : nand02 port map ( Y=>gen_11_cmp_BSCmp_op2_5, A0=>nx6537, A1=>
      nx6543);
   ix6538 : nor02_2x port map ( Y=>nx6537, A0=>nx4396, A1=>nx4392);
   ix4397 : nor03_2x port map ( Y=>nx4396, A0=>gen_11_cmp_mReg_4, A1=>
      nx10292, A2=>nx11330);
   ix4393 : nor03_2x port map ( Y=>nx4392, A0=>nx6532, A1=>nx11336, A2=>
      nx11346);
   ix6544 : nor02_2x port map ( Y=>nx6543, A0=>nx4388, A1=>nx4386);
   ix4389 : nor03_2x port map ( Y=>nx4388, A0=>nx6547, A1=>nx10288, A2=>
      nx11354);
   gen_11_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_11_cmp_mReg_5, QB=>
      nx6547, D=>window_11_5, CLK=>start, R=>rst);
   ix4387 : nor03_2x port map ( Y=>nx4386, A0=>gen_11_cmp_mReg_5, A1=>
      nx10796, A2=>nx11362);
   ix4423 : nand02 port map ( Y=>gen_11_cmp_BSCmp_op2_6, A0=>nx6553, A1=>
      nx6557);
   ix6554 : nor02_2x port map ( Y=>nx6553, A0=>nx4418, A1=>nx4414);
   ix4419 : nor03_2x port map ( Y=>nx4418, A0=>gen_11_cmp_mReg_5, A1=>
      nx10294, A2=>nx11330);
   ix4415 : nor03_2x port map ( Y=>nx4414, A0=>nx6547, A1=>nx11336, A2=>
      nx11346);
   ix6558 : nor02_2x port map ( Y=>nx6557, A0=>nx4410, A1=>nx4408);
   ix4411 : nor03_2x port map ( Y=>nx4410, A0=>nx6561, A1=>nx10288, A2=>
      nx11354);
   gen_11_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_11_cmp_mReg_6, QB=>
      nx6561, D=>window_11_6, CLK=>start, R=>rst);
   ix4409 : nor03_2x port map ( Y=>nx4408, A0=>gen_11_cmp_mReg_6, A1=>
      nx10796, A2=>nx11362);
   ix4445 : nand02 port map ( Y=>gen_11_cmp_BSCmp_op2_7, A0=>nx6567, A1=>
      nx6572);
   ix6568 : nor02_2x port map ( Y=>nx6567, A0=>nx4440, A1=>nx4436);
   ix4441 : nor03_2x port map ( Y=>nx4440, A0=>gen_11_cmp_mReg_6, A1=>
      nx10294, A2=>nx11332);
   ix4437 : nor03_2x port map ( Y=>nx4436, A0=>nx6561, A1=>nx11338, A2=>
      nx11348);
   ix6573 : nor02_2x port map ( Y=>nx6572, A0=>nx4432, A1=>nx4430);
   ix4433 : nor03_2x port map ( Y=>nx4432, A0=>nx6575, A1=>nx10288, A2=>
      nx11356);
   gen_11_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_11_cmp_mReg_7, QB=>
      nx6575, D=>window_11_7, CLK=>start, R=>rst);
   ix4431 : nor03_2x port map ( Y=>nx4430, A0=>gen_11_cmp_mReg_7, A1=>
      nx10796, A2=>nx11364);
   ix4467 : nand02 port map ( Y=>gen_11_cmp_BSCmp_op2_8, A0=>nx6579, A1=>
      nx6585);
   ix6580 : nor02_2x port map ( Y=>nx6579, A0=>nx4462, A1=>nx4458);
   ix4463 : nor03_2x port map ( Y=>nx4462, A0=>gen_11_cmp_mReg_7, A1=>
      nx10294, A2=>nx11332);
   ix4459 : nor03_2x port map ( Y=>nx4458, A0=>nx6575, A1=>nx11338, A2=>
      nx11348);
   ix6586 : nor02_2x port map ( Y=>nx6585, A0=>nx4454, A1=>nx4452);
   ix4455 : nor03_2x port map ( Y=>nx4454, A0=>nx6589, A1=>nx10288, A2=>
      nx11356);
   gen_11_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_11_cmp_mReg_8, QB=>
      nx6589, D=>window_11_8, CLK=>start, R=>rst);
   ix4453 : nor03_2x port map ( Y=>nx4452, A0=>gen_11_cmp_mReg_8, A1=>
      nx10798, A2=>nx11364);
   ix4489 : nand02 port map ( Y=>gen_11_cmp_BSCmp_op2_9, A0=>nx6595, A1=>
      nx6601);
   ix6596 : nor02_2x port map ( Y=>nx6595, A0=>nx4484, A1=>nx4480);
   ix4485 : nor03_2x port map ( Y=>nx4484, A0=>gen_11_cmp_mReg_8, A1=>
      nx10294, A2=>nx11332);
   ix4481 : nor03_2x port map ( Y=>nx4480, A0=>nx6589, A1=>nx11338, A2=>
      nx11348);
   ix6602 : nor02_2x port map ( Y=>nx6601, A0=>nx4476, A1=>nx4474);
   ix4477 : nor03_2x port map ( Y=>nx4476, A0=>nx6604, A1=>nx10288, A2=>
      nx11356);
   gen_11_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_11_cmp_mReg_9, QB=>
      nx6604, D=>window_11_9, CLK=>start, R=>rst);
   ix4475 : nor03_2x port map ( Y=>nx4474, A0=>gen_11_cmp_mReg_9, A1=>
      nx10798, A2=>nx11364);
   ix4511 : nand02 port map ( Y=>gen_11_cmp_BSCmp_op2_10, A0=>nx6609, A1=>
      nx6615);
   ix6610 : nor02_2x port map ( Y=>nx6609, A0=>nx4506, A1=>nx4502);
   ix4507 : nor03_2x port map ( Y=>nx4506, A0=>gen_11_cmp_mReg_9, A1=>
      nx10294, A2=>nx11332);
   ix4503 : nor03_2x port map ( Y=>nx4502, A0=>nx6604, A1=>nx11338, A2=>
      nx11348);
   ix6616 : nor02_2x port map ( Y=>nx6615, A0=>nx4498, A1=>nx4496);
   ix4499 : nor03_2x port map ( Y=>nx4498, A0=>nx6619, A1=>nx10288, A2=>
      nx11356);
   gen_11_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_11_cmp_mReg_10, QB=>
      nx6619, D=>window_11_10, CLK=>start, R=>rst);
   ix4497 : nor03_2x port map ( Y=>nx4496, A0=>gen_11_cmp_mReg_10, A1=>
      nx10798, A2=>nx11364);
   ix4533 : nand02 port map ( Y=>gen_11_cmp_BSCmp_op2_11, A0=>nx6625, A1=>
      nx6631);
   ix6626 : nor02_2x port map ( Y=>nx6625, A0=>nx4528, A1=>nx4524);
   ix4529 : nor03_2x port map ( Y=>nx4528, A0=>gen_11_cmp_mReg_10, A1=>
      nx10294, A2=>nx11332);
   ix4525 : nor03_2x port map ( Y=>nx4524, A0=>nx6619, A1=>nx11338, A2=>
      nx11348);
   ix6632 : nor02_2x port map ( Y=>nx6631, A0=>nx4520, A1=>nx4518);
   ix4521 : nor03_2x port map ( Y=>nx4520, A0=>nx6634, A1=>nx10288, A2=>
      nx11356);
   gen_11_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_11_cmp_mReg_11, QB=>
      nx6634, D=>window_11_11, CLK=>start, R=>rst);
   ix4519 : nor03_2x port map ( Y=>nx4518, A0=>gen_11_cmp_mReg_11, A1=>
      nx10798, A2=>nx11364);
   ix4555 : nand02 port map ( Y=>gen_11_cmp_BSCmp_op2_12, A0=>nx6641, A1=>
      nx6647);
   ix6642 : nor02_2x port map ( Y=>nx6641, A0=>nx4550, A1=>nx4546);
   ix4551 : nor03_2x port map ( Y=>nx4550, A0=>gen_11_cmp_mReg_11, A1=>
      nx10294, A2=>nx11332);
   ix4547 : nor03_2x port map ( Y=>nx4546, A0=>nx6634, A1=>nx11338, A2=>
      nx11348);
   ix6648 : nor02_2x port map ( Y=>nx6647, A0=>nx4542, A1=>nx4540);
   ix4543 : nor03_2x port map ( Y=>nx4542, A0=>nx6651, A1=>nx10290, A2=>
      nx11356);
   gen_11_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_11_cmp_mReg_12, QB=>
      nx6651, D=>window_11_12, CLK=>start, R=>rst);
   ix4541 : nor03_2x port map ( Y=>nx4540, A0=>gen_11_cmp_mReg_12, A1=>
      nx10798, A2=>nx11364);
   ix4577 : nand02 port map ( Y=>gen_11_cmp_BSCmp_op2_13, A0=>nx6655, A1=>
      nx6661);
   ix6656 : nor02_2x port map ( Y=>nx6655, A0=>nx4572, A1=>nx4568);
   ix4573 : nor03_2x port map ( Y=>nx4572, A0=>gen_11_cmp_mReg_12, A1=>
      nx10296, A2=>nx11334);
   ix4569 : nor03_2x port map ( Y=>nx4568, A0=>nx6651, A1=>nx11338, A2=>
      nx11350);
   ix6662 : nor02_2x port map ( Y=>nx6661, A0=>nx4564, A1=>nx4562);
   ix4565 : nor03_2x port map ( Y=>nx4564, A0=>nx6665, A1=>nx10290, A2=>
      nx11358);
   gen_11_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_11_cmp_mReg_13, QB=>
      nx6665, D=>window_11_13, CLK=>start, R=>rst);
   ix4563 : nor03_2x port map ( Y=>nx4562, A0=>gen_11_cmp_mReg_13, A1=>
      nx10798, A2=>nx11366);
   ix4599 : nand02 port map ( Y=>gen_11_cmp_BSCmp_op2_14, A0=>nx6669, A1=>
      nx6675);
   ix6670 : nor02_2x port map ( Y=>nx6669, A0=>nx4594, A1=>nx4590);
   ix4595 : nor03_2x port map ( Y=>nx4594, A0=>gen_11_cmp_mReg_13, A1=>
      nx10296, A2=>nx11334);
   ix4591 : nor03_2x port map ( Y=>nx4590, A0=>nx6665, A1=>nx11340, A2=>
      nx11350);
   ix6676 : nor02_2x port map ( Y=>nx6675, A0=>nx4586, A1=>nx4584);
   ix4587 : nor03_2x port map ( Y=>nx4586, A0=>nx6678, A1=>nx10290, A2=>
      nx11358);
   gen_11_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_11_cmp_mReg_14, QB=>
      nx6678, D=>window_11_14, CLK=>start, R=>rst);
   ix4585 : nor03_2x port map ( Y=>nx4584, A0=>gen_11_cmp_mReg_14, A1=>
      nx10798, A2=>nx11366);
   ix4621 : nand02 port map ( Y=>gen_11_cmp_BSCmp_op2_15, A0=>nx6685, A1=>
      nx6691);
   ix6686 : nor02_2x port map ( Y=>nx6685, A0=>nx4616, A1=>nx4612);
   ix4617 : nor03_2x port map ( Y=>nx4616, A0=>gen_11_cmp_mReg_14, A1=>
      nx10296, A2=>nx11334);
   ix4613 : nor03_2x port map ( Y=>nx4612, A0=>nx6678, A1=>nx11340, A2=>
      nx11350);
   ix6692 : nor02_2x port map ( Y=>nx6691, A0=>nx4608, A1=>nx4606);
   ix4609 : nor03_2x port map ( Y=>nx4608, A0=>nx6695, A1=>nx10290, A2=>
      nx11358);
   gen_11_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_11_cmp_mReg_15, QB=>
      nx6695, D=>window_11_15, CLK=>start, R=>rst);
   ix4607 : nor03_2x port map ( Y=>nx4606, A0=>gen_11_cmp_mReg_15, A1=>
      nx10800, A2=>nx11366);
   ix4631 : nand02 port map ( Y=>gen_11_cmp_BSCmp_op2_16, A0=>nx6699, A1=>
      nx6691);
   ix6700 : nor02_2x port map ( Y=>nx6699, A0=>nx4626, A1=>nx4622);
   ix4627 : nor03_2x port map ( Y=>nx4626, A0=>gen_11_cmp_mReg_15, A1=>
      nx10296, A2=>nx11334);
   ix4623 : nor03_2x port map ( Y=>nx4622, A0=>nx6695, A1=>nx11340, A2=>
      nx11350);
   ix4699 : nand02 port map ( Y=>gen_12_cmp_BSCmp_op2_1, A0=>nx6707, A1=>
      nx6727);
   ix6708 : nor02_2x port map ( Y=>nx6707, A0=>nx4694, A1=>nx4690);
   ix4695 : nor03_2x port map ( Y=>nx4694, A0=>gen_12_cmp_mReg_0, A1=>
      nx10280, A2=>nx11370);
   gen_12_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_12_cmp_mReg_0, QB=>
      nx6713, D=>window_12_0, CLK=>start, R=>rst);
   ix6718 : inv01 port map ( Y=>nx6717, A=>gen_12_cmp_pMux_0);
   ix4691 : nor03_2x port map ( Y=>nx4690, A0=>nx6713, A1=>nx11376, A2=>
      nx11386);
   ix6726 : inv02 port map ( Y=>nx6725, A=>gen_12_cmp_pMux_2);
   ix6728 : nor02_2x port map ( Y=>nx6727, A0=>nx4680, A1=>nx4678);
   ix4681 : nor03_2x port map ( Y=>nx4680, A0=>nx6731, A1=>nx10274, A2=>
      nx11394);
   gen_12_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_12_cmp_mReg_1, QB=>
      nx6731, D=>window_12_1, CLK=>start, R=>rst);
   ix4679 : nor03_2x port map ( Y=>nx4678, A0=>gen_12_cmp_mReg_1, A1=>
      nx10802, A2=>nx11402);
   ix4639 : nor03_2x port map ( Y=>nx4638, A0=>nx10280, A1=>nx6725, A2=>
      gen_12_cmp_pMux_0);
   ix4721 : nand02 port map ( Y=>gen_12_cmp_BSCmp_op2_2, A0=>nx6742, A1=>
      nx6747);
   ix6743 : nor02_2x port map ( Y=>nx6742, A0=>nx4716, A1=>nx4712);
   ix4717 : nor03_2x port map ( Y=>nx4716, A0=>gen_12_cmp_mReg_1, A1=>
      nx10280, A2=>nx11370);
   ix4713 : nor03_2x port map ( Y=>nx4712, A0=>nx6731, A1=>nx11376, A2=>
      nx11386);
   ix6748 : nor02_2x port map ( Y=>nx6747, A0=>nx4708, A1=>nx4706);
   ix4709 : nor03_2x port map ( Y=>nx4708, A0=>nx6751, A1=>nx10274, A2=>
      nx11394);
   gen_12_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_12_cmp_mReg_2, QB=>
      nx6751, D=>window_12_2, CLK=>start, R=>rst);
   ix4707 : nor03_2x port map ( Y=>nx4706, A0=>gen_12_cmp_mReg_2, A1=>
      nx10802, A2=>nx11402);
   ix4743 : nand02 port map ( Y=>gen_12_cmp_BSCmp_op2_3, A0=>nx6757, A1=>
      nx6763);
   ix6758 : nor02_2x port map ( Y=>nx6757, A0=>nx4738, A1=>nx4734);
   ix4739 : nor03_2x port map ( Y=>nx4738, A0=>gen_12_cmp_mReg_2, A1=>
      nx10280, A2=>nx11370);
   ix4735 : nor03_2x port map ( Y=>nx4734, A0=>nx6751, A1=>nx11376, A2=>
      nx11386);
   ix6764 : nor02_2x port map ( Y=>nx6763, A0=>nx4730, A1=>nx4728);
   ix4731 : nor03_2x port map ( Y=>nx4730, A0=>nx6766, A1=>nx10274, A2=>
      nx11394);
   gen_12_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_12_cmp_mReg_3, QB=>
      nx6766, D=>window_12_3, CLK=>start, R=>rst);
   ix4729 : nor03_2x port map ( Y=>nx4728, A0=>gen_12_cmp_mReg_3, A1=>
      nx10802, A2=>nx11402);
   ix4765 : nand02 port map ( Y=>gen_12_cmp_BSCmp_op2_4, A0=>nx6773, A1=>
      nx6779);
   ix6774 : nor02_2x port map ( Y=>nx6773, A0=>nx4760, A1=>nx4756);
   ix4761 : nor03_2x port map ( Y=>nx4760, A0=>gen_12_cmp_mReg_3, A1=>
      nx10280, A2=>nx11370);
   ix4757 : nor03_2x port map ( Y=>nx4756, A0=>nx6766, A1=>nx11376, A2=>
      nx11386);
   ix6780 : nor02_2x port map ( Y=>nx6779, A0=>nx4752, A1=>nx4750);
   ix4753 : nor03_2x port map ( Y=>nx4752, A0=>nx6783, A1=>nx10274, A2=>
      nx11394);
   gen_12_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_12_cmp_mReg_4, QB=>
      nx6783, D=>window_12_4, CLK=>start, R=>rst);
   ix4751 : nor03_2x port map ( Y=>nx4750, A0=>gen_12_cmp_mReg_4, A1=>
      nx10802, A2=>nx11402);
   ix4787 : nand02 port map ( Y=>gen_12_cmp_BSCmp_op2_5, A0=>nx6787, A1=>
      nx6793);
   ix6788 : nor02_2x port map ( Y=>nx6787, A0=>nx4782, A1=>nx4778);
   ix4783 : nor03_2x port map ( Y=>nx4782, A0=>gen_12_cmp_mReg_4, A1=>
      nx10280, A2=>nx11370);
   ix4779 : nor03_2x port map ( Y=>nx4778, A0=>nx6783, A1=>nx11376, A2=>
      nx11386);
   ix6794 : nor02_2x port map ( Y=>nx6793, A0=>nx4774, A1=>nx4772);
   ix4775 : nor03_2x port map ( Y=>nx4774, A0=>nx6797, A1=>nx10276, A2=>
      nx11394);
   gen_12_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_12_cmp_mReg_5, QB=>
      nx6797, D=>window_12_5, CLK=>start, R=>rst);
   ix4773 : nor03_2x port map ( Y=>nx4772, A0=>gen_12_cmp_mReg_5, A1=>
      nx10802, A2=>nx11402);
   ix4809 : nand02 port map ( Y=>gen_12_cmp_BSCmp_op2_6, A0=>nx6801, A1=>
      nx6807);
   ix6802 : nor02_2x port map ( Y=>nx6801, A0=>nx4804, A1=>nx4800);
   ix4805 : nor03_2x port map ( Y=>nx4804, A0=>gen_12_cmp_mReg_5, A1=>
      nx10282, A2=>nx11370);
   ix4801 : nor03_2x port map ( Y=>nx4800, A0=>nx6797, A1=>nx11376, A2=>
      nx11386);
   ix6808 : nor02_2x port map ( Y=>nx6807, A0=>nx4796, A1=>nx4794);
   ix4797 : nor03_2x port map ( Y=>nx4796, A0=>nx6810, A1=>nx10276, A2=>
      nx11394);
   gen_12_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_12_cmp_mReg_6, QB=>
      nx6810, D=>window_12_6, CLK=>start, R=>rst);
   ix4795 : nor03_2x port map ( Y=>nx4794, A0=>gen_12_cmp_mReg_6, A1=>
      nx10802, A2=>nx11402);
   ix4831 : nand02 port map ( Y=>gen_12_cmp_BSCmp_op2_7, A0=>nx6817, A1=>
      nx6823);
   ix6818 : nor02_2x port map ( Y=>nx6817, A0=>nx4826, A1=>nx4822);
   ix4827 : nor03_2x port map ( Y=>nx4826, A0=>gen_12_cmp_mReg_6, A1=>
      nx10282, A2=>nx11372);
   ix4823 : nor03_2x port map ( Y=>nx4822, A0=>nx6810, A1=>nx11378, A2=>
      nx11388);
   ix6824 : nor02_2x port map ( Y=>nx6823, A0=>nx4818, A1=>nx4816);
   ix4819 : nor03_2x port map ( Y=>nx4818, A0=>nx6827, A1=>nx10276, A2=>
      nx11396);
   gen_12_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_12_cmp_mReg_7, QB=>
      nx6827, D=>window_12_7, CLK=>start, R=>rst);
   ix4817 : nor03_2x port map ( Y=>nx4816, A0=>gen_12_cmp_mReg_7, A1=>
      nx10802, A2=>nx11404);
   ix4853 : nand02 port map ( Y=>gen_12_cmp_BSCmp_op2_8, A0=>nx6831, A1=>
      nx6837);
   ix6832 : nor02_2x port map ( Y=>nx6831, A0=>nx4848, A1=>nx4844);
   ix4849 : nor03_2x port map ( Y=>nx4848, A0=>gen_12_cmp_mReg_7, A1=>
      nx10282, A2=>nx11372);
   ix4845 : nor03_2x port map ( Y=>nx4844, A0=>nx6827, A1=>nx11378, A2=>
      nx11388);
   ix6838 : nor02_2x port map ( Y=>nx6837, A0=>nx4840, A1=>nx4838);
   ix4841 : nor03_2x port map ( Y=>nx4840, A0=>nx6841, A1=>nx10276, A2=>
      nx11396);
   gen_12_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_12_cmp_mReg_8, QB=>
      nx6841, D=>window_12_8, CLK=>start, R=>rst);
   ix4839 : nor03_2x port map ( Y=>nx4838, A0=>gen_12_cmp_mReg_8, A1=>
      nx10804, A2=>nx11404);
   ix4875 : nand02 port map ( Y=>gen_12_cmp_BSCmp_op2_9, A0=>nx6845, A1=>
      nx6851);
   ix6846 : nor02_2x port map ( Y=>nx6845, A0=>nx4870, A1=>nx4866);
   ix4871 : nor03_2x port map ( Y=>nx4870, A0=>gen_12_cmp_mReg_8, A1=>
      nx10282, A2=>nx11372);
   ix4867 : nor03_2x port map ( Y=>nx4866, A0=>nx6841, A1=>nx11378, A2=>
      nx11388);
   ix6852 : nor02_2x port map ( Y=>nx6851, A0=>nx4862, A1=>nx4860);
   ix4863 : nor03_2x port map ( Y=>nx4862, A0=>nx6854, A1=>nx10276, A2=>
      nx11396);
   gen_12_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_12_cmp_mReg_9, QB=>
      nx6854, D=>window_12_9, CLK=>start, R=>rst);
   ix4861 : nor03_2x port map ( Y=>nx4860, A0=>gen_12_cmp_mReg_9, A1=>
      nx10804, A2=>nx11404);
   ix4897 : nand02 port map ( Y=>gen_12_cmp_BSCmp_op2_10, A0=>nx6861, A1=>
      nx6867);
   ix6862 : nor02_2x port map ( Y=>nx6861, A0=>nx4892, A1=>nx4888);
   ix4893 : nor03_2x port map ( Y=>nx4892, A0=>gen_12_cmp_mReg_9, A1=>
      nx10282, A2=>nx11372);
   ix4889 : nor03_2x port map ( Y=>nx4888, A0=>nx6854, A1=>nx11378, A2=>
      nx11388);
   ix6868 : nor02_2x port map ( Y=>nx6867, A0=>nx4884, A1=>nx4882);
   ix4885 : nor03_2x port map ( Y=>nx4884, A0=>nx6871, A1=>nx10276, A2=>
      nx11396);
   gen_12_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_12_cmp_mReg_10, QB=>
      nx6871, D=>window_12_10, CLK=>start, R=>rst);
   ix4883 : nor03_2x port map ( Y=>nx4882, A0=>gen_12_cmp_mReg_10, A1=>
      nx10804, A2=>nx11404);
   ix4919 : nand02 port map ( Y=>gen_12_cmp_BSCmp_op2_11, A0=>nx6875, A1=>
      nx6881);
   ix6876 : nor02_2x port map ( Y=>nx6875, A0=>nx4914, A1=>nx4910);
   ix4915 : nor03_2x port map ( Y=>nx4914, A0=>gen_12_cmp_mReg_10, A1=>
      nx10282, A2=>nx11372);
   ix4911 : nor03_2x port map ( Y=>nx4910, A0=>nx6871, A1=>nx11378, A2=>
      nx11388);
   ix6882 : nor02_2x port map ( Y=>nx6881, A0=>nx4906, A1=>nx4904);
   ix4907 : nor03_2x port map ( Y=>nx4906, A0=>nx6885, A1=>nx10276, A2=>
      nx11396);
   gen_12_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_12_cmp_mReg_11, QB=>
      nx6885, D=>window_12_11, CLK=>start, R=>rst);
   ix4905 : nor03_2x port map ( Y=>nx4904, A0=>gen_12_cmp_mReg_11, A1=>
      nx10804, A2=>nx11404);
   ix4941 : nand02 port map ( Y=>gen_12_cmp_BSCmp_op2_12, A0=>nx6889, A1=>
      nx6895);
   ix6890 : nor02_2x port map ( Y=>nx6889, A0=>nx4936, A1=>nx4932);
   ix4937 : nor03_2x port map ( Y=>nx4936, A0=>gen_12_cmp_mReg_11, A1=>
      nx10282, A2=>nx11372);
   ix4933 : nor03_2x port map ( Y=>nx4932, A0=>nx6885, A1=>nx11378, A2=>
      nx11388);
   ix6896 : nor02_2x port map ( Y=>nx6895, A0=>nx4928, A1=>nx4926);
   ix4929 : nor03_2x port map ( Y=>nx4928, A0=>nx6898, A1=>nx10278, A2=>
      nx11396);
   gen_12_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_12_cmp_mReg_12, QB=>
      nx6898, D=>window_12_12, CLK=>start, R=>rst);
   ix4927 : nor03_2x port map ( Y=>nx4926, A0=>gen_12_cmp_mReg_12, A1=>
      nx10804, A2=>nx11404);
   ix4963 : nand02 port map ( Y=>gen_12_cmp_BSCmp_op2_13, A0=>nx6905, A1=>
      nx6911);
   ix6906 : nor02_2x port map ( Y=>nx6905, A0=>nx4958, A1=>nx4954);
   ix4959 : nor03_2x port map ( Y=>nx4958, A0=>gen_12_cmp_mReg_12, A1=>
      nx10284, A2=>nx11374);
   ix4955 : nor03_2x port map ( Y=>nx4954, A0=>nx6898, A1=>nx11378, A2=>
      nx11390);
   ix6912 : nor02_2x port map ( Y=>nx6911, A0=>nx4950, A1=>nx4948);
   ix4951 : nor03_2x port map ( Y=>nx4950, A0=>nx6915, A1=>nx10278, A2=>
      nx11398);
   gen_12_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_12_cmp_mReg_13, QB=>
      nx6915, D=>window_12_13, CLK=>start, R=>rst);
   ix4949 : nor03_2x port map ( Y=>nx4948, A0=>gen_12_cmp_mReg_13, A1=>
      nx10804, A2=>nx11406);
   ix4985 : nand02 port map ( Y=>gen_12_cmp_BSCmp_op2_14, A0=>nx6919, A1=>
      nx6925);
   ix6920 : nor02_2x port map ( Y=>nx6919, A0=>nx4980, A1=>nx4976);
   ix4981 : nor03_2x port map ( Y=>nx4980, A0=>gen_12_cmp_mReg_13, A1=>
      nx10284, A2=>nx11374);
   ix4977 : nor03_2x port map ( Y=>nx4976, A0=>nx6915, A1=>nx11380, A2=>
      nx11390);
   ix6926 : nor02_2x port map ( Y=>nx6925, A0=>nx4972, A1=>nx4970);
   ix4973 : nor03_2x port map ( Y=>nx4972, A0=>nx6929, A1=>nx10278, A2=>
      nx11398);
   gen_12_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_12_cmp_mReg_14, QB=>
      nx6929, D=>window_12_14, CLK=>start, R=>rst);
   ix4971 : nor03_2x port map ( Y=>nx4970, A0=>gen_12_cmp_mReg_14, A1=>
      nx10804, A2=>nx11406);
   ix5007 : nand02 port map ( Y=>gen_12_cmp_BSCmp_op2_15, A0=>nx6933, A1=>
      nx6939);
   ix6934 : nor02_2x port map ( Y=>nx6933, A0=>nx5002, A1=>nx4998);
   ix5003 : nor03_2x port map ( Y=>nx5002, A0=>gen_12_cmp_mReg_14, A1=>
      nx10284, A2=>nx11374);
   ix4999 : nor03_2x port map ( Y=>nx4998, A0=>nx6929, A1=>nx11380, A2=>
      nx11390);
   ix6940 : nor02_2x port map ( Y=>nx6939, A0=>nx4994, A1=>nx4992);
   ix4995 : nor03_2x port map ( Y=>nx4994, A0=>nx6943, A1=>nx10278, A2=>
      nx11398);
   gen_12_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_12_cmp_mReg_15, QB=>
      nx6943, D=>window_12_15, CLK=>start, R=>rst);
   ix4993 : nor03_2x port map ( Y=>nx4992, A0=>gen_12_cmp_mReg_15, A1=>
      nx10806, A2=>nx11406);
   ix5017 : nand02 port map ( Y=>gen_12_cmp_BSCmp_op2_16, A0=>nx6949, A1=>
      nx6939);
   ix6950 : nor02_2x port map ( Y=>nx6949, A0=>nx5012, A1=>nx5008);
   ix5013 : nor03_2x port map ( Y=>nx5012, A0=>gen_12_cmp_mReg_15, A1=>
      nx10284, A2=>nx11374);
   ix5009 : nor03_2x port map ( Y=>nx5008, A0=>nx6943, A1=>nx11380, A2=>
      nx11390);
   ix5085 : nand02 port map ( Y=>gen_13_cmp_BSCmp_op2_1, A0=>nx6957, A1=>
      nx6975);
   ix6958 : nor02_2x port map ( Y=>nx6957, A0=>nx5080, A1=>nx5076);
   ix5081 : nor03_2x port map ( Y=>nx5080, A0=>gen_13_cmp_mReg_0, A1=>
      nx10268, A2=>nx11410);
   gen_13_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_13_cmp_mReg_0, QB=>
      nx6961, D=>window_13_0, CLK=>start, R=>rst);
   ix6966 : inv01 port map ( Y=>nx6965, A=>gen_13_cmp_pMux_0);
   ix5077 : nor03_2x port map ( Y=>nx5076, A0=>nx6961, A1=>nx11416, A2=>
      nx11426);
   ix6974 : inv02 port map ( Y=>nx6973, A=>gen_13_cmp_pMux_2);
   ix6976 : nor02_2x port map ( Y=>nx6975, A0=>nx5066, A1=>nx5064);
   ix5067 : nor03_2x port map ( Y=>nx5066, A0=>nx6979, A1=>nx10262, A2=>
      nx11434);
   gen_13_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_13_cmp_mReg_1, QB=>
      nx6979, D=>window_13_1, CLK=>start, R=>rst);
   ix5065 : nor03_2x port map ( Y=>nx5064, A0=>gen_13_cmp_mReg_1, A1=>
      nx10808, A2=>nx11442);
   ix5025 : nor03_2x port map ( Y=>nx5024, A0=>nx10268, A1=>nx6973, A2=>
      gen_13_cmp_pMux_0);
   ix5107 : nand02 port map ( Y=>gen_13_cmp_BSCmp_op2_2, A0=>nx6990, A1=>
      nx6995);
   ix6991 : nor02_2x port map ( Y=>nx6990, A0=>nx5102, A1=>nx5098);
   ix5103 : nor03_2x port map ( Y=>nx5102, A0=>gen_13_cmp_mReg_1, A1=>
      nx10268, A2=>nx11410);
   ix5099 : nor03_2x port map ( Y=>nx5098, A0=>nx6979, A1=>nx11416, A2=>
      nx11426);
   ix6996 : nor02_2x port map ( Y=>nx6995, A0=>nx5094, A1=>nx5092);
   ix5095 : nor03_2x port map ( Y=>nx5094, A0=>nx6999, A1=>nx10262, A2=>
      nx11434);
   gen_13_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_13_cmp_mReg_2, QB=>
      nx6999, D=>window_13_2, CLK=>start, R=>rst);
   ix5093 : nor03_2x port map ( Y=>nx5092, A0=>gen_13_cmp_mReg_2, A1=>
      nx10808, A2=>nx11442);
   ix5129 : nand02 port map ( Y=>gen_13_cmp_BSCmp_op2_3, A0=>nx7003, A1=>
      nx7009);
   ix7004 : nor02_2x port map ( Y=>nx7003, A0=>nx5124, A1=>nx5120);
   ix5125 : nor03_2x port map ( Y=>nx5124, A0=>gen_13_cmp_mReg_2, A1=>
      nx10268, A2=>nx11410);
   ix5121 : nor03_2x port map ( Y=>nx5120, A0=>nx6999, A1=>nx11416, A2=>
      nx11426);
   ix7010 : nor02_2x port map ( Y=>nx7009, A0=>nx5116, A1=>nx5114);
   ix5117 : nor03_2x port map ( Y=>nx5116, A0=>nx7013, A1=>nx10262, A2=>
      nx11434);
   gen_13_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_13_cmp_mReg_3, QB=>
      nx7013, D=>window_13_3, CLK=>start, R=>rst);
   ix5115 : nor03_2x port map ( Y=>nx5114, A0=>gen_13_cmp_mReg_3, A1=>
      nx10808, A2=>nx11442);
   ix5151 : nand02 port map ( Y=>gen_13_cmp_BSCmp_op2_4, A0=>nx7018, A1=>
      nx7023);
   ix7019 : nor02_2x port map ( Y=>nx7018, A0=>nx5146, A1=>nx5142);
   ix5147 : nor03_2x port map ( Y=>nx5146, A0=>gen_13_cmp_mReg_3, A1=>
      nx10268, A2=>nx11410);
   ix5143 : nor03_2x port map ( Y=>nx5142, A0=>nx7013, A1=>nx11416, A2=>
      nx11426);
   ix7024 : nor02_2x port map ( Y=>nx7023, A0=>nx5138, A1=>nx5136);
   ix5139 : nor03_2x port map ( Y=>nx5138, A0=>nx7027, A1=>nx10262, A2=>
      nx11434);
   gen_13_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_13_cmp_mReg_4, QB=>
      nx7027, D=>window_13_4, CLK=>start, R=>rst);
   ix5137 : nor03_2x port map ( Y=>nx5136, A0=>gen_13_cmp_mReg_4, A1=>
      nx10808, A2=>nx11442);
   ix5173 : nand02 port map ( Y=>gen_13_cmp_BSCmp_op2_5, A0=>nx7033, A1=>
      nx7039);
   ix7034 : nor02_2x port map ( Y=>nx7033, A0=>nx5168, A1=>nx5164);
   ix5169 : nor03_2x port map ( Y=>nx5168, A0=>gen_13_cmp_mReg_4, A1=>
      nx10268, A2=>nx11410);
   ix5165 : nor03_2x port map ( Y=>nx5164, A0=>nx7027, A1=>nx11416, A2=>
      nx11426);
   ix7040 : nor02_2x port map ( Y=>nx7039, A0=>nx5160, A1=>nx5158);
   ix5161 : nor03_2x port map ( Y=>nx5160, A0=>nx7042, A1=>nx10264, A2=>
      nx11434);
   gen_13_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_13_cmp_mReg_5, QB=>
      nx7042, D=>window_13_5, CLK=>start, R=>rst);
   ix5159 : nor03_2x port map ( Y=>nx5158, A0=>gen_13_cmp_mReg_5, A1=>
      nx10808, A2=>nx11442);
   ix5195 : nand02 port map ( Y=>gen_13_cmp_BSCmp_op2_6, A0=>nx7049, A1=>
      nx7055);
   ix7050 : nor02_2x port map ( Y=>nx7049, A0=>nx5190, A1=>nx5186);
   ix5191 : nor03_2x port map ( Y=>nx5190, A0=>gen_13_cmp_mReg_5, A1=>
      nx10270, A2=>nx11410);
   ix5187 : nor03_2x port map ( Y=>nx5186, A0=>nx7042, A1=>nx11416, A2=>
      nx11426);
   ix7056 : nor02_2x port map ( Y=>nx7055, A0=>nx5182, A1=>nx5180);
   ix5183 : nor03_2x port map ( Y=>nx5182, A0=>nx7059, A1=>nx10264, A2=>
      nx11434);
   gen_13_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_13_cmp_mReg_6, QB=>
      nx7059, D=>window_13_6, CLK=>start, R=>rst);
   ix5181 : nor03_2x port map ( Y=>nx5180, A0=>gen_13_cmp_mReg_6, A1=>
      nx10808, A2=>nx11442);
   ix5217 : nand02 port map ( Y=>gen_13_cmp_BSCmp_op2_7, A0=>nx7063, A1=>
      nx7069);
   ix7064 : nor02_2x port map ( Y=>nx7063, A0=>nx5212, A1=>nx5208);
   ix5213 : nor03_2x port map ( Y=>nx5212, A0=>gen_13_cmp_mReg_6, A1=>
      nx10270, A2=>nx11412);
   ix5209 : nor03_2x port map ( Y=>nx5208, A0=>nx7059, A1=>nx11418, A2=>
      nx11428);
   ix7070 : nor02_2x port map ( Y=>nx7069, A0=>nx5204, A1=>nx5202);
   ix5205 : nor03_2x port map ( Y=>nx5204, A0=>nx7073, A1=>nx10264, A2=>
      nx11436);
   gen_13_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_13_cmp_mReg_7, QB=>
      nx7073, D=>window_13_7, CLK=>start, R=>rst);
   ix5203 : nor03_2x port map ( Y=>nx5202, A0=>gen_13_cmp_mReg_7, A1=>
      nx10808, A2=>nx11444);
   ix5239 : nand02 port map ( Y=>gen_13_cmp_BSCmp_op2_8, A0=>nx7077, A1=>
      nx7083);
   ix7078 : nor02_2x port map ( Y=>nx7077, A0=>nx5234, A1=>nx5230);
   ix5235 : nor03_2x port map ( Y=>nx5234, A0=>gen_13_cmp_mReg_7, A1=>
      nx10270, A2=>nx11412);
   ix5231 : nor03_2x port map ( Y=>nx5230, A0=>nx7073, A1=>nx11418, A2=>
      nx11428);
   ix7084 : nor02_2x port map ( Y=>nx7083, A0=>nx5226, A1=>nx5224);
   ix5227 : nor03_2x port map ( Y=>nx5226, A0=>nx7086, A1=>nx10264, A2=>
      nx11436);
   gen_13_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_13_cmp_mReg_8, QB=>
      nx7086, D=>window_13_8, CLK=>start, R=>rst);
   ix5225 : nor03_2x port map ( Y=>nx5224, A0=>gen_13_cmp_mReg_8, A1=>
      nx10810, A2=>nx11444);
   ix5261 : nand02 port map ( Y=>gen_13_cmp_BSCmp_op2_9, A0=>nx7093, A1=>
      nx7099);
   ix7094 : nor02_2x port map ( Y=>nx7093, A0=>nx5256, A1=>nx5252);
   ix5257 : nor03_2x port map ( Y=>nx5256, A0=>gen_13_cmp_mReg_8, A1=>
      nx10270, A2=>nx11412);
   ix5253 : nor03_2x port map ( Y=>nx5252, A0=>nx7086, A1=>nx11418, A2=>
      nx11428);
   ix7100 : nor02_2x port map ( Y=>nx7099, A0=>nx5248, A1=>nx5246);
   ix5249 : nor03_2x port map ( Y=>nx5248, A0=>nx7103, A1=>nx10264, A2=>
      nx11436);
   gen_13_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_13_cmp_mReg_9, QB=>
      nx7103, D=>window_13_9, CLK=>start, R=>rst);
   ix5247 : nor03_2x port map ( Y=>nx5246, A0=>gen_13_cmp_mReg_9, A1=>
      nx10810, A2=>nx11444);
   ix5283 : nand02 port map ( Y=>gen_13_cmp_BSCmp_op2_10, A0=>nx7107, A1=>
      nx7113);
   ix7108 : nor02_2x port map ( Y=>nx7107, A0=>nx5278, A1=>nx5274);
   ix5279 : nor03_2x port map ( Y=>nx5278, A0=>gen_13_cmp_mReg_9, A1=>
      nx10270, A2=>nx11412);
   ix5275 : nor03_2x port map ( Y=>nx5274, A0=>nx7103, A1=>nx11418, A2=>
      nx11428);
   ix7114 : nor02_2x port map ( Y=>nx7113, A0=>nx5270, A1=>nx5268);
   ix5271 : nor03_2x port map ( Y=>nx5270, A0=>nx7117, A1=>nx10264, A2=>
      nx11436);
   gen_13_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_13_cmp_mReg_10, QB=>
      nx7117, D=>window_13_10, CLK=>start, R=>rst);
   ix5269 : nor03_2x port map ( Y=>nx5268, A0=>gen_13_cmp_mReg_10, A1=>
      nx10810, A2=>nx11444);
   ix5305 : nand02 port map ( Y=>gen_13_cmp_BSCmp_op2_11, A0=>nx7121, A1=>
      nx7127);
   ix7122 : nor02_2x port map ( Y=>nx7121, A0=>nx5300, A1=>nx5296);
   ix5301 : nor03_2x port map ( Y=>nx5300, A0=>gen_13_cmp_mReg_10, A1=>
      nx10270, A2=>nx11412);
   ix5297 : nor03_2x port map ( Y=>nx5296, A0=>nx7117, A1=>nx11418, A2=>
      nx11428);
   ix7128 : nor02_2x port map ( Y=>nx7127, A0=>nx5292, A1=>nx5290);
   ix5293 : nor03_2x port map ( Y=>nx5292, A0=>nx7130, A1=>nx10264, A2=>
      nx11436);
   gen_13_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_13_cmp_mReg_11, QB=>
      nx7130, D=>window_13_11, CLK=>start, R=>rst);
   ix5291 : nor03_2x port map ( Y=>nx5290, A0=>gen_13_cmp_mReg_11, A1=>
      nx10810, A2=>nx11444);
   ix5327 : nand02 port map ( Y=>gen_13_cmp_BSCmp_op2_12, A0=>nx7137, A1=>
      nx7143);
   ix7138 : nor02_2x port map ( Y=>nx7137, A0=>nx5322, A1=>nx5318);
   ix5323 : nor03_2x port map ( Y=>nx5322, A0=>gen_13_cmp_mReg_11, A1=>
      nx10270, A2=>nx11412);
   ix5319 : nor03_2x port map ( Y=>nx5318, A0=>nx7130, A1=>nx11418, A2=>
      nx11428);
   ix7144 : nor02_2x port map ( Y=>nx7143, A0=>nx5314, A1=>nx5312);
   ix5315 : nor03_2x port map ( Y=>nx5314, A0=>nx7147, A1=>nx10266, A2=>
      nx11436);
   gen_13_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_13_cmp_mReg_12, QB=>
      nx7147, D=>window_13_12, CLK=>start, R=>rst);
   ix5313 : nor03_2x port map ( Y=>nx5312, A0=>gen_13_cmp_mReg_12, A1=>
      nx10810, A2=>nx11444);
   ix5349 : nand02 port map ( Y=>gen_13_cmp_BSCmp_op2_13, A0=>nx7151, A1=>
      nx7157);
   ix7152 : nor02_2x port map ( Y=>nx7151, A0=>nx5344, A1=>nx5340);
   ix5345 : nor03_2x port map ( Y=>nx5344, A0=>gen_13_cmp_mReg_12, A1=>
      nx10272, A2=>nx11414);
   ix5341 : nor03_2x port map ( Y=>nx5340, A0=>nx7147, A1=>nx11418, A2=>
      nx11430);
   ix7158 : nor02_2x port map ( Y=>nx7157, A0=>nx5336, A1=>nx5334);
   ix5337 : nor03_2x port map ( Y=>nx5336, A0=>nx7161, A1=>nx10266, A2=>
      nx11438);
   gen_13_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_13_cmp_mReg_13, QB=>
      nx7161, D=>window_13_13, CLK=>start, R=>rst);
   ix5335 : nor03_2x port map ( Y=>nx5334, A0=>gen_13_cmp_mReg_13, A1=>
      nx10810, A2=>nx11446);
   ix5371 : nand02 port map ( Y=>gen_13_cmp_BSCmp_op2_14, A0=>nx7165, A1=>
      nx7171);
   ix7166 : nor02_2x port map ( Y=>nx7165, A0=>nx5366, A1=>nx5362);
   ix5367 : nor03_2x port map ( Y=>nx5366, A0=>gen_13_cmp_mReg_13, A1=>
      nx10272, A2=>nx11414);
   ix5363 : nor03_2x port map ( Y=>nx5362, A0=>nx7161, A1=>nx11420, A2=>
      nx11430);
   ix7172 : nor02_2x port map ( Y=>nx7171, A0=>nx5358, A1=>nx5356);
   ix5359 : nor03_2x port map ( Y=>nx5358, A0=>nx7174, A1=>nx10266, A2=>
      nx11438);
   gen_13_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_13_cmp_mReg_14, QB=>
      nx7174, D=>window_13_14, CLK=>start, R=>rst);
   ix5357 : nor03_2x port map ( Y=>nx5356, A0=>gen_13_cmp_mReg_14, A1=>
      nx10810, A2=>nx11446);
   ix5393 : nand02 port map ( Y=>gen_13_cmp_BSCmp_op2_15, A0=>nx7181, A1=>
      nx7187);
   ix7182 : nor02_2x port map ( Y=>nx7181, A0=>nx5388, A1=>nx5384);
   ix5389 : nor03_2x port map ( Y=>nx5388, A0=>gen_13_cmp_mReg_14, A1=>
      nx10272, A2=>nx11414);
   ix5385 : nor03_2x port map ( Y=>nx5384, A0=>nx7174, A1=>nx11420, A2=>
      nx11430);
   ix7188 : nor02_2x port map ( Y=>nx7187, A0=>nx5380, A1=>nx5378);
   ix5381 : nor03_2x port map ( Y=>nx5380, A0=>nx7191, A1=>nx10266, A2=>
      nx11438);
   gen_13_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_13_cmp_mReg_15, QB=>
      nx7191, D=>window_13_15, CLK=>start, R=>rst);
   ix5379 : nor03_2x port map ( Y=>nx5378, A0=>gen_13_cmp_mReg_15, A1=>
      nx10812, A2=>nx11446);
   ix5403 : nand02 port map ( Y=>gen_13_cmp_BSCmp_op2_16, A0=>nx7195, A1=>
      nx7187);
   ix7196 : nor02_2x port map ( Y=>nx7195, A0=>nx5398, A1=>nx5394);
   ix5399 : nor03_2x port map ( Y=>nx5398, A0=>gen_13_cmp_mReg_15, A1=>
      nx10272, A2=>nx11414);
   ix5395 : nor03_2x port map ( Y=>nx5394, A0=>nx7191, A1=>nx11420, A2=>
      nx11430);
   ix5471 : nand02 port map ( Y=>gen_14_cmp_BSCmp_op2_1, A0=>nx7203, A1=>
      nx7223);
   ix7204 : nor02_2x port map ( Y=>nx7203, A0=>nx5466, A1=>nx5462);
   ix5467 : nor03_2x port map ( Y=>nx5466, A0=>gen_14_cmp_mReg_0, A1=>
      nx10256, A2=>nx11450);
   gen_14_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_14_cmp_mReg_0, QB=>
      nx7209, D=>window_14_0, CLK=>start, R=>rst);
   ix7214 : inv01 port map ( Y=>nx7213, A=>gen_14_cmp_pMux_0);
   ix5463 : nor03_2x port map ( Y=>nx5462, A0=>nx7209, A1=>nx11456, A2=>
      nx11466);
   ix7222 : inv02 port map ( Y=>nx7221, A=>gen_14_cmp_pMux_2);
   ix7224 : nor02_2x port map ( Y=>nx7223, A0=>nx5452, A1=>nx5450);
   ix5453 : nor03_2x port map ( Y=>nx5452, A0=>nx7227, A1=>nx10250, A2=>
      nx11474);
   gen_14_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_14_cmp_mReg_1, QB=>
      nx7227, D=>window_14_1, CLK=>start, R=>rst);
   ix5451 : nor03_2x port map ( Y=>nx5450, A0=>gen_14_cmp_mReg_1, A1=>
      nx10814, A2=>nx11482);
   ix5411 : nor03_2x port map ( Y=>nx5410, A0=>nx10256, A1=>nx7221, A2=>
      gen_14_cmp_pMux_0);
   ix5493 : nand02 port map ( Y=>gen_14_cmp_BSCmp_op2_2, A0=>nx7238, A1=>
      nx7243);
   ix7239 : nor02_2x port map ( Y=>nx7238, A0=>nx5488, A1=>nx5484);
   ix5489 : nor03_2x port map ( Y=>nx5488, A0=>gen_14_cmp_mReg_1, A1=>
      nx10256, A2=>nx11450);
   ix5485 : nor03_2x port map ( Y=>nx5484, A0=>nx7227, A1=>nx11456, A2=>
      nx11466);
   ix7244 : nor02_2x port map ( Y=>nx7243, A0=>nx5480, A1=>nx5478);
   ix5481 : nor03_2x port map ( Y=>nx5480, A0=>nx7247, A1=>nx10250, A2=>
      nx11474);
   gen_14_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_14_cmp_mReg_2, QB=>
      nx7247, D=>window_14_2, CLK=>start, R=>rst);
   ix5479 : nor03_2x port map ( Y=>nx5478, A0=>gen_14_cmp_mReg_2, A1=>
      nx10814, A2=>nx11482);
   ix5515 : nand02 port map ( Y=>gen_14_cmp_BSCmp_op2_3, A0=>nx7253, A1=>
      nx7259);
   ix7254 : nor02_2x port map ( Y=>nx7253, A0=>nx5510, A1=>nx5506);
   ix5511 : nor03_2x port map ( Y=>nx5510, A0=>gen_14_cmp_mReg_2, A1=>
      nx10256, A2=>nx11450);
   ix5507 : nor03_2x port map ( Y=>nx5506, A0=>nx7247, A1=>nx11456, A2=>
      nx11466);
   ix7260 : nor02_2x port map ( Y=>nx7259, A0=>nx5502, A1=>nx5500);
   ix5503 : nor03_2x port map ( Y=>nx5502, A0=>nx7262, A1=>nx10250, A2=>
      nx11474);
   gen_14_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_14_cmp_mReg_3, QB=>
      nx7262, D=>window_14_3, CLK=>start, R=>rst);
   ix5501 : nor03_2x port map ( Y=>nx5500, A0=>gen_14_cmp_mReg_3, A1=>
      nx10814, A2=>nx11482);
   ix5537 : nand02 port map ( Y=>gen_14_cmp_BSCmp_op2_4, A0=>nx7269, A1=>
      nx7275);
   ix7270 : nor02_2x port map ( Y=>nx7269, A0=>nx5532, A1=>nx5528);
   ix5533 : nor03_2x port map ( Y=>nx5532, A0=>gen_14_cmp_mReg_3, A1=>
      nx10256, A2=>nx11450);
   ix5529 : nor03_2x port map ( Y=>nx5528, A0=>nx7262, A1=>nx11456, A2=>
      nx11466);
   ix7276 : nor02_2x port map ( Y=>nx7275, A0=>nx5524, A1=>nx5522);
   ix5525 : nor03_2x port map ( Y=>nx5524, A0=>nx7279, A1=>nx10250, A2=>
      nx11474);
   gen_14_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_14_cmp_mReg_4, QB=>
      nx7279, D=>window_14_4, CLK=>start, R=>rst);
   ix5523 : nor03_2x port map ( Y=>nx5522, A0=>gen_14_cmp_mReg_4, A1=>
      nx10814, A2=>nx11482);
   ix5559 : nand02 port map ( Y=>gen_14_cmp_BSCmp_op2_5, A0=>nx7283, A1=>
      nx7289);
   ix7284 : nor02_2x port map ( Y=>nx7283, A0=>nx5554, A1=>nx5550);
   ix5555 : nor03_2x port map ( Y=>nx5554, A0=>gen_14_cmp_mReg_4, A1=>
      nx10256, A2=>nx11450);
   ix5551 : nor03_2x port map ( Y=>nx5550, A0=>nx7279, A1=>nx11456, A2=>
      nx11466);
   ix7290 : nor02_2x port map ( Y=>nx7289, A0=>nx5546, A1=>nx5544);
   ix5547 : nor03_2x port map ( Y=>nx5546, A0=>nx7293, A1=>nx10252, A2=>
      nx11474);
   gen_14_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_14_cmp_mReg_5, QB=>
      nx7293, D=>window_14_5, CLK=>start, R=>rst);
   ix5545 : nor03_2x port map ( Y=>nx5544, A0=>gen_14_cmp_mReg_5, A1=>
      nx10814, A2=>nx11482);
   ix5581 : nand02 port map ( Y=>gen_14_cmp_BSCmp_op2_6, A0=>nx7297, A1=>
      nx7303);
   ix7298 : nor02_2x port map ( Y=>nx7297, A0=>nx5576, A1=>nx5572);
   ix5577 : nor03_2x port map ( Y=>nx5576, A0=>gen_14_cmp_mReg_5, A1=>
      nx10258, A2=>nx11450);
   ix5573 : nor03_2x port map ( Y=>nx5572, A0=>nx7293, A1=>nx11456, A2=>
      nx11466);
   ix7304 : nor02_2x port map ( Y=>nx7303, A0=>nx5568, A1=>nx5566);
   ix5569 : nor03_2x port map ( Y=>nx5568, A0=>nx7306, A1=>nx10252, A2=>
      nx11474);
   gen_14_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_14_cmp_mReg_6, QB=>
      nx7306, D=>window_14_6, CLK=>start, R=>rst);
   ix5567 : nor03_2x port map ( Y=>nx5566, A0=>gen_14_cmp_mReg_6, A1=>
      nx10814, A2=>nx11482);
   ix5603 : nand02 port map ( Y=>gen_14_cmp_BSCmp_op2_7, A0=>nx7313, A1=>
      nx7319);
   ix7314 : nor02_2x port map ( Y=>nx7313, A0=>nx5598, A1=>nx5594);
   ix5599 : nor03_2x port map ( Y=>nx5598, A0=>gen_14_cmp_mReg_6, A1=>
      nx10258, A2=>nx11452);
   ix5595 : nor03_2x port map ( Y=>nx5594, A0=>nx7306, A1=>nx11458, A2=>
      nx11468);
   ix7320 : nor02_2x port map ( Y=>nx7319, A0=>nx5590, A1=>nx5588);
   ix5591 : nor03_2x port map ( Y=>nx5590, A0=>nx7323, A1=>nx10252, A2=>
      nx11476);
   gen_14_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_14_cmp_mReg_7, QB=>
      nx7323, D=>window_14_7, CLK=>start, R=>rst);
   ix5589 : nor03_2x port map ( Y=>nx5588, A0=>gen_14_cmp_mReg_7, A1=>
      nx10814, A2=>nx11484);
   ix5625 : nand02 port map ( Y=>gen_14_cmp_BSCmp_op2_8, A0=>nx7329, A1=>
      nx7335);
   ix7330 : nor02_2x port map ( Y=>nx7329, A0=>nx5620, A1=>nx5616);
   ix5621 : nor03_2x port map ( Y=>nx5620, A0=>gen_14_cmp_mReg_7, A1=>
      nx10258, A2=>nx11452);
   ix5617 : nor03_2x port map ( Y=>nx5616, A0=>nx7323, A1=>nx11458, A2=>
      nx11468);
   ix7336 : nor02_2x port map ( Y=>nx7335, A0=>nx5612, A1=>nx5610);
   ix5613 : nor03_2x port map ( Y=>nx5612, A0=>nx7339, A1=>nx10252, A2=>
      nx11476);
   gen_14_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_14_cmp_mReg_8, QB=>
      nx7339, D=>window_14_8, CLK=>start, R=>rst);
   ix5611 : nor03_2x port map ( Y=>nx5610, A0=>gen_14_cmp_mReg_8, A1=>
      nx10816, A2=>nx11484);
   ix5647 : nand02 port map ( Y=>gen_14_cmp_BSCmp_op2_9, A0=>nx7344, A1=>
      nx7348);
   ix7345 : nor02_2x port map ( Y=>nx7344, A0=>nx5642, A1=>nx5638);
   ix5643 : nor03_2x port map ( Y=>nx5642, A0=>gen_14_cmp_mReg_8, A1=>
      nx10258, A2=>nx11452);
   ix5639 : nor03_2x port map ( Y=>nx5638, A0=>nx7339, A1=>nx11458, A2=>
      nx11468);
   ix7349 : nor02_2x port map ( Y=>nx7348, A0=>nx5634, A1=>nx5632);
   ix5635 : nor03_2x port map ( Y=>nx5634, A0=>nx7351, A1=>nx10252, A2=>
      nx11476);
   gen_14_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_14_cmp_mReg_9, QB=>
      nx7351, D=>window_14_9, CLK=>start, R=>rst);
   ix5633 : nor03_2x port map ( Y=>nx5632, A0=>gen_14_cmp_mReg_9, A1=>
      nx10816, A2=>nx11484);
   ix5669 : nand02 port map ( Y=>gen_14_cmp_BSCmp_op2_10, A0=>nx7357, A1=>
      nx7363);
   ix7358 : nor02_2x port map ( Y=>nx7357, A0=>nx5664, A1=>nx5660);
   ix5665 : nor03_2x port map ( Y=>nx5664, A0=>gen_14_cmp_mReg_9, A1=>
      nx10258, A2=>nx11452);
   ix5661 : nor03_2x port map ( Y=>nx5660, A0=>nx7351, A1=>nx11458, A2=>
      nx11468);
   ix7364 : nor02_2x port map ( Y=>nx7363, A0=>nx5656, A1=>nx5654);
   ix5657 : nor03_2x port map ( Y=>nx5656, A0=>nx7367, A1=>nx10252, A2=>
      nx11476);
   gen_14_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_14_cmp_mReg_10, QB=>
      nx7367, D=>window_14_10, CLK=>start, R=>rst);
   ix5655 : nor03_2x port map ( Y=>nx5654, A0=>gen_14_cmp_mReg_10, A1=>
      nx10816, A2=>nx11484);
   ix5691 : nand02 port map ( Y=>gen_14_cmp_BSCmp_op2_11, A0=>nx7373, A1=>
      nx7377);
   ix7374 : nor02_2x port map ( Y=>nx7373, A0=>nx5686, A1=>nx5682);
   ix5687 : nor03_2x port map ( Y=>nx5686, A0=>gen_14_cmp_mReg_10, A1=>
      nx10258, A2=>nx11452);
   ix5683 : nor03_2x port map ( Y=>nx5682, A0=>nx7367, A1=>nx11458, A2=>
      nx11468);
   ix7378 : nor02_2x port map ( Y=>nx7377, A0=>nx5678, A1=>nx5676);
   ix5679 : nor03_2x port map ( Y=>nx5678, A0=>nx7381, A1=>nx10252, A2=>
      nx11476);
   gen_14_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_14_cmp_mReg_11, QB=>
      nx7381, D=>window_14_11, CLK=>start, R=>rst);
   ix5677 : nor03_2x port map ( Y=>nx5676, A0=>gen_14_cmp_mReg_11, A1=>
      nx10816, A2=>nx11484);
   ix5713 : nand02 port map ( Y=>gen_14_cmp_BSCmp_op2_12, A0=>nx7387, A1=>
      nx7393);
   ix7388 : nor02_2x port map ( Y=>nx7387, A0=>nx5708, A1=>nx5704);
   ix5709 : nor03_2x port map ( Y=>nx5708, A0=>gen_14_cmp_mReg_11, A1=>
      nx10258, A2=>nx11452);
   ix5705 : nor03_2x port map ( Y=>nx5704, A0=>nx7381, A1=>nx11458, A2=>
      nx11468);
   ix7394 : nor02_2x port map ( Y=>nx7393, A0=>nx5700, A1=>nx5698);
   ix5701 : nor03_2x port map ( Y=>nx5700, A0=>nx7397, A1=>nx10254, A2=>
      nx11476);
   gen_14_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_14_cmp_mReg_12, QB=>
      nx7397, D=>window_14_12, CLK=>start, R=>rst);
   ix5699 : nor03_2x port map ( Y=>nx5698, A0=>gen_14_cmp_mReg_12, A1=>
      nx10816, A2=>nx11484);
   ix5735 : nand02 port map ( Y=>gen_14_cmp_BSCmp_op2_13, A0=>nx7403, A1=>
      nx7407);
   ix7404 : nor02_2x port map ( Y=>nx7403, A0=>nx5730, A1=>nx5726);
   ix5731 : nor03_2x port map ( Y=>nx5730, A0=>gen_14_cmp_mReg_12, A1=>
      nx10260, A2=>nx11454);
   ix5727 : nor03_2x port map ( Y=>nx5726, A0=>nx7397, A1=>nx11458, A2=>
      nx11470);
   ix7408 : nor02_2x port map ( Y=>nx7407, A0=>nx5722, A1=>nx5720);
   ix5723 : nor03_2x port map ( Y=>nx5722, A0=>nx7411, A1=>nx10254, A2=>
      nx11478);
   gen_14_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_14_cmp_mReg_13, QB=>
      nx7411, D=>window_14_13, CLK=>start, R=>rst);
   ix5721 : nor03_2x port map ( Y=>nx5720, A0=>gen_14_cmp_mReg_13, A1=>
      nx10816, A2=>nx11486);
   ix5757 : nand02 port map ( Y=>gen_14_cmp_BSCmp_op2_14, A0=>nx7417, A1=>
      nx7423);
   ix7418 : nor02_2x port map ( Y=>nx7417, A0=>nx5752, A1=>nx5748);
   ix5753 : nor03_2x port map ( Y=>nx5752, A0=>gen_14_cmp_mReg_13, A1=>
      nx10260, A2=>nx11454);
   ix5749 : nor03_2x port map ( Y=>nx5748, A0=>nx7411, A1=>nx11460, A2=>
      nx11470);
   ix7424 : nor02_2x port map ( Y=>nx7423, A0=>nx5744, A1=>nx5742);
   ix5745 : nor03_2x port map ( Y=>nx5744, A0=>nx7426, A1=>nx10254, A2=>
      nx11478);
   gen_14_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_14_cmp_mReg_14, QB=>
      nx7426, D=>window_14_14, CLK=>start, R=>rst);
   ix5743 : nor03_2x port map ( Y=>nx5742, A0=>gen_14_cmp_mReg_14, A1=>
      nx10816, A2=>nx11486);
   ix5779 : nand02 port map ( Y=>gen_14_cmp_BSCmp_op2_15, A0=>nx7431, A1=>
      nx7437);
   ix7432 : nor02_2x port map ( Y=>nx7431, A0=>nx5774, A1=>nx5770);
   ix5775 : nor03_2x port map ( Y=>nx5774, A0=>gen_14_cmp_mReg_14, A1=>
      nx10260, A2=>nx11454);
   ix5771 : nor03_2x port map ( Y=>nx5770, A0=>nx7426, A1=>nx11460, A2=>
      nx11470);
   ix7438 : nor02_2x port map ( Y=>nx7437, A0=>nx5766, A1=>nx5764);
   ix5767 : nor03_2x port map ( Y=>nx5766, A0=>nx7441, A1=>nx10254, A2=>
      nx11478);
   gen_14_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_14_cmp_mReg_15, QB=>
      nx7441, D=>window_14_15, CLK=>start, R=>rst);
   ix5765 : nor03_2x port map ( Y=>nx5764, A0=>gen_14_cmp_mReg_15, A1=>
      nx10818, A2=>nx11486);
   ix5789 : nand02 port map ( Y=>gen_14_cmp_BSCmp_op2_16, A0=>nx7447, A1=>
      nx7437);
   ix7448 : nor02_2x port map ( Y=>nx7447, A0=>nx5784, A1=>nx5780);
   ix5785 : nor03_2x port map ( Y=>nx5784, A0=>gen_14_cmp_mReg_15, A1=>
      nx10260, A2=>nx11454);
   ix5781 : nor03_2x port map ( Y=>nx5780, A0=>nx7441, A1=>nx11460, A2=>
      nx11470);
   ix5857 : nand02 port map ( Y=>gen_15_cmp_BSCmp_op2_1, A0=>nx7453, A1=>
      nx7473);
   ix7454 : nor02_2x port map ( Y=>nx7453, A0=>nx5852, A1=>nx5848);
   ix5853 : nor03_2x port map ( Y=>nx5852, A0=>gen_15_cmp_mReg_0, A1=>
      nx10244, A2=>nx11490);
   gen_15_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_15_cmp_mReg_0, QB=>
      nx7459, D=>window_15_0, CLK=>start, R=>rst);
   ix7464 : inv01 port map ( Y=>nx7463, A=>gen_15_cmp_pMux_0);
   ix5849 : nor03_2x port map ( Y=>nx5848, A0=>nx7459, A1=>nx11496, A2=>
      nx11506);
   ix7472 : inv02 port map ( Y=>nx7471, A=>gen_15_cmp_pMux_2);
   ix7474 : nor02_2x port map ( Y=>nx7473, A0=>nx5838, A1=>nx5836);
   ix5839 : nor03_2x port map ( Y=>nx5838, A0=>nx7477, A1=>nx10238, A2=>
      nx11514);
   gen_15_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_15_cmp_mReg_1, QB=>
      nx7477, D=>window_15_1, CLK=>start, R=>rst);
   ix5837 : nor03_2x port map ( Y=>nx5836, A0=>gen_15_cmp_mReg_1, A1=>
      nx10820, A2=>nx11522);
   ix5797 : nor03_2x port map ( Y=>nx5796, A0=>nx10244, A1=>nx7471, A2=>
      gen_15_cmp_pMux_0);
   ix5879 : nand02 port map ( Y=>gen_15_cmp_BSCmp_op2_2, A0=>nx7489, A1=>
      nx7493);
   ix7490 : nor02_2x port map ( Y=>nx7489, A0=>nx5874, A1=>nx5870);
   ix5875 : nor03_2x port map ( Y=>nx5874, A0=>gen_15_cmp_mReg_1, A1=>
      nx10244, A2=>nx11490);
   ix5871 : nor03_2x port map ( Y=>nx5870, A0=>nx7477, A1=>nx11496, A2=>
      nx11506);
   ix7494 : nor02_2x port map ( Y=>nx7493, A0=>nx5866, A1=>nx5864);
   ix5867 : nor03_2x port map ( Y=>nx5866, A0=>nx7497, A1=>nx10238, A2=>
      nx11514);
   gen_15_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_15_cmp_mReg_2, QB=>
      nx7497, D=>window_15_2, CLK=>start, R=>rst);
   ix5865 : nor03_2x port map ( Y=>nx5864, A0=>gen_15_cmp_mReg_2, A1=>
      nx10820, A2=>nx11522);
   ix5901 : nand02 port map ( Y=>gen_15_cmp_BSCmp_op2_3, A0=>nx7503, A1=>
      nx7507);
   ix7504 : nor02_2x port map ( Y=>nx7503, A0=>nx5896, A1=>nx5892);
   ix5897 : nor03_2x port map ( Y=>nx5896, A0=>gen_15_cmp_mReg_2, A1=>
      nx10244, A2=>nx11490);
   ix5893 : nor03_2x port map ( Y=>nx5892, A0=>nx7497, A1=>nx11496, A2=>
      nx11506);
   ix7508 : nor02_2x port map ( Y=>nx7507, A0=>nx5888, A1=>nx5886);
   ix5889 : nor03_2x port map ( Y=>nx5888, A0=>nx7511, A1=>nx10238, A2=>
      nx11514);
   gen_15_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_15_cmp_mReg_3, QB=>
      nx7511, D=>window_15_3, CLK=>start, R=>rst);
   ix5887 : nor03_2x port map ( Y=>nx5886, A0=>gen_15_cmp_mReg_3, A1=>
      nx10820, A2=>nx11522);
   ix5923 : nand02 port map ( Y=>gen_15_cmp_BSCmp_op2_4, A0=>nx7515, A1=>
      nx7521);
   ix7516 : nor02_2x port map ( Y=>nx7515, A0=>nx5918, A1=>nx5914);
   ix5919 : nor03_2x port map ( Y=>nx5918, A0=>gen_15_cmp_mReg_3, A1=>
      nx10244, A2=>nx11490);
   ix5915 : nor03_2x port map ( Y=>nx5914, A0=>nx7511, A1=>nx11496, A2=>
      nx11506);
   ix7522 : nor02_2x port map ( Y=>nx7521, A0=>nx5910, A1=>nx5908);
   ix5911 : nor03_2x port map ( Y=>nx5910, A0=>nx7525, A1=>nx10238, A2=>
      nx11514);
   gen_15_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_15_cmp_mReg_4, QB=>
      nx7525, D=>window_15_4, CLK=>start, R=>rst);
   ix5909 : nor03_2x port map ( Y=>nx5908, A0=>gen_15_cmp_mReg_4, A1=>
      nx10820, A2=>nx11522);
   ix5945 : nand02 port map ( Y=>gen_15_cmp_BSCmp_op2_5, A0=>nx7529, A1=>
      nx7535);
   ix7530 : nor02_2x port map ( Y=>nx7529, A0=>nx5940, A1=>nx5936);
   ix5941 : nor03_2x port map ( Y=>nx5940, A0=>gen_15_cmp_mReg_4, A1=>
      nx10244, A2=>nx11490);
   ix5937 : nor03_2x port map ( Y=>nx5936, A0=>nx7525, A1=>nx11496, A2=>
      nx11506);
   ix7536 : nor02_2x port map ( Y=>nx7535, A0=>nx5932, A1=>nx5930);
   ix5933 : nor03_2x port map ( Y=>nx5932, A0=>nx7538, A1=>nx10240, A2=>
      nx11514);
   gen_15_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_15_cmp_mReg_5, QB=>
      nx7538, D=>window_15_5, CLK=>start, R=>rst);
   ix5931 : nor03_2x port map ( Y=>nx5930, A0=>gen_15_cmp_mReg_5, A1=>
      nx10820, A2=>nx11522);
   ix5967 : nand02 port map ( Y=>gen_15_cmp_BSCmp_op2_6, A0=>nx7545, A1=>
      nx7551);
   ix7546 : nor02_2x port map ( Y=>nx7545, A0=>nx5962, A1=>nx5958);
   ix5963 : nor03_2x port map ( Y=>nx5962, A0=>gen_15_cmp_mReg_5, A1=>
      nx10246, A2=>nx11490);
   ix5959 : nor03_2x port map ( Y=>nx5958, A0=>nx7538, A1=>nx11496, A2=>
      nx11506);
   ix7552 : nor02_2x port map ( Y=>nx7551, A0=>nx5954, A1=>nx5952);
   ix5955 : nor03_2x port map ( Y=>nx5954, A0=>nx7555, A1=>nx10240, A2=>
      nx11514);
   gen_15_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_15_cmp_mReg_6, QB=>
      nx7555, D=>window_15_6, CLK=>start, R=>rst);
   ix5953 : nor03_2x port map ( Y=>nx5952, A0=>gen_15_cmp_mReg_6, A1=>
      nx10820, A2=>nx11522);
   ix5989 : nand02 port map ( Y=>gen_15_cmp_BSCmp_op2_7, A0=>nx7559, A1=>
      nx7565);
   ix7560 : nor02_2x port map ( Y=>nx7559, A0=>nx5984, A1=>nx5980);
   ix5985 : nor03_2x port map ( Y=>nx5984, A0=>gen_15_cmp_mReg_6, A1=>
      nx10246, A2=>nx11492);
   ix5981 : nor03_2x port map ( Y=>nx5980, A0=>nx7555, A1=>nx11498, A2=>
      nx11508);
   ix7566 : nor02_2x port map ( Y=>nx7565, A0=>nx5976, A1=>nx5974);
   ix5977 : nor03_2x port map ( Y=>nx5976, A0=>nx7569, A1=>nx10240, A2=>
      nx11516);
   gen_15_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_15_cmp_mReg_7, QB=>
      nx7569, D=>window_15_7, CLK=>start, R=>rst);
   ix5975 : nor03_2x port map ( Y=>nx5974, A0=>gen_15_cmp_mReg_7, A1=>
      nx10820, A2=>nx11524);
   ix6011 : nand02 port map ( Y=>gen_15_cmp_BSCmp_op2_8, A0=>nx7573, A1=>
      nx7579);
   ix7574 : nor02_2x port map ( Y=>nx7573, A0=>nx6006, A1=>nx6002);
   ix6007 : nor03_2x port map ( Y=>nx6006, A0=>gen_15_cmp_mReg_7, A1=>
      nx10246, A2=>nx11492);
   ix6003 : nor03_2x port map ( Y=>nx6002, A0=>nx7569, A1=>nx11498, A2=>
      nx11508);
   ix7580 : nor02_2x port map ( Y=>nx7579, A0=>nx5998, A1=>nx5996);
   ix5999 : nor03_2x port map ( Y=>nx5998, A0=>nx7582, A1=>nx10240, A2=>
      nx11516);
   gen_15_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_15_cmp_mReg_8, QB=>
      nx7582, D=>window_15_8, CLK=>start, R=>rst);
   ix5997 : nor03_2x port map ( Y=>nx5996, A0=>gen_15_cmp_mReg_8, A1=>
      nx10822, A2=>nx11524);
   ix6033 : nand02 port map ( Y=>gen_15_cmp_BSCmp_op2_9, A0=>nx7589, A1=>
      nx7595);
   ix7590 : nor02_2x port map ( Y=>nx7589, A0=>nx6028, A1=>nx6024);
   ix6029 : nor03_2x port map ( Y=>nx6028, A0=>gen_15_cmp_mReg_8, A1=>
      nx10246, A2=>nx11492);
   ix6025 : nor03_2x port map ( Y=>nx6024, A0=>nx7582, A1=>nx11498, A2=>
      nx11508);
   ix7596 : nor02_2x port map ( Y=>nx7595, A0=>nx6020, A1=>nx6018);
   ix6021 : nor03_2x port map ( Y=>nx6020, A0=>nx7599, A1=>nx10240, A2=>
      nx11516);
   gen_15_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_15_cmp_mReg_9, QB=>
      nx7599, D=>window_15_9, CLK=>start, R=>rst);
   ix6019 : nor03_2x port map ( Y=>nx6018, A0=>gen_15_cmp_mReg_9, A1=>
      nx10822, A2=>nx11524);
   ix6055 : nand02 port map ( Y=>gen_15_cmp_BSCmp_op2_10, A0=>nx7603, A1=>
      nx7609);
   ix7604 : nor02_2x port map ( Y=>nx7603, A0=>nx6050, A1=>nx6046);
   ix6051 : nor03_2x port map ( Y=>nx6050, A0=>gen_15_cmp_mReg_9, A1=>
      nx10246, A2=>nx11492);
   ix6047 : nor03_2x port map ( Y=>nx6046, A0=>nx7599, A1=>nx11498, A2=>
      nx11508);
   ix7610 : nor02_2x port map ( Y=>nx7609, A0=>nx6042, A1=>nx6040);
   ix6043 : nor03_2x port map ( Y=>nx6042, A0=>nx7613, A1=>nx10240, A2=>
      nx11516);
   gen_15_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_15_cmp_mReg_10, QB=>
      nx7613, D=>window_15_10, CLK=>start, R=>rst);
   ix6041 : nor03_2x port map ( Y=>nx6040, A0=>gen_15_cmp_mReg_10, A1=>
      nx10822, A2=>nx11524);
   ix6077 : nand02 port map ( Y=>gen_15_cmp_BSCmp_op2_11, A0=>nx7617, A1=>
      nx7623);
   ix7618 : nor02_2x port map ( Y=>nx7617, A0=>nx6072, A1=>nx6068);
   ix6073 : nor03_2x port map ( Y=>nx6072, A0=>gen_15_cmp_mReg_10, A1=>
      nx10246, A2=>nx11492);
   ix6069 : nor03_2x port map ( Y=>nx6068, A0=>nx7613, A1=>nx11498, A2=>
      nx11508);
   ix7624 : nor02_2x port map ( Y=>nx7623, A0=>nx6064, A1=>nx6062);
   ix6065 : nor03_2x port map ( Y=>nx6064, A0=>nx7626, A1=>nx10240, A2=>
      nx11516);
   gen_15_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_15_cmp_mReg_11, QB=>
      nx7626, D=>window_15_11, CLK=>start, R=>rst);
   ix6063 : nor03_2x port map ( Y=>nx6062, A0=>gen_15_cmp_mReg_11, A1=>
      nx10822, A2=>nx11524);
   ix6099 : nand02 port map ( Y=>gen_15_cmp_BSCmp_op2_12, A0=>nx7633, A1=>
      nx7639);
   ix7634 : nor02_2x port map ( Y=>nx7633, A0=>nx6094, A1=>nx6090);
   ix6095 : nor03_2x port map ( Y=>nx6094, A0=>gen_15_cmp_mReg_11, A1=>
      nx10246, A2=>nx11492);
   ix6091 : nor03_2x port map ( Y=>nx6090, A0=>nx7626, A1=>nx11498, A2=>
      nx11508);
   ix7640 : nor02_2x port map ( Y=>nx7639, A0=>nx6086, A1=>nx6084);
   ix6087 : nor03_2x port map ( Y=>nx6086, A0=>nx7643, A1=>nx10242, A2=>
      nx11516);
   gen_15_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_15_cmp_mReg_12, QB=>
      nx7643, D=>window_15_12, CLK=>start, R=>rst);
   ix6085 : nor03_2x port map ( Y=>nx6084, A0=>gen_15_cmp_mReg_12, A1=>
      nx10822, A2=>nx11524);
   ix6121 : nand02 port map ( Y=>gen_15_cmp_BSCmp_op2_13, A0=>nx7647, A1=>
      nx7653);
   ix7648 : nor02_2x port map ( Y=>nx7647, A0=>nx6116, A1=>nx6112);
   ix6117 : nor03_2x port map ( Y=>nx6116, A0=>gen_15_cmp_mReg_12, A1=>
      nx10248, A2=>nx11494);
   ix6113 : nor03_2x port map ( Y=>nx6112, A0=>nx7643, A1=>nx11498, A2=>
      nx11510);
   ix7654 : nor02_2x port map ( Y=>nx7653, A0=>nx6108, A1=>nx6106);
   ix6109 : nor03_2x port map ( Y=>nx6108, A0=>nx7657, A1=>nx10242, A2=>
      nx11518);
   gen_15_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_15_cmp_mReg_13, QB=>
      nx7657, D=>window_15_13, CLK=>start, R=>rst);
   ix6107 : nor03_2x port map ( Y=>nx6106, A0=>gen_15_cmp_mReg_13, A1=>
      nx10822, A2=>nx11526);
   ix6143 : nand02 port map ( Y=>gen_15_cmp_BSCmp_op2_14, A0=>nx7661, A1=>
      nx7667);
   ix7662 : nor02_2x port map ( Y=>nx7661, A0=>nx6138, A1=>nx6134);
   ix6139 : nor03_2x port map ( Y=>nx6138, A0=>gen_15_cmp_mReg_13, A1=>
      nx10248, A2=>nx11494);
   ix6135 : nor03_2x port map ( Y=>nx6134, A0=>nx7657, A1=>nx11500, A2=>
      nx11510);
   ix7668 : nor02_2x port map ( Y=>nx7667, A0=>nx6130, A1=>nx6128);
   ix6131 : nor03_2x port map ( Y=>nx6130, A0=>nx7670, A1=>nx10242, A2=>
      nx11518);
   gen_15_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_15_cmp_mReg_14, QB=>
      nx7670, D=>window_15_14, CLK=>start, R=>rst);
   ix6129 : nor03_2x port map ( Y=>nx6128, A0=>gen_15_cmp_mReg_14, A1=>
      nx10822, A2=>nx11526);
   ix6165 : nand02 port map ( Y=>gen_15_cmp_BSCmp_op2_15, A0=>nx7677, A1=>
      nx7683);
   ix7678 : nor02_2x port map ( Y=>nx7677, A0=>nx6160, A1=>nx6156);
   ix6161 : nor03_2x port map ( Y=>nx6160, A0=>gen_15_cmp_mReg_14, A1=>
      nx10248, A2=>nx11494);
   ix6157 : nor03_2x port map ( Y=>nx6156, A0=>nx7670, A1=>nx11500, A2=>
      nx11510);
   ix7684 : nor02_2x port map ( Y=>nx7683, A0=>nx6152, A1=>nx6150);
   ix6153 : nor03_2x port map ( Y=>nx6152, A0=>nx7687, A1=>nx10242, A2=>
      nx11518);
   gen_15_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_15_cmp_mReg_15, QB=>
      nx7687, D=>window_15_15, CLK=>start, R=>rst);
   ix6151 : nor03_2x port map ( Y=>nx6150, A0=>gen_15_cmp_mReg_15, A1=>
      nx10824, A2=>nx11526);
   ix6175 : nand02 port map ( Y=>gen_15_cmp_BSCmp_op2_16, A0=>nx7691, A1=>
      nx7683);
   ix7692 : nor02_2x port map ( Y=>nx7691, A0=>nx6170, A1=>nx6166);
   ix6171 : nor03_2x port map ( Y=>nx6170, A0=>gen_15_cmp_mReg_15, A1=>
      nx10248, A2=>nx11494);
   ix6167 : nor03_2x port map ( Y=>nx6166, A0=>nx7687, A1=>nx11500, A2=>
      nx11510);
   ix6243 : nand02 port map ( Y=>gen_16_cmp_BSCmp_op2_1, A0=>nx7699, A1=>
      nx7719);
   ix7700 : nor02_2x port map ( Y=>nx7699, A0=>nx6238, A1=>nx6234);
   ix6239 : nor03_2x port map ( Y=>nx6238, A0=>gen_16_cmp_mReg_0, A1=>
      nx10232, A2=>nx11530);
   gen_16_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_16_cmp_mReg_0, QB=>
      nx7705, D=>window_16_0, CLK=>start, R=>rst);
   ix7710 : inv01 port map ( Y=>nx7709, A=>gen_16_cmp_pMux_0);
   ix6235 : nor03_2x port map ( Y=>nx6234, A0=>nx7705, A1=>nx11536, A2=>
      nx11546);
   ix7718 : inv02 port map ( Y=>nx7717, A=>gen_16_cmp_pMux_2);
   ix7720 : nor02_2x port map ( Y=>nx7719, A0=>nx6224, A1=>nx6222);
   ix6225 : nor03_2x port map ( Y=>nx6224, A0=>nx7723, A1=>nx10226, A2=>
      nx11554);
   gen_16_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_16_cmp_mReg_1, QB=>
      nx7723, D=>window_16_1, CLK=>start, R=>rst);
   ix6223 : nor03_2x port map ( Y=>nx6222, A0=>gen_16_cmp_mReg_1, A1=>
      nx10826, A2=>nx11562);
   ix6183 : nor03_2x port map ( Y=>nx6182, A0=>nx10232, A1=>nx7717, A2=>
      gen_16_cmp_pMux_0);
   ix6265 : nand02 port map ( Y=>gen_16_cmp_BSCmp_op2_2, A0=>nx7733, A1=>
      nx7737);
   ix7734 : nor02_2x port map ( Y=>nx7733, A0=>nx6260, A1=>nx6256);
   ix6261 : nor03_2x port map ( Y=>nx6260, A0=>gen_16_cmp_mReg_1, A1=>
      nx10232, A2=>nx11530);
   ix6257 : nor03_2x port map ( Y=>nx6256, A0=>nx7723, A1=>nx11536, A2=>
      nx11546);
   ix7738 : nor02_2x port map ( Y=>nx7737, A0=>nx6252, A1=>nx6250);
   ix6253 : nor03_2x port map ( Y=>nx6252, A0=>nx7741, A1=>nx10226, A2=>
      nx11554);
   gen_16_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_16_cmp_mReg_2, QB=>
      nx7741, D=>window_16_2, CLK=>start, R=>rst);
   ix6251 : nor03_2x port map ( Y=>nx6250, A0=>gen_16_cmp_mReg_2, A1=>
      nx10826, A2=>nx11562);
   ix6287 : nand02 port map ( Y=>gen_16_cmp_BSCmp_op2_3, A0=>nx7747, A1=>
      nx7753);
   ix7748 : nor02_2x port map ( Y=>nx7747, A0=>nx6282, A1=>nx6278);
   ix6283 : nor03_2x port map ( Y=>nx6282, A0=>gen_16_cmp_mReg_2, A1=>
      nx10232, A2=>nx11530);
   ix6279 : nor03_2x port map ( Y=>nx6278, A0=>nx7741, A1=>nx11536, A2=>
      nx11546);
   ix7754 : nor02_2x port map ( Y=>nx7753, A0=>nx6274, A1=>nx6272);
   ix6275 : nor03_2x port map ( Y=>nx6274, A0=>nx7757, A1=>nx10226, A2=>
      nx11554);
   gen_16_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_16_cmp_mReg_3, QB=>
      nx7757, D=>window_16_3, CLK=>start, R=>rst);
   ix6273 : nor03_2x port map ( Y=>nx6272, A0=>gen_16_cmp_mReg_3, A1=>
      nx10826, A2=>nx11562);
   ix6309 : nand02 port map ( Y=>gen_16_cmp_BSCmp_op2_4, A0=>nx7762, A1=>
      nx7767);
   ix7763 : nor02_2x port map ( Y=>nx7762, A0=>nx6304, A1=>nx6300);
   ix6305 : nor03_2x port map ( Y=>nx6304, A0=>gen_16_cmp_mReg_3, A1=>
      nx10232, A2=>nx11530);
   ix6301 : nor03_2x port map ( Y=>nx6300, A0=>nx7757, A1=>nx11536, A2=>
      nx11546);
   ix7768 : nor02_2x port map ( Y=>nx7767, A0=>nx6296, A1=>nx6294);
   ix6297 : nor03_2x port map ( Y=>nx6296, A0=>nx7771, A1=>nx10226, A2=>
      nx11554);
   gen_16_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_16_cmp_mReg_4, QB=>
      nx7771, D=>window_16_4, CLK=>start, R=>rst);
   ix6295 : nor03_2x port map ( Y=>nx6294, A0=>gen_16_cmp_mReg_4, A1=>
      nx10826, A2=>nx11562);
   ix6331 : nand02 port map ( Y=>gen_16_cmp_BSCmp_op2_5, A0=>nx7775, A1=>
      nx7781);
   ix7776 : nor02_2x port map ( Y=>nx7775, A0=>nx6326, A1=>nx6322);
   ix6327 : nor03_2x port map ( Y=>nx6326, A0=>gen_16_cmp_mReg_4, A1=>
      nx10232, A2=>nx11530);
   ix6323 : nor03_2x port map ( Y=>nx6322, A0=>nx7771, A1=>nx11536, A2=>
      nx11546);
   ix7782 : nor02_2x port map ( Y=>nx7781, A0=>nx6318, A1=>nx6316);
   ix6319 : nor03_2x port map ( Y=>nx6318, A0=>nx7785, A1=>nx10228, A2=>
      nx11554);
   gen_16_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_16_cmp_mReg_5, QB=>
      nx7785, D=>window_16_5, CLK=>start, R=>rst);
   ix6317 : nor03_2x port map ( Y=>nx6316, A0=>gen_16_cmp_mReg_5, A1=>
      nx10826, A2=>nx11562);
   ix6353 : nand02 port map ( Y=>gen_16_cmp_BSCmp_op2_6, A0=>nx7790, A1=>
      nx7795);
   ix7791 : nor02_2x port map ( Y=>nx7790, A0=>nx6348, A1=>nx6344);
   ix6349 : nor03_2x port map ( Y=>nx6348, A0=>gen_16_cmp_mReg_5, A1=>
      nx10234, A2=>nx11530);
   ix6345 : nor03_2x port map ( Y=>nx6344, A0=>nx7785, A1=>nx11536, A2=>
      nx11546);
   ix7796 : nor02_2x port map ( Y=>nx7795, A0=>nx6340, A1=>nx6338);
   ix6341 : nor03_2x port map ( Y=>nx6340, A0=>nx7799, A1=>nx10228, A2=>
      nx11554);
   gen_16_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_16_cmp_mReg_6, QB=>
      nx7799, D=>window_16_6, CLK=>start, R=>rst);
   ix6339 : nor03_2x port map ( Y=>nx6338, A0=>gen_16_cmp_mReg_6, A1=>
      nx10826, A2=>nx11562);
   ix6375 : nand02 port map ( Y=>gen_16_cmp_BSCmp_op2_7, A0=>nx7805, A1=>
      nx7811);
   ix7806 : nor02_2x port map ( Y=>nx7805, A0=>nx6370, A1=>nx6366);
   ix6371 : nor03_2x port map ( Y=>nx6370, A0=>gen_16_cmp_mReg_6, A1=>
      nx10234, A2=>nx11532);
   ix6367 : nor03_2x port map ( Y=>nx6366, A0=>nx7799, A1=>nx11538, A2=>
      nx11548);
   ix7812 : nor02_2x port map ( Y=>nx7811, A0=>nx6362, A1=>nx6360);
   ix6363 : nor03_2x port map ( Y=>nx6362, A0=>nx7814, A1=>nx10228, A2=>
      nx11556);
   gen_16_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_16_cmp_mReg_7, QB=>
      nx7814, D=>window_16_7, CLK=>start, R=>rst);
   ix6361 : nor03_2x port map ( Y=>nx6360, A0=>gen_16_cmp_mReg_7, A1=>
      nx10826, A2=>nx11564);
   ix6397 : nand02 port map ( Y=>gen_16_cmp_BSCmp_op2_8, A0=>nx7821, A1=>
      nx7827);
   ix7822 : nor02_2x port map ( Y=>nx7821, A0=>nx6392, A1=>nx6388);
   ix6393 : nor03_2x port map ( Y=>nx6392, A0=>gen_16_cmp_mReg_7, A1=>
      nx10234, A2=>nx11532);
   ix6389 : nor03_2x port map ( Y=>nx6388, A0=>nx7814, A1=>nx11538, A2=>
      nx11548);
   ix7828 : nor02_2x port map ( Y=>nx7827, A0=>nx6384, A1=>nx6382);
   ix6385 : nor03_2x port map ( Y=>nx6384, A0=>nx7831, A1=>nx10228, A2=>
      nx11556);
   gen_16_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_16_cmp_mReg_8, QB=>
      nx7831, D=>window_16_8, CLK=>start, R=>rst);
   ix6383 : nor03_2x port map ( Y=>nx6382, A0=>gen_16_cmp_mReg_8, A1=>
      nx10828, A2=>nx11564);
   ix6419 : nand02 port map ( Y=>gen_16_cmp_BSCmp_op2_9, A0=>nx7835, A1=>
      nx7841);
   ix7836 : nor02_2x port map ( Y=>nx7835, A0=>nx6414, A1=>nx6410);
   ix6415 : nor03_2x port map ( Y=>nx6414, A0=>gen_16_cmp_mReg_8, A1=>
      nx10234, A2=>nx11532);
   ix6411 : nor03_2x port map ( Y=>nx6410, A0=>nx7831, A1=>nx11538, A2=>
      nx11548);
   ix7842 : nor02_2x port map ( Y=>nx7841, A0=>nx6406, A1=>nx6404);
   ix6407 : nor03_2x port map ( Y=>nx6406, A0=>nx7845, A1=>nx10228, A2=>
      nx11556);
   gen_16_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_16_cmp_mReg_9, QB=>
      nx7845, D=>window_16_9, CLK=>start, R=>rst);
   ix6405 : nor03_2x port map ( Y=>nx6404, A0=>gen_16_cmp_mReg_9, A1=>
      nx10828, A2=>nx11564);
   ix6441 : nand02 port map ( Y=>gen_16_cmp_BSCmp_op2_10, A0=>nx7849, A1=>
      nx7855);
   ix7850 : nor02_2x port map ( Y=>nx7849, A0=>nx6436, A1=>nx6432);
   ix6437 : nor03_2x port map ( Y=>nx6436, A0=>gen_16_cmp_mReg_9, A1=>
      nx10234, A2=>nx11532);
   ix6433 : nor03_2x port map ( Y=>nx6432, A0=>nx7845, A1=>nx11538, A2=>
      nx11548);
   ix7856 : nor02_2x port map ( Y=>nx7855, A0=>nx6428, A1=>nx6426);
   ix6429 : nor03_2x port map ( Y=>nx6428, A0=>nx7858, A1=>nx10228, A2=>
      nx11556);
   gen_16_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_16_cmp_mReg_10, QB=>
      nx7858, D=>window_16_10, CLK=>start, R=>rst);
   ix6427 : nor03_2x port map ( Y=>nx6426, A0=>gen_16_cmp_mReg_10, A1=>
      nx10828, A2=>nx11564);
   ix6463 : nand02 port map ( Y=>gen_16_cmp_BSCmp_op2_11, A0=>nx7865, A1=>
      nx7871);
   ix7866 : nor02_2x port map ( Y=>nx7865, A0=>nx6458, A1=>nx6454);
   ix6459 : nor03_2x port map ( Y=>nx6458, A0=>gen_16_cmp_mReg_10, A1=>
      nx10234, A2=>nx11532);
   ix6455 : nor03_2x port map ( Y=>nx6454, A0=>nx7858, A1=>nx11538, A2=>
      nx11548);
   ix7872 : nor02_2x port map ( Y=>nx7871, A0=>nx6450, A1=>nx6448);
   ix6451 : nor03_2x port map ( Y=>nx6450, A0=>nx7875, A1=>nx10228, A2=>
      nx11556);
   gen_16_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_16_cmp_mReg_11, QB=>
      nx7875, D=>window_16_11, CLK=>start, R=>rst);
   ix6449 : nor03_2x port map ( Y=>nx6448, A0=>gen_16_cmp_mReg_11, A1=>
      nx10828, A2=>nx11564);
   ix6485 : nand02 port map ( Y=>gen_16_cmp_BSCmp_op2_12, A0=>nx7879, A1=>
      nx7885);
   ix7880 : nor02_2x port map ( Y=>nx7879, A0=>nx6480, A1=>nx6476);
   ix6481 : nor03_2x port map ( Y=>nx6480, A0=>gen_16_cmp_mReg_11, A1=>
      nx10234, A2=>nx11532);
   ix6477 : nor03_2x port map ( Y=>nx6476, A0=>nx7875, A1=>nx11538, A2=>
      nx11548);
   ix7886 : nor02_2x port map ( Y=>nx7885, A0=>nx6472, A1=>nx6470);
   ix6473 : nor03_2x port map ( Y=>nx6472, A0=>nx7889, A1=>nx10230, A2=>
      nx11556);
   gen_16_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_16_cmp_mReg_12, QB=>
      nx7889, D=>window_16_12, CLK=>start, R=>rst);
   ix6471 : nor03_2x port map ( Y=>nx6470, A0=>gen_16_cmp_mReg_12, A1=>
      nx10828, A2=>nx11564);
   ix6507 : nand02 port map ( Y=>gen_16_cmp_BSCmp_op2_13, A0=>nx7893, A1=>
      nx7899);
   ix7894 : nor02_2x port map ( Y=>nx7893, A0=>nx6502, A1=>nx6498);
   ix6503 : nor03_2x port map ( Y=>nx6502, A0=>gen_16_cmp_mReg_12, A1=>
      nx10236, A2=>nx11534);
   ix6499 : nor03_2x port map ( Y=>nx6498, A0=>nx7889, A1=>nx11538, A2=>
      nx11550);
   ix7900 : nor02_2x port map ( Y=>nx7899, A0=>nx6494, A1=>nx6492);
   ix6495 : nor03_2x port map ( Y=>nx6494, A0=>nx7902, A1=>nx10230, A2=>
      nx11558);
   gen_16_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_16_cmp_mReg_13, QB=>
      nx7902, D=>window_16_13, CLK=>start, R=>rst);
   ix6493 : nor03_2x port map ( Y=>nx6492, A0=>gen_16_cmp_mReg_13, A1=>
      nx10828, A2=>nx11566);
   ix6529 : nand02 port map ( Y=>gen_16_cmp_BSCmp_op2_14, A0=>nx7909, A1=>
      nx7915);
   ix7910 : nor02_2x port map ( Y=>nx7909, A0=>nx6524, A1=>nx6520);
   ix6525 : nor03_2x port map ( Y=>nx6524, A0=>gen_16_cmp_mReg_13, A1=>
      nx10236, A2=>nx11534);
   ix6521 : nor03_2x port map ( Y=>nx6520, A0=>nx7902, A1=>nx11540, A2=>
      nx11550);
   ix7916 : nor02_2x port map ( Y=>nx7915, A0=>nx6516, A1=>nx6514);
   ix6517 : nor03_2x port map ( Y=>nx6516, A0=>nx7919, A1=>nx10230, A2=>
      nx11558);
   gen_16_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_16_cmp_mReg_14, QB=>
      nx7919, D=>window_16_14, CLK=>start, R=>rst);
   ix6515 : nor03_2x port map ( Y=>nx6514, A0=>gen_16_cmp_mReg_14, A1=>
      nx10828, A2=>nx11566);
   ix6551 : nand02 port map ( Y=>gen_16_cmp_BSCmp_op2_15, A0=>nx7923, A1=>
      nx7929);
   ix7924 : nor02_2x port map ( Y=>nx7923, A0=>nx6546, A1=>nx6542);
   ix6547 : nor03_2x port map ( Y=>nx6546, A0=>gen_16_cmp_mReg_14, A1=>
      nx10236, A2=>nx11534);
   ix6543 : nor03_2x port map ( Y=>nx6542, A0=>nx7919, A1=>nx11540, A2=>
      nx11550);
   ix7930 : nor02_2x port map ( Y=>nx7929, A0=>nx6538, A1=>nx6536);
   ix6539 : nor03_2x port map ( Y=>nx6538, A0=>nx7933, A1=>nx10230, A2=>
      nx11558);
   gen_16_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_16_cmp_mReg_15, QB=>
      nx7933, D=>window_16_15, CLK=>start, R=>rst);
   ix6537 : nor03_2x port map ( Y=>nx6536, A0=>gen_16_cmp_mReg_15, A1=>
      nx10830, A2=>nx11566);
   ix6561 : nand02 port map ( Y=>gen_16_cmp_BSCmp_op2_16, A0=>nx7937, A1=>
      nx7929);
   ix7938 : nor02_2x port map ( Y=>nx7937, A0=>nx6556, A1=>nx6552);
   ix6557 : nor03_2x port map ( Y=>nx6556, A0=>gen_16_cmp_mReg_15, A1=>
      nx10236, A2=>nx11534);
   ix6553 : nor03_2x port map ( Y=>nx6552, A0=>nx7933, A1=>nx11540, A2=>
      nx11550);
   ix6629 : nand02 port map ( Y=>gen_17_cmp_BSCmp_op2_1, A0=>nx7944, A1=>
      nx7963);
   ix7945 : nor02_2x port map ( Y=>nx7944, A0=>nx6624, A1=>nx6620);
   ix6625 : nor03_2x port map ( Y=>nx6624, A0=>gen_17_cmp_mReg_0, A1=>
      nx10220, A2=>nx11570);
   gen_17_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_17_cmp_mReg_0, QB=>
      nx7949, D=>window_17_0, CLK=>start, R=>rst);
   ix7954 : inv01 port map ( Y=>nx7953, A=>gen_17_cmp_pMux_0);
   ix6621 : nor03_2x port map ( Y=>nx6620, A0=>nx7949, A1=>nx11576, A2=>
      nx11586);
   ix7962 : inv02 port map ( Y=>nx7961, A=>gen_17_cmp_pMux_2);
   ix7964 : nor02_2x port map ( Y=>nx7963, A0=>nx6610, A1=>nx6608);
   ix6611 : nor03_2x port map ( Y=>nx6610, A0=>nx7966, A1=>nx10214, A2=>
      nx11594);
   gen_17_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_17_cmp_mReg_1, QB=>
      nx7966, D=>window_17_1, CLK=>start, R=>rst);
   ix6609 : nor03_2x port map ( Y=>nx6608, A0=>gen_17_cmp_mReg_1, A1=>
      nx10832, A2=>nx11602);
   ix6569 : nor03_2x port map ( Y=>nx6568, A0=>nx10220, A1=>nx7961, A2=>
      gen_17_cmp_pMux_0);
   ix6651 : nand02 port map ( Y=>gen_17_cmp_BSCmp_op2_2, A0=>nx7979, A1=>
      nx7985);
   ix7980 : nor02_2x port map ( Y=>nx7979, A0=>nx6646, A1=>nx6642);
   ix6647 : nor03_2x port map ( Y=>nx6646, A0=>gen_17_cmp_mReg_1, A1=>
      nx10220, A2=>nx11570);
   ix6643 : nor03_2x port map ( Y=>nx6642, A0=>nx7966, A1=>nx11576, A2=>
      nx11586);
   ix7986 : nor02_2x port map ( Y=>nx7985, A0=>nx6638, A1=>nx6636);
   ix6639 : nor03_2x port map ( Y=>nx6638, A0=>nx7988, A1=>nx10214, A2=>
      nx11594);
   gen_17_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_17_cmp_mReg_2, QB=>
      nx7988, D=>window_17_2, CLK=>start, R=>rst);
   ix6637 : nor03_2x port map ( Y=>nx6636, A0=>gen_17_cmp_mReg_2, A1=>
      nx10832, A2=>nx11602);
   ix6673 : nand02 port map ( Y=>gen_17_cmp_BSCmp_op2_3, A0=>nx7993, A1=>
      nx7999);
   ix7994 : nor02_2x port map ( Y=>nx7993, A0=>nx6668, A1=>nx6664);
   ix6669 : nor03_2x port map ( Y=>nx6668, A0=>gen_17_cmp_mReg_2, A1=>
      nx10220, A2=>nx11570);
   ix6665 : nor03_2x port map ( Y=>nx6664, A0=>nx7988, A1=>nx11576, A2=>
      nx11586);
   ix8000 : nor02_2x port map ( Y=>nx7999, A0=>nx6660, A1=>nx6658);
   ix6661 : nor03_2x port map ( Y=>nx6660, A0=>nx8003, A1=>nx10214, A2=>
      nx11594);
   gen_17_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_17_cmp_mReg_3, QB=>
      nx8003, D=>window_17_3, CLK=>start, R=>rst);
   ix6659 : nor03_2x port map ( Y=>nx6658, A0=>gen_17_cmp_mReg_3, A1=>
      nx10832, A2=>nx11602);
   ix6695 : nand02 port map ( Y=>gen_17_cmp_BSCmp_op2_4, A0=>nx8009, A1=>
      nx8013);
   ix8010 : nor02_2x port map ( Y=>nx8009, A0=>nx6690, A1=>nx6686);
   ix6691 : nor03_2x port map ( Y=>nx6690, A0=>gen_17_cmp_mReg_3, A1=>
      nx10220, A2=>nx11570);
   ix6687 : nor03_2x port map ( Y=>nx6686, A0=>nx8003, A1=>nx11576, A2=>
      nx11586);
   ix8014 : nor02_2x port map ( Y=>nx8013, A0=>nx6682, A1=>nx6680);
   ix6683 : nor03_2x port map ( Y=>nx6682, A0=>nx8017, A1=>nx10214, A2=>
      nx11594);
   gen_17_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_17_cmp_mReg_4, QB=>
      nx8017, D=>window_17_4, CLK=>start, R=>rst);
   ix6681 : nor03_2x port map ( Y=>nx6680, A0=>gen_17_cmp_mReg_4, A1=>
      nx10832, A2=>nx11602);
   ix6717 : nand02 port map ( Y=>gen_17_cmp_BSCmp_op2_5, A0=>nx8023, A1=>
      nx8029);
   ix8024 : nor02_2x port map ( Y=>nx8023, A0=>nx6712, A1=>nx6708);
   ix6713 : nor03_2x port map ( Y=>nx6712, A0=>gen_17_cmp_mReg_4, A1=>
      nx10220, A2=>nx11570);
   ix6709 : nor03_2x port map ( Y=>nx6708, A0=>nx8017, A1=>nx11576, A2=>
      nx11586);
   ix8030 : nor02_2x port map ( Y=>nx8029, A0=>nx6704, A1=>nx6702);
   ix6705 : nor03_2x port map ( Y=>nx6704, A0=>nx8032, A1=>nx10216, A2=>
      nx11594);
   gen_17_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_17_cmp_mReg_5, QB=>
      nx8032, D=>window_17_5, CLK=>start, R=>rst);
   ix6703 : nor03_2x port map ( Y=>nx6702, A0=>gen_17_cmp_mReg_5, A1=>
      nx10832, A2=>nx11602);
   ix6739 : nand02 port map ( Y=>gen_17_cmp_BSCmp_op2_6, A0=>nx8037, A1=>
      nx8043);
   ix8038 : nor02_2x port map ( Y=>nx8037, A0=>nx6734, A1=>nx6730);
   ix6735 : nor03_2x port map ( Y=>nx6734, A0=>gen_17_cmp_mReg_5, A1=>
      nx10222, A2=>nx11570);
   ix6731 : nor03_2x port map ( Y=>nx6730, A0=>nx8032, A1=>nx11576, A2=>
      nx11586);
   ix8044 : nor02_2x port map ( Y=>nx8043, A0=>nx6726, A1=>nx6724);
   ix6727 : nor03_2x port map ( Y=>nx6726, A0=>nx8047, A1=>nx10216, A2=>
      nx11594);
   gen_17_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_17_cmp_mReg_6, QB=>
      nx8047, D=>window_17_6, CLK=>start, R=>rst);
   ix6725 : nor03_2x port map ( Y=>nx6724, A0=>gen_17_cmp_mReg_6, A1=>
      nx10832, A2=>nx11602);
   ix6761 : nand02 port map ( Y=>gen_17_cmp_BSCmp_op2_7, A0=>nx8053, A1=>
      nx8057);
   ix8054 : nor02_2x port map ( Y=>nx8053, A0=>nx6756, A1=>nx6752);
   ix6757 : nor03_2x port map ( Y=>nx6756, A0=>gen_17_cmp_mReg_6, A1=>
      nx10222, A2=>nx11572);
   ix6753 : nor03_2x port map ( Y=>nx6752, A0=>nx8047, A1=>nx11578, A2=>
      nx11588);
   ix8058 : nor02_2x port map ( Y=>nx8057, A0=>nx6748, A1=>nx6746);
   ix6749 : nor03_2x port map ( Y=>nx6748, A0=>nx8061, A1=>nx10216, A2=>
      nx11596);
   gen_17_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_17_cmp_mReg_7, QB=>
      nx8061, D=>window_17_7, CLK=>start, R=>rst);
   ix6747 : nor03_2x port map ( Y=>nx6746, A0=>gen_17_cmp_mReg_7, A1=>
      nx10832, A2=>nx11604);
   ix6783 : nand02 port map ( Y=>gen_17_cmp_BSCmp_op2_8, A0=>nx8067, A1=>
      nx8073);
   ix8068 : nor02_2x port map ( Y=>nx8067, A0=>nx6778, A1=>nx6774);
   ix6779 : nor03_2x port map ( Y=>nx6778, A0=>gen_17_cmp_mReg_7, A1=>
      nx10222, A2=>nx11572);
   ix6775 : nor03_2x port map ( Y=>nx6774, A0=>nx8061, A1=>nx11578, A2=>
      nx11588);
   ix8074 : nor02_2x port map ( Y=>nx8073, A0=>nx6770, A1=>nx6768);
   ix6771 : nor03_2x port map ( Y=>nx6770, A0=>nx8076, A1=>nx10216, A2=>
      nx11596);
   gen_17_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_17_cmp_mReg_8, QB=>
      nx8076, D=>window_17_8, CLK=>start, R=>rst);
   ix6769 : nor03_2x port map ( Y=>nx6768, A0=>gen_17_cmp_mReg_8, A1=>
      nx10834, A2=>nx11604);
   ix6805 : nand02 port map ( Y=>gen_17_cmp_BSCmp_op2_9, A0=>nx8081, A1=>
      nx8087);
   ix8082 : nor02_2x port map ( Y=>nx8081, A0=>nx6800, A1=>nx6796);
   ix6801 : nor03_2x port map ( Y=>nx6800, A0=>gen_17_cmp_mReg_8, A1=>
      nx10222, A2=>nx11572);
   ix6797 : nor03_2x port map ( Y=>nx6796, A0=>nx8076, A1=>nx11578, A2=>
      nx11588);
   ix8088 : nor02_2x port map ( Y=>nx8087, A0=>nx6792, A1=>nx6790);
   ix6793 : nor03_2x port map ( Y=>nx6792, A0=>nx8091, A1=>nx10216, A2=>
      nx11596);
   gen_17_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_17_cmp_mReg_9, QB=>
      nx8091, D=>window_17_9, CLK=>start, R=>rst);
   ix6791 : nor03_2x port map ( Y=>nx6790, A0=>gen_17_cmp_mReg_9, A1=>
      nx10834, A2=>nx11604);
   ix6827 : nand02 port map ( Y=>gen_17_cmp_BSCmp_op2_10, A0=>nx8097, A1=>
      nx8101);
   ix8098 : nor02_2x port map ( Y=>nx8097, A0=>nx6822, A1=>nx6818);
   ix6823 : nor03_2x port map ( Y=>nx6822, A0=>gen_17_cmp_mReg_9, A1=>
      nx10222, A2=>nx11572);
   ix6819 : nor03_2x port map ( Y=>nx6818, A0=>nx8091, A1=>nx11578, A2=>
      nx11588);
   ix8102 : nor02_2x port map ( Y=>nx8101, A0=>nx6814, A1=>nx6812);
   ix6815 : nor03_2x port map ( Y=>nx6814, A0=>nx8105, A1=>nx10216, A2=>
      nx11596);
   gen_17_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_17_cmp_mReg_10, QB=>
      nx8105, D=>window_17_10, CLK=>start, R=>rst);
   ix6813 : nor03_2x port map ( Y=>nx6812, A0=>gen_17_cmp_mReg_10, A1=>
      nx10834, A2=>nx11604);
   ix6849 : nand02 port map ( Y=>gen_17_cmp_BSCmp_op2_11, A0=>nx8111, A1=>
      nx8116);
   ix8112 : nor02_2x port map ( Y=>nx8111, A0=>nx6844, A1=>nx6840);
   ix6845 : nor03_2x port map ( Y=>nx6844, A0=>gen_17_cmp_mReg_10, A1=>
      nx10222, A2=>nx11572);
   ix6841 : nor03_2x port map ( Y=>nx6840, A0=>nx8105, A1=>nx11578, A2=>
      nx11588);
   ix8117 : nor02_2x port map ( Y=>nx8116, A0=>nx6836, A1=>nx6834);
   ix6837 : nor03_2x port map ( Y=>nx6836, A0=>nx8119, A1=>nx10216, A2=>
      nx11596);
   gen_17_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_17_cmp_mReg_11, QB=>
      nx8119, D=>window_17_11, CLK=>start, R=>rst);
   ix6835 : nor03_2x port map ( Y=>nx6834, A0=>gen_17_cmp_mReg_11, A1=>
      nx10834, A2=>nx11604);
   ix6871 : nand02 port map ( Y=>gen_17_cmp_BSCmp_op2_12, A0=>nx8123, A1=>
      nx8129);
   ix8124 : nor02_2x port map ( Y=>nx8123, A0=>nx6866, A1=>nx6862);
   ix6867 : nor03_2x port map ( Y=>nx6866, A0=>gen_17_cmp_mReg_11, A1=>
      nx10222, A2=>nx11572);
   ix6863 : nor03_2x port map ( Y=>nx6862, A0=>nx8119, A1=>nx11578, A2=>
      nx11588);
   ix8130 : nor02_2x port map ( Y=>nx8129, A0=>nx6858, A1=>nx6856);
   ix6859 : nor03_2x port map ( Y=>nx6858, A0=>nx8133, A1=>nx10218, A2=>
      nx11596);
   gen_17_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_17_cmp_mReg_12, QB=>
      nx8133, D=>window_17_12, CLK=>start, R=>rst);
   ix6857 : nor03_2x port map ( Y=>nx6856, A0=>gen_17_cmp_mReg_12, A1=>
      nx10834, A2=>nx11604);
   ix6893 : nand02 port map ( Y=>gen_17_cmp_BSCmp_op2_13, A0=>nx8139, A1=>
      nx8145);
   ix8140 : nor02_2x port map ( Y=>nx8139, A0=>nx6888, A1=>nx6884);
   ix6889 : nor03_2x port map ( Y=>nx6888, A0=>gen_17_cmp_mReg_12, A1=>
      nx10224, A2=>nx11574);
   ix6885 : nor03_2x port map ( Y=>nx6884, A0=>nx8133, A1=>nx11578, A2=>
      nx11590);
   ix8146 : nor02_2x port map ( Y=>nx8145, A0=>nx6880, A1=>nx6878);
   ix6881 : nor03_2x port map ( Y=>nx6880, A0=>nx8148, A1=>nx10218, A2=>
      nx11598);
   gen_17_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_17_cmp_mReg_13, QB=>
      nx8148, D=>window_17_13, CLK=>start, R=>rst);
   ix6879 : nor03_2x port map ( Y=>nx6878, A0=>gen_17_cmp_mReg_13, A1=>
      nx10834, A2=>nx11606);
   ix6915 : nand02 port map ( Y=>gen_17_cmp_BSCmp_op2_14, A0=>nx8153, A1=>
      nx8159);
   ix8154 : nor02_2x port map ( Y=>nx8153, A0=>nx6910, A1=>nx6906);
   ix6911 : nor03_2x port map ( Y=>nx6910, A0=>gen_17_cmp_mReg_13, A1=>
      nx10224, A2=>nx11574);
   ix6907 : nor03_2x port map ( Y=>nx6906, A0=>nx8148, A1=>nx11580, A2=>
      nx11590);
   ix8160 : nor02_2x port map ( Y=>nx8159, A0=>nx6902, A1=>nx6900);
   ix6903 : nor03_2x port map ( Y=>nx6902, A0=>nx8163, A1=>nx10218, A2=>
      nx11598);
   gen_17_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_17_cmp_mReg_14, QB=>
      nx8163, D=>window_17_14, CLK=>start, R=>rst);
   ix6901 : nor03_2x port map ( Y=>nx6900, A0=>gen_17_cmp_mReg_14, A1=>
      nx10834, A2=>nx11606);
   ix6937 : nand02 port map ( Y=>gen_17_cmp_BSCmp_op2_15, A0=>nx8169, A1=>
      nx8175);
   ix8170 : nor02_2x port map ( Y=>nx8169, A0=>nx6932, A1=>nx6928);
   ix6933 : nor03_2x port map ( Y=>nx6932, A0=>gen_17_cmp_mReg_14, A1=>
      nx10224, A2=>nx11574);
   ix6929 : nor03_2x port map ( Y=>nx6928, A0=>nx8163, A1=>nx11580, A2=>
      nx11590);
   ix8176 : nor02_2x port map ( Y=>nx8175, A0=>nx6924, A1=>nx6922);
   ix6925 : nor03_2x port map ( Y=>nx6924, A0=>nx8178, A1=>nx10218, A2=>
      nx11598);
   gen_17_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_17_cmp_mReg_15, QB=>
      nx8178, D=>window_17_15, CLK=>start, R=>rst);
   ix6923 : nor03_2x port map ( Y=>nx6922, A0=>gen_17_cmp_mReg_15, A1=>
      nx10836, A2=>nx11606);
   ix6947 : nand02 port map ( Y=>gen_17_cmp_BSCmp_op2_16, A0=>nx8185, A1=>
      nx8175);
   ix8186 : nor02_2x port map ( Y=>nx8185, A0=>nx6942, A1=>nx6938);
   ix6943 : nor03_2x port map ( Y=>nx6942, A0=>gen_17_cmp_mReg_15, A1=>
      nx10224, A2=>nx11574);
   ix6939 : nor03_2x port map ( Y=>nx6938, A0=>nx8178, A1=>nx11580, A2=>
      nx11590);
   ix7015 : nand02 port map ( Y=>gen_18_cmp_BSCmp_op2_1, A0=>nx8191, A1=>
      nx8211);
   ix8192 : nor02_2x port map ( Y=>nx8191, A0=>nx7010, A1=>nx7006);
   ix7011 : nor03_2x port map ( Y=>nx7010, A0=>gen_18_cmp_mReg_0, A1=>
      nx10208, A2=>nx11610);
   gen_18_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_18_cmp_mReg_0, QB=>
      nx8197, D=>window_18_0, CLK=>start, R=>rst);
   ix8202 : inv01 port map ( Y=>nx8200, A=>gen_18_cmp_pMux_0);
   ix7007 : nor03_2x port map ( Y=>nx7006, A0=>nx8197, A1=>nx11616, A2=>
      nx11626);
   ix8210 : inv02 port map ( Y=>nx8209, A=>gen_18_cmp_pMux_2);
   ix8212 : nor02_2x port map ( Y=>nx8211, A0=>nx6996, A1=>nx6994);
   ix6997 : nor03_2x port map ( Y=>nx6996, A0=>nx8215, A1=>nx10202, A2=>
      nx11634);
   gen_18_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_18_cmp_mReg_1, QB=>
      nx8215, D=>window_18_1, CLK=>start, R=>rst);
   ix6995 : nor03_2x port map ( Y=>nx6994, A0=>gen_18_cmp_mReg_1, A1=>
      nx10838, A2=>nx11642);
   ix6955 : nor03_2x port map ( Y=>nx6954, A0=>nx10208, A1=>nx8209, A2=>
      gen_18_cmp_pMux_0);
   ix7037 : nand02 port map ( Y=>gen_18_cmp_BSCmp_op2_2, A0=>nx8225, A1=>
      nx8231);
   ix8226 : nor02_2x port map ( Y=>nx8225, A0=>nx7032, A1=>nx7028);
   ix7033 : nor03_2x port map ( Y=>nx7032, A0=>gen_18_cmp_mReg_1, A1=>
      nx10208, A2=>nx11610);
   ix7029 : nor03_2x port map ( Y=>nx7028, A0=>nx8215, A1=>nx11616, A2=>
      nx11626);
   ix8232 : nor02_2x port map ( Y=>nx8231, A0=>nx7024, A1=>nx7022);
   ix7025 : nor03_2x port map ( Y=>nx7024, A0=>nx8235, A1=>nx10202, A2=>
      nx11634);
   gen_18_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_18_cmp_mReg_2, QB=>
      nx8235, D=>window_18_2, CLK=>start, R=>rst);
   ix7023 : nor03_2x port map ( Y=>nx7022, A0=>gen_18_cmp_mReg_2, A1=>
      nx10838, A2=>nx11642);
   ix7059 : nand02 port map ( Y=>gen_18_cmp_BSCmp_op2_3, A0=>nx8241, A1=>
      nx8245);
   ix8242 : nor02_2x port map ( Y=>nx8241, A0=>nx7054, A1=>nx7050);
   ix7055 : nor03_2x port map ( Y=>nx7054, A0=>gen_18_cmp_mReg_2, A1=>
      nx10208, A2=>nx11610);
   ix7051 : nor03_2x port map ( Y=>nx7050, A0=>nx8235, A1=>nx11616, A2=>
      nx11626);
   ix8246 : nor02_2x port map ( Y=>nx8245, A0=>nx7046, A1=>nx7044);
   ix7047 : nor03_2x port map ( Y=>nx7046, A0=>nx8249, A1=>nx10202, A2=>
      nx11634);
   gen_18_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_18_cmp_mReg_3, QB=>
      nx8249, D=>window_18_3, CLK=>start, R=>rst);
   ix7045 : nor03_2x port map ( Y=>nx7044, A0=>gen_18_cmp_mReg_3, A1=>
      nx10838, A2=>nx11642);
   ix7081 : nand02 port map ( Y=>gen_18_cmp_BSCmp_op2_4, A0=>nx8255, A1=>
      nx8261);
   ix8256 : nor02_2x port map ( Y=>nx8255, A0=>nx7076, A1=>nx7072);
   ix7077 : nor03_2x port map ( Y=>nx7076, A0=>gen_18_cmp_mReg_3, A1=>
      nx10208, A2=>nx11610);
   ix7073 : nor03_2x port map ( Y=>nx7072, A0=>nx8249, A1=>nx11616, A2=>
      nx11626);
   ix8262 : nor02_2x port map ( Y=>nx8261, A0=>nx7068, A1=>nx7066);
   ix7069 : nor03_2x port map ( Y=>nx7068, A0=>nx8264, A1=>nx10202, A2=>
      nx11634);
   gen_18_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_18_cmp_mReg_4, QB=>
      nx8264, D=>window_18_4, CLK=>start, R=>rst);
   ix7067 : nor03_2x port map ( Y=>nx7066, A0=>gen_18_cmp_mReg_4, A1=>
      nx10838, A2=>nx11642);
   ix7103 : nand02 port map ( Y=>gen_18_cmp_BSCmp_op2_5, A0=>nx8269, A1=>
      nx8275);
   ix8270 : nor02_2x port map ( Y=>nx8269, A0=>nx7098, A1=>nx7094);
   ix7099 : nor03_2x port map ( Y=>nx7098, A0=>gen_18_cmp_mReg_4, A1=>
      nx10208, A2=>nx11610);
   ix7095 : nor03_2x port map ( Y=>nx7094, A0=>nx8264, A1=>nx11616, A2=>
      nx11626);
   ix8276 : nor02_2x port map ( Y=>nx8275, A0=>nx7090, A1=>nx7088);
   ix7091 : nor03_2x port map ( Y=>nx7090, A0=>nx8279, A1=>nx10204, A2=>
      nx11634);
   gen_18_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_18_cmp_mReg_5, QB=>
      nx8279, D=>window_18_5, CLK=>start, R=>rst);
   ix7089 : nor03_2x port map ( Y=>nx7088, A0=>gen_18_cmp_mReg_5, A1=>
      nx10838, A2=>nx11642);
   ix7125 : nand02 port map ( Y=>gen_18_cmp_BSCmp_op2_6, A0=>nx8285, A1=>
      nx8289);
   ix8286 : nor02_2x port map ( Y=>nx8285, A0=>nx7120, A1=>nx7116);
   ix7121 : nor03_2x port map ( Y=>nx7120, A0=>gen_18_cmp_mReg_5, A1=>
      nx10210, A2=>nx11610);
   ix7117 : nor03_2x port map ( Y=>nx7116, A0=>nx8279, A1=>nx11616, A2=>
      nx11626);
   ix8290 : nor02_2x port map ( Y=>nx8289, A0=>nx7112, A1=>nx7110);
   ix7113 : nor03_2x port map ( Y=>nx7112, A0=>nx8293, A1=>nx10204, A2=>
      nx11634);
   gen_18_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_18_cmp_mReg_6, QB=>
      nx8293, D=>window_18_6, CLK=>start, R=>rst);
   ix7111 : nor03_2x port map ( Y=>nx7110, A0=>gen_18_cmp_mReg_6, A1=>
      nx10838, A2=>nx11642);
   ix7147 : nand02 port map ( Y=>gen_18_cmp_BSCmp_op2_7, A0=>nx8299, A1=>
      nx8305);
   ix8300 : nor02_2x port map ( Y=>nx8299, A0=>nx7142, A1=>nx7138);
   ix7143 : nor03_2x port map ( Y=>nx7142, A0=>gen_18_cmp_mReg_6, A1=>
      nx10210, A2=>nx11612);
   ix7139 : nor03_2x port map ( Y=>nx7138, A0=>nx8293, A1=>nx11618, A2=>
      nx11628);
   ix8306 : nor02_2x port map ( Y=>nx8305, A0=>nx7134, A1=>nx7132);
   ix7135 : nor03_2x port map ( Y=>nx7134, A0=>nx8308, A1=>nx10204, A2=>
      nx11636);
   gen_18_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_18_cmp_mReg_7, QB=>
      nx8308, D=>window_18_7, CLK=>start, R=>rst);
   ix7133 : nor03_2x port map ( Y=>nx7132, A0=>gen_18_cmp_mReg_7, A1=>
      nx10838, A2=>nx11644);
   ix7169 : nand02 port map ( Y=>gen_18_cmp_BSCmp_op2_8, A0=>nx8313, A1=>
      nx8319);
   ix8314 : nor02_2x port map ( Y=>nx8313, A0=>nx7164, A1=>nx7160);
   ix7165 : nor03_2x port map ( Y=>nx7164, A0=>gen_18_cmp_mReg_7, A1=>
      nx10210, A2=>nx11612);
   ix7161 : nor03_2x port map ( Y=>nx7160, A0=>nx8308, A1=>nx11618, A2=>
      nx11628);
   ix8320 : nor02_2x port map ( Y=>nx8319, A0=>nx7156, A1=>nx7154);
   ix7157 : nor03_2x port map ( Y=>nx7156, A0=>nx8323, A1=>nx10204, A2=>
      nx11636);
   gen_18_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_18_cmp_mReg_8, QB=>
      nx8323, D=>window_18_8, CLK=>start, R=>rst);
   ix7155 : nor03_2x port map ( Y=>nx7154, A0=>gen_18_cmp_mReg_8, A1=>
      nx10840, A2=>nx11644);
   ix7191 : nand02 port map ( Y=>gen_18_cmp_BSCmp_op2_9, A0=>nx8329, A1=>
      nx8333);
   ix8330 : nor02_2x port map ( Y=>nx8329, A0=>nx7186, A1=>nx7182);
   ix7187 : nor03_2x port map ( Y=>nx7186, A0=>gen_18_cmp_mReg_8, A1=>
      nx10210, A2=>nx11612);
   ix7183 : nor03_2x port map ( Y=>nx7182, A0=>nx8323, A1=>nx11618, A2=>
      nx11628);
   ix8334 : nor02_2x port map ( Y=>nx8333, A0=>nx7178, A1=>nx7176);
   ix7179 : nor03_2x port map ( Y=>nx7178, A0=>nx8337, A1=>nx10204, A2=>
      nx11636);
   gen_18_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_18_cmp_mReg_9, QB=>
      nx8337, D=>window_18_9, CLK=>start, R=>rst);
   ix7177 : nor03_2x port map ( Y=>nx7176, A0=>gen_18_cmp_mReg_9, A1=>
      nx10840, A2=>nx11644);
   ix7213 : nand02 port map ( Y=>gen_18_cmp_BSCmp_op2_10, A0=>nx8343, A1=>
      nx8349);
   ix8344 : nor02_2x port map ( Y=>nx8343, A0=>nx7208, A1=>nx7204);
   ix7209 : nor03_2x port map ( Y=>nx7208, A0=>gen_18_cmp_mReg_9, A1=>
      nx10210, A2=>nx11612);
   ix7205 : nor03_2x port map ( Y=>nx7204, A0=>nx8337, A1=>nx11618, A2=>
      nx11628);
   ix8350 : nor02_2x port map ( Y=>nx8349, A0=>nx7200, A1=>nx7198);
   ix7201 : nor03_2x port map ( Y=>nx7200, A0=>nx8352, A1=>nx10204, A2=>
      nx11636);
   gen_18_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_18_cmp_mReg_10, QB=>
      nx8352, D=>window_18_10, CLK=>start, R=>rst);
   ix7199 : nor03_2x port map ( Y=>nx7198, A0=>gen_18_cmp_mReg_10, A1=>
      nx10840, A2=>nx11644);
   ix7235 : nand02 port map ( Y=>gen_18_cmp_BSCmp_op2_11, A0=>nx8357, A1=>
      nx8363);
   ix8358 : nor02_2x port map ( Y=>nx8357, A0=>nx7230, A1=>nx7226);
   ix7231 : nor03_2x port map ( Y=>nx7230, A0=>gen_18_cmp_mReg_10, A1=>
      nx10210, A2=>nx11612);
   ix7227 : nor03_2x port map ( Y=>nx7226, A0=>nx8352, A1=>nx11618, A2=>
      nx11628);
   ix8364 : nor02_2x port map ( Y=>nx8363, A0=>nx7222, A1=>nx7220);
   ix7223 : nor03_2x port map ( Y=>nx7222, A0=>nx8367, A1=>nx10204, A2=>
      nx11636);
   gen_18_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_18_cmp_mReg_11, QB=>
      nx8367, D=>window_18_11, CLK=>start, R=>rst);
   ix7221 : nor03_2x port map ( Y=>nx7220, A0=>gen_18_cmp_mReg_11, A1=>
      nx10840, A2=>nx11644);
   ix7257 : nand02 port map ( Y=>gen_18_cmp_BSCmp_op2_12, A0=>nx8373, A1=>
      nx8377);
   ix8374 : nor02_2x port map ( Y=>nx8373, A0=>nx7252, A1=>nx7248);
   ix7253 : nor03_2x port map ( Y=>nx7252, A0=>gen_18_cmp_mReg_11, A1=>
      nx10210, A2=>nx11612);
   ix7249 : nor03_2x port map ( Y=>nx7248, A0=>nx8367, A1=>nx11618, A2=>
      nx11628);
   ix8378 : nor02_2x port map ( Y=>nx8377, A0=>nx7244, A1=>nx7242);
   ix7245 : nor03_2x port map ( Y=>nx7244, A0=>nx8381, A1=>nx10206, A2=>
      nx11636);
   gen_18_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_18_cmp_mReg_12, QB=>
      nx8381, D=>window_18_12, CLK=>start, R=>rst);
   ix7243 : nor03_2x port map ( Y=>nx7242, A0=>gen_18_cmp_mReg_12, A1=>
      nx10840, A2=>nx11644);
   ix7279 : nand02 port map ( Y=>gen_18_cmp_BSCmp_op2_13, A0=>nx8387, A1=>
      nx8393);
   ix8388 : nor02_2x port map ( Y=>nx8387, A0=>nx7274, A1=>nx7270);
   ix7275 : nor03_2x port map ( Y=>nx7274, A0=>gen_18_cmp_mReg_12, A1=>
      nx10212, A2=>nx11614);
   ix7271 : nor03_2x port map ( Y=>nx7270, A0=>nx8381, A1=>nx11618, A2=>
      nx11630);
   ix8394 : nor02_2x port map ( Y=>nx8393, A0=>nx7266, A1=>nx7264);
   ix7267 : nor03_2x port map ( Y=>nx7266, A0=>nx8396, A1=>nx10206, A2=>
      nx11638);
   gen_18_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_18_cmp_mReg_13, QB=>
      nx8396, D=>window_18_13, CLK=>start, R=>rst);
   ix7265 : nor03_2x port map ( Y=>nx7264, A0=>gen_18_cmp_mReg_13, A1=>
      nx10840, A2=>nx11646);
   ix7301 : nand02 port map ( Y=>gen_18_cmp_BSCmp_op2_14, A0=>nx8401, A1=>
      nx8407);
   ix8402 : nor02_2x port map ( Y=>nx8401, A0=>nx7296, A1=>nx7292);
   ix7297 : nor03_2x port map ( Y=>nx7296, A0=>gen_18_cmp_mReg_13, A1=>
      nx10212, A2=>nx11614);
   ix7293 : nor03_2x port map ( Y=>nx7292, A0=>nx8396, A1=>nx11620, A2=>
      nx11630);
   ix8408 : nor02_2x port map ( Y=>nx8407, A0=>nx7288, A1=>nx7286);
   ix7289 : nor03_2x port map ( Y=>nx7288, A0=>nx8411, A1=>nx10206, A2=>
      nx11638);
   gen_18_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_18_cmp_mReg_14, QB=>
      nx8411, D=>window_18_14, CLK=>start, R=>rst);
   ix7287 : nor03_2x port map ( Y=>nx7286, A0=>gen_18_cmp_mReg_14, A1=>
      nx10840, A2=>nx11646);
   ix7323 : nand02 port map ( Y=>gen_18_cmp_BSCmp_op2_15, A0=>nx8417, A1=>
      nx8421);
   ix8418 : nor02_2x port map ( Y=>nx8417, A0=>nx7318, A1=>nx7314);
   ix7319 : nor03_2x port map ( Y=>nx7318, A0=>gen_18_cmp_mReg_14, A1=>
      nx10212, A2=>nx11614);
   ix7315 : nor03_2x port map ( Y=>nx7314, A0=>nx8411, A1=>nx11620, A2=>
      nx11630);
   ix8422 : nor02_2x port map ( Y=>nx8421, A0=>nx7310, A1=>nx7308);
   ix7311 : nor03_2x port map ( Y=>nx7310, A0=>nx8425, A1=>nx10206, A2=>
      nx11638);
   gen_18_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_18_cmp_mReg_15, QB=>
      nx8425, D=>window_18_15, CLK=>start, R=>rst);
   ix7309 : nor03_2x port map ( Y=>nx7308, A0=>gen_18_cmp_mReg_15, A1=>
      nx10842, A2=>nx11646);
   ix7333 : nand02 port map ( Y=>gen_18_cmp_BSCmp_op2_16, A0=>nx8431, A1=>
      nx8421);
   ix8432 : nor02_2x port map ( Y=>nx8431, A0=>nx7328, A1=>nx7324);
   ix7329 : nor03_2x port map ( Y=>nx7328, A0=>gen_18_cmp_mReg_15, A1=>
      nx10212, A2=>nx11614);
   ix7325 : nor03_2x port map ( Y=>nx7324, A0=>nx8425, A1=>nx11620, A2=>
      nx11630);
   ix7401 : nand02 port map ( Y=>gen_19_cmp_BSCmp_op2_1, A0=>nx8439, A1=>
      nx8457);
   ix8440 : nor02_2x port map ( Y=>nx8439, A0=>nx7396, A1=>nx7392);
   ix7397 : nor03_2x port map ( Y=>nx7396, A0=>gen_19_cmp_mReg_0, A1=>
      nx10196, A2=>nx11650);
   gen_19_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_19_cmp_mReg_0, QB=>
      nx8443, D=>window_19_0, CLK=>start, R=>rst);
   ix8448 : inv01 port map ( Y=>nx8447, A=>gen_19_cmp_pMux_0);
   ix7393 : nor03_2x port map ( Y=>nx7392, A0=>nx8443, A1=>nx11656, A2=>
      nx11666);
   ix8456 : inv02 port map ( Y=>nx8455, A=>gen_19_cmp_pMux_2);
   ix8458 : nor02_2x port map ( Y=>nx8457, A0=>nx7382, A1=>nx7380);
   ix7383 : nor03_2x port map ( Y=>nx7382, A0=>nx8461, A1=>nx10190, A2=>
      nx11674);
   gen_19_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_19_cmp_mReg_1, QB=>
      nx8461, D=>window_19_1, CLK=>start, R=>rst);
   ix7381 : nor03_2x port map ( Y=>nx7380, A0=>gen_19_cmp_mReg_1, A1=>
      nx10844, A2=>nx11682);
   ix7341 : nor03_2x port map ( Y=>nx7340, A0=>nx10196, A1=>nx8455, A2=>
      gen_19_cmp_pMux_0);
   ix7423 : nand02 port map ( Y=>gen_19_cmp_BSCmp_op2_2, A0=>nx8473, A1=>
      nx8477);
   ix8474 : nor02_2x port map ( Y=>nx8473, A0=>nx7418, A1=>nx7414);
   ix7419 : nor03_2x port map ( Y=>nx7418, A0=>gen_19_cmp_mReg_1, A1=>
      nx10196, A2=>nx11650);
   ix7415 : nor03_2x port map ( Y=>nx7414, A0=>nx8461, A1=>nx11656, A2=>
      nx11666);
   ix8478 : nor02_2x port map ( Y=>nx8477, A0=>nx7410, A1=>nx7408);
   ix7411 : nor03_2x port map ( Y=>nx7410, A0=>nx8481, A1=>nx10190, A2=>
      nx11674);
   gen_19_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_19_cmp_mReg_2, QB=>
      nx8481, D=>window_19_2, CLK=>start, R=>rst);
   ix7409 : nor03_2x port map ( Y=>nx7408, A0=>gen_19_cmp_mReg_2, A1=>
      nx10844, A2=>nx11682);
   ix7445 : nand02 port map ( Y=>gen_19_cmp_BSCmp_op2_3, A0=>nx8487, A1=>
      nx8493);
   ix8488 : nor02_2x port map ( Y=>nx8487, A0=>nx7440, A1=>nx7436);
   ix7441 : nor03_2x port map ( Y=>nx7440, A0=>gen_19_cmp_mReg_2, A1=>
      nx10196, A2=>nx11650);
   ix7437 : nor03_2x port map ( Y=>nx7436, A0=>nx8481, A1=>nx11656, A2=>
      nx11666);
   ix8494 : nor02_2x port map ( Y=>nx8493, A0=>nx7432, A1=>nx7430);
   ix7433 : nor03_2x port map ( Y=>nx7432, A0=>nx8497, A1=>nx10190, A2=>
      nx11674);
   gen_19_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_19_cmp_mReg_3, QB=>
      nx8497, D=>window_19_3, CLK=>start, R=>rst);
   ix7431 : nor03_2x port map ( Y=>nx7430, A0=>gen_19_cmp_mReg_3, A1=>
      nx10844, A2=>nx11682);
   ix7467 : nand02 port map ( Y=>gen_19_cmp_BSCmp_op2_4, A0=>nx8502, A1=>
      nx8506);
   ix8503 : nor02_2x port map ( Y=>nx8502, A0=>nx7462, A1=>nx7458);
   ix7463 : nor03_2x port map ( Y=>nx7462, A0=>gen_19_cmp_mReg_3, A1=>
      nx10196, A2=>nx11650);
   ix7459 : nor03_2x port map ( Y=>nx7458, A0=>nx8497, A1=>nx11656, A2=>
      nx11666);
   ix8507 : nor02_2x port map ( Y=>nx8506, A0=>nx7454, A1=>nx7452);
   ix7455 : nor03_2x port map ( Y=>nx7454, A0=>nx8509, A1=>nx10190, A2=>
      nx11674);
   gen_19_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_19_cmp_mReg_4, QB=>
      nx8509, D=>window_19_4, CLK=>start, R=>rst);
   ix7453 : nor03_2x port map ( Y=>nx7452, A0=>gen_19_cmp_mReg_4, A1=>
      nx10844, A2=>nx11682);
   ix7489 : nand02 port map ( Y=>gen_19_cmp_BSCmp_op2_5, A0=>nx8515, A1=>
      nx8521);
   ix8516 : nor02_2x port map ( Y=>nx8515, A0=>nx7484, A1=>nx7480);
   ix7485 : nor03_2x port map ( Y=>nx7484, A0=>gen_19_cmp_mReg_4, A1=>
      nx10196, A2=>nx11650);
   ix7481 : nor03_2x port map ( Y=>nx7480, A0=>nx8509, A1=>nx11656, A2=>
      nx11666);
   ix8522 : nor02_2x port map ( Y=>nx8521, A0=>nx7476, A1=>nx7474);
   ix7477 : nor03_2x port map ( Y=>nx7476, A0=>nx8525, A1=>nx10192, A2=>
      nx11674);
   gen_19_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_19_cmp_mReg_5, QB=>
      nx8525, D=>window_19_5, CLK=>start, R=>rst);
   ix7475 : nor03_2x port map ( Y=>nx7474, A0=>gen_19_cmp_mReg_5, A1=>
      nx10844, A2=>nx11682);
   ix7511 : nand02 port map ( Y=>gen_19_cmp_BSCmp_op2_6, A0=>nx8531, A1=>
      nx8535);
   ix8532 : nor02_2x port map ( Y=>nx8531, A0=>nx7506, A1=>nx7502);
   ix7507 : nor03_2x port map ( Y=>nx7506, A0=>gen_19_cmp_mReg_5, A1=>
      nx10198, A2=>nx11650);
   ix7503 : nor03_2x port map ( Y=>nx7502, A0=>nx8525, A1=>nx11656, A2=>
      nx11666);
   ix8536 : nor02_2x port map ( Y=>nx8535, A0=>nx7498, A1=>nx7496);
   ix7499 : nor03_2x port map ( Y=>nx7498, A0=>nx8539, A1=>nx10192, A2=>
      nx11674);
   gen_19_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_19_cmp_mReg_6, QB=>
      nx8539, D=>window_19_6, CLK=>start, R=>rst);
   ix7497 : nor03_2x port map ( Y=>nx7496, A0=>gen_19_cmp_mReg_6, A1=>
      nx10844, A2=>nx11682);
   ix7533 : nand02 port map ( Y=>gen_19_cmp_BSCmp_op2_7, A0=>nx8545, A1=>
      nx8551);
   ix8546 : nor02_2x port map ( Y=>nx8545, A0=>nx7528, A1=>nx7524);
   ix7529 : nor03_2x port map ( Y=>nx7528, A0=>gen_19_cmp_mReg_6, A1=>
      nx10198, A2=>nx11652);
   ix7525 : nor03_2x port map ( Y=>nx7524, A0=>nx8539, A1=>nx11658, A2=>
      nx11668);
   ix8552 : nor02_2x port map ( Y=>nx8551, A0=>nx7520, A1=>nx7518);
   ix7521 : nor03_2x port map ( Y=>nx7520, A0=>nx8555, A1=>nx10192, A2=>
      nx11676);
   gen_19_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_19_cmp_mReg_7, QB=>
      nx8555, D=>window_19_7, CLK=>start, R=>rst);
   ix7519 : nor03_2x port map ( Y=>nx7518, A0=>gen_19_cmp_mReg_7, A1=>
      nx10844, A2=>nx11684);
   ix7555 : nand02 port map ( Y=>gen_19_cmp_BSCmp_op2_8, A0=>nx8561, A1=>
      nx8565);
   ix8562 : nor02_2x port map ( Y=>nx8561, A0=>nx7550, A1=>nx7546);
   ix7551 : nor03_2x port map ( Y=>nx7550, A0=>gen_19_cmp_mReg_7, A1=>
      nx10198, A2=>nx11652);
   ix7547 : nor03_2x port map ( Y=>nx7546, A0=>nx8555, A1=>nx11658, A2=>
      nx11668);
   ix8566 : nor02_2x port map ( Y=>nx8565, A0=>nx7542, A1=>nx7540);
   ix7543 : nor03_2x port map ( Y=>nx7542, A0=>nx8569, A1=>nx10192, A2=>
      nx11676);
   gen_19_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_19_cmp_mReg_8, QB=>
      nx8569, D=>window_19_8, CLK=>start, R=>rst);
   ix7541 : nor03_2x port map ( Y=>nx7540, A0=>gen_19_cmp_mReg_8, A1=>
      nx10846, A2=>nx11684);
   ix7577 : nand02 port map ( Y=>gen_19_cmp_BSCmp_op2_9, A0=>nx8575, A1=>
      nx8581);
   ix8576 : nor02_2x port map ( Y=>nx8575, A0=>nx7572, A1=>nx7568);
   ix7573 : nor03_2x port map ( Y=>nx7572, A0=>gen_19_cmp_mReg_8, A1=>
      nx10198, A2=>nx11652);
   ix7569 : nor03_2x port map ( Y=>nx7568, A0=>nx8569, A1=>nx11658, A2=>
      nx11668);
   ix8582 : nor02_2x port map ( Y=>nx8581, A0=>nx7564, A1=>nx7562);
   ix7565 : nor03_2x port map ( Y=>nx7564, A0=>nx8584, A1=>nx10192, A2=>
      nx11676);
   gen_19_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_19_cmp_mReg_9, QB=>
      nx8584, D=>window_19_9, CLK=>start, R=>rst);
   ix7563 : nor03_2x port map ( Y=>nx7562, A0=>gen_19_cmp_mReg_9, A1=>
      nx10846, A2=>nx11684);
   ix7599 : nand02 port map ( Y=>gen_19_cmp_BSCmp_op2_10, A0=>nx8589, A1=>
      nx8595);
   ix8590 : nor02_2x port map ( Y=>nx8589, A0=>nx7594, A1=>nx7590);
   ix7595 : nor03_2x port map ( Y=>nx7594, A0=>gen_19_cmp_mReg_9, A1=>
      nx10198, A2=>nx11652);
   ix7591 : nor03_2x port map ( Y=>nx7590, A0=>nx8584, A1=>nx11658, A2=>
      nx11668);
   ix8596 : nor02_2x port map ( Y=>nx8595, A0=>nx7586, A1=>nx7584);
   ix7587 : nor03_2x port map ( Y=>nx7586, A0=>nx8599, A1=>nx10192, A2=>
      nx11676);
   gen_19_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_19_cmp_mReg_10, QB=>
      nx8599, D=>window_19_10, CLK=>start, R=>rst);
   ix7585 : nor03_2x port map ( Y=>nx7584, A0=>gen_19_cmp_mReg_10, A1=>
      nx10846, A2=>nx11684);
   ix7621 : nand02 port map ( Y=>gen_19_cmp_BSCmp_op2_11, A0=>nx8605, A1=>
      nx8609);
   ix8606 : nor02_2x port map ( Y=>nx8605, A0=>nx7616, A1=>nx7612);
   ix7617 : nor03_2x port map ( Y=>nx7616, A0=>gen_19_cmp_mReg_10, A1=>
      nx10198, A2=>nx11652);
   ix7613 : nor03_2x port map ( Y=>nx7612, A0=>nx8599, A1=>nx11658, A2=>
      nx11668);
   ix8610 : nor02_2x port map ( Y=>nx8609, A0=>nx7608, A1=>nx7606);
   ix7609 : nor03_2x port map ( Y=>nx7608, A0=>nx8613, A1=>nx10192, A2=>
      nx11676);
   gen_19_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_19_cmp_mReg_11, QB=>
      nx8613, D=>window_19_11, CLK=>start, R=>rst);
   ix7607 : nor03_2x port map ( Y=>nx7606, A0=>gen_19_cmp_mReg_11, A1=>
      nx10846, A2=>nx11684);
   ix7643 : nand02 port map ( Y=>gen_19_cmp_BSCmp_op2_12, A0=>nx8619, A1=>
      nx8625);
   ix8620 : nor02_2x port map ( Y=>nx8619, A0=>nx7638, A1=>nx7634);
   ix7639 : nor03_2x port map ( Y=>nx7638, A0=>gen_19_cmp_mReg_11, A1=>
      nx10198, A2=>nx11652);
   ix7635 : nor03_2x port map ( Y=>nx7634, A0=>nx8613, A1=>nx11658, A2=>
      nx11668);
   ix8626 : nor02_2x port map ( Y=>nx8625, A0=>nx7630, A1=>nx7628);
   ix7631 : nor03_2x port map ( Y=>nx7630, A0=>nx8628, A1=>nx10194, A2=>
      nx11676);
   gen_19_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_19_cmp_mReg_12, QB=>
      nx8628, D=>window_19_12, CLK=>start, R=>rst);
   ix7629 : nor03_2x port map ( Y=>nx7628, A0=>gen_19_cmp_mReg_12, A1=>
      nx10846, A2=>nx11684);
   ix7665 : nand02 port map ( Y=>gen_19_cmp_BSCmp_op2_13, A0=>nx8633, A1=>
      nx8639);
   ix8634 : nor02_2x port map ( Y=>nx8633, A0=>nx7660, A1=>nx7656);
   ix7661 : nor03_2x port map ( Y=>nx7660, A0=>gen_19_cmp_mReg_12, A1=>
      nx10200, A2=>nx11654);
   ix7657 : nor03_2x port map ( Y=>nx7656, A0=>nx8628, A1=>nx11658, A2=>
      nx11670);
   ix8640 : nor02_2x port map ( Y=>nx8639, A0=>nx7652, A1=>nx7650);
   ix7653 : nor03_2x port map ( Y=>nx7652, A0=>nx8643, A1=>nx10194, A2=>
      nx11678);
   gen_19_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_19_cmp_mReg_13, QB=>
      nx8643, D=>window_19_13, CLK=>start, R=>rst);
   ix7651 : nor03_2x port map ( Y=>nx7650, A0=>gen_19_cmp_mReg_13, A1=>
      nx10846, A2=>nx11686);
   ix7687 : nand02 port map ( Y=>gen_19_cmp_BSCmp_op2_14, A0=>nx8649, A1=>
      nx8653);
   ix8650 : nor02_2x port map ( Y=>nx8649, A0=>nx7682, A1=>nx7678);
   ix7683 : nor03_2x port map ( Y=>nx7682, A0=>gen_19_cmp_mReg_13, A1=>
      nx10200, A2=>nx11654);
   ix7679 : nor03_2x port map ( Y=>nx7678, A0=>nx8643, A1=>nx11660, A2=>
      nx11670);
   ix8654 : nor02_2x port map ( Y=>nx8653, A0=>nx7674, A1=>nx7672);
   ix7675 : nor03_2x port map ( Y=>nx7674, A0=>nx8657, A1=>nx10194, A2=>
      nx11678);
   gen_19_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_19_cmp_mReg_14, QB=>
      nx8657, D=>window_19_14, CLK=>start, R=>rst);
   ix7673 : nor03_2x port map ( Y=>nx7672, A0=>gen_19_cmp_mReg_14, A1=>
      nx10846, A2=>nx11686);
   ix7709 : nand02 port map ( Y=>gen_19_cmp_BSCmp_op2_15, A0=>nx8663, A1=>
      nx8669);
   ix8664 : nor02_2x port map ( Y=>nx8663, A0=>nx7704, A1=>nx7700);
   ix7705 : nor03_2x port map ( Y=>nx7704, A0=>gen_19_cmp_mReg_14, A1=>
      nx10200, A2=>nx11654);
   ix7701 : nor03_2x port map ( Y=>nx7700, A0=>nx8657, A1=>nx11660, A2=>
      nx11670);
   ix8670 : nor02_2x port map ( Y=>nx8669, A0=>nx7696, A1=>nx7694);
   ix7697 : nor03_2x port map ( Y=>nx7696, A0=>nx8672, A1=>nx10194, A2=>
      nx11678);
   gen_19_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_19_cmp_mReg_15, QB=>
      nx8672, D=>window_19_15, CLK=>start, R=>rst);
   ix7695 : nor03_2x port map ( Y=>nx7694, A0=>gen_19_cmp_mReg_15, A1=>
      nx10848, A2=>nx11686);
   ix7719 : nand02 port map ( Y=>gen_19_cmp_BSCmp_op2_16, A0=>nx8677, A1=>
      nx8669);
   ix8678 : nor02_2x port map ( Y=>nx8677, A0=>nx7714, A1=>nx7710);
   ix7715 : nor03_2x port map ( Y=>nx7714, A0=>gen_19_cmp_mReg_15, A1=>
      nx10200, A2=>nx11654);
   ix7711 : nor03_2x port map ( Y=>nx7710, A0=>nx8672, A1=>nx11660, A2=>
      nx11670);
   ix7787 : nand02 port map ( Y=>gen_20_cmp_BSCmp_op2_1, A0=>nx8685, A1=>
      nx8703);
   ix8686 : nor02_2x port map ( Y=>nx8685, A0=>nx7782, A1=>nx7778);
   ix7783 : nor03_2x port map ( Y=>nx7782, A0=>gen_20_cmp_mReg_0, A1=>
      nx10184, A2=>nx11690);
   gen_20_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_20_cmp_mReg_0, QB=>
      nx8691, D=>window_20_0, CLK=>start, R=>rst);
   ix8695 : inv01 port map ( Y=>nx8694, A=>gen_20_cmp_pMux_0);
   ix7779 : nor03_2x port map ( Y=>nx7778, A0=>nx8691, A1=>nx11696, A2=>
      nx11706);
   ix8702 : inv02 port map ( Y=>nx8701, A=>gen_20_cmp_pMux_2);
   ix8704 : nor02_2x port map ( Y=>nx8703, A0=>nx7768, A1=>nx7766);
   ix7769 : nor03_2x port map ( Y=>nx7768, A0=>nx8707, A1=>nx10178, A2=>
      nx11714);
   gen_20_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_20_cmp_mReg_1, QB=>
      nx8707, D=>window_20_1, CLK=>start, R=>rst);
   ix7767 : nor03_2x port map ( Y=>nx7766, A0=>gen_20_cmp_mReg_1, A1=>
      nx10850, A2=>nx11722);
   ix7727 : nor03_2x port map ( Y=>nx7726, A0=>nx10184, A1=>nx8701, A2=>
      gen_20_cmp_pMux_0);
   ix7809 : nand02 port map ( Y=>gen_20_cmp_BSCmp_op2_2, A0=>nx8718, A1=>
      nx8725);
   ix8720 : nor02_2x port map ( Y=>nx8718, A0=>nx7804, A1=>nx7800);
   ix7805 : nor03_2x port map ( Y=>nx7804, A0=>gen_20_cmp_mReg_1, A1=>
      nx10184, A2=>nx11690);
   ix7801 : nor03_2x port map ( Y=>nx7800, A0=>nx8707, A1=>nx11696, A2=>
      nx11706);
   ix8726 : nor02_2x port map ( Y=>nx8725, A0=>nx7796, A1=>nx7794);
   ix7797 : nor03_2x port map ( Y=>nx7796, A0=>nx8729, A1=>nx10178, A2=>
      nx11714);
   gen_20_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_20_cmp_mReg_2, QB=>
      nx8729, D=>window_20_2, CLK=>start, R=>rst);
   ix7795 : nor03_2x port map ( Y=>nx7794, A0=>gen_20_cmp_mReg_2, A1=>
      nx10850, A2=>nx11722);
   ix7831 : nand02 port map ( Y=>gen_20_cmp_BSCmp_op2_3, A0=>nx8735, A1=>
      nx8739);
   ix8736 : nor02_2x port map ( Y=>nx8735, A0=>nx7826, A1=>nx7822);
   ix7827 : nor03_2x port map ( Y=>nx7826, A0=>gen_20_cmp_mReg_2, A1=>
      nx10184, A2=>nx11690);
   ix7823 : nor03_2x port map ( Y=>nx7822, A0=>nx8729, A1=>nx11696, A2=>
      nx11706);
   ix8740 : nor02_2x port map ( Y=>nx8739, A0=>nx7818, A1=>nx7816);
   ix7819 : nor03_2x port map ( Y=>nx7818, A0=>nx8743, A1=>nx10178, A2=>
      nx11714);
   gen_20_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_20_cmp_mReg_3, QB=>
      nx8743, D=>window_20_3, CLK=>start, R=>rst);
   ix7817 : nor03_2x port map ( Y=>nx7816, A0=>gen_20_cmp_mReg_3, A1=>
      nx10850, A2=>nx11722);
   ix7853 : nand02 port map ( Y=>gen_20_cmp_BSCmp_op2_4, A0=>nx8749, A1=>
      nx8753);
   ix8750 : nor02_2x port map ( Y=>nx8749, A0=>nx7848, A1=>nx7844);
   ix7849 : nor03_2x port map ( Y=>nx7848, A0=>gen_20_cmp_mReg_3, A1=>
      nx10184, A2=>nx11690);
   ix7845 : nor03_2x port map ( Y=>nx7844, A0=>nx8743, A1=>nx11696, A2=>
      nx11706);
   ix8754 : nor02_2x port map ( Y=>nx8753, A0=>nx7840, A1=>nx7838);
   ix7841 : nor03_2x port map ( Y=>nx7840, A0=>nx8757, A1=>nx10178, A2=>
      nx11714);
   gen_20_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_20_cmp_mReg_4, QB=>
      nx8757, D=>window_20_4, CLK=>start, R=>rst);
   ix7839 : nor03_2x port map ( Y=>nx7838, A0=>gen_20_cmp_mReg_4, A1=>
      nx10850, A2=>nx11722);
   ix7875 : nand02 port map ( Y=>gen_20_cmp_BSCmp_op2_5, A0=>nx8761, A1=>
      nx8767);
   ix8762 : nor02_2x port map ( Y=>nx8761, A0=>nx7870, A1=>nx7866);
   ix7871 : nor03_2x port map ( Y=>nx7870, A0=>gen_20_cmp_mReg_4, A1=>
      nx10184, A2=>nx11690);
   ix7867 : nor03_2x port map ( Y=>nx7866, A0=>nx8757, A1=>nx11696, A2=>
      nx11706);
   ix8768 : nor02_2x port map ( Y=>nx8767, A0=>nx7862, A1=>nx7860);
   ix7863 : nor03_2x port map ( Y=>nx7862, A0=>nx8771, A1=>nx10180, A2=>
      nx11714);
   gen_20_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_20_cmp_mReg_5, QB=>
      nx8771, D=>window_20_5, CLK=>start, R=>rst);
   ix7861 : nor03_2x port map ( Y=>nx7860, A0=>gen_20_cmp_mReg_5, A1=>
      nx10850, A2=>nx11722);
   ix7897 : nand02 port map ( Y=>gen_20_cmp_BSCmp_op2_6, A0=>nx8775, A1=>
      nx8781);
   ix8776 : nor02_2x port map ( Y=>nx8775, A0=>nx7892, A1=>nx7888);
   ix7893 : nor03_2x port map ( Y=>nx7892, A0=>gen_20_cmp_mReg_5, A1=>
      nx10186, A2=>nx11690);
   ix7889 : nor03_2x port map ( Y=>nx7888, A0=>nx8771, A1=>nx11696, A2=>
      nx11706);
   ix8782 : nor02_2x port map ( Y=>nx8781, A0=>nx7884, A1=>nx7882);
   ix7885 : nor03_2x port map ( Y=>nx7884, A0=>nx8784, A1=>nx10180, A2=>
      nx11714);
   gen_20_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_20_cmp_mReg_6, QB=>
      nx8784, D=>window_20_6, CLK=>start, R=>rst);
   ix7883 : nor03_2x port map ( Y=>nx7882, A0=>gen_20_cmp_mReg_6, A1=>
      nx10850, A2=>nx11722);
   ix7919 : nand02 port map ( Y=>gen_20_cmp_BSCmp_op2_7, A0=>nx8791, A1=>
      nx8797);
   ix8792 : nor02_2x port map ( Y=>nx8791, A0=>nx7914, A1=>nx7910);
   ix7915 : nor03_2x port map ( Y=>nx7914, A0=>gen_20_cmp_mReg_6, A1=>
      nx10186, A2=>nx11692);
   ix7911 : nor03_2x port map ( Y=>nx7910, A0=>nx8784, A1=>nx11698, A2=>
      nx11708);
   ix8798 : nor02_2x port map ( Y=>nx8797, A0=>nx7906, A1=>nx7904);
   ix7907 : nor03_2x port map ( Y=>nx7906, A0=>nx8801, A1=>nx10180, A2=>
      nx11716);
   gen_20_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_20_cmp_mReg_7, QB=>
      nx8801, D=>window_20_7, CLK=>start, R=>rst);
   ix7905 : nor03_2x port map ( Y=>nx7904, A0=>gen_20_cmp_mReg_7, A1=>
      nx10850, A2=>nx11724);
   ix7941 : nand02 port map ( Y=>gen_20_cmp_BSCmp_op2_8, A0=>nx8805, A1=>
      nx8811);
   ix8806 : nor02_2x port map ( Y=>nx8805, A0=>nx7936, A1=>nx7932);
   ix7937 : nor03_2x port map ( Y=>nx7936, A0=>gen_20_cmp_mReg_7, A1=>
      nx10186, A2=>nx11692);
   ix7933 : nor03_2x port map ( Y=>nx7932, A0=>nx8801, A1=>nx11698, A2=>
      nx11708);
   ix8812 : nor02_2x port map ( Y=>nx8811, A0=>nx7928, A1=>nx7926);
   ix7929 : nor03_2x port map ( Y=>nx7928, A0=>nx8815, A1=>nx10180, A2=>
      nx11716);
   gen_20_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_20_cmp_mReg_8, QB=>
      nx8815, D=>window_20_8, CLK=>start, R=>rst);
   ix7927 : nor03_2x port map ( Y=>nx7926, A0=>gen_20_cmp_mReg_8, A1=>
      nx10852, A2=>nx11724);
   ix7963 : nand02 port map ( Y=>gen_20_cmp_BSCmp_op2_9, A0=>nx8819, A1=>
      nx8825);
   ix8820 : nor02_2x port map ( Y=>nx8819, A0=>nx7958, A1=>nx7954);
   ix7959 : nor03_2x port map ( Y=>nx7958, A0=>gen_20_cmp_mReg_8, A1=>
      nx10186, A2=>nx11692);
   ix7955 : nor03_2x port map ( Y=>nx7954, A0=>nx8815, A1=>nx11698, A2=>
      nx11708);
   ix8826 : nor02_2x port map ( Y=>nx8825, A0=>nx7950, A1=>nx7948);
   ix7951 : nor03_2x port map ( Y=>nx7950, A0=>nx8828, A1=>nx10180, A2=>
      nx11716);
   gen_20_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_20_cmp_mReg_9, QB=>
      nx8828, D=>window_20_9, CLK=>start, R=>rst);
   ix7949 : nor03_2x port map ( Y=>nx7948, A0=>gen_20_cmp_mReg_9, A1=>
      nx10852, A2=>nx11724);
   ix7985 : nand02 port map ( Y=>gen_20_cmp_BSCmp_op2_10, A0=>nx8835, A1=>
      nx8841);
   ix8836 : nor02_2x port map ( Y=>nx8835, A0=>nx7980, A1=>nx7976);
   ix7981 : nor03_2x port map ( Y=>nx7980, A0=>gen_20_cmp_mReg_9, A1=>
      nx10186, A2=>nx11692);
   ix7977 : nor03_2x port map ( Y=>nx7976, A0=>nx8828, A1=>nx11698, A2=>
      nx11708);
   ix8842 : nor02_2x port map ( Y=>nx8841, A0=>nx7972, A1=>nx7970);
   ix7973 : nor03_2x port map ( Y=>nx7972, A0=>nx8845, A1=>nx10180, A2=>
      nx11716);
   gen_20_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_20_cmp_mReg_10, QB=>
      nx8845, D=>window_20_10, CLK=>start, R=>rst);
   ix7971 : nor03_2x port map ( Y=>nx7970, A0=>gen_20_cmp_mReg_10, A1=>
      nx10852, A2=>nx11724);
   ix8007 : nand02 port map ( Y=>gen_20_cmp_BSCmp_op2_11, A0=>nx8849, A1=>
      nx8855);
   ix8850 : nor02_2x port map ( Y=>nx8849, A0=>nx8002, A1=>nx7998);
   ix8003 : nor03_2x port map ( Y=>nx8002, A0=>gen_20_cmp_mReg_10, A1=>
      nx10186, A2=>nx11692);
   ix7999 : nor03_2x port map ( Y=>nx7998, A0=>nx8845, A1=>nx11698, A2=>
      nx11708);
   ix8856 : nor02_2x port map ( Y=>nx8855, A0=>nx7994, A1=>nx7992);
   ix7995 : nor03_2x port map ( Y=>nx7994, A0=>nx8859, A1=>nx10180, A2=>
      nx11716);
   gen_20_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_20_cmp_mReg_11, QB=>
      nx8859, D=>window_20_11, CLK=>start, R=>rst);
   ix7993 : nor03_2x port map ( Y=>nx7992, A0=>gen_20_cmp_mReg_11, A1=>
      nx10852, A2=>nx11724);
   ix8029 : nand02 port map ( Y=>gen_20_cmp_BSCmp_op2_12, A0=>nx8863, A1=>
      nx8869);
   ix8864 : nor02_2x port map ( Y=>nx8863, A0=>nx8024, A1=>nx8020);
   ix8025 : nor03_2x port map ( Y=>nx8024, A0=>gen_20_cmp_mReg_11, A1=>
      nx10186, A2=>nx11692);
   ix8021 : nor03_2x port map ( Y=>nx8020, A0=>nx8859, A1=>nx11698, A2=>
      nx11708);
   ix8870 : nor02_2x port map ( Y=>nx8869, A0=>nx8016, A1=>nx8014);
   ix8017 : nor03_2x port map ( Y=>nx8016, A0=>nx8873, A1=>nx10182, A2=>
      nx11716);
   gen_20_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_20_cmp_mReg_12, QB=>
      nx8873, D=>window_20_12, CLK=>start, R=>rst);
   ix8015 : nor03_2x port map ( Y=>nx8014, A0=>gen_20_cmp_mReg_12, A1=>
      nx10852, A2=>nx11724);
   ix8051 : nand02 port map ( Y=>gen_20_cmp_BSCmp_op2_13, A0=>nx8879, A1=>
      nx8885);
   ix8880 : nor02_2x port map ( Y=>nx8879, A0=>nx8046, A1=>nx8042);
   ix8047 : nor03_2x port map ( Y=>nx8046, A0=>gen_20_cmp_mReg_12, A1=>
      nx10188, A2=>nx11694);
   ix8043 : nor03_2x port map ( Y=>nx8042, A0=>nx8873, A1=>nx11698, A2=>
      nx11710);
   ix8886 : nor02_2x port map ( Y=>nx8885, A0=>nx8038, A1=>nx8036);
   ix8039 : nor03_2x port map ( Y=>nx8038, A0=>nx8888, A1=>nx10182, A2=>
      nx11718);
   gen_20_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_20_cmp_mReg_13, QB=>
      nx8888, D=>window_20_13, CLK=>start, R=>rst);
   ix8037 : nor03_2x port map ( Y=>nx8036, A0=>gen_20_cmp_mReg_13, A1=>
      nx10852, A2=>nx11726);
   ix8073 : nand02 port map ( Y=>gen_20_cmp_BSCmp_op2_14, A0=>nx8892, A1=>
      nx8897);
   ix8893 : nor02_2x port map ( Y=>nx8892, A0=>nx8068, A1=>nx8064);
   ix8069 : nor03_2x port map ( Y=>nx8068, A0=>gen_20_cmp_mReg_13, A1=>
      nx10188, A2=>nx11694);
   ix8065 : nor03_2x port map ( Y=>nx8064, A0=>nx8888, A1=>nx11700, A2=>
      nx11710);
   ix8898 : nor02_2x port map ( Y=>nx8897, A0=>nx8060, A1=>nx8058);
   ix8061 : nor03_2x port map ( Y=>nx8060, A0=>nx8901, A1=>nx10182, A2=>
      nx11718);
   gen_20_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_20_cmp_mReg_14, QB=>
      nx8901, D=>window_20_14, CLK=>start, R=>rst);
   ix8059 : nor03_2x port map ( Y=>nx8058, A0=>gen_20_cmp_mReg_14, A1=>
      nx10852, A2=>nx11726);
   ix8095 : nand02 port map ( Y=>gen_20_cmp_BSCmp_op2_15, A0=>nx8907, A1=>
      nx8913);
   ix8908 : nor02_2x port map ( Y=>nx8907, A0=>nx8090, A1=>nx8086);
   ix8091 : nor03_2x port map ( Y=>nx8090, A0=>gen_20_cmp_mReg_14, A1=>
      nx10188, A2=>nx11694);
   ix8087 : nor03_2x port map ( Y=>nx8086, A0=>nx8901, A1=>nx11700, A2=>
      nx11710);
   ix8914 : nor02_2x port map ( Y=>nx8913, A0=>nx8082, A1=>nx8080);
   ix8083 : nor03_2x port map ( Y=>nx8082, A0=>nx8917, A1=>nx10182, A2=>
      nx11718);
   gen_20_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_20_cmp_mReg_15, QB=>
      nx8917, D=>window_20_15, CLK=>start, R=>rst);
   ix8081 : nor03_2x port map ( Y=>nx8080, A0=>gen_20_cmp_mReg_15, A1=>
      nx10854, A2=>nx11726);
   ix8105 : nand02 port map ( Y=>gen_20_cmp_BSCmp_op2_16, A0=>nx8921, A1=>
      nx8913);
   ix8922 : nor02_2x port map ( Y=>nx8921, A0=>nx8100, A1=>nx8096);
   ix8101 : nor03_2x port map ( Y=>nx8100, A0=>gen_20_cmp_mReg_15, A1=>
      nx10188, A2=>nx11694);
   ix8097 : nor03_2x port map ( Y=>nx8096, A0=>nx8917, A1=>nx11700, A2=>
      nx11710);
   ix8173 : nand02 port map ( Y=>gen_21_cmp_BSCmp_op2_1, A0=>nx8929, A1=>
      nx8947);
   ix8930 : nor02_2x port map ( Y=>nx8929, A0=>nx8168, A1=>nx8164);
   ix8169 : nor03_2x port map ( Y=>nx8168, A0=>gen_21_cmp_mReg_0, A1=>
      nx10172, A2=>nx11730);
   gen_21_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_21_cmp_mReg_0, QB=>
      nx8933, D=>window_21_0, CLK=>start, R=>rst);
   ix8938 : inv01 port map ( Y=>nx8937, A=>gen_21_cmp_pMux_0);
   ix8165 : nor03_2x port map ( Y=>nx8164, A0=>nx8933, A1=>nx11736, A2=>
      nx11746);
   ix8946 : inv02 port map ( Y=>nx8945, A=>gen_21_cmp_pMux_2);
   ix8948 : nor02_2x port map ( Y=>nx8947, A0=>nx8154, A1=>nx8152);
   ix8155 : nor03_2x port map ( Y=>nx8154, A0=>nx8950, A1=>nx10166, A2=>
      nx11754);
   gen_21_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_21_cmp_mReg_1, QB=>
      nx8950, D=>window_21_1, CLK=>start, R=>rst);
   ix8153 : nor03_2x port map ( Y=>nx8152, A0=>gen_21_cmp_mReg_1, A1=>
      nx10856, A2=>nx11762);
   ix8113 : nor03_2x port map ( Y=>nx8112, A0=>nx10172, A1=>nx8945, A2=>
      gen_21_cmp_pMux_0);
   ix8195 : nand02 port map ( Y=>gen_21_cmp_BSCmp_op2_2, A0=>nx8963, A1=>
      nx8969);
   ix8964 : nor02_2x port map ( Y=>nx8963, A0=>nx8190, A1=>nx8186);
   ix8191 : nor03_2x port map ( Y=>nx8190, A0=>gen_21_cmp_mReg_1, A1=>
      nx10172, A2=>nx11730);
   ix8187 : nor03_2x port map ( Y=>nx8186, A0=>nx8950, A1=>nx11736, A2=>
      nx11746);
   ix8970 : nor02_2x port map ( Y=>nx8969, A0=>nx8182, A1=>nx8180);
   ix8183 : nor03_2x port map ( Y=>nx8182, A0=>nx8972, A1=>nx10166, A2=>
      nx11754);
   gen_21_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_21_cmp_mReg_2, QB=>
      nx8972, D=>window_21_2, CLK=>start, R=>rst);
   ix8181 : nor03_2x port map ( Y=>nx8180, A0=>gen_21_cmp_mReg_2, A1=>
      nx10856, A2=>nx11762);
   ix8217 : nand02 port map ( Y=>gen_21_cmp_BSCmp_op2_3, A0=>nx8979, A1=>
      nx8985);
   ix8980 : nor02_2x port map ( Y=>nx8979, A0=>nx8212, A1=>nx8208);
   ix8213 : nor03_2x port map ( Y=>nx8212, A0=>gen_21_cmp_mReg_2, A1=>
      nx10172, A2=>nx11730);
   ix8209 : nor03_2x port map ( Y=>nx8208, A0=>nx8972, A1=>nx11736, A2=>
      nx11746);
   ix8986 : nor02_2x port map ( Y=>nx8985, A0=>nx8204, A1=>nx8202);
   ix8205 : nor03_2x port map ( Y=>nx8204, A0=>nx8989, A1=>nx10166, A2=>
      nx11754);
   gen_21_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_21_cmp_mReg_3, QB=>
      nx8989, D=>window_21_3, CLK=>start, R=>rst);
   ix8203 : nor03_2x port map ( Y=>nx8202, A0=>gen_21_cmp_mReg_3, A1=>
      nx10856, A2=>nx11762);
   ix8239 : nand02 port map ( Y=>gen_21_cmp_BSCmp_op2_4, A0=>nx8993, A1=>
      nx8999);
   ix8994 : nor02_2x port map ( Y=>nx8993, A0=>nx8234, A1=>nx8230);
   ix8235 : nor03_2x port map ( Y=>nx8234, A0=>gen_21_cmp_mReg_3, A1=>
      nx10172, A2=>nx11730);
   ix8231 : nor03_2x port map ( Y=>nx8230, A0=>nx8989, A1=>nx11736, A2=>
      nx11746);
   ix9000 : nor02_2x port map ( Y=>nx8999, A0=>nx8226, A1=>nx8224);
   ix8227 : nor03_2x port map ( Y=>nx8226, A0=>nx9003, A1=>nx10166, A2=>
      nx11754);
   gen_21_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_21_cmp_mReg_4, QB=>
      nx9003, D=>window_21_4, CLK=>start, R=>rst);
   ix8225 : nor03_2x port map ( Y=>nx8224, A0=>gen_21_cmp_mReg_4, A1=>
      nx10856, A2=>nx11762);
   ix8261 : nand02 port map ( Y=>gen_21_cmp_BSCmp_op2_5, A0=>nx9007, A1=>
      nx9013);
   ix9008 : nor02_2x port map ( Y=>nx9007, A0=>nx8256, A1=>nx8252);
   ix8257 : nor03_2x port map ( Y=>nx8256, A0=>gen_21_cmp_mReg_4, A1=>
      nx10172, A2=>nx11730);
   ix8253 : nor03_2x port map ( Y=>nx8252, A0=>nx9003, A1=>nx11736, A2=>
      nx11746);
   ix9014 : nor02_2x port map ( Y=>nx9013, A0=>nx8248, A1=>nx8246);
   ix8249 : nor03_2x port map ( Y=>nx8248, A0=>nx9016, A1=>nx10168, A2=>
      nx11754);
   gen_21_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_21_cmp_mReg_5, QB=>
      nx9016, D=>window_21_5, CLK=>start, R=>rst);
   ix8247 : nor03_2x port map ( Y=>nx8246, A0=>gen_21_cmp_mReg_5, A1=>
      nx10856, A2=>nx11762);
   ix8283 : nand02 port map ( Y=>gen_21_cmp_BSCmp_op2_6, A0=>nx9023, A1=>
      nx9029);
   ix9024 : nor02_2x port map ( Y=>nx9023, A0=>nx8278, A1=>nx8274);
   ix8279 : nor03_2x port map ( Y=>nx8278, A0=>gen_21_cmp_mReg_5, A1=>
      nx10174, A2=>nx11730);
   ix8275 : nor03_2x port map ( Y=>nx8274, A0=>nx9016, A1=>nx11736, A2=>
      nx11746);
   ix9030 : nor02_2x port map ( Y=>nx9029, A0=>nx8270, A1=>nx8268);
   ix8271 : nor03_2x port map ( Y=>nx8270, A0=>nx9033, A1=>nx10168, A2=>
      nx11754);
   gen_21_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_21_cmp_mReg_6, QB=>
      nx9033, D=>window_21_6, CLK=>start, R=>rst);
   ix8269 : nor03_2x port map ( Y=>nx8268, A0=>gen_21_cmp_mReg_6, A1=>
      nx10856, A2=>nx11762);
   ix8305 : nand02 port map ( Y=>gen_21_cmp_BSCmp_op2_7, A0=>nx9037, A1=>
      nx9043);
   ix9038 : nor02_2x port map ( Y=>nx9037, A0=>nx8300, A1=>nx8296);
   ix8301 : nor03_2x port map ( Y=>nx8300, A0=>gen_21_cmp_mReg_6, A1=>
      nx10174, A2=>nx11732);
   ix8297 : nor03_2x port map ( Y=>nx8296, A0=>nx9033, A1=>nx11738, A2=>
      nx11748);
   ix9044 : nor02_2x port map ( Y=>nx9043, A0=>nx8292, A1=>nx8290);
   ix8293 : nor03_2x port map ( Y=>nx8292, A0=>nx9047, A1=>nx10168, A2=>
      nx11756);
   gen_21_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_21_cmp_mReg_7, QB=>
      nx9047, D=>window_21_7, CLK=>start, R=>rst);
   ix8291 : nor03_2x port map ( Y=>nx8290, A0=>gen_21_cmp_mReg_7, A1=>
      nx10856, A2=>nx11764);
   ix8327 : nand02 port map ( Y=>gen_21_cmp_BSCmp_op2_8, A0=>nx9051, A1=>
      nx9057);
   ix9052 : nor02_2x port map ( Y=>nx9051, A0=>nx8322, A1=>nx8318);
   ix8323 : nor03_2x port map ( Y=>nx8322, A0=>gen_21_cmp_mReg_7, A1=>
      nx10174, A2=>nx11732);
   ix8319 : nor03_2x port map ( Y=>nx8318, A0=>nx9047, A1=>nx11738, A2=>
      nx11748);
   ix9058 : nor02_2x port map ( Y=>nx9057, A0=>nx8314, A1=>nx8312);
   ix8315 : nor03_2x port map ( Y=>nx8314, A0=>nx9060, A1=>nx10168, A2=>
      nx11756);
   gen_21_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_21_cmp_mReg_8, QB=>
      nx9060, D=>window_21_8, CLK=>start, R=>rst);
   ix8313 : nor03_2x port map ( Y=>nx8312, A0=>gen_21_cmp_mReg_8, A1=>
      nx10858, A2=>nx11764);
   ix8349 : nand02 port map ( Y=>gen_21_cmp_BSCmp_op2_9, A0=>nx9067, A1=>
      nx9073);
   ix9068 : nor02_2x port map ( Y=>nx9067, A0=>nx8344, A1=>nx8340);
   ix8345 : nor03_2x port map ( Y=>nx8344, A0=>gen_21_cmp_mReg_8, A1=>
      nx10174, A2=>nx11732);
   ix8341 : nor03_2x port map ( Y=>nx8340, A0=>nx9060, A1=>nx11738, A2=>
      nx11748);
   ix9074 : nor02_2x port map ( Y=>nx9073, A0=>nx8336, A1=>nx8334);
   ix8337 : nor03_2x port map ( Y=>nx8336, A0=>nx9077, A1=>nx10168, A2=>
      nx11756);
   gen_21_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_21_cmp_mReg_9, QB=>
      nx9077, D=>window_21_9, CLK=>start, R=>rst);
   ix8335 : nor03_2x port map ( Y=>nx8334, A0=>gen_21_cmp_mReg_9, A1=>
      nx10858, A2=>nx11764);
   ix8371 : nand02 port map ( Y=>gen_21_cmp_BSCmp_op2_10, A0=>nx9081, A1=>
      nx9087);
   ix9082 : nor02_2x port map ( Y=>nx9081, A0=>nx8366, A1=>nx8362);
   ix8367 : nor03_2x port map ( Y=>nx8366, A0=>gen_21_cmp_mReg_9, A1=>
      nx10174, A2=>nx11732);
   ix8363 : nor03_2x port map ( Y=>nx8362, A0=>nx9077, A1=>nx11738, A2=>
      nx11748);
   ix9088 : nor02_2x port map ( Y=>nx9087, A0=>nx8358, A1=>nx8356);
   ix8359 : nor03_2x port map ( Y=>nx8358, A0=>nx9091, A1=>nx10168, A2=>
      nx11756);
   gen_21_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_21_cmp_mReg_10, QB=>
      nx9091, D=>window_21_10, CLK=>start, R=>rst);
   ix8357 : nor03_2x port map ( Y=>nx8356, A0=>gen_21_cmp_mReg_10, A1=>
      nx10858, A2=>nx11764);
   ix8393 : nand02 port map ( Y=>gen_21_cmp_BSCmp_op2_11, A0=>nx9095, A1=>
      nx9101);
   ix9096 : nor02_2x port map ( Y=>nx9095, A0=>nx8388, A1=>nx8384);
   ix8389 : nor03_2x port map ( Y=>nx8388, A0=>gen_21_cmp_mReg_10, A1=>
      nx10174, A2=>nx11732);
   ix8385 : nor03_2x port map ( Y=>nx8384, A0=>nx9091, A1=>nx11738, A2=>
      nx11748);
   ix9102 : nor02_2x port map ( Y=>nx9101, A0=>nx8380, A1=>nx8378);
   ix8381 : nor03_2x port map ( Y=>nx8380, A0=>nx9104, A1=>nx10168, A2=>
      nx11756);
   gen_21_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_21_cmp_mReg_11, QB=>
      nx9104, D=>window_21_11, CLK=>start, R=>rst);
   ix8379 : nor03_2x port map ( Y=>nx8378, A0=>gen_21_cmp_mReg_11, A1=>
      nx10858, A2=>nx11764);
   ix8415 : nand02 port map ( Y=>gen_21_cmp_BSCmp_op2_12, A0=>nx9111, A1=>
      nx9117);
   ix9112 : nor02_2x port map ( Y=>nx9111, A0=>nx8410, A1=>nx8406);
   ix8411 : nor03_2x port map ( Y=>nx8410, A0=>gen_21_cmp_mReg_11, A1=>
      nx10174, A2=>nx11732);
   ix8407 : nor03_2x port map ( Y=>nx8406, A0=>nx9104, A1=>nx11738, A2=>
      nx11748);
   ix9118 : nor02_2x port map ( Y=>nx9117, A0=>nx8402, A1=>nx8400);
   ix8403 : nor03_2x port map ( Y=>nx8402, A0=>nx9121, A1=>nx10170, A2=>
      nx11756);
   gen_21_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_21_cmp_mReg_12, QB=>
      nx9121, D=>window_21_12, CLK=>start, R=>rst);
   ix8401 : nor03_2x port map ( Y=>nx8400, A0=>gen_21_cmp_mReg_12, A1=>
      nx10858, A2=>nx11764);
   ix8437 : nand02 port map ( Y=>gen_21_cmp_BSCmp_op2_13, A0=>nx9125, A1=>
      nx9131);
   ix9126 : nor02_2x port map ( Y=>nx9125, A0=>nx8432, A1=>nx8428);
   ix8433 : nor03_2x port map ( Y=>nx8432, A0=>gen_21_cmp_mReg_12, A1=>
      nx10176, A2=>nx11734);
   ix8429 : nor03_2x port map ( Y=>nx8428, A0=>nx9121, A1=>nx11738, A2=>
      nx11750);
   ix9132 : nor02_2x port map ( Y=>nx9131, A0=>nx8424, A1=>nx8422);
   ix8425 : nor03_2x port map ( Y=>nx8424, A0=>nx9135, A1=>nx10170, A2=>
      nx11758);
   gen_21_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_21_cmp_mReg_13, QB=>
      nx9135, D=>window_21_13, CLK=>start, R=>rst);
   ix8423 : nor03_2x port map ( Y=>nx8422, A0=>gen_21_cmp_mReg_13, A1=>
      nx10858, A2=>nx11766);
   ix8459 : nand02 port map ( Y=>gen_21_cmp_BSCmp_op2_14, A0=>nx9139, A1=>
      nx9145);
   ix9140 : nor02_2x port map ( Y=>nx9139, A0=>nx8454, A1=>nx8450);
   ix8455 : nor03_2x port map ( Y=>nx8454, A0=>gen_21_cmp_mReg_13, A1=>
      nx10176, A2=>nx11734);
   ix8451 : nor03_2x port map ( Y=>nx8450, A0=>nx9135, A1=>nx11740, A2=>
      nx11750);
   ix9146 : nor02_2x port map ( Y=>nx9145, A0=>nx8446, A1=>nx8444);
   ix8447 : nor03_2x port map ( Y=>nx8446, A0=>nx9148, A1=>nx10170, A2=>
      nx11758);
   gen_21_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_21_cmp_mReg_14, QB=>
      nx9148, D=>window_21_14, CLK=>start, R=>rst);
   ix8445 : nor03_2x port map ( Y=>nx8444, A0=>gen_21_cmp_mReg_14, A1=>
      nx10858, A2=>nx11766);
   ix8481 : nand02 port map ( Y=>gen_21_cmp_BSCmp_op2_15, A0=>nx9155, A1=>
      nx9161);
   ix9156 : nor02_2x port map ( Y=>nx9155, A0=>nx8476, A1=>nx8472);
   ix8477 : nor03_2x port map ( Y=>nx8476, A0=>gen_21_cmp_mReg_14, A1=>
      nx10176, A2=>nx11734);
   ix8473 : nor03_2x port map ( Y=>nx8472, A0=>nx9148, A1=>nx11740, A2=>
      nx11750);
   ix9162 : nor02_2x port map ( Y=>nx9161, A0=>nx8468, A1=>nx8466);
   ix8469 : nor03_2x port map ( Y=>nx8468, A0=>nx9165, A1=>nx10170, A2=>
      nx11758);
   gen_21_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_21_cmp_mReg_15, QB=>
      nx9165, D=>window_21_15, CLK=>start, R=>rst);
   ix8467 : nor03_2x port map ( Y=>nx8466, A0=>gen_21_cmp_mReg_15, A1=>
      nx10860, A2=>nx11766);
   ix8491 : nand02 port map ( Y=>gen_21_cmp_BSCmp_op2_16, A0=>nx9169, A1=>
      nx9161);
   ix9170 : nor02_2x port map ( Y=>nx9169, A0=>nx8486, A1=>nx8482);
   ix8487 : nor03_2x port map ( Y=>nx8486, A0=>gen_21_cmp_mReg_15, A1=>
      nx10176, A2=>nx11734);
   ix8483 : nor03_2x port map ( Y=>nx8482, A0=>nx9165, A1=>nx11740, A2=>
      nx11750);
   ix8559 : nand02 port map ( Y=>gen_22_cmp_BSCmp_op2_1, A0=>nx9177, A1=>
      nx9197);
   ix9178 : nor02_2x port map ( Y=>nx9177, A0=>nx8554, A1=>nx8550);
   ix8555 : nor03_2x port map ( Y=>nx8554, A0=>gen_22_cmp_mReg_0, A1=>
      nx10160, A2=>nx11770);
   gen_22_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_22_cmp_mReg_0, QB=>
      nx9183, D=>window_22_0, CLK=>start, R=>rst);
   ix9188 : inv01 port map ( Y=>nx9187, A=>gen_22_cmp_pMux_0);
   ix8551 : nor03_2x port map ( Y=>nx8550, A0=>nx9183, A1=>nx11776, A2=>
      nx11786);
   ix9196 : inv02 port map ( Y=>nx9195, A=>gen_22_cmp_pMux_2);
   ix9198 : nor02_2x port map ( Y=>nx9197, A0=>nx8540, A1=>nx8538);
   ix8541 : nor03_2x port map ( Y=>nx8540, A0=>nx9201, A1=>nx10154, A2=>
      nx11794);
   gen_22_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_22_cmp_mReg_1, QB=>
      nx9201, D=>window_22_1, CLK=>start, R=>rst);
   ix8539 : nor03_2x port map ( Y=>nx8538, A0=>gen_22_cmp_mReg_1, A1=>
      nx10862, A2=>nx11802);
   ix8499 : nor03_2x port map ( Y=>nx8498, A0=>nx10160, A1=>nx9195, A2=>
      gen_22_cmp_pMux_0);
   ix8581 : nand02 port map ( Y=>gen_22_cmp_BSCmp_op2_2, A0=>nx9212, A1=>
      nx9217);
   ix9213 : nor02_2x port map ( Y=>nx9212, A0=>nx8576, A1=>nx8572);
   ix8577 : nor03_2x port map ( Y=>nx8576, A0=>gen_22_cmp_mReg_1, A1=>
      nx10160, A2=>nx11770);
   ix8573 : nor03_2x port map ( Y=>nx8572, A0=>nx9201, A1=>nx11776, A2=>
      nx11786);
   ix9218 : nor02_2x port map ( Y=>nx9217, A0=>nx8568, A1=>nx8566);
   ix8569 : nor03_2x port map ( Y=>nx8568, A0=>nx9221, A1=>nx10154, A2=>
      nx11794);
   gen_22_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_22_cmp_mReg_2, QB=>
      nx9221, D=>window_22_2, CLK=>start, R=>rst);
   ix8567 : nor03_2x port map ( Y=>nx8566, A0=>gen_22_cmp_mReg_2, A1=>
      nx10862, A2=>nx11802);
   ix8603 : nand02 port map ( Y=>gen_22_cmp_BSCmp_op2_3, A0=>nx9227, A1=>
      nx9233);
   ix9228 : nor02_2x port map ( Y=>nx9227, A0=>nx8598, A1=>nx8594);
   ix8599 : nor03_2x port map ( Y=>nx8598, A0=>gen_22_cmp_mReg_2, A1=>
      nx10160, A2=>nx11770);
   ix8595 : nor03_2x port map ( Y=>nx8594, A0=>nx9221, A1=>nx11776, A2=>
      nx11786);
   ix9234 : nor02_2x port map ( Y=>nx9233, A0=>nx8590, A1=>nx8588);
   ix8591 : nor03_2x port map ( Y=>nx8590, A0=>nx9236, A1=>nx10154, A2=>
      nx11794);
   gen_22_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_22_cmp_mReg_3, QB=>
      nx9236, D=>window_22_3, CLK=>start, R=>rst);
   ix8589 : nor03_2x port map ( Y=>nx8588, A0=>gen_22_cmp_mReg_3, A1=>
      nx10862, A2=>nx11802);
   ix8625 : nand02 port map ( Y=>gen_22_cmp_BSCmp_op2_4, A0=>nx9243, A1=>
      nx9249);
   ix9244 : nor02_2x port map ( Y=>nx9243, A0=>nx8620, A1=>nx8616);
   ix8621 : nor03_2x port map ( Y=>nx8620, A0=>gen_22_cmp_mReg_3, A1=>
      nx10160, A2=>nx11770);
   ix8617 : nor03_2x port map ( Y=>nx8616, A0=>nx9236, A1=>nx11776, A2=>
      nx11786);
   ix9250 : nor02_2x port map ( Y=>nx9249, A0=>nx8612, A1=>nx8610);
   ix8613 : nor03_2x port map ( Y=>nx8612, A0=>nx9253, A1=>nx10154, A2=>
      nx11794);
   gen_22_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_22_cmp_mReg_4, QB=>
      nx9253, D=>window_22_4, CLK=>start, R=>rst);
   ix8611 : nor03_2x port map ( Y=>nx8610, A0=>gen_22_cmp_mReg_4, A1=>
      nx10862, A2=>nx11802);
   ix8647 : nand02 port map ( Y=>gen_22_cmp_BSCmp_op2_5, A0=>nx9259, A1=>
      nx9265);
   ix9260 : nor02_2x port map ( Y=>nx9259, A0=>nx8642, A1=>nx8638);
   ix8643 : nor03_2x port map ( Y=>nx8642, A0=>gen_22_cmp_mReg_4, A1=>
      nx10160, A2=>nx11770);
   ix8639 : nor03_2x port map ( Y=>nx8638, A0=>nx9253, A1=>nx11776, A2=>
      nx11786);
   ix9266 : nor02_2x port map ( Y=>nx9265, A0=>nx8634, A1=>nx8632);
   ix8635 : nor03_2x port map ( Y=>nx8634, A0=>nx9269, A1=>nx10156, A2=>
      nx11794);
   gen_22_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_22_cmp_mReg_5, QB=>
      nx9269, D=>window_22_5, CLK=>start, R=>rst);
   ix8633 : nor03_2x port map ( Y=>nx8632, A0=>gen_22_cmp_mReg_5, A1=>
      nx10862, A2=>nx11802);
   ix8669 : nand02 port map ( Y=>gen_22_cmp_BSCmp_op2_6, A0=>nx9274, A1=>
      nx9278);
   ix9275 : nor02_2x port map ( Y=>nx9274, A0=>nx8664, A1=>nx8660);
   ix8665 : nor03_2x port map ( Y=>nx8664, A0=>gen_22_cmp_mReg_5, A1=>
      nx10162, A2=>nx11770);
   ix8661 : nor03_2x port map ( Y=>nx8660, A0=>nx9269, A1=>nx11776, A2=>
      nx11786);
   ix9279 : nor02_2x port map ( Y=>nx9278, A0=>nx8656, A1=>nx8654);
   ix8657 : nor03_2x port map ( Y=>nx8656, A0=>nx9281, A1=>nx10156, A2=>
      nx11794);
   gen_22_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_22_cmp_mReg_6, QB=>
      nx9281, D=>window_22_6, CLK=>start, R=>rst);
   ix8655 : nor03_2x port map ( Y=>nx8654, A0=>gen_22_cmp_mReg_6, A1=>
      nx10862, A2=>nx11802);
   ix8691 : nand02 port map ( Y=>gen_22_cmp_BSCmp_op2_7, A0=>nx9287, A1=>
      nx9293);
   ix9288 : nor02_2x port map ( Y=>nx9287, A0=>nx8686, A1=>nx8682);
   ix8687 : nor03_2x port map ( Y=>nx8686, A0=>gen_22_cmp_mReg_6, A1=>
      nx10162, A2=>nx11772);
   ix8683 : nor03_2x port map ( Y=>nx8682, A0=>nx9281, A1=>nx11778, A2=>
      nx11788);
   ix9294 : nor02_2x port map ( Y=>nx9293, A0=>nx8678, A1=>nx8676);
   ix8679 : nor03_2x port map ( Y=>nx8678, A0=>nx9297, A1=>nx10156, A2=>
      nx11796);
   gen_22_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_22_cmp_mReg_7, QB=>
      nx9297, D=>window_22_7, CLK=>start, R=>rst);
   ix8677 : nor03_2x port map ( Y=>nx8676, A0=>gen_22_cmp_mReg_7, A1=>
      nx10862, A2=>nx11804);
   ix8713 : nand02 port map ( Y=>gen_22_cmp_BSCmp_op2_8, A0=>nx9303, A1=>
      nx9307);
   ix9304 : nor02_2x port map ( Y=>nx9303, A0=>nx8708, A1=>nx8704);
   ix8709 : nor03_2x port map ( Y=>nx8708, A0=>gen_22_cmp_mReg_7, A1=>
      nx10162, A2=>nx11772);
   ix8705 : nor03_2x port map ( Y=>nx8704, A0=>nx9297, A1=>nx11778, A2=>
      nx11788);
   ix9308 : nor02_2x port map ( Y=>nx9307, A0=>nx8700, A1=>nx8698);
   ix8701 : nor03_2x port map ( Y=>nx8700, A0=>nx9311, A1=>nx10156, A2=>
      nx11796);
   gen_22_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_22_cmp_mReg_8, QB=>
      nx9311, D=>window_22_8, CLK=>start, R=>rst);
   ix8699 : nor03_2x port map ( Y=>nx8698, A0=>gen_22_cmp_mReg_8, A1=>
      nx10864, A2=>nx11804);
   ix8735 : nand02 port map ( Y=>gen_22_cmp_BSCmp_op2_9, A0=>nx9317, A1=>
      nx9323);
   ix9318 : nor02_2x port map ( Y=>nx9317, A0=>nx8730, A1=>nx8726);
   ix8731 : nor03_2x port map ( Y=>nx8730, A0=>gen_22_cmp_mReg_8, A1=>
      nx10162, A2=>nx11772);
   ix8727 : nor03_2x port map ( Y=>nx8726, A0=>nx9311, A1=>nx11778, A2=>
      nx11788);
   ix9324 : nor02_2x port map ( Y=>nx9323, A0=>nx8722, A1=>nx8720);
   ix8723 : nor03_2x port map ( Y=>nx8722, A0=>nx9327, A1=>nx10156, A2=>
      nx11796);
   gen_22_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_22_cmp_mReg_9, QB=>
      nx9327, D=>window_22_9, CLK=>start, R=>rst);
   ix8721 : nor03_2x port map ( Y=>nx8720, A0=>gen_22_cmp_mReg_9, A1=>
      nx10864, A2=>nx11804);
   ix8757 : nand02 port map ( Y=>gen_22_cmp_BSCmp_op2_10, A0=>nx9333, A1=>
      nx9337);
   ix9334 : nor02_2x port map ( Y=>nx9333, A0=>nx8752, A1=>nx8748);
   ix8753 : nor03_2x port map ( Y=>nx8752, A0=>gen_22_cmp_mReg_9, A1=>
      nx10162, A2=>nx11772);
   ix8749 : nor03_2x port map ( Y=>nx8748, A0=>nx9327, A1=>nx11778, A2=>
      nx11788);
   ix9338 : nor02_2x port map ( Y=>nx9337, A0=>nx8744, A1=>nx8742);
   ix8745 : nor03_2x port map ( Y=>nx8744, A0=>nx9341, A1=>nx10156, A2=>
      nx11796);
   gen_22_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_22_cmp_mReg_10, QB=>
      nx9341, D=>window_22_10, CLK=>start, R=>rst);
   ix8743 : nor03_2x port map ( Y=>nx8742, A0=>gen_22_cmp_mReg_10, A1=>
      nx10864, A2=>nx11804);
   ix8779 : nand02 port map ( Y=>gen_22_cmp_BSCmp_op2_11, A0=>nx9347, A1=>
      nx9353);
   ix9348 : nor02_2x port map ( Y=>nx9347, A0=>nx8774, A1=>nx8770);
   ix8775 : nor03_2x port map ( Y=>nx8774, A0=>gen_22_cmp_mReg_10, A1=>
      nx10162, A2=>nx11772);
   ix8771 : nor03_2x port map ( Y=>nx8770, A0=>nx9341, A1=>nx11778, A2=>
      nx11788);
   ix9354 : nor02_2x port map ( Y=>nx9353, A0=>nx8766, A1=>nx8764);
   ix8767 : nor03_2x port map ( Y=>nx8766, A0=>nx9356, A1=>nx10156, A2=>
      nx11796);
   gen_22_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_22_cmp_mReg_11, QB=>
      nx9356, D=>window_22_11, CLK=>start, R=>rst);
   ix8765 : nor03_2x port map ( Y=>nx8764, A0=>gen_22_cmp_mReg_11, A1=>
      nx10864, A2=>nx11804);
   ix8801 : nand02 port map ( Y=>gen_22_cmp_BSCmp_op2_12, A0=>nx9361, A1=>
      nx9367);
   ix9362 : nor02_2x port map ( Y=>nx9361, A0=>nx8796, A1=>nx8792);
   ix8797 : nor03_2x port map ( Y=>nx8796, A0=>gen_22_cmp_mReg_11, A1=>
      nx10162, A2=>nx11772);
   ix8793 : nor03_2x port map ( Y=>nx8792, A0=>nx9356, A1=>nx11778, A2=>
      nx11788);
   ix9368 : nor02_2x port map ( Y=>nx9367, A0=>nx8788, A1=>nx8786);
   ix8789 : nor03_2x port map ( Y=>nx8788, A0=>nx9371, A1=>nx10158, A2=>
      nx11796);
   gen_22_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_22_cmp_mReg_12, QB=>
      nx9371, D=>window_22_12, CLK=>start, R=>rst);
   ix8787 : nor03_2x port map ( Y=>nx8786, A0=>gen_22_cmp_mReg_12, A1=>
      nx10864, A2=>nx11804);
   ix8823 : nand02 port map ( Y=>gen_22_cmp_BSCmp_op2_13, A0=>nx9377, A1=>
      nx9381);
   ix9378 : nor02_2x port map ( Y=>nx9377, A0=>nx8818, A1=>nx8814);
   ix8819 : nor03_2x port map ( Y=>nx8818, A0=>gen_22_cmp_mReg_12, A1=>
      nx10164, A2=>nx11774);
   ix8815 : nor03_2x port map ( Y=>nx8814, A0=>nx9371, A1=>nx11778, A2=>
      nx11790);
   ix9382 : nor02_2x port map ( Y=>nx9381, A0=>nx8810, A1=>nx8808);
   ix8811 : nor03_2x port map ( Y=>nx8810, A0=>nx9385, A1=>nx10158, A2=>
      nx11798);
   gen_22_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_22_cmp_mReg_13, QB=>
      nx9385, D=>window_22_13, CLK=>start, R=>rst);
   ix8809 : nor03_2x port map ( Y=>nx8808, A0=>gen_22_cmp_mReg_13, A1=>
      nx10864, A2=>nx11806);
   ix8845 : nand02 port map ( Y=>gen_22_cmp_BSCmp_op2_14, A0=>nx9391, A1=>
      nx9397);
   ix9392 : nor02_2x port map ( Y=>nx9391, A0=>nx8840, A1=>nx8836);
   ix8841 : nor03_2x port map ( Y=>nx8840, A0=>gen_22_cmp_mReg_13, A1=>
      nx10164, A2=>nx11774);
   ix8837 : nor03_2x port map ( Y=>nx8836, A0=>nx9385, A1=>nx11780, A2=>
      nx11790);
   ix9398 : nor02_2x port map ( Y=>nx9397, A0=>nx8832, A1=>nx8830);
   ix8833 : nor03_2x port map ( Y=>nx8832, A0=>nx9400, A1=>nx10158, A2=>
      nx11798);
   gen_22_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_22_cmp_mReg_14, QB=>
      nx9400, D=>window_22_14, CLK=>start, R=>rst);
   ix8831 : nor03_2x port map ( Y=>nx8830, A0=>gen_22_cmp_mReg_14, A1=>
      nx10864, A2=>nx11806);
   ix8867 : nand02 port map ( Y=>gen_22_cmp_BSCmp_op2_15, A0=>nx9405, A1=>
      nx9411);
   ix9406 : nor02_2x port map ( Y=>nx9405, A0=>nx8862, A1=>nx8858);
   ix8863 : nor03_2x port map ( Y=>nx8862, A0=>gen_22_cmp_mReg_14, A1=>
      nx10164, A2=>nx11774);
   ix8859 : nor03_2x port map ( Y=>nx8858, A0=>nx9400, A1=>nx11780, A2=>
      nx11790);
   ix9412 : nor02_2x port map ( Y=>nx9411, A0=>nx8854, A1=>nx8852);
   ix8855 : nor03_2x port map ( Y=>nx8854, A0=>nx9415, A1=>nx10158, A2=>
      nx11798);
   gen_22_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_22_cmp_mReg_15, QB=>
      nx9415, D=>window_22_15, CLK=>start, R=>rst);
   ix8853 : nor03_2x port map ( Y=>nx8852, A0=>gen_22_cmp_mReg_15, A1=>
      nx10866, A2=>nx11806);
   ix8877 : nand02 port map ( Y=>gen_22_cmp_BSCmp_op2_16, A0=>nx9421, A1=>
      nx9411);
   ix9422 : nor02_2x port map ( Y=>nx9421, A0=>nx8872, A1=>nx8868);
   ix8873 : nor03_2x port map ( Y=>nx8872, A0=>gen_22_cmp_mReg_15, A1=>
      nx10164, A2=>nx11774);
   ix8869 : nor03_2x port map ( Y=>nx8868, A0=>nx9415, A1=>nx11780, A2=>
      nx11790);
   ix8945 : nand02 port map ( Y=>gen_23_cmp_BSCmp_op2_1, A0=>nx9427, A1=>
      nx9447);
   ix9428 : nor02_2x port map ( Y=>nx9427, A0=>nx8940, A1=>nx8936);
   ix8941 : nor03_2x port map ( Y=>nx8940, A0=>gen_23_cmp_mReg_0, A1=>
      nx10148, A2=>nx11810);
   gen_23_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_23_cmp_mReg_0, QB=>
      nx9433, D=>window_23_0, CLK=>start, R=>rst);
   ix9438 : inv01 port map ( Y=>nx9437, A=>gen_23_cmp_pMux_0);
   ix8937 : nor03_2x port map ( Y=>nx8936, A0=>nx9433, A1=>nx11816, A2=>
      nx11826);
   ix9446 : inv02 port map ( Y=>nx9445, A=>gen_23_cmp_pMux_2);
   ix9448 : nor02_2x port map ( Y=>nx9447, A0=>nx8926, A1=>nx8924);
   ix8927 : nor03_2x port map ( Y=>nx8926, A0=>nx9451, A1=>nx10142, A2=>
      nx11834);
   gen_23_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_23_cmp_mReg_1, QB=>
      nx9451, D=>window_23_1, CLK=>start, R=>rst);
   ix8925 : nor03_2x port map ( Y=>nx8924, A0=>gen_23_cmp_mReg_1, A1=>
      nx10868, A2=>nx11842);
   ix8885 : nor03_2x port map ( Y=>nx8884, A0=>nx10148, A1=>nx9445, A2=>
      gen_23_cmp_pMux_0);
   ix8967 : nand02 port map ( Y=>gen_23_cmp_BSCmp_op2_2, A0=>nx9463, A1=>
      nx9467);
   ix9464 : nor02_2x port map ( Y=>nx9463, A0=>nx8962, A1=>nx8958);
   ix8963 : nor03_2x port map ( Y=>nx8962, A0=>gen_23_cmp_mReg_1, A1=>
      nx10148, A2=>nx11810);
   ix8959 : nor03_2x port map ( Y=>nx8958, A0=>nx9451, A1=>nx11816, A2=>
      nx11826);
   ix9468 : nor02_2x port map ( Y=>nx9467, A0=>nx8954, A1=>nx8952);
   ix8955 : nor03_2x port map ( Y=>nx8954, A0=>nx9471, A1=>nx10142, A2=>
      nx11834);
   gen_23_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_23_cmp_mReg_2, QB=>
      nx9471, D=>window_23_2, CLK=>start, R=>rst);
   ix8953 : nor03_2x port map ( Y=>nx8952, A0=>gen_23_cmp_mReg_2, A1=>
      nx10868, A2=>nx11842);
   ix8989 : nand02 port map ( Y=>gen_23_cmp_BSCmp_op2_3, A0=>nx9477, A1=>
      nx9481);
   ix9478 : nor02_2x port map ( Y=>nx9477, A0=>nx8984, A1=>nx8980);
   ix8985 : nor03_2x port map ( Y=>nx8984, A0=>gen_23_cmp_mReg_2, A1=>
      nx10148, A2=>nx11810);
   ix8981 : nor03_2x port map ( Y=>nx8980, A0=>nx9471, A1=>nx11816, A2=>
      nx11826);
   ix9482 : nor02_2x port map ( Y=>nx9481, A0=>nx8976, A1=>nx8974);
   ix8977 : nor03_2x port map ( Y=>nx8976, A0=>nx9485, A1=>nx10142, A2=>
      nx11834);
   gen_23_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_23_cmp_mReg_3, QB=>
      nx9485, D=>window_23_3, CLK=>start, R=>rst);
   ix8975 : nor03_2x port map ( Y=>nx8974, A0=>gen_23_cmp_mReg_3, A1=>
      nx10868, A2=>nx11842);
   ix9011 : nand02 port map ( Y=>gen_23_cmp_BSCmp_op2_4, A0=>nx9489, A1=>
      nx9495);
   ix9490 : nor02_2x port map ( Y=>nx9489, A0=>nx9006, A1=>nx9002);
   ix9007 : nor03_2x port map ( Y=>nx9006, A0=>gen_23_cmp_mReg_3, A1=>
      nx10148, A2=>nx11810);
   ix9003 : nor03_2x port map ( Y=>nx9002, A0=>nx9485, A1=>nx11816, A2=>
      nx11826);
   ix9496 : nor02_2x port map ( Y=>nx9495, A0=>nx8998, A1=>nx8996);
   ix8999 : nor03_2x port map ( Y=>nx8998, A0=>nx9499, A1=>nx10142, A2=>
      nx11834);
   gen_23_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_23_cmp_mReg_4, QB=>
      nx9499, D=>window_23_4, CLK=>start, R=>rst);
   ix8997 : nor03_2x port map ( Y=>nx8996, A0=>gen_23_cmp_mReg_4, A1=>
      nx10868, A2=>nx11842);
   ix9033 : nand02 port map ( Y=>gen_23_cmp_BSCmp_op2_5, A0=>nx9503, A1=>
      nx9509);
   ix9504 : nor02_2x port map ( Y=>nx9503, A0=>nx9028, A1=>nx9024);
   ix9029 : nor03_2x port map ( Y=>nx9028, A0=>gen_23_cmp_mReg_4, A1=>
      nx10148, A2=>nx11810);
   ix9025 : nor03_2x port map ( Y=>nx9024, A0=>nx9499, A1=>nx11816, A2=>
      nx11826);
   ix9510 : nor02_2x port map ( Y=>nx9509, A0=>nx9020, A1=>nx9018);
   ix9021 : nor03_2x port map ( Y=>nx9020, A0=>nx9512, A1=>nx10144, A2=>
      nx11834);
   gen_23_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_23_cmp_mReg_5, QB=>
      nx9512, D=>window_23_5, CLK=>start, R=>rst);
   ix9019 : nor03_2x port map ( Y=>nx9018, A0=>gen_23_cmp_mReg_5, A1=>
      nx10868, A2=>nx11842);
   ix9055 : nand02 port map ( Y=>gen_23_cmp_BSCmp_op2_6, A0=>nx9519, A1=>
      nx9525);
   ix9520 : nor02_2x port map ( Y=>nx9519, A0=>nx9050, A1=>nx9046);
   ix9051 : nor03_2x port map ( Y=>nx9050, A0=>gen_23_cmp_mReg_5, A1=>
      nx10150, A2=>nx11810);
   ix9047 : nor03_2x port map ( Y=>nx9046, A0=>nx9512, A1=>nx11816, A2=>
      nx11826);
   ix9526 : nor02_2x port map ( Y=>nx9525, A0=>nx9042, A1=>nx9040);
   ix9043 : nor03_2x port map ( Y=>nx9042, A0=>nx9529, A1=>nx10144, A2=>
      nx11834);
   gen_23_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_23_cmp_mReg_6, QB=>
      nx9529, D=>window_23_6, CLK=>start, R=>rst);
   ix9041 : nor03_2x port map ( Y=>nx9040, A0=>gen_23_cmp_mReg_6, A1=>
      nx10868, A2=>nx11842);
   ix9077 : nand02 port map ( Y=>gen_23_cmp_BSCmp_op2_7, A0=>nx9533, A1=>
      nx9539);
   ix9534 : nor02_2x port map ( Y=>nx9533, A0=>nx9072, A1=>nx9068);
   ix9073 : nor03_2x port map ( Y=>nx9072, A0=>gen_23_cmp_mReg_6, A1=>
      nx10150, A2=>nx11812);
   ix9069 : nor03_2x port map ( Y=>nx9068, A0=>nx9529, A1=>nx11818, A2=>
      nx11828);
   ix9540 : nor02_2x port map ( Y=>nx9539, A0=>nx9064, A1=>nx9062);
   ix9065 : nor03_2x port map ( Y=>nx9064, A0=>nx9543, A1=>nx10144, A2=>
      nx11836);
   gen_23_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_23_cmp_mReg_7, QB=>
      nx9543, D=>window_23_7, CLK=>start, R=>rst);
   ix9063 : nor03_2x port map ( Y=>nx9062, A0=>gen_23_cmp_mReg_7, A1=>
      nx10868, A2=>nx11844);
   ix9099 : nand02 port map ( Y=>gen_23_cmp_BSCmp_op2_8, A0=>nx9547, A1=>
      nx9553);
   ix9548 : nor02_2x port map ( Y=>nx9547, A0=>nx9094, A1=>nx9090);
   ix9095 : nor03_2x port map ( Y=>nx9094, A0=>gen_23_cmp_mReg_7, A1=>
      nx10150, A2=>nx11812);
   ix9091 : nor03_2x port map ( Y=>nx9090, A0=>nx9543, A1=>nx11818, A2=>
      nx11828);
   ix9554 : nor02_2x port map ( Y=>nx9553, A0=>nx9086, A1=>nx9084);
   ix9087 : nor03_2x port map ( Y=>nx9086, A0=>nx9556, A1=>nx10144, A2=>
      nx11836);
   gen_23_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_23_cmp_mReg_8, QB=>
      nx9556, D=>window_23_8, CLK=>start, R=>rst);
   ix9085 : nor03_2x port map ( Y=>nx9084, A0=>gen_23_cmp_mReg_8, A1=>
      nx10870, A2=>nx11844);
   ix9121 : nand02 port map ( Y=>gen_23_cmp_BSCmp_op2_9, A0=>nx9563, A1=>
      nx9569);
   ix9564 : nor02_2x port map ( Y=>nx9563, A0=>nx9116, A1=>nx9112);
   ix9117 : nor03_2x port map ( Y=>nx9116, A0=>gen_23_cmp_mReg_8, A1=>
      nx10150, A2=>nx11812);
   ix9113 : nor03_2x port map ( Y=>nx9112, A0=>nx9556, A1=>nx11818, A2=>
      nx11828);
   ix9570 : nor02_2x port map ( Y=>nx9569, A0=>nx9108, A1=>nx9106);
   ix9109 : nor03_2x port map ( Y=>nx9108, A0=>nx9573, A1=>nx10144, A2=>
      nx11836);
   gen_23_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_23_cmp_mReg_9, QB=>
      nx9573, D=>window_23_9, CLK=>start, R=>rst);
   ix9107 : nor03_2x port map ( Y=>nx9106, A0=>gen_23_cmp_mReg_9, A1=>
      nx10870, A2=>nx11844);
   ix9143 : nand02 port map ( Y=>gen_23_cmp_BSCmp_op2_10, A0=>nx9577, A1=>
      nx9583);
   ix9578 : nor02_2x port map ( Y=>nx9577, A0=>nx9138, A1=>nx9134);
   ix9139 : nor03_2x port map ( Y=>nx9138, A0=>gen_23_cmp_mReg_9, A1=>
      nx10150, A2=>nx11812);
   ix9135 : nor03_2x port map ( Y=>nx9134, A0=>nx9573, A1=>nx11818, A2=>
      nx11828);
   ix9584 : nor02_2x port map ( Y=>nx9583, A0=>nx9130, A1=>nx9128);
   ix9131 : nor03_2x port map ( Y=>nx9130, A0=>nx9587, A1=>nx10144, A2=>
      nx11836);
   gen_23_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_23_cmp_mReg_10, QB=>
      nx9587, D=>window_23_10, CLK=>start, R=>rst);
   ix9129 : nor03_2x port map ( Y=>nx9128, A0=>gen_23_cmp_mReg_10, A1=>
      nx10870, A2=>nx11844);
   ix9165 : nand02 port map ( Y=>gen_23_cmp_BSCmp_op2_11, A0=>nx9591, A1=>
      nx9597);
   ix9592 : nor02_2x port map ( Y=>nx9591, A0=>nx9160, A1=>nx9156);
   ix9161 : nor03_2x port map ( Y=>nx9160, A0=>gen_23_cmp_mReg_10, A1=>
      nx10150, A2=>nx11812);
   ix9157 : nor03_2x port map ( Y=>nx9156, A0=>nx9587, A1=>nx11818, A2=>
      nx11828);
   ix9598 : nor02_2x port map ( Y=>nx9597, A0=>nx9152, A1=>nx9150);
   ix9153 : nor03_2x port map ( Y=>nx9152, A0=>nx9600, A1=>nx10144, A2=>
      nx11836);
   gen_23_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_23_cmp_mReg_11, QB=>
      nx9600, D=>window_23_11, CLK=>start, R=>rst);
   ix9151 : nor03_2x port map ( Y=>nx9150, A0=>gen_23_cmp_mReg_11, A1=>
      nx10870, A2=>nx11844);
   ix9187 : nand02 port map ( Y=>gen_23_cmp_BSCmp_op2_12, A0=>nx9607, A1=>
      nx9613);
   ix9608 : nor02_2x port map ( Y=>nx9607, A0=>nx9182, A1=>nx9178);
   ix9183 : nor03_2x port map ( Y=>nx9182, A0=>gen_23_cmp_mReg_11, A1=>
      nx10150, A2=>nx11812);
   ix9179 : nor03_2x port map ( Y=>nx9178, A0=>nx9600, A1=>nx11818, A2=>
      nx11828);
   ix9614 : nor02_2x port map ( Y=>nx9613, A0=>nx9174, A1=>nx9172);
   ix9175 : nor03_2x port map ( Y=>nx9174, A0=>nx9617, A1=>nx10146, A2=>
      nx11836);
   gen_23_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_23_cmp_mReg_12, QB=>
      nx9617, D=>window_23_12, CLK=>start, R=>rst);
   ix9173 : nor03_2x port map ( Y=>nx9172, A0=>gen_23_cmp_mReg_12, A1=>
      nx10870, A2=>nx11844);
   ix9209 : nand02 port map ( Y=>gen_23_cmp_BSCmp_op2_13, A0=>nx9621, A1=>
      nx9627);
   ix9622 : nor02_2x port map ( Y=>nx9621, A0=>nx9204, A1=>nx9200);
   ix9205 : nor03_2x port map ( Y=>nx9204, A0=>gen_23_cmp_mReg_12, A1=>
      nx10152, A2=>nx11814);
   ix9201 : nor03_2x port map ( Y=>nx9200, A0=>nx9617, A1=>nx11818, A2=>
      nx11830);
   ix9628 : nor02_2x port map ( Y=>nx9627, A0=>nx9196, A1=>nx9194);
   ix9197 : nor03_2x port map ( Y=>nx9196, A0=>nx9631, A1=>nx10146, A2=>
      nx11838);
   gen_23_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_23_cmp_mReg_13, QB=>
      nx9631, D=>window_23_13, CLK=>start, R=>rst);
   ix9195 : nor03_2x port map ( Y=>nx9194, A0=>gen_23_cmp_mReg_13, A1=>
      nx10870, A2=>nx11846);
   ix9231 : nand02 port map ( Y=>gen_23_cmp_BSCmp_op2_14, A0=>nx9635, A1=>
      nx9641);
   ix9636 : nor02_2x port map ( Y=>nx9635, A0=>nx9226, A1=>nx9222);
   ix9227 : nor03_2x port map ( Y=>nx9226, A0=>gen_23_cmp_mReg_13, A1=>
      nx10152, A2=>nx11814);
   ix9223 : nor03_2x port map ( Y=>nx9222, A0=>nx9631, A1=>nx11820, A2=>
      nx11830);
   ix9642 : nor02_2x port map ( Y=>nx9641, A0=>nx9218, A1=>nx9216);
   ix9219 : nor03_2x port map ( Y=>nx9218, A0=>nx9645, A1=>nx10146, A2=>
      nx11838);
   gen_23_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_23_cmp_mReg_14, QB=>
      nx9645, D=>window_23_14, CLK=>start, R=>rst);
   ix9217 : nor03_2x port map ( Y=>nx9216, A0=>gen_23_cmp_mReg_14, A1=>
      nx10870, A2=>nx11846);
   ix9253 : nand02 port map ( Y=>gen_23_cmp_BSCmp_op2_15, A0=>nx9651, A1=>
      nx9655);
   ix9652 : nor02_2x port map ( Y=>nx9651, A0=>nx9248, A1=>nx9244);
   ix9249 : nor03_2x port map ( Y=>nx9248, A0=>gen_23_cmp_mReg_14, A1=>
      nx10152, A2=>nx11814);
   ix9245 : nor03_2x port map ( Y=>nx9244, A0=>nx9645, A1=>nx11820, A2=>
      nx11830);
   ix9656 : nor02_2x port map ( Y=>nx9655, A0=>nx9240, A1=>nx9238);
   ix9241 : nor03_2x port map ( Y=>nx9240, A0=>nx9658, A1=>nx10146, A2=>
      nx11838);
   gen_23_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_23_cmp_mReg_15, QB=>
      nx9658, D=>window_23_15, CLK=>start, R=>rst);
   ix9239 : nor03_2x port map ( Y=>nx9238, A0=>gen_23_cmp_mReg_15, A1=>
      nx10872, A2=>nx11846);
   ix9263 : nand02 port map ( Y=>gen_23_cmp_BSCmp_op2_16, A0=>nx9663, A1=>
      nx9655);
   ix9664 : nor02_2x port map ( Y=>nx9663, A0=>nx9258, A1=>nx9254);
   ix9259 : nor03_2x port map ( Y=>nx9258, A0=>gen_23_cmp_mReg_15, A1=>
      nx10152, A2=>nx11814);
   ix9255 : nor03_2x port map ( Y=>nx9254, A0=>nx9658, A1=>nx11820, A2=>
      nx11830);
   ix9331 : nand02 port map ( Y=>gen_24_cmp_BSCmp_op2_1, A0=>nx9669, A1=>
      nx9685);
   ix9670 : nor02_2x port map ( Y=>nx9669, A0=>nx9326, A1=>nx9322);
   ix9327 : nor03_2x port map ( Y=>nx9326, A0=>gen_24_cmp_mReg_0, A1=>
      nx10136, A2=>nx11850);
   gen_24_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_24_cmp_mReg_0, QB=>
      nx9673, D=>window_24_0, CLK=>start, R=>rst);
   ix9677 : inv01 port map ( Y=>nx9676, A=>gen_24_cmp_pMux_0);
   ix9323 : nor03_2x port map ( Y=>nx9322, A0=>nx9673, A1=>nx11856, A2=>
      nx11866);
   ix9684 : inv02 port map ( Y=>nx9683, A=>gen_24_cmp_pMux_2);
   ix9686 : nor02_2x port map ( Y=>nx9685, A0=>nx9312, A1=>nx9310);
   ix9313 : nor03_2x port map ( Y=>nx9312, A0=>nx9688, A1=>nx10130, A2=>
      nx11874);
   gen_24_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_24_cmp_mReg_1, QB=>
      nx9688, D=>window_24_1, CLK=>start, R=>rst);
   ix9311 : nor03_2x port map ( Y=>nx9310, A0=>gen_24_cmp_mReg_1, A1=>
      nx10874, A2=>nx11882);
   ix9271 : nor03_2x port map ( Y=>nx9270, A0=>nx10136, A1=>nx9683, A2=>
      gen_24_cmp_pMux_0);
   ix9353 : nand02 port map ( Y=>gen_24_cmp_BSCmp_op2_2, A0=>nx9698, A1=>
      nx9702);
   ix9699 : nor02_2x port map ( Y=>nx9698, A0=>nx9348, A1=>nx9344);
   ix9349 : nor03_2x port map ( Y=>nx9348, A0=>gen_24_cmp_mReg_1, A1=>
      nx10136, A2=>nx11850);
   ix9345 : nor03_2x port map ( Y=>nx9344, A0=>nx9688, A1=>nx11856, A2=>
      nx11866);
   ix9703 : nor02_2x port map ( Y=>nx9702, A0=>nx9340, A1=>nx9338);
   ix9341 : nor03_2x port map ( Y=>nx9340, A0=>nx9705, A1=>nx10130, A2=>
      nx11874);
   gen_24_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_24_cmp_mReg_2, QB=>
      nx9705, D=>window_24_2, CLK=>start, R=>rst);
   ix9339 : nor03_2x port map ( Y=>nx9338, A0=>gen_24_cmp_mReg_2, A1=>
      nx10874, A2=>nx11882);
   ix9375 : nand02 port map ( Y=>gen_24_cmp_BSCmp_op2_3, A0=>nx9709, A1=>
      nx9713);
   ix9710 : nor02_2x port map ( Y=>nx9709, A0=>nx9370, A1=>nx9366);
   ix9371 : nor03_2x port map ( Y=>nx9370, A0=>gen_24_cmp_mReg_2, A1=>
      nx10136, A2=>nx11850);
   ix9367 : nor03_2x port map ( Y=>nx9366, A0=>nx9705, A1=>nx11856, A2=>
      nx11866);
   ix9714 : nor02_2x port map ( Y=>nx9713, A0=>nx9362, A1=>nx9360);
   ix9363 : nor03_2x port map ( Y=>nx9362, A0=>nx9716, A1=>nx10130, A2=>
      nx11874);
   gen_24_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_24_cmp_mReg_3, QB=>
      nx9716, D=>window_24_3, CLK=>start, R=>rst);
   ix9361 : nor03_2x port map ( Y=>nx9360, A0=>gen_24_cmp_mReg_3, A1=>
      nx10874, A2=>nx11882);
   ix9397 : nand02 port map ( Y=>gen_24_cmp_BSCmp_op2_4, A0=>nx9720, A1=>
      nx9724);
   ix9721 : nor02_2x port map ( Y=>nx9720, A0=>nx9392, A1=>nx9388);
   ix9393 : nor03_2x port map ( Y=>nx9392, A0=>gen_24_cmp_mReg_3, A1=>
      nx10136, A2=>nx11850);
   ix9389 : nor03_2x port map ( Y=>nx9388, A0=>nx9716, A1=>nx11856, A2=>
      nx11866);
   ix9725 : nor02_2x port map ( Y=>nx9724, A0=>nx9384, A1=>nx9382);
   ix9385 : nor03_2x port map ( Y=>nx9384, A0=>nx9727, A1=>nx10130, A2=>
      nx11874);
   gen_24_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_24_cmp_mReg_4, QB=>
      nx9727, D=>window_24_4, CLK=>start, R=>rst);
   ix9383 : nor03_2x port map ( Y=>nx9382, A0=>gen_24_cmp_mReg_4, A1=>
      nx10874, A2=>nx11882);
   ix9419 : nand02 port map ( Y=>gen_24_cmp_BSCmp_op2_5, A0=>nx9731, A1=>
      nx9735);
   ix9732 : nor02_2x port map ( Y=>nx9731, A0=>nx9414, A1=>nx9410);
   ix9415 : nor03_2x port map ( Y=>nx9414, A0=>gen_24_cmp_mReg_4, A1=>
      nx10136, A2=>nx11850);
   ix9411 : nor03_2x port map ( Y=>nx9410, A0=>nx9727, A1=>nx11856, A2=>
      nx11866);
   ix9736 : nor02_2x port map ( Y=>nx9735, A0=>nx9406, A1=>nx9404);
   ix9407 : nor03_2x port map ( Y=>nx9406, A0=>nx9738, A1=>nx10132, A2=>
      nx11874);
   gen_24_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_24_cmp_mReg_5, QB=>
      nx9738, D=>window_24_5, CLK=>start, R=>rst);
   ix9405 : nor03_2x port map ( Y=>nx9404, A0=>gen_24_cmp_mReg_5, A1=>
      nx10874, A2=>nx11882);
   ix9441 : nand02 port map ( Y=>gen_24_cmp_BSCmp_op2_6, A0=>nx9742, A1=>
      nx9746);
   ix9743 : nor02_2x port map ( Y=>nx9742, A0=>nx9436, A1=>nx9432);
   ix9437 : nor03_2x port map ( Y=>nx9436, A0=>gen_24_cmp_mReg_5, A1=>
      nx10138, A2=>nx11850);
   ix9433 : nor03_2x port map ( Y=>nx9432, A0=>nx9738, A1=>nx11856, A2=>
      nx11866);
   ix9747 : nor02_2x port map ( Y=>nx9746, A0=>nx9428, A1=>nx9426);
   ix9429 : nor03_2x port map ( Y=>nx9428, A0=>nx9749, A1=>nx10132, A2=>
      nx11874);
   gen_24_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_24_cmp_mReg_6, QB=>
      nx9749, D=>window_24_6, CLK=>start, R=>rst);
   ix9427 : nor03_2x port map ( Y=>nx9426, A0=>gen_24_cmp_mReg_6, A1=>
      nx10874, A2=>nx11882);
   ix9463 : nand02 port map ( Y=>gen_24_cmp_BSCmp_op2_7, A0=>nx9753, A1=>
      nx9757);
   ix9754 : nor02_2x port map ( Y=>nx9753, A0=>nx9458, A1=>nx9454);
   ix9459 : nor03_2x port map ( Y=>nx9458, A0=>gen_24_cmp_mReg_6, A1=>
      nx10138, A2=>nx11852);
   ix9455 : nor03_2x port map ( Y=>nx9454, A0=>nx9749, A1=>nx11858, A2=>
      nx11868);
   ix9758 : nor02_2x port map ( Y=>nx9757, A0=>nx9450, A1=>nx9448);
   ix9451 : nor03_2x port map ( Y=>nx9450, A0=>nx9760, A1=>nx10132, A2=>
      nx11876);
   gen_24_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_24_cmp_mReg_7, QB=>
      nx9760, D=>window_24_7, CLK=>start, R=>rst);
   ix9449 : nor03_2x port map ( Y=>nx9448, A0=>gen_24_cmp_mReg_7, A1=>
      nx10874, A2=>nx11884);
   ix9485 : nand02 port map ( Y=>gen_24_cmp_BSCmp_op2_8, A0=>nx9764, A1=>
      nx9768);
   ix9765 : nor02_2x port map ( Y=>nx9764, A0=>nx9480, A1=>nx9476);
   ix9481 : nor03_2x port map ( Y=>nx9480, A0=>gen_24_cmp_mReg_7, A1=>
      nx10138, A2=>nx11852);
   ix9477 : nor03_2x port map ( Y=>nx9476, A0=>nx9760, A1=>nx11858, A2=>
      nx11868);
   ix9769 : nor02_2x port map ( Y=>nx9768, A0=>nx9472, A1=>nx9470);
   ix9473 : nor03_2x port map ( Y=>nx9472, A0=>nx9771, A1=>nx10132, A2=>
      nx11876);
   gen_24_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_24_cmp_mReg_8, QB=>
      nx9771, D=>window_24_8, CLK=>start, R=>rst);
   ix9471 : nor03_2x port map ( Y=>nx9470, A0=>gen_24_cmp_mReg_8, A1=>
      nx10876, A2=>nx11884);
   ix9507 : nand02 port map ( Y=>gen_24_cmp_BSCmp_op2_9, A0=>nx9775, A1=>
      nx9779);
   ix9776 : nor02_2x port map ( Y=>nx9775, A0=>nx9502, A1=>nx9498);
   ix9503 : nor03_2x port map ( Y=>nx9502, A0=>gen_24_cmp_mReg_8, A1=>
      nx10138, A2=>nx11852);
   ix9499 : nor03_2x port map ( Y=>nx9498, A0=>nx9771, A1=>nx11858, A2=>
      nx11868);
   ix9780 : nor02_2x port map ( Y=>nx9779, A0=>nx9494, A1=>nx9492);
   ix9495 : nor03_2x port map ( Y=>nx9494, A0=>nx9782, A1=>nx10132, A2=>
      nx11876);
   gen_24_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_24_cmp_mReg_9, QB=>
      nx9782, D=>window_24_9, CLK=>start, R=>rst);
   ix9493 : nor03_2x port map ( Y=>nx9492, A0=>gen_24_cmp_mReg_9, A1=>
      nx10876, A2=>nx11884);
   ix9529 : nand02 port map ( Y=>gen_24_cmp_BSCmp_op2_10, A0=>nx9786, A1=>
      nx9790);
   ix9787 : nor02_2x port map ( Y=>nx9786, A0=>nx9524, A1=>nx9520);
   ix9525 : nor03_2x port map ( Y=>nx9524, A0=>gen_24_cmp_mReg_9, A1=>
      nx10138, A2=>nx11852);
   ix9521 : nor03_2x port map ( Y=>nx9520, A0=>nx9782, A1=>nx11858, A2=>
      nx11868);
   ix9791 : nor02_2x port map ( Y=>nx9790, A0=>nx9516, A1=>nx9514);
   ix9517 : nor03_2x port map ( Y=>nx9516, A0=>nx9793, A1=>nx10132, A2=>
      nx11876);
   gen_24_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_24_cmp_mReg_10, QB=>
      nx9793, D=>window_24_10, CLK=>start, R=>rst);
   ix9515 : nor03_2x port map ( Y=>nx9514, A0=>gen_24_cmp_mReg_10, A1=>
      nx10876, A2=>nx11884);
   ix9551 : nand02 port map ( Y=>gen_24_cmp_BSCmp_op2_11, A0=>nx9797, A1=>
      nx9801);
   ix9798 : nor02_2x port map ( Y=>nx9797, A0=>nx9546, A1=>nx9542);
   ix9547 : nor03_2x port map ( Y=>nx9546, A0=>gen_24_cmp_mReg_10, A1=>
      nx10138, A2=>nx11852);
   ix9543 : nor03_2x port map ( Y=>nx9542, A0=>nx9793, A1=>nx11858, A2=>
      nx11868);
   ix9802 : nor02_2x port map ( Y=>nx9801, A0=>nx9538, A1=>nx9536);
   ix9539 : nor03_2x port map ( Y=>nx9538, A0=>nx9804, A1=>nx10132, A2=>
      nx11876);
   gen_24_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_24_cmp_mReg_11, QB=>
      nx9804, D=>window_24_11, CLK=>start, R=>rst);
   ix9537 : nor03_2x port map ( Y=>nx9536, A0=>gen_24_cmp_mReg_11, A1=>
      nx10876, A2=>nx11884);
   ix9573 : nand02 port map ( Y=>gen_24_cmp_BSCmp_op2_12, A0=>nx9808, A1=>
      nx9812);
   ix9809 : nor02_2x port map ( Y=>nx9808, A0=>nx9568, A1=>nx9564);
   ix9569 : nor03_2x port map ( Y=>nx9568, A0=>gen_24_cmp_mReg_11, A1=>
      nx10138, A2=>nx11852);
   ix9565 : nor03_2x port map ( Y=>nx9564, A0=>nx9804, A1=>nx11858, A2=>
      nx11868);
   ix9813 : nor02_2x port map ( Y=>nx9812, A0=>nx9560, A1=>nx9558);
   ix9561 : nor03_2x port map ( Y=>nx9560, A0=>nx9815, A1=>nx10134, A2=>
      nx11876);
   gen_24_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_24_cmp_mReg_12, QB=>
      nx9815, D=>window_24_12, CLK=>start, R=>rst);
   ix9559 : nor03_2x port map ( Y=>nx9558, A0=>gen_24_cmp_mReg_12, A1=>
      nx10876, A2=>nx11884);
   ix9595 : nand02 port map ( Y=>gen_24_cmp_BSCmp_op2_13, A0=>nx9819, A1=>
      nx9823);
   ix9820 : nor02_2x port map ( Y=>nx9819, A0=>nx9590, A1=>nx9586);
   ix9591 : nor03_2x port map ( Y=>nx9590, A0=>gen_24_cmp_mReg_12, A1=>
      nx10140, A2=>nx11854);
   ix9587 : nor03_2x port map ( Y=>nx9586, A0=>nx9815, A1=>nx11858, A2=>
      nx11870);
   ix9824 : nor02_2x port map ( Y=>nx9823, A0=>nx9582, A1=>nx9580);
   ix9583 : nor03_2x port map ( Y=>nx9582, A0=>nx9826, A1=>nx10134, A2=>
      nx11878);
   gen_24_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_24_cmp_mReg_13, QB=>
      nx9826, D=>window_24_13, CLK=>start, R=>rst);
   ix9581 : nor03_2x port map ( Y=>nx9580, A0=>gen_24_cmp_mReg_13, A1=>
      nx10876, A2=>nx11886);
   ix9617 : nand02 port map ( Y=>gen_24_cmp_BSCmp_op2_14, A0=>nx9830, A1=>
      nx9834);
   ix9831 : nor02_2x port map ( Y=>nx9830, A0=>nx9612, A1=>nx9608);
   ix9613 : nor03_2x port map ( Y=>nx9612, A0=>gen_24_cmp_mReg_13, A1=>
      nx10140, A2=>nx11854);
   ix9609 : nor03_2x port map ( Y=>nx9608, A0=>nx9826, A1=>nx11860, A2=>
      nx11870);
   ix9835 : nor02_2x port map ( Y=>nx9834, A0=>nx9604, A1=>nx9602);
   ix9605 : nor03_2x port map ( Y=>nx9604, A0=>nx9837, A1=>nx10134, A2=>
      nx11878);
   gen_24_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_24_cmp_mReg_14, QB=>
      nx9837, D=>window_24_14, CLK=>start, R=>rst);
   ix9603 : nor03_2x port map ( Y=>nx9602, A0=>gen_24_cmp_mReg_14, A1=>
      nx10876, A2=>nx11886);
   ix9639 : nand02 port map ( Y=>gen_24_cmp_BSCmp_op2_15, A0=>nx9841, A1=>
      nx9845);
   ix9842 : nor02_2x port map ( Y=>nx9841, A0=>nx9634, A1=>nx9630);
   ix9635 : nor03_2x port map ( Y=>nx9634, A0=>gen_24_cmp_mReg_14, A1=>
      nx10140, A2=>nx11854);
   ix9631 : nor03_2x port map ( Y=>nx9630, A0=>nx9837, A1=>nx11860, A2=>
      nx11870);
   ix9846 : nor02_2x port map ( Y=>nx9845, A0=>nx9626, A1=>nx9624);
   ix9627 : nor03_2x port map ( Y=>nx9626, A0=>nx9848, A1=>nx10134, A2=>
      nx11878);
   gen_24_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_24_cmp_mReg_15, QB=>
      nx9848, D=>window_24_15, CLK=>start, R=>rst);
   ix9625 : nor03_2x port map ( Y=>nx9624, A0=>gen_24_cmp_mReg_15, A1=>
      nx10878, A2=>nx11886);
   ix9649 : nand02 port map ( Y=>gen_24_cmp_BSCmp_op2_16, A0=>nx9852, A1=>
      nx9845);
   ix9853 : nor02_2x port map ( Y=>nx9852, A0=>nx9644, A1=>nx9640);
   ix9645 : nor03_2x port map ( Y=>nx9644, A0=>gen_24_cmp_mReg_15, A1=>
      nx10140, A2=>nx11854);
   ix9641 : nor03_2x port map ( Y=>nx9640, A0=>nx9848, A1=>nx11860, A2=>
      nx11870);
   ix19 : nor02_2x port map ( Y=>gen_0_cmp_BSCmp_carryIn, A0=>nx3769, A1=>
      nx9857);
   ix9858 : nor02_2x port map ( Y=>nx9857, A0=>nx10900, A1=>nx3761);
   ix39 : nand02 port map ( Y=>gen_0_cmp_BSCmp_op2_0, A0=>nx9860, A1=>nx9864
   );
   ix9861 : nor02_2x port map ( Y=>nx9860, A0=>nx34, A1=>nx26);
   ix35 : nor03_2x port map ( Y=>nx34, A0=>nx3757, A1=>nx10422, A2=>nx10918
   );
   ix27 : nor03_2x port map ( Y=>nx26, A0=>gen_0_cmp_mReg_0, A1=>nx10734, A2
      =>nx10926);
   ix9865 : nand03 port map ( Y=>nx9864, A0=>nx10900, A1=>nx10422, A2=>
      nx3761);
   ix405 : nor02_2x port map ( Y=>gen_1_cmp_BSCmp_carryIn, A0=>nx4013, A1=>
      nx9867);
   ix9868 : nor02_2x port map ( Y=>nx9867, A0=>nx10940, A1=>nx4005);
   ix425 : nand02 port map ( Y=>gen_1_cmp_BSCmp_op2_0, A0=>nx9870, A1=>
      nx9874);
   ix9871 : nor02_2x port map ( Y=>nx9870, A0=>nx420, A1=>nx412);
   ix421 : nor03_2x port map ( Y=>nx420, A0=>nx4001, A1=>nx10410, A2=>
      nx10958);
   ix413 : nor03_2x port map ( Y=>nx412, A0=>gen_1_cmp_mReg_0, A1=>nx10740, 
      A2=>nx10966);
   ix9875 : nand03 port map ( Y=>nx9874, A0=>nx10940, A1=>nx10410, A2=>
      nx4005);
   ix791 : nor02_2x port map ( Y=>gen_2_cmp_BSCmp_carryIn, A0=>nx4260, A1=>
      nx9877);
   ix9878 : nor02_2x port map ( Y=>nx9877, A0=>nx10980, A1=>nx4253);
   ix811 : nand02 port map ( Y=>gen_2_cmp_BSCmp_op2_0, A0=>nx9880, A1=>
      nx9884);
   ix9881 : nor02_2x port map ( Y=>nx9880, A0=>nx806, A1=>nx798);
   ix807 : nor03_2x port map ( Y=>nx806, A0=>nx4249, A1=>nx10398, A2=>
      nx10998);
   ix799 : nor03_2x port map ( Y=>nx798, A0=>gen_2_cmp_mReg_0, A1=>nx10746, 
      A2=>nx11006);
   ix9885 : nand03 port map ( Y=>nx9884, A0=>nx10980, A1=>nx10398, A2=>
      nx4253);
   ix1177 : nor02_2x port map ( Y=>gen_3_cmp_BSCmp_carryIn, A0=>nx4509, A1=>
      nx9887);
   ix9888 : nor02_2x port map ( Y=>nx9887, A0=>nx11020, A1=>nx4501);
   ix1197 : nand02 port map ( Y=>gen_3_cmp_BSCmp_op2_0, A0=>nx9890, A1=>
      nx9894);
   ix9891 : nor02_2x port map ( Y=>nx9890, A0=>nx1192, A1=>nx1184);
   ix1193 : nor03_2x port map ( Y=>nx1192, A0=>nx4497, A1=>nx10386, A2=>
      nx11038);
   ix1185 : nor03_2x port map ( Y=>nx1184, A0=>gen_3_cmp_mReg_0, A1=>nx10752, 
      A2=>nx11046);
   ix9895 : nand03 port map ( Y=>nx9894, A0=>nx11020, A1=>nx10386, A2=>
      nx4501);
   ix1563 : nor02_2x port map ( Y=>gen_4_cmp_BSCmp_carryIn, A0=>nx4757, A1=>
      nx9897);
   ix9898 : nor02_2x port map ( Y=>nx9897, A0=>nx11060, A1=>nx4748);
   ix1583 : nand02 port map ( Y=>gen_4_cmp_BSCmp_op2_0, A0=>nx9900, A1=>
      nx9904);
   ix9901 : nor02_2x port map ( Y=>nx9900, A0=>nx1578, A1=>nx1570);
   ix1579 : nor03_2x port map ( Y=>nx1578, A0=>nx4745, A1=>nx10374, A2=>
      nx11078);
   ix1571 : nor03_2x port map ( Y=>nx1570, A0=>gen_4_cmp_mReg_0, A1=>nx10758, 
      A2=>nx11086);
   ix9905 : nand03 port map ( Y=>nx9904, A0=>nx11060, A1=>nx10374, A2=>
      nx4748);
   ix1949 : nor02_2x port map ( Y=>gen_5_cmp_BSCmp_carryIn, A0=>nx5003, A1=>
      nx9907);
   ix9908 : nor02_2x port map ( Y=>nx9907, A0=>nx11100, A1=>nx4995);
   ix1969 : nand02 port map ( Y=>gen_5_cmp_BSCmp_op2_0, A0=>nx9910, A1=>
      nx9914);
   ix9911 : nor02_2x port map ( Y=>nx9910, A0=>nx1964, A1=>nx1956);
   ix1965 : nor03_2x port map ( Y=>nx1964, A0=>nx4991, A1=>nx10362, A2=>
      nx11118);
   ix1957 : nor03_2x port map ( Y=>nx1956, A0=>gen_5_cmp_mReg_0, A1=>nx10764, 
      A2=>nx11126);
   ix9915 : nand03 port map ( Y=>nx9914, A0=>nx11100, A1=>nx10362, A2=>
      nx4995);
   ix2335 : nor02_2x port map ( Y=>gen_6_cmp_BSCmp_carryIn, A0=>nx5253, A1=>
      nx9917);
   ix9918 : nor02_2x port map ( Y=>nx9917, A0=>nx11140, A1=>nx5244);
   ix2355 : nand02 port map ( Y=>gen_6_cmp_BSCmp_op2_0, A0=>nx9920, A1=>
      nx9924);
   ix9921 : nor02_2x port map ( Y=>nx9920, A0=>nx2350, A1=>nx2342);
   ix2351 : nor03_2x port map ( Y=>nx2350, A0=>nx5241, A1=>nx10350, A2=>
      nx11158);
   ix2343 : nor03_2x port map ( Y=>nx2342, A0=>gen_6_cmp_mReg_0, A1=>nx10770, 
      A2=>nx11166);
   ix9925 : nand03 port map ( Y=>nx9924, A0=>nx11140, A1=>nx10350, A2=>
      nx5244);
   ix2721 : nor02_2x port map ( Y=>gen_7_cmp_BSCmp_carryIn, A0=>nx5499, A1=>
      nx9927);
   ix9928 : nor02_2x port map ( Y=>nx9927, A0=>nx11180, A1=>nx5491);
   ix2741 : nand02 port map ( Y=>gen_7_cmp_BSCmp_op2_0, A0=>nx9930, A1=>
      nx9934);
   ix9931 : nor02_2x port map ( Y=>nx9930, A0=>nx2736, A1=>nx2728);
   ix2737 : nor03_2x port map ( Y=>nx2736, A0=>nx5487, A1=>nx10338, A2=>
      nx11198);
   ix2729 : nor03_2x port map ( Y=>nx2728, A0=>gen_7_cmp_mReg_0, A1=>nx10776, 
      A2=>nx11206);
   ix9935 : nand03 port map ( Y=>nx9934, A0=>nx11180, A1=>nx10338, A2=>
      nx5491);
   ix3107 : nor02_2x port map ( Y=>gen_8_cmp_BSCmp_carryIn, A0=>nx5743, A1=>
      nx9937);
   ix9938 : nor02_2x port map ( Y=>nx9937, A0=>nx11220, A1=>nx5735);
   ix3127 : nand02 port map ( Y=>gen_8_cmp_BSCmp_op2_0, A0=>nx9940, A1=>
      nx9944);
   ix9941 : nor02_2x port map ( Y=>nx9940, A0=>nx3122, A1=>nx3114);
   ix3123 : nor03_2x port map ( Y=>nx3122, A0=>nx5731, A1=>nx10326, A2=>
      nx11238);
   ix3115 : nor03_2x port map ( Y=>nx3114, A0=>gen_8_cmp_mReg_0, A1=>nx10782, 
      A2=>nx11246);
   ix9945 : nand03 port map ( Y=>nx9944, A0=>nx11220, A1=>nx10326, A2=>
      nx5735);
   ix3493 : nor02_2x port map ( Y=>gen_9_cmp_BSCmp_carryIn, A0=>nx5987, A1=>
      nx9947);
   ix9948 : nor02_2x port map ( Y=>nx9947, A0=>nx11260, A1=>nx5979);
   ix3513 : nand02 port map ( Y=>gen_9_cmp_BSCmp_op2_0, A0=>nx9950, A1=>
      nx9954);
   ix9951 : nor02_2x port map ( Y=>nx9950, A0=>nx3508, A1=>nx3500);
   ix3509 : nor03_2x port map ( Y=>nx3508, A0=>nx5975, A1=>nx10314, A2=>
      nx11278);
   ix3501 : nor03_2x port map ( Y=>nx3500, A0=>gen_9_cmp_mReg_0, A1=>nx10788, 
      A2=>nx11286);
   ix9955 : nand03 port map ( Y=>nx9954, A0=>nx11260, A1=>nx10314, A2=>
      nx5979);
   ix3879 : nor02_2x port map ( Y=>gen_10_cmp_BSCmp_carryIn, A0=>nx6233, A1
      =>nx9957);
   ix9958 : nor02_2x port map ( Y=>nx9957, A0=>nx11300, A1=>nx6225);
   ix3899 : nand02 port map ( Y=>gen_10_cmp_BSCmp_op2_0, A0=>nx9960, A1=>
      nx9964);
   ix9961 : nor02_2x port map ( Y=>nx9960, A0=>nx3894, A1=>nx3886);
   ix3895 : nor03_2x port map ( Y=>nx3894, A0=>nx6221, A1=>nx10302, A2=>
      nx11318);
   ix3887 : nor03_2x port map ( Y=>nx3886, A0=>gen_10_cmp_mReg_0, A1=>
      nx10794, A2=>nx11326);
   ix9965 : nand03 port map ( Y=>nx9964, A0=>nx11300, A1=>nx10302, A2=>
      nx6225);
   ix4265 : nor02_2x port map ( Y=>gen_11_cmp_BSCmp_carryIn, A0=>nx6477, A1
      =>nx9967);
   ix9968 : nor02_2x port map ( Y=>nx9967, A0=>nx11340, A1=>nx6468);
   ix4285 : nand02 port map ( Y=>gen_11_cmp_BSCmp_op2_0, A0=>nx9970, A1=>
      nx9974);
   ix9971 : nor02_2x port map ( Y=>nx9970, A0=>nx4280, A1=>nx4272);
   ix4281 : nor03_2x port map ( Y=>nx4280, A0=>nx6465, A1=>nx10290, A2=>
      nx11358);
   ix4273 : nor03_2x port map ( Y=>nx4272, A0=>gen_11_cmp_mReg_0, A1=>
      nx10800, A2=>nx11366);
   ix9975 : nand03 port map ( Y=>nx9974, A0=>nx11340, A1=>nx10290, A2=>
      nx6468);
   ix4651 : nor02_2x port map ( Y=>gen_12_cmp_BSCmp_carryIn, A0=>nx6725, A1
      =>nx9977);
   ix9978 : nor02_2x port map ( Y=>nx9977, A0=>nx11380, A1=>nx6717);
   ix4671 : nand02 port map ( Y=>gen_12_cmp_BSCmp_op2_0, A0=>nx9980, A1=>
      nx9984);
   ix9981 : nor02_2x port map ( Y=>nx9980, A0=>nx4666, A1=>nx4658);
   ix4667 : nor03_2x port map ( Y=>nx4666, A0=>nx6713, A1=>nx10278, A2=>
      nx11398);
   ix4659 : nor03_2x port map ( Y=>nx4658, A0=>gen_12_cmp_mReg_0, A1=>
      nx10806, A2=>nx11406);
   ix9985 : nand03 port map ( Y=>nx9984, A0=>nx11380, A1=>nx10278, A2=>
      nx6717);
   ix5037 : nor02_2x port map ( Y=>gen_13_cmp_BSCmp_carryIn, A0=>nx6973, A1
      =>nx9987);
   ix9988 : nor02_2x port map ( Y=>nx9987, A0=>nx11420, A1=>nx6965);
   ix5057 : nand02 port map ( Y=>gen_13_cmp_BSCmp_op2_0, A0=>nx9990, A1=>
      nx9994);
   ix9991 : nor02_2x port map ( Y=>nx9990, A0=>nx5052, A1=>nx5044);
   ix5053 : nor03_2x port map ( Y=>nx5052, A0=>nx6961, A1=>nx10266, A2=>
      nx11438);
   ix5045 : nor03_2x port map ( Y=>nx5044, A0=>gen_13_cmp_mReg_0, A1=>
      nx10812, A2=>nx11446);
   ix9995 : nand03 port map ( Y=>nx9994, A0=>nx11420, A1=>nx10266, A2=>
      nx6965);
   ix5423 : nor02_2x port map ( Y=>gen_14_cmp_BSCmp_carryIn, A0=>nx7221, A1
      =>nx9997);
   ix9998 : nor02_2x port map ( Y=>nx9997, A0=>nx11460, A1=>nx7213);
   ix5443 : nand02 port map ( Y=>gen_14_cmp_BSCmp_op2_0, A0=>nx10000, A1=>
      nx10004);
   ix10001 : nor02_2x port map ( Y=>nx10000, A0=>nx5438, A1=>nx5430);
   ix5439 : nor03_2x port map ( Y=>nx5438, A0=>nx7209, A1=>nx10254, A2=>
      nx11478);
   ix5431 : nor03_2x port map ( Y=>nx5430, A0=>gen_14_cmp_mReg_0, A1=>
      nx10818, A2=>nx11486);
   ix10005 : nand03 port map ( Y=>nx10004, A0=>nx11460, A1=>nx10254, A2=>
      nx7213);
   ix5809 : nor02_2x port map ( Y=>gen_15_cmp_BSCmp_carryIn, A0=>nx7471, A1
      =>nx10007);
   ix10008 : nor02_2x port map ( Y=>nx10007, A0=>nx11500, A1=>nx7463);
   ix5829 : nand02 port map ( Y=>gen_15_cmp_BSCmp_op2_0, A0=>nx10010, A1=>
      nx10014);
   ix10011 : nor02_2x port map ( Y=>nx10010, A0=>nx5824, A1=>nx5816);
   ix5825 : nor03_2x port map ( Y=>nx5824, A0=>nx7459, A1=>nx10242, A2=>
      nx11518);
   ix5817 : nor03_2x port map ( Y=>nx5816, A0=>gen_15_cmp_mReg_0, A1=>
      nx10824, A2=>nx11526);
   ix10015 : nand03 port map ( Y=>nx10014, A0=>nx11500, A1=>nx10242, A2=>
      nx7463);
   ix6195 : nor02_2x port map ( Y=>gen_16_cmp_BSCmp_carryIn, A0=>nx7717, A1
      =>nx10017);
   ix10018 : nor02_2x port map ( Y=>nx10017, A0=>nx11540, A1=>nx7709);
   ix6215 : nand02 port map ( Y=>gen_16_cmp_BSCmp_op2_0, A0=>nx10020, A1=>
      nx10024);
   ix10021 : nor02_2x port map ( Y=>nx10020, A0=>nx6210, A1=>nx6202);
   ix6211 : nor03_2x port map ( Y=>nx6210, A0=>nx7705, A1=>nx10230, A2=>
      nx11558);
   ix6203 : nor03_2x port map ( Y=>nx6202, A0=>gen_16_cmp_mReg_0, A1=>
      nx10830, A2=>nx11566);
   ix10025 : nand03 port map ( Y=>nx10024, A0=>nx11540, A1=>nx10230, A2=>
      nx7709);
   ix6581 : nor02_2x port map ( Y=>gen_17_cmp_BSCmp_carryIn, A0=>nx7961, A1
      =>nx10027);
   ix10028 : nor02_2x port map ( Y=>nx10027, A0=>nx11580, A1=>nx7953);
   ix6601 : nand02 port map ( Y=>gen_17_cmp_BSCmp_op2_0, A0=>nx10030, A1=>
      nx10034);
   ix10031 : nor02_2x port map ( Y=>nx10030, A0=>nx6596, A1=>nx6588);
   ix6597 : nor03_2x port map ( Y=>nx6596, A0=>nx7949, A1=>nx10218, A2=>
      nx11598);
   ix6589 : nor03_2x port map ( Y=>nx6588, A0=>gen_17_cmp_mReg_0, A1=>
      nx10836, A2=>nx11606);
   ix10035 : nand03 port map ( Y=>nx10034, A0=>nx11580, A1=>nx10218, A2=>
      nx7953);
   ix6967 : nor02_2x port map ( Y=>gen_18_cmp_BSCmp_carryIn, A0=>nx8209, A1
      =>nx10037);
   ix10038 : nor02_2x port map ( Y=>nx10037, A0=>nx11620, A1=>nx8200);
   ix6987 : nand02 port map ( Y=>gen_18_cmp_BSCmp_op2_0, A0=>nx10040, A1=>
      nx10044);
   ix10041 : nor02_2x port map ( Y=>nx10040, A0=>nx6982, A1=>nx6974);
   ix6983 : nor03_2x port map ( Y=>nx6982, A0=>nx8197, A1=>nx10206, A2=>
      nx11638);
   ix6975 : nor03_2x port map ( Y=>nx6974, A0=>gen_18_cmp_mReg_0, A1=>
      nx10842, A2=>nx11646);
   ix10045 : nand03 port map ( Y=>nx10044, A0=>nx11620, A1=>nx10206, A2=>
      nx8200);
   ix7353 : nor02_2x port map ( Y=>gen_19_cmp_BSCmp_carryIn, A0=>nx8455, A1
      =>nx10047);
   ix10048 : nor02_2x port map ( Y=>nx10047, A0=>nx11660, A1=>nx8447);
   ix7373 : nand02 port map ( Y=>gen_19_cmp_BSCmp_op2_0, A0=>nx10050, A1=>
      nx10054);
   ix10051 : nor02_2x port map ( Y=>nx10050, A0=>nx7368, A1=>nx7360);
   ix7369 : nor03_2x port map ( Y=>nx7368, A0=>nx8443, A1=>nx10194, A2=>
      nx11678);
   ix7361 : nor03_2x port map ( Y=>nx7360, A0=>gen_19_cmp_mReg_0, A1=>
      nx10848, A2=>nx11686);
   ix10055 : nand03 port map ( Y=>nx10054, A0=>nx11660, A1=>nx10194, A2=>
      nx8447);
   ix7739 : nor02_2x port map ( Y=>gen_20_cmp_BSCmp_carryIn, A0=>nx8701, A1
      =>nx10057);
   ix10058 : nor02_2x port map ( Y=>nx10057, A0=>nx11700, A1=>nx8694);
   ix7759 : nand02 port map ( Y=>gen_20_cmp_BSCmp_op2_0, A0=>nx10060, A1=>
      nx10064);
   ix10061 : nor02_2x port map ( Y=>nx10060, A0=>nx7754, A1=>nx7746);
   ix7755 : nor03_2x port map ( Y=>nx7754, A0=>nx8691, A1=>nx10182, A2=>
      nx11718);
   ix7747 : nor03_2x port map ( Y=>nx7746, A0=>gen_20_cmp_mReg_0, A1=>
      nx10854, A2=>nx11726);
   ix10065 : nand03 port map ( Y=>nx10064, A0=>nx11700, A1=>nx10182, A2=>
      nx8694);
   ix8125 : nor02_2x port map ( Y=>gen_21_cmp_BSCmp_carryIn, A0=>nx8945, A1
      =>nx10067);
   ix10068 : nor02_2x port map ( Y=>nx10067, A0=>nx11740, A1=>nx8937);
   ix8145 : nand02 port map ( Y=>gen_21_cmp_BSCmp_op2_0, A0=>nx10070, A1=>
      nx10074);
   ix10071 : nor02_2x port map ( Y=>nx10070, A0=>nx8140, A1=>nx8132);
   ix8141 : nor03_2x port map ( Y=>nx8140, A0=>nx8933, A1=>nx10170, A2=>
      nx11758);
   ix8133 : nor03_2x port map ( Y=>nx8132, A0=>gen_21_cmp_mReg_0, A1=>
      nx10860, A2=>nx11766);
   ix10075 : nand03 port map ( Y=>nx10074, A0=>nx11740, A1=>nx10170, A2=>
      nx8937);
   ix8511 : nor02_2x port map ( Y=>gen_22_cmp_BSCmp_carryIn, A0=>nx9195, A1
      =>nx10077);
   ix10078 : nor02_2x port map ( Y=>nx10077, A0=>nx11780, A1=>nx9187);
   ix8531 : nand02 port map ( Y=>gen_22_cmp_BSCmp_op2_0, A0=>nx10080, A1=>
      nx10084);
   ix10081 : nor02_2x port map ( Y=>nx10080, A0=>nx8526, A1=>nx8518);
   ix8527 : nor03_2x port map ( Y=>nx8526, A0=>nx9183, A1=>nx10158, A2=>
      nx11798);
   ix8519 : nor03_2x port map ( Y=>nx8518, A0=>gen_22_cmp_mReg_0, A1=>
      nx10866, A2=>nx11806);
   ix10085 : nand03 port map ( Y=>nx10084, A0=>nx11780, A1=>nx10158, A2=>
      nx9187);
   ix8897 : nor02_2x port map ( Y=>gen_23_cmp_BSCmp_carryIn, A0=>nx9445, A1
      =>nx10087);
   ix10088 : nor02_2x port map ( Y=>nx10087, A0=>nx11820, A1=>nx9437);
   ix8917 : nand02 port map ( Y=>gen_23_cmp_BSCmp_op2_0, A0=>nx10090, A1=>
      nx10094);
   ix10091 : nor02_2x port map ( Y=>nx10090, A0=>nx8912, A1=>nx8904);
   ix8913 : nor03_2x port map ( Y=>nx8912, A0=>nx9433, A1=>nx10146, A2=>
      nx11838);
   ix8905 : nor03_2x port map ( Y=>nx8904, A0=>gen_23_cmp_mReg_0, A1=>
      nx10872, A2=>nx11846);
   ix10095 : nand03 port map ( Y=>nx10094, A0=>nx11820, A1=>nx10146, A2=>
      nx9437);
   ix9283 : nor02_2x port map ( Y=>gen_24_cmp_BSCmp_carryIn, A0=>nx9683, A1
      =>nx10097);
   ix10098 : nor02_2x port map ( Y=>nx10097, A0=>nx11860, A1=>nx9676);
   ix9303 : nand02 port map ( Y=>gen_24_cmp_BSCmp_op2_0, A0=>nx10100, A1=>
      nx10104);
   ix10101 : nor02_2x port map ( Y=>nx10100, A0=>nx9298, A1=>nx9290);
   ix9299 : nor03_2x port map ( Y=>nx9298, A0=>nx9673, A1=>nx10134, A2=>
      nx11878);
   ix9291 : nor03_2x port map ( Y=>nx9290, A0=>gen_24_cmp_mReg_0, A1=>
      nx10878, A2=>nx11886);
   ix10105 : nand03 port map ( Y=>nx10104, A0=>nx11860, A1=>nx10134, A2=>
      nx9676);
   ix9695 : nor02_2x port map ( Y=>working, A0=>nx10107, A1=>nx11934);
   firtStartLachCmp_reg_Q_0 : dffr port map ( Q=>OPEN, QB=>nx10107, D=>
      nx9650, CLK=>start, R=>rst);
   ix10119 : inv01 port map ( Y=>nx10120, A=>nx3745);
   ix10121 : inv01 port map ( Y=>nx10122, A=>clk);
   ix10123 : inv01 port map ( Y=>nx10124, A=>clk);
   ix10125 : inv01 port map ( Y=>nx10126, A=>clk);
   ix10127 : inv01 port map ( Y=>nx10128, A=>clk);
   ix10129 : inv04 port map ( Y=>nx10130, A=>nx9683);
   ix10131 : inv04 port map ( Y=>nx10132, A=>nx9683);
   ix10133 : inv04 port map ( Y=>nx10134, A=>nx9683);
   ix10135 : inv04 port map ( Y=>nx10136, A=>nx11860);
   ix10137 : inv04 port map ( Y=>nx10138, A=>nx11860);
   ix10139 : inv04 port map ( Y=>nx10140, A=>nx11862);
   ix10141 : inv04 port map ( Y=>nx10142, A=>nx9445);
   ix10143 : inv04 port map ( Y=>nx10144, A=>nx9445);
   ix10145 : inv04 port map ( Y=>nx10146, A=>nx9445);
   ix10147 : inv04 port map ( Y=>nx10148, A=>nx11820);
   ix10149 : inv04 port map ( Y=>nx10150, A=>nx11820);
   ix10151 : inv04 port map ( Y=>nx10152, A=>nx11822);
   ix10153 : inv04 port map ( Y=>nx10154, A=>nx9195);
   ix10155 : inv04 port map ( Y=>nx10156, A=>nx9195);
   ix10157 : inv04 port map ( Y=>nx10158, A=>nx9195);
   ix10159 : inv04 port map ( Y=>nx10160, A=>nx11780);
   ix10161 : inv04 port map ( Y=>nx10162, A=>nx11780);
   ix10163 : inv04 port map ( Y=>nx10164, A=>nx11782);
   ix10165 : inv04 port map ( Y=>nx10166, A=>nx8945);
   ix10167 : inv04 port map ( Y=>nx10168, A=>nx8945);
   ix10169 : inv04 port map ( Y=>nx10170, A=>nx8945);
   ix10171 : inv04 port map ( Y=>nx10172, A=>nx11740);
   ix10173 : inv04 port map ( Y=>nx10174, A=>nx11740);
   ix10175 : inv04 port map ( Y=>nx10176, A=>nx11742);
   ix10177 : inv04 port map ( Y=>nx10178, A=>nx8701);
   ix10179 : inv04 port map ( Y=>nx10180, A=>nx8701);
   ix10181 : inv04 port map ( Y=>nx10182, A=>nx8701);
   ix10183 : inv04 port map ( Y=>nx10184, A=>nx11700);
   ix10185 : inv04 port map ( Y=>nx10186, A=>nx11700);
   ix10187 : inv04 port map ( Y=>nx10188, A=>nx11702);
   ix10189 : inv04 port map ( Y=>nx10190, A=>nx8455);
   ix10191 : inv04 port map ( Y=>nx10192, A=>nx8455);
   ix10193 : inv04 port map ( Y=>nx10194, A=>nx8455);
   ix10195 : inv04 port map ( Y=>nx10196, A=>nx11660);
   ix10197 : inv04 port map ( Y=>nx10198, A=>nx11660);
   ix10199 : inv04 port map ( Y=>nx10200, A=>nx11662);
   ix10201 : inv04 port map ( Y=>nx10202, A=>nx8209);
   ix10203 : inv04 port map ( Y=>nx10204, A=>nx8209);
   ix10205 : inv04 port map ( Y=>nx10206, A=>nx8209);
   ix10207 : inv04 port map ( Y=>nx10208, A=>nx11620);
   ix10209 : inv04 port map ( Y=>nx10210, A=>nx11620);
   ix10211 : inv04 port map ( Y=>nx10212, A=>nx11622);
   ix10213 : inv04 port map ( Y=>nx10214, A=>nx7961);
   ix10215 : inv04 port map ( Y=>nx10216, A=>nx7961);
   ix10217 : inv04 port map ( Y=>nx10218, A=>nx7961);
   ix10219 : inv04 port map ( Y=>nx10220, A=>nx11580);
   ix10221 : inv04 port map ( Y=>nx10222, A=>nx11580);
   ix10223 : inv04 port map ( Y=>nx10224, A=>nx11582);
   ix10225 : inv04 port map ( Y=>nx10226, A=>nx7717);
   ix10227 : inv04 port map ( Y=>nx10228, A=>nx7717);
   ix10229 : inv04 port map ( Y=>nx10230, A=>nx7717);
   ix10231 : inv04 port map ( Y=>nx10232, A=>nx11540);
   ix10233 : inv04 port map ( Y=>nx10234, A=>nx11540);
   ix10235 : inv04 port map ( Y=>nx10236, A=>nx11542);
   ix10237 : inv04 port map ( Y=>nx10238, A=>nx7471);
   ix10239 : inv04 port map ( Y=>nx10240, A=>nx7471);
   ix10241 : inv04 port map ( Y=>nx10242, A=>nx7471);
   ix10243 : inv04 port map ( Y=>nx10244, A=>nx11500);
   ix10245 : inv04 port map ( Y=>nx10246, A=>nx11500);
   ix10247 : inv04 port map ( Y=>nx10248, A=>nx11502);
   ix10249 : inv04 port map ( Y=>nx10250, A=>nx7221);
   ix10251 : inv04 port map ( Y=>nx10252, A=>nx7221);
   ix10253 : inv04 port map ( Y=>nx10254, A=>nx7221);
   ix10255 : inv04 port map ( Y=>nx10256, A=>nx11460);
   ix10257 : inv04 port map ( Y=>nx10258, A=>nx11460);
   ix10259 : inv04 port map ( Y=>nx10260, A=>nx11462);
   ix10261 : inv04 port map ( Y=>nx10262, A=>nx6973);
   ix10263 : inv04 port map ( Y=>nx10264, A=>nx6973);
   ix10265 : inv04 port map ( Y=>nx10266, A=>nx6973);
   ix10267 : inv04 port map ( Y=>nx10268, A=>nx11420);
   ix10269 : inv04 port map ( Y=>nx10270, A=>nx11420);
   ix10271 : inv04 port map ( Y=>nx10272, A=>nx11422);
   ix10273 : inv04 port map ( Y=>nx10274, A=>nx6725);
   ix10275 : inv04 port map ( Y=>nx10276, A=>nx6725);
   ix10277 : inv04 port map ( Y=>nx10278, A=>nx6725);
   ix10279 : inv04 port map ( Y=>nx10280, A=>nx11380);
   ix10281 : inv04 port map ( Y=>nx10282, A=>nx11380);
   ix10283 : inv04 port map ( Y=>nx10284, A=>nx11382);
   ix10285 : inv04 port map ( Y=>nx10286, A=>nx6477);
   ix10287 : inv04 port map ( Y=>nx10288, A=>nx6477);
   ix10289 : inv04 port map ( Y=>nx10290, A=>nx6477);
   ix10291 : inv04 port map ( Y=>nx10292, A=>nx11340);
   ix10293 : inv04 port map ( Y=>nx10294, A=>nx11340);
   ix10295 : inv04 port map ( Y=>nx10296, A=>nx11342);
   ix10297 : inv04 port map ( Y=>nx10298, A=>nx6233);
   ix10299 : inv04 port map ( Y=>nx10300, A=>nx6233);
   ix10301 : inv04 port map ( Y=>nx10302, A=>nx6233);
   ix10303 : inv04 port map ( Y=>nx10304, A=>nx11300);
   ix10305 : inv04 port map ( Y=>nx10306, A=>nx11300);
   ix10307 : inv04 port map ( Y=>nx10308, A=>nx11302);
   ix10309 : inv04 port map ( Y=>nx10310, A=>nx5987);
   ix10311 : inv04 port map ( Y=>nx10312, A=>nx5987);
   ix10313 : inv04 port map ( Y=>nx10314, A=>nx5987);
   ix10315 : inv04 port map ( Y=>nx10316, A=>nx11260);
   ix10317 : inv04 port map ( Y=>nx10318, A=>nx11260);
   ix10319 : inv04 port map ( Y=>nx10320, A=>nx11262);
   ix10321 : inv04 port map ( Y=>nx10322, A=>nx5743);
   ix10323 : inv04 port map ( Y=>nx10324, A=>nx5743);
   ix10325 : inv04 port map ( Y=>nx10326, A=>nx5743);
   ix10327 : inv04 port map ( Y=>nx10328, A=>nx11220);
   ix10329 : inv04 port map ( Y=>nx10330, A=>nx11220);
   ix10331 : inv04 port map ( Y=>nx10332, A=>nx11222);
   ix10333 : inv04 port map ( Y=>nx10334, A=>nx5499);
   ix10335 : inv04 port map ( Y=>nx10336, A=>nx5499);
   ix10337 : inv04 port map ( Y=>nx10338, A=>nx5499);
   ix10339 : inv04 port map ( Y=>nx10340, A=>nx11180);
   ix10341 : inv04 port map ( Y=>nx10342, A=>nx11180);
   ix10343 : inv04 port map ( Y=>nx10344, A=>nx11182);
   ix10345 : inv04 port map ( Y=>nx10346, A=>nx5253);
   ix10347 : inv04 port map ( Y=>nx10348, A=>nx5253);
   ix10349 : inv04 port map ( Y=>nx10350, A=>nx5253);
   ix10351 : inv04 port map ( Y=>nx10352, A=>nx11140);
   ix10353 : inv04 port map ( Y=>nx10354, A=>nx11140);
   ix10355 : inv04 port map ( Y=>nx10356, A=>nx11142);
   ix10357 : inv04 port map ( Y=>nx10358, A=>nx5003);
   ix10359 : inv04 port map ( Y=>nx10360, A=>nx5003);
   ix10361 : inv04 port map ( Y=>nx10362, A=>nx5003);
   ix10363 : inv04 port map ( Y=>nx10364, A=>nx11100);
   ix10365 : inv04 port map ( Y=>nx10366, A=>nx11100);
   ix10367 : inv04 port map ( Y=>nx10368, A=>nx11102);
   ix10369 : inv04 port map ( Y=>nx10370, A=>nx4757);
   ix10371 : inv04 port map ( Y=>nx10372, A=>nx4757);
   ix10373 : inv04 port map ( Y=>nx10374, A=>nx4757);
   ix10375 : inv04 port map ( Y=>nx10376, A=>nx11060);
   ix10377 : inv04 port map ( Y=>nx10378, A=>nx11060);
   ix10379 : inv04 port map ( Y=>nx10380, A=>nx11062);
   ix10381 : inv04 port map ( Y=>nx10382, A=>nx4509);
   ix10383 : inv04 port map ( Y=>nx10384, A=>nx4509);
   ix10385 : inv04 port map ( Y=>nx10386, A=>nx4509);
   ix10387 : inv04 port map ( Y=>nx10388, A=>nx11020);
   ix10389 : inv04 port map ( Y=>nx10390, A=>nx11020);
   ix10391 : inv04 port map ( Y=>nx10392, A=>nx11022);
   ix10393 : inv04 port map ( Y=>nx10394, A=>nx4260);
   ix10395 : inv04 port map ( Y=>nx10396, A=>nx4260);
   ix10397 : inv04 port map ( Y=>nx10398, A=>nx4260);
   ix10399 : inv04 port map ( Y=>nx10400, A=>nx10980);
   ix10401 : inv04 port map ( Y=>nx10402, A=>nx10980);
   ix10403 : inv04 port map ( Y=>nx10404, A=>nx10982);
   ix10405 : inv04 port map ( Y=>nx10406, A=>nx4013);
   ix10407 : inv04 port map ( Y=>nx10408, A=>nx4013);
   ix10409 : inv04 port map ( Y=>nx10410, A=>nx4013);
   ix10411 : inv04 port map ( Y=>nx10412, A=>nx10940);
   ix10413 : inv04 port map ( Y=>nx10414, A=>nx10940);
   ix10415 : inv04 port map ( Y=>nx10416, A=>nx10942);
   ix10417 : inv04 port map ( Y=>nx10418, A=>nx3769);
   ix10419 : inv04 port map ( Y=>nx10420, A=>nx3769);
   ix10421 : inv04 port map ( Y=>nx10422, A=>nx3769);
   ix10423 : inv04 port map ( Y=>nx10424, A=>nx10900);
   ix10425 : inv04 port map ( Y=>nx10426, A=>nx10900);
   ix10427 : inv04 port map ( Y=>nx10428, A=>nx10902);
   ix10429 : inv01 port map ( Y=>nx10430, A=>gen_24_cmp_BSCmp_op2_16);
   ix10431 : inv02 port map ( Y=>nx10432, A=>nx10430);
   ix10433 : inv02 port map ( Y=>nx10434, A=>nx10430);
   ix10435 : inv02 port map ( Y=>nx10436, A=>nx10430);
   ix10437 : inv02 port map ( Y=>nx10438, A=>nx10430);
   ix10439 : inv02 port map ( Y=>nx10440, A=>nx10430);
   ix10441 : inv01 port map ( Y=>nx10442, A=>gen_23_cmp_BSCmp_op2_16);
   ix10443 : inv02 port map ( Y=>nx10444, A=>nx10442);
   ix10445 : inv02 port map ( Y=>nx10446, A=>nx10442);
   ix10447 : inv02 port map ( Y=>nx10448, A=>nx10442);
   ix10449 : inv02 port map ( Y=>nx10450, A=>nx10442);
   ix10451 : inv02 port map ( Y=>nx10452, A=>nx10442);
   ix10453 : inv01 port map ( Y=>nx10454, A=>gen_22_cmp_BSCmp_op2_16);
   ix10455 : inv02 port map ( Y=>nx10456, A=>nx10454);
   ix10457 : inv02 port map ( Y=>nx10458, A=>nx10454);
   ix10459 : inv02 port map ( Y=>nx10460, A=>nx10454);
   ix10461 : inv02 port map ( Y=>nx10462, A=>nx10454);
   ix10463 : inv02 port map ( Y=>nx10464, A=>nx10454);
   ix10465 : inv01 port map ( Y=>nx10466, A=>gen_21_cmp_BSCmp_op2_16);
   ix10467 : inv02 port map ( Y=>nx10468, A=>nx10466);
   ix10469 : inv02 port map ( Y=>nx10470, A=>nx10466);
   ix10471 : inv02 port map ( Y=>nx10472, A=>nx10466);
   ix10473 : inv02 port map ( Y=>nx10474, A=>nx10466);
   ix10475 : inv02 port map ( Y=>nx10476, A=>nx10466);
   ix10477 : inv01 port map ( Y=>nx10478, A=>gen_20_cmp_BSCmp_op2_16);
   ix10479 : inv02 port map ( Y=>nx10480, A=>nx10478);
   ix10481 : inv02 port map ( Y=>nx10482, A=>nx10478);
   ix10483 : inv02 port map ( Y=>nx10484, A=>nx10478);
   ix10485 : inv02 port map ( Y=>nx10486, A=>nx10478);
   ix10487 : inv02 port map ( Y=>nx10488, A=>nx10478);
   ix10489 : inv01 port map ( Y=>nx10490, A=>gen_19_cmp_BSCmp_op2_16);
   ix10491 : inv02 port map ( Y=>nx10492, A=>nx10490);
   ix10493 : inv02 port map ( Y=>nx10494, A=>nx10490);
   ix10495 : inv02 port map ( Y=>nx10496, A=>nx10490);
   ix10497 : inv02 port map ( Y=>nx10498, A=>nx10490);
   ix10499 : inv02 port map ( Y=>nx10500, A=>nx10490);
   ix10501 : inv01 port map ( Y=>nx10502, A=>gen_18_cmp_BSCmp_op2_16);
   ix10503 : inv02 port map ( Y=>nx10504, A=>nx10502);
   ix10505 : inv02 port map ( Y=>nx10506, A=>nx10502);
   ix10507 : inv02 port map ( Y=>nx10508, A=>nx10502);
   ix10509 : inv02 port map ( Y=>nx10510, A=>nx10502);
   ix10511 : inv02 port map ( Y=>nx10512, A=>nx10502);
   ix10513 : inv01 port map ( Y=>nx10514, A=>gen_17_cmp_BSCmp_op2_16);
   ix10515 : inv02 port map ( Y=>nx10516, A=>nx10514);
   ix10517 : inv02 port map ( Y=>nx10518, A=>nx10514);
   ix10519 : inv02 port map ( Y=>nx10520, A=>nx10514);
   ix10521 : inv02 port map ( Y=>nx10522, A=>nx10514);
   ix10523 : inv02 port map ( Y=>nx10524, A=>nx10514);
   ix10525 : inv01 port map ( Y=>nx10526, A=>gen_16_cmp_BSCmp_op2_16);
   ix10527 : inv02 port map ( Y=>nx10528, A=>nx10526);
   ix10529 : inv02 port map ( Y=>nx10530, A=>nx10526);
   ix10531 : inv02 port map ( Y=>nx10532, A=>nx10526);
   ix10533 : inv02 port map ( Y=>nx10534, A=>nx10526);
   ix10535 : inv02 port map ( Y=>nx10536, A=>nx10526);
   ix10537 : inv01 port map ( Y=>nx10538, A=>gen_15_cmp_BSCmp_op2_16);
   ix10539 : inv02 port map ( Y=>nx10540, A=>nx10538);
   ix10541 : inv02 port map ( Y=>nx10542, A=>nx10538);
   ix10543 : inv02 port map ( Y=>nx10544, A=>nx10538);
   ix10545 : inv02 port map ( Y=>nx10546, A=>nx10538);
   ix10547 : inv02 port map ( Y=>nx10548, A=>nx10538);
   ix10549 : inv01 port map ( Y=>nx10550, A=>gen_14_cmp_BSCmp_op2_16);
   ix10551 : inv02 port map ( Y=>nx10552, A=>nx10550);
   ix10553 : inv02 port map ( Y=>nx10554, A=>nx10550);
   ix10555 : inv02 port map ( Y=>nx10556, A=>nx10550);
   ix10557 : inv02 port map ( Y=>nx10558, A=>nx10550);
   ix10559 : inv02 port map ( Y=>nx10560, A=>nx10550);
   ix10561 : inv01 port map ( Y=>nx10562, A=>gen_13_cmp_BSCmp_op2_16);
   ix10563 : inv02 port map ( Y=>nx10564, A=>nx10562);
   ix10565 : inv02 port map ( Y=>nx10566, A=>nx10562);
   ix10567 : inv02 port map ( Y=>nx10568, A=>nx10562);
   ix10569 : inv02 port map ( Y=>nx10570, A=>nx10562);
   ix10571 : inv02 port map ( Y=>nx10572, A=>nx10562);
   ix10573 : inv01 port map ( Y=>nx10574, A=>gen_12_cmp_BSCmp_op2_16);
   ix10575 : inv02 port map ( Y=>nx10576, A=>nx10574);
   ix10577 : inv02 port map ( Y=>nx10578, A=>nx10574);
   ix10579 : inv02 port map ( Y=>nx10580, A=>nx10574);
   ix10581 : inv02 port map ( Y=>nx10582, A=>nx10574);
   ix10583 : inv02 port map ( Y=>nx10584, A=>nx10574);
   ix10585 : inv01 port map ( Y=>nx10586, A=>gen_11_cmp_BSCmp_op2_16);
   ix10587 : inv02 port map ( Y=>nx10588, A=>nx10586);
   ix10589 : inv02 port map ( Y=>nx10590, A=>nx10586);
   ix10591 : inv02 port map ( Y=>nx10592, A=>nx10586);
   ix10593 : inv02 port map ( Y=>nx10594, A=>nx10586);
   ix10595 : inv02 port map ( Y=>nx10596, A=>nx10586);
   ix10597 : inv01 port map ( Y=>nx10598, A=>gen_10_cmp_BSCmp_op2_16);
   ix10599 : inv02 port map ( Y=>nx10600, A=>nx10598);
   ix10601 : inv02 port map ( Y=>nx10602, A=>nx10598);
   ix10603 : inv02 port map ( Y=>nx10604, A=>nx10598);
   ix10605 : inv02 port map ( Y=>nx10606, A=>nx10598);
   ix10607 : inv02 port map ( Y=>nx10608, A=>nx10598);
   ix10609 : inv01 port map ( Y=>nx10610, A=>gen_9_cmp_BSCmp_op2_16);
   ix10611 : inv02 port map ( Y=>nx10612, A=>nx10610);
   ix10613 : inv02 port map ( Y=>nx10614, A=>nx10610);
   ix10615 : inv02 port map ( Y=>nx10616, A=>nx10610);
   ix10617 : inv02 port map ( Y=>nx10618, A=>nx10610);
   ix10619 : inv02 port map ( Y=>nx10620, A=>nx10610);
   ix10621 : inv01 port map ( Y=>nx10622, A=>gen_8_cmp_BSCmp_op2_16);
   ix10623 : inv02 port map ( Y=>nx10624, A=>nx10622);
   ix10625 : inv02 port map ( Y=>nx10626, A=>nx10622);
   ix10627 : inv02 port map ( Y=>nx10628, A=>nx10622);
   ix10629 : inv02 port map ( Y=>nx10630, A=>nx10622);
   ix10631 : inv02 port map ( Y=>nx10632, A=>nx10622);
   ix10633 : inv01 port map ( Y=>nx10634, A=>gen_7_cmp_BSCmp_op2_16);
   ix10635 : inv02 port map ( Y=>nx10636, A=>nx10634);
   ix10637 : inv02 port map ( Y=>nx10638, A=>nx10634);
   ix10639 : inv02 port map ( Y=>nx10640, A=>nx10634);
   ix10641 : inv02 port map ( Y=>nx10642, A=>nx10634);
   ix10643 : inv02 port map ( Y=>nx10644, A=>nx10634);
   ix10645 : inv01 port map ( Y=>nx10646, A=>gen_6_cmp_BSCmp_op2_16);
   ix10647 : inv02 port map ( Y=>nx10648, A=>nx10646);
   ix10649 : inv02 port map ( Y=>nx10650, A=>nx10646);
   ix10651 : inv02 port map ( Y=>nx10652, A=>nx10646);
   ix10653 : inv02 port map ( Y=>nx10654, A=>nx10646);
   ix10655 : inv02 port map ( Y=>nx10656, A=>nx10646);
   ix10657 : inv01 port map ( Y=>nx10658, A=>gen_5_cmp_BSCmp_op2_16);
   ix10659 : inv02 port map ( Y=>nx10660, A=>nx10658);
   ix10661 : inv02 port map ( Y=>nx10662, A=>nx10658);
   ix10663 : inv02 port map ( Y=>nx10664, A=>nx10658);
   ix10665 : inv02 port map ( Y=>nx10666, A=>nx10658);
   ix10667 : inv02 port map ( Y=>nx10668, A=>nx10658);
   ix10669 : inv01 port map ( Y=>nx10670, A=>gen_4_cmp_BSCmp_op2_16);
   ix10671 : inv02 port map ( Y=>nx10672, A=>nx10670);
   ix10673 : inv02 port map ( Y=>nx10674, A=>nx10670);
   ix10675 : inv02 port map ( Y=>nx10676, A=>nx10670);
   ix10677 : inv02 port map ( Y=>nx10678, A=>nx10670);
   ix10679 : inv02 port map ( Y=>nx10680, A=>nx10670);
   ix10681 : inv01 port map ( Y=>nx10682, A=>gen_3_cmp_BSCmp_op2_16);
   ix10683 : inv02 port map ( Y=>nx10684, A=>nx10682);
   ix10685 : inv02 port map ( Y=>nx10686, A=>nx10682);
   ix10687 : inv02 port map ( Y=>nx10688, A=>nx10682);
   ix10689 : inv02 port map ( Y=>nx10690, A=>nx10682);
   ix10691 : inv02 port map ( Y=>nx10692, A=>nx10682);
   ix10693 : inv01 port map ( Y=>nx10694, A=>gen_2_cmp_BSCmp_op2_16);
   ix10695 : inv02 port map ( Y=>nx10696, A=>nx10694);
   ix10697 : inv02 port map ( Y=>nx10698, A=>nx10694);
   ix10699 : inv02 port map ( Y=>nx10700, A=>nx10694);
   ix10701 : inv02 port map ( Y=>nx10702, A=>nx10694);
   ix10703 : inv02 port map ( Y=>nx10704, A=>nx10694);
   ix10705 : inv01 port map ( Y=>nx10706, A=>gen_1_cmp_BSCmp_op2_16);
   ix10707 : inv02 port map ( Y=>nx10708, A=>nx10706);
   ix10709 : inv02 port map ( Y=>nx10710, A=>nx10706);
   ix10711 : inv02 port map ( Y=>nx10712, A=>nx10706);
   ix10713 : inv02 port map ( Y=>nx10714, A=>nx10706);
   ix10715 : inv02 port map ( Y=>nx10716, A=>nx10706);
   ix10717 : inv01 port map ( Y=>nx10718, A=>gen_0_cmp_BSCmp_op2_16);
   ix10719 : inv02 port map ( Y=>nx10720, A=>nx10718);
   ix10721 : inv02 port map ( Y=>nx10722, A=>nx10718);
   ix10723 : inv02 port map ( Y=>nx10724, A=>nx10718);
   ix10725 : inv02 port map ( Y=>nx10726, A=>nx10718);
   ix10727 : inv02 port map ( Y=>nx10728, A=>nx10718);
   ix10729 : buf02 port map ( Y=>nx10730, A=>nx6);
   ix10731 : buf02 port map ( Y=>nx10732, A=>nx6);
   ix10733 : buf02 port map ( Y=>nx10734, A=>nx6);
   ix10735 : buf02 port map ( Y=>nx10736, A=>nx392);
   ix10737 : buf02 port map ( Y=>nx10738, A=>nx392);
   ix10739 : buf02 port map ( Y=>nx10740, A=>nx392);
   ix10741 : buf02 port map ( Y=>nx10742, A=>nx778);
   ix10743 : buf02 port map ( Y=>nx10744, A=>nx778);
   ix10745 : buf02 port map ( Y=>nx10746, A=>nx778);
   ix10747 : buf02 port map ( Y=>nx10748, A=>nx1164);
   ix10749 : buf02 port map ( Y=>nx10750, A=>nx1164);
   ix10751 : buf02 port map ( Y=>nx10752, A=>nx1164);
   ix10753 : buf02 port map ( Y=>nx10754, A=>nx1550);
   ix10755 : buf02 port map ( Y=>nx10756, A=>nx1550);
   ix10757 : buf02 port map ( Y=>nx10758, A=>nx1550);
   ix10759 : buf02 port map ( Y=>nx10760, A=>nx1936);
   ix10761 : buf02 port map ( Y=>nx10762, A=>nx1936);
   ix10763 : buf02 port map ( Y=>nx10764, A=>nx1936);
   ix10765 : buf02 port map ( Y=>nx10766, A=>nx2322);
   ix10767 : buf02 port map ( Y=>nx10768, A=>nx2322);
   ix10769 : buf02 port map ( Y=>nx10770, A=>nx2322);
   ix10771 : buf02 port map ( Y=>nx10772, A=>nx2708);
   ix10773 : buf02 port map ( Y=>nx10774, A=>nx2708);
   ix10775 : buf02 port map ( Y=>nx10776, A=>nx2708);
   ix10777 : buf02 port map ( Y=>nx10778, A=>nx3094);
   ix10779 : buf02 port map ( Y=>nx10780, A=>nx3094);
   ix10781 : buf02 port map ( Y=>nx10782, A=>nx3094);
   ix10783 : buf02 port map ( Y=>nx10784, A=>nx3480);
   ix10785 : buf02 port map ( Y=>nx10786, A=>nx3480);
   ix10787 : buf02 port map ( Y=>nx10788, A=>nx3480);
   ix10789 : buf02 port map ( Y=>nx10790, A=>nx3866);
   ix10791 : buf02 port map ( Y=>nx10792, A=>nx3866);
   ix10793 : buf02 port map ( Y=>nx10794, A=>nx3866);
   ix10795 : buf02 port map ( Y=>nx10796, A=>nx4252);
   ix10797 : buf02 port map ( Y=>nx10798, A=>nx4252);
   ix10799 : buf02 port map ( Y=>nx10800, A=>nx4252);
   ix10801 : buf02 port map ( Y=>nx10802, A=>nx4638);
   ix10803 : buf02 port map ( Y=>nx10804, A=>nx4638);
   ix10805 : buf02 port map ( Y=>nx10806, A=>nx4638);
   ix10807 : buf02 port map ( Y=>nx10808, A=>nx5024);
   ix10809 : buf02 port map ( Y=>nx10810, A=>nx5024);
   ix10811 : buf02 port map ( Y=>nx10812, A=>nx5024);
   ix10813 : buf02 port map ( Y=>nx10814, A=>nx5410);
   ix10815 : buf02 port map ( Y=>nx10816, A=>nx5410);
   ix10817 : buf02 port map ( Y=>nx10818, A=>nx5410);
   ix10819 : buf02 port map ( Y=>nx10820, A=>nx5796);
   ix10821 : buf02 port map ( Y=>nx10822, A=>nx5796);
   ix10823 : buf02 port map ( Y=>nx10824, A=>nx5796);
   ix10825 : buf02 port map ( Y=>nx10826, A=>nx6182);
   ix10827 : buf02 port map ( Y=>nx10828, A=>nx6182);
   ix10829 : buf02 port map ( Y=>nx10830, A=>nx6182);
   ix10831 : buf02 port map ( Y=>nx10832, A=>nx6568);
   ix10833 : buf02 port map ( Y=>nx10834, A=>nx6568);
   ix10835 : buf02 port map ( Y=>nx10836, A=>nx6568);
   ix10837 : buf02 port map ( Y=>nx10838, A=>nx6954);
   ix10839 : buf02 port map ( Y=>nx10840, A=>nx6954);
   ix10841 : buf02 port map ( Y=>nx10842, A=>nx6954);
   ix10843 : buf02 port map ( Y=>nx10844, A=>nx7340);
   ix10845 : buf02 port map ( Y=>nx10846, A=>nx7340);
   ix10847 : buf02 port map ( Y=>nx10848, A=>nx7340);
   ix10849 : buf02 port map ( Y=>nx10850, A=>nx7726);
   ix10851 : buf02 port map ( Y=>nx10852, A=>nx7726);
   ix10853 : buf02 port map ( Y=>nx10854, A=>nx7726);
   ix10855 : buf02 port map ( Y=>nx10856, A=>nx8112);
   ix10857 : buf02 port map ( Y=>nx10858, A=>nx8112);
   ix10859 : buf02 port map ( Y=>nx10860, A=>nx8112);
   ix10861 : buf02 port map ( Y=>nx10862, A=>nx8498);
   ix10863 : buf02 port map ( Y=>nx10864, A=>nx8498);
   ix10865 : buf02 port map ( Y=>nx10866, A=>nx8498);
   ix10867 : buf02 port map ( Y=>nx10868, A=>nx8884);
   ix10869 : buf02 port map ( Y=>nx10870, A=>nx8884);
   ix10871 : buf02 port map ( Y=>nx10872, A=>nx8884);
   ix10873 : buf02 port map ( Y=>nx10874, A=>nx9270);
   ix10875 : buf02 port map ( Y=>nx10876, A=>nx9270);
   ix10877 : buf02 port map ( Y=>nx10878, A=>nx9270);
   ix10879 : inv02 port map ( Y=>nx10880, A=>done);
   ix10881 : inv02 port map ( Y=>nx10882, A=>nx11934);
   ix10883 : inv02 port map ( Y=>nx10884, A=>nx11934);
   ix10885 : inv02 port map ( Y=>nx10886, A=>nx11934);
   ix10889 : inv02 port map ( Y=>nx10890, A=>nx10888);
   ix10891 : inv02 port map ( Y=>nx10892, A=>nx10888);
   ix10893 : inv02 port map ( Y=>nx10894, A=>nx10888);
   ix10895 : inv04 port map ( Y=>nx10896, A=>gen_0_cmp_pMux_1);
   ix10897 : inv04 port map ( Y=>nx10898, A=>gen_0_cmp_pMux_1);
   ix10899 : inv04 port map ( Y=>nx10900, A=>gen_0_cmp_pMux_1);
   ix10901 : inv04 port map ( Y=>nx10902, A=>gen_0_cmp_pMux_1);
   ix10905 : inv02 port map ( Y=>nx10906, A=>nx10904);
   ix10907 : inv02 port map ( Y=>nx10908, A=>nx10904);
   ix10909 : inv02 port map ( Y=>nx10910, A=>nx10904);
   ix10913 : inv02 port map ( Y=>nx10914, A=>nx10912);
   ix10915 : inv02 port map ( Y=>nx10916, A=>nx10912);
   ix10917 : inv02 port map ( Y=>nx10918, A=>nx10912);
   ix10921 : inv02 port map ( Y=>nx10922, A=>nx10920);
   ix10923 : inv02 port map ( Y=>nx10924, A=>nx10920);
   ix10925 : inv02 port map ( Y=>nx10926, A=>nx10920);
   ix10929 : inv02 port map ( Y=>nx10930, A=>nx10928);
   ix10931 : inv02 port map ( Y=>nx10932, A=>nx10928);
   ix10933 : inv02 port map ( Y=>nx10934, A=>nx10928);
   ix10935 : inv04 port map ( Y=>nx10936, A=>gen_1_cmp_pMux_1);
   ix10937 : inv04 port map ( Y=>nx10938, A=>gen_1_cmp_pMux_1);
   ix10939 : inv04 port map ( Y=>nx10940, A=>gen_1_cmp_pMux_1);
   ix10941 : inv04 port map ( Y=>nx10942, A=>gen_1_cmp_pMux_1);
   ix10945 : inv02 port map ( Y=>nx10946, A=>nx10944);
   ix10947 : inv02 port map ( Y=>nx10948, A=>nx10944);
   ix10949 : inv02 port map ( Y=>nx10950, A=>nx10944);
   ix10953 : inv02 port map ( Y=>nx10954, A=>nx10952);
   ix10955 : inv02 port map ( Y=>nx10956, A=>nx10952);
   ix10957 : inv02 port map ( Y=>nx10958, A=>nx10952);
   ix10961 : inv02 port map ( Y=>nx10962, A=>nx10960);
   ix10963 : inv02 port map ( Y=>nx10964, A=>nx10960);
   ix10965 : inv02 port map ( Y=>nx10966, A=>nx10960);
   ix10969 : inv02 port map ( Y=>nx10970, A=>nx10968);
   ix10971 : inv02 port map ( Y=>nx10972, A=>nx10968);
   ix10973 : inv02 port map ( Y=>nx10974, A=>nx10968);
   ix10975 : inv04 port map ( Y=>nx10976, A=>gen_2_cmp_pMux_1);
   ix10977 : inv04 port map ( Y=>nx10978, A=>gen_2_cmp_pMux_1);
   ix10979 : inv04 port map ( Y=>nx10980, A=>gen_2_cmp_pMux_1);
   ix10981 : inv04 port map ( Y=>nx10982, A=>gen_2_cmp_pMux_1);
   ix10985 : inv02 port map ( Y=>nx10986, A=>nx10984);
   ix10987 : inv02 port map ( Y=>nx10988, A=>nx10984);
   ix10989 : inv02 port map ( Y=>nx10990, A=>nx10984);
   ix10993 : inv02 port map ( Y=>nx10994, A=>nx10992);
   ix10995 : inv02 port map ( Y=>nx10996, A=>nx10992);
   ix10997 : inv02 port map ( Y=>nx10998, A=>nx10992);
   ix11001 : inv02 port map ( Y=>nx11002, A=>nx11000);
   ix11003 : inv02 port map ( Y=>nx11004, A=>nx11000);
   ix11005 : inv02 port map ( Y=>nx11006, A=>nx11000);
   ix11009 : inv02 port map ( Y=>nx11010, A=>nx11008);
   ix11011 : inv02 port map ( Y=>nx11012, A=>nx11008);
   ix11013 : inv02 port map ( Y=>nx11014, A=>nx11008);
   ix11015 : inv04 port map ( Y=>nx11016, A=>gen_3_cmp_pMux_1);
   ix11017 : inv04 port map ( Y=>nx11018, A=>gen_3_cmp_pMux_1);
   ix11019 : inv04 port map ( Y=>nx11020, A=>gen_3_cmp_pMux_1);
   ix11021 : inv04 port map ( Y=>nx11022, A=>gen_3_cmp_pMux_1);
   ix11025 : inv02 port map ( Y=>nx11026, A=>nx11024);
   ix11027 : inv02 port map ( Y=>nx11028, A=>nx11024);
   ix11029 : inv02 port map ( Y=>nx11030, A=>nx11024);
   ix11033 : inv02 port map ( Y=>nx11034, A=>nx11032);
   ix11035 : inv02 port map ( Y=>nx11036, A=>nx11032);
   ix11037 : inv02 port map ( Y=>nx11038, A=>nx11032);
   ix11041 : inv02 port map ( Y=>nx11042, A=>nx11040);
   ix11043 : inv02 port map ( Y=>nx11044, A=>nx11040);
   ix11045 : inv02 port map ( Y=>nx11046, A=>nx11040);
   ix11049 : inv02 port map ( Y=>nx11050, A=>nx11048);
   ix11051 : inv02 port map ( Y=>nx11052, A=>nx11048);
   ix11053 : inv02 port map ( Y=>nx11054, A=>nx11048);
   ix11055 : inv04 port map ( Y=>nx11056, A=>gen_4_cmp_pMux_1);
   ix11057 : inv04 port map ( Y=>nx11058, A=>gen_4_cmp_pMux_1);
   ix11059 : inv04 port map ( Y=>nx11060, A=>gen_4_cmp_pMux_1);
   ix11061 : inv04 port map ( Y=>nx11062, A=>gen_4_cmp_pMux_1);
   ix11065 : inv02 port map ( Y=>nx11066, A=>nx11064);
   ix11067 : inv02 port map ( Y=>nx11068, A=>nx11064);
   ix11069 : inv02 port map ( Y=>nx11070, A=>nx11064);
   ix11073 : inv02 port map ( Y=>nx11074, A=>nx11072);
   ix11075 : inv02 port map ( Y=>nx11076, A=>nx11072);
   ix11077 : inv02 port map ( Y=>nx11078, A=>nx11072);
   ix11081 : inv02 port map ( Y=>nx11082, A=>nx11080);
   ix11083 : inv02 port map ( Y=>nx11084, A=>nx11080);
   ix11085 : inv02 port map ( Y=>nx11086, A=>nx11080);
   ix11089 : inv02 port map ( Y=>nx11090, A=>nx11088);
   ix11091 : inv02 port map ( Y=>nx11092, A=>nx11088);
   ix11093 : inv02 port map ( Y=>nx11094, A=>nx11088);
   ix11095 : inv04 port map ( Y=>nx11096, A=>gen_5_cmp_pMux_1);
   ix11097 : inv04 port map ( Y=>nx11098, A=>gen_5_cmp_pMux_1);
   ix11099 : inv04 port map ( Y=>nx11100, A=>gen_5_cmp_pMux_1);
   ix11101 : inv04 port map ( Y=>nx11102, A=>gen_5_cmp_pMux_1);
   ix11105 : inv02 port map ( Y=>nx11106, A=>nx11104);
   ix11107 : inv02 port map ( Y=>nx11108, A=>nx11104);
   ix11109 : inv02 port map ( Y=>nx11110, A=>nx11104);
   ix11113 : inv02 port map ( Y=>nx11114, A=>nx11112);
   ix11115 : inv02 port map ( Y=>nx11116, A=>nx11112);
   ix11117 : inv02 port map ( Y=>nx11118, A=>nx11112);
   ix11121 : inv02 port map ( Y=>nx11122, A=>nx11120);
   ix11123 : inv02 port map ( Y=>nx11124, A=>nx11120);
   ix11125 : inv02 port map ( Y=>nx11126, A=>nx11120);
   ix11129 : inv02 port map ( Y=>nx11130, A=>nx11128);
   ix11131 : inv02 port map ( Y=>nx11132, A=>nx11128);
   ix11133 : inv02 port map ( Y=>nx11134, A=>nx11128);
   ix11135 : inv04 port map ( Y=>nx11136, A=>gen_6_cmp_pMux_1);
   ix11137 : inv04 port map ( Y=>nx11138, A=>gen_6_cmp_pMux_1);
   ix11139 : inv04 port map ( Y=>nx11140, A=>gen_6_cmp_pMux_1);
   ix11141 : inv04 port map ( Y=>nx11142, A=>gen_6_cmp_pMux_1);
   ix11145 : inv02 port map ( Y=>nx11146, A=>nx11144);
   ix11147 : inv02 port map ( Y=>nx11148, A=>nx11144);
   ix11149 : inv02 port map ( Y=>nx11150, A=>nx11144);
   ix11153 : inv02 port map ( Y=>nx11154, A=>nx11152);
   ix11155 : inv02 port map ( Y=>nx11156, A=>nx11152);
   ix11157 : inv02 port map ( Y=>nx11158, A=>nx11152);
   ix11161 : inv02 port map ( Y=>nx11162, A=>nx11160);
   ix11163 : inv02 port map ( Y=>nx11164, A=>nx11160);
   ix11165 : inv02 port map ( Y=>nx11166, A=>nx11160);
   ix11169 : inv02 port map ( Y=>nx11170, A=>nx11168);
   ix11171 : inv02 port map ( Y=>nx11172, A=>nx11168);
   ix11173 : inv02 port map ( Y=>nx11174, A=>nx11168);
   ix11175 : inv04 port map ( Y=>nx11176, A=>gen_7_cmp_pMux_1);
   ix11177 : inv04 port map ( Y=>nx11178, A=>gen_7_cmp_pMux_1);
   ix11179 : inv04 port map ( Y=>nx11180, A=>gen_7_cmp_pMux_1);
   ix11181 : inv04 port map ( Y=>nx11182, A=>gen_7_cmp_pMux_1);
   ix11185 : inv02 port map ( Y=>nx11186, A=>nx11184);
   ix11187 : inv02 port map ( Y=>nx11188, A=>nx11184);
   ix11189 : inv02 port map ( Y=>nx11190, A=>nx11184);
   ix11193 : inv02 port map ( Y=>nx11194, A=>nx11192);
   ix11195 : inv02 port map ( Y=>nx11196, A=>nx11192);
   ix11197 : inv02 port map ( Y=>nx11198, A=>nx11192);
   ix11201 : inv02 port map ( Y=>nx11202, A=>nx11200);
   ix11203 : inv02 port map ( Y=>nx11204, A=>nx11200);
   ix11205 : inv02 port map ( Y=>nx11206, A=>nx11200);
   ix11209 : inv02 port map ( Y=>nx11210, A=>nx11208);
   ix11211 : inv02 port map ( Y=>nx11212, A=>nx11208);
   ix11213 : inv02 port map ( Y=>nx11214, A=>nx11208);
   ix11215 : inv04 port map ( Y=>nx11216, A=>gen_8_cmp_pMux_1);
   ix11217 : inv04 port map ( Y=>nx11218, A=>gen_8_cmp_pMux_1);
   ix11219 : inv04 port map ( Y=>nx11220, A=>gen_8_cmp_pMux_1);
   ix11221 : inv04 port map ( Y=>nx11222, A=>gen_8_cmp_pMux_1);
   ix11225 : inv02 port map ( Y=>nx11226, A=>nx11224);
   ix11227 : inv02 port map ( Y=>nx11228, A=>nx11224);
   ix11229 : inv02 port map ( Y=>nx11230, A=>nx11224);
   ix11233 : inv02 port map ( Y=>nx11234, A=>nx11232);
   ix11235 : inv02 port map ( Y=>nx11236, A=>nx11232);
   ix11237 : inv02 port map ( Y=>nx11238, A=>nx11232);
   ix11241 : inv02 port map ( Y=>nx11242, A=>nx11240);
   ix11243 : inv02 port map ( Y=>nx11244, A=>nx11240);
   ix11245 : inv02 port map ( Y=>nx11246, A=>nx11240);
   ix11249 : inv02 port map ( Y=>nx11250, A=>nx11248);
   ix11251 : inv02 port map ( Y=>nx11252, A=>nx11248);
   ix11253 : inv02 port map ( Y=>nx11254, A=>nx11248);
   ix11255 : inv04 port map ( Y=>nx11256, A=>gen_9_cmp_pMux_1);
   ix11257 : inv04 port map ( Y=>nx11258, A=>gen_9_cmp_pMux_1);
   ix11259 : inv04 port map ( Y=>nx11260, A=>gen_9_cmp_pMux_1);
   ix11261 : inv04 port map ( Y=>nx11262, A=>gen_9_cmp_pMux_1);
   ix11265 : inv02 port map ( Y=>nx11266, A=>nx11264);
   ix11267 : inv02 port map ( Y=>nx11268, A=>nx11264);
   ix11269 : inv02 port map ( Y=>nx11270, A=>nx11264);
   ix11273 : inv02 port map ( Y=>nx11274, A=>nx11272);
   ix11275 : inv02 port map ( Y=>nx11276, A=>nx11272);
   ix11277 : inv02 port map ( Y=>nx11278, A=>nx11272);
   ix11281 : inv02 port map ( Y=>nx11282, A=>nx11280);
   ix11283 : inv02 port map ( Y=>nx11284, A=>nx11280);
   ix11285 : inv02 port map ( Y=>nx11286, A=>nx11280);
   ix11289 : inv02 port map ( Y=>nx11290, A=>nx11288);
   ix11291 : inv02 port map ( Y=>nx11292, A=>nx11288);
   ix11293 : inv02 port map ( Y=>nx11294, A=>nx11288);
   ix11295 : inv04 port map ( Y=>nx11296, A=>gen_10_cmp_pMux_1);
   ix11297 : inv04 port map ( Y=>nx11298, A=>gen_10_cmp_pMux_1);
   ix11299 : inv04 port map ( Y=>nx11300, A=>gen_10_cmp_pMux_1);
   ix11301 : inv04 port map ( Y=>nx11302, A=>gen_10_cmp_pMux_1);
   ix11305 : inv02 port map ( Y=>nx11306, A=>nx11304);
   ix11307 : inv02 port map ( Y=>nx11308, A=>nx11304);
   ix11309 : inv02 port map ( Y=>nx11310, A=>nx11304);
   ix11313 : inv02 port map ( Y=>nx11314, A=>nx11312);
   ix11315 : inv02 port map ( Y=>nx11316, A=>nx11312);
   ix11317 : inv02 port map ( Y=>nx11318, A=>nx11312);
   ix11321 : inv02 port map ( Y=>nx11322, A=>nx11320);
   ix11323 : inv02 port map ( Y=>nx11324, A=>nx11320);
   ix11325 : inv02 port map ( Y=>nx11326, A=>nx11320);
   ix11329 : inv02 port map ( Y=>nx11330, A=>nx11328);
   ix11331 : inv02 port map ( Y=>nx11332, A=>nx11328);
   ix11333 : inv02 port map ( Y=>nx11334, A=>nx11328);
   ix11335 : inv04 port map ( Y=>nx11336, A=>gen_11_cmp_pMux_1);
   ix11337 : inv04 port map ( Y=>nx11338, A=>gen_11_cmp_pMux_1);
   ix11339 : inv04 port map ( Y=>nx11340, A=>gen_11_cmp_pMux_1);
   ix11341 : inv04 port map ( Y=>nx11342, A=>gen_11_cmp_pMux_1);
   ix11345 : inv02 port map ( Y=>nx11346, A=>nx11344);
   ix11347 : inv02 port map ( Y=>nx11348, A=>nx11344);
   ix11349 : inv02 port map ( Y=>nx11350, A=>nx11344);
   ix11353 : inv02 port map ( Y=>nx11354, A=>nx11352);
   ix11355 : inv02 port map ( Y=>nx11356, A=>nx11352);
   ix11357 : inv02 port map ( Y=>nx11358, A=>nx11352);
   ix11361 : inv02 port map ( Y=>nx11362, A=>nx11360);
   ix11363 : inv02 port map ( Y=>nx11364, A=>nx11360);
   ix11365 : inv02 port map ( Y=>nx11366, A=>nx11360);
   ix11369 : inv02 port map ( Y=>nx11370, A=>nx11368);
   ix11371 : inv02 port map ( Y=>nx11372, A=>nx11368);
   ix11373 : inv02 port map ( Y=>nx11374, A=>nx11368);
   ix11375 : inv04 port map ( Y=>nx11376, A=>gen_12_cmp_pMux_1);
   ix11377 : inv04 port map ( Y=>nx11378, A=>gen_12_cmp_pMux_1);
   ix11379 : inv04 port map ( Y=>nx11380, A=>gen_12_cmp_pMux_1);
   ix11381 : inv04 port map ( Y=>nx11382, A=>gen_12_cmp_pMux_1);
   ix11385 : inv02 port map ( Y=>nx11386, A=>nx11384);
   ix11387 : inv02 port map ( Y=>nx11388, A=>nx11384);
   ix11389 : inv02 port map ( Y=>nx11390, A=>nx11384);
   ix11393 : inv02 port map ( Y=>nx11394, A=>nx11392);
   ix11395 : inv02 port map ( Y=>nx11396, A=>nx11392);
   ix11397 : inv02 port map ( Y=>nx11398, A=>nx11392);
   ix11401 : inv02 port map ( Y=>nx11402, A=>nx11400);
   ix11403 : inv02 port map ( Y=>nx11404, A=>nx11400);
   ix11405 : inv02 port map ( Y=>nx11406, A=>nx11400);
   ix11409 : inv02 port map ( Y=>nx11410, A=>nx11408);
   ix11411 : inv02 port map ( Y=>nx11412, A=>nx11408);
   ix11413 : inv02 port map ( Y=>nx11414, A=>nx11408);
   ix11415 : inv04 port map ( Y=>nx11416, A=>gen_13_cmp_pMux_1);
   ix11417 : inv04 port map ( Y=>nx11418, A=>gen_13_cmp_pMux_1);
   ix11419 : inv04 port map ( Y=>nx11420, A=>gen_13_cmp_pMux_1);
   ix11421 : inv04 port map ( Y=>nx11422, A=>gen_13_cmp_pMux_1);
   ix11425 : inv02 port map ( Y=>nx11426, A=>nx11424);
   ix11427 : inv02 port map ( Y=>nx11428, A=>nx11424);
   ix11429 : inv02 port map ( Y=>nx11430, A=>nx11424);
   ix11433 : inv02 port map ( Y=>nx11434, A=>nx11432);
   ix11435 : inv02 port map ( Y=>nx11436, A=>nx11432);
   ix11437 : inv02 port map ( Y=>nx11438, A=>nx11432);
   ix11441 : inv02 port map ( Y=>nx11442, A=>nx11440);
   ix11443 : inv02 port map ( Y=>nx11444, A=>nx11440);
   ix11445 : inv02 port map ( Y=>nx11446, A=>nx11440);
   ix11449 : inv02 port map ( Y=>nx11450, A=>nx11448);
   ix11451 : inv02 port map ( Y=>nx11452, A=>nx11448);
   ix11453 : inv02 port map ( Y=>nx11454, A=>nx11448);
   ix11455 : inv04 port map ( Y=>nx11456, A=>gen_14_cmp_pMux_1);
   ix11457 : inv04 port map ( Y=>nx11458, A=>gen_14_cmp_pMux_1);
   ix11459 : inv04 port map ( Y=>nx11460, A=>gen_14_cmp_pMux_1);
   ix11461 : inv04 port map ( Y=>nx11462, A=>gen_14_cmp_pMux_1);
   ix11465 : inv02 port map ( Y=>nx11466, A=>nx11464);
   ix11467 : inv02 port map ( Y=>nx11468, A=>nx11464);
   ix11469 : inv02 port map ( Y=>nx11470, A=>nx11464);
   ix11473 : inv02 port map ( Y=>nx11474, A=>nx11472);
   ix11475 : inv02 port map ( Y=>nx11476, A=>nx11472);
   ix11477 : inv02 port map ( Y=>nx11478, A=>nx11472);
   ix11481 : inv02 port map ( Y=>nx11482, A=>nx11480);
   ix11483 : inv02 port map ( Y=>nx11484, A=>nx11480);
   ix11485 : inv02 port map ( Y=>nx11486, A=>nx11480);
   ix11489 : inv02 port map ( Y=>nx11490, A=>nx11488);
   ix11491 : inv02 port map ( Y=>nx11492, A=>nx11488);
   ix11493 : inv02 port map ( Y=>nx11494, A=>nx11488);
   ix11495 : inv04 port map ( Y=>nx11496, A=>gen_15_cmp_pMux_1);
   ix11497 : inv04 port map ( Y=>nx11498, A=>gen_15_cmp_pMux_1);
   ix11499 : inv04 port map ( Y=>nx11500, A=>gen_15_cmp_pMux_1);
   ix11501 : inv04 port map ( Y=>nx11502, A=>gen_15_cmp_pMux_1);
   ix11505 : inv02 port map ( Y=>nx11506, A=>nx11504);
   ix11507 : inv02 port map ( Y=>nx11508, A=>nx11504);
   ix11509 : inv02 port map ( Y=>nx11510, A=>nx11504);
   ix11513 : inv02 port map ( Y=>nx11514, A=>nx11512);
   ix11515 : inv02 port map ( Y=>nx11516, A=>nx11512);
   ix11517 : inv02 port map ( Y=>nx11518, A=>nx11512);
   ix11521 : inv02 port map ( Y=>nx11522, A=>nx11520);
   ix11523 : inv02 port map ( Y=>nx11524, A=>nx11520);
   ix11525 : inv02 port map ( Y=>nx11526, A=>nx11520);
   ix11529 : inv02 port map ( Y=>nx11530, A=>nx11528);
   ix11531 : inv02 port map ( Y=>nx11532, A=>nx11528);
   ix11533 : inv02 port map ( Y=>nx11534, A=>nx11528);
   ix11535 : inv04 port map ( Y=>nx11536, A=>gen_16_cmp_pMux_1);
   ix11537 : inv04 port map ( Y=>nx11538, A=>gen_16_cmp_pMux_1);
   ix11539 : inv04 port map ( Y=>nx11540, A=>gen_16_cmp_pMux_1);
   ix11541 : inv04 port map ( Y=>nx11542, A=>gen_16_cmp_pMux_1);
   ix11545 : inv02 port map ( Y=>nx11546, A=>nx11544);
   ix11547 : inv02 port map ( Y=>nx11548, A=>nx11544);
   ix11549 : inv02 port map ( Y=>nx11550, A=>nx11544);
   ix11553 : inv02 port map ( Y=>nx11554, A=>nx11552);
   ix11555 : inv02 port map ( Y=>nx11556, A=>nx11552);
   ix11557 : inv02 port map ( Y=>nx11558, A=>nx11552);
   ix11561 : inv02 port map ( Y=>nx11562, A=>nx11560);
   ix11563 : inv02 port map ( Y=>nx11564, A=>nx11560);
   ix11565 : inv02 port map ( Y=>nx11566, A=>nx11560);
   ix11569 : inv02 port map ( Y=>nx11570, A=>nx11568);
   ix11571 : inv02 port map ( Y=>nx11572, A=>nx11568);
   ix11573 : inv02 port map ( Y=>nx11574, A=>nx11568);
   ix11575 : inv04 port map ( Y=>nx11576, A=>gen_17_cmp_pMux_1);
   ix11577 : inv04 port map ( Y=>nx11578, A=>gen_17_cmp_pMux_1);
   ix11579 : inv04 port map ( Y=>nx11580, A=>gen_17_cmp_pMux_1);
   ix11581 : inv04 port map ( Y=>nx11582, A=>gen_17_cmp_pMux_1);
   ix11585 : inv02 port map ( Y=>nx11586, A=>nx11584);
   ix11587 : inv02 port map ( Y=>nx11588, A=>nx11584);
   ix11589 : inv02 port map ( Y=>nx11590, A=>nx11584);
   ix11593 : inv02 port map ( Y=>nx11594, A=>nx11592);
   ix11595 : inv02 port map ( Y=>nx11596, A=>nx11592);
   ix11597 : inv02 port map ( Y=>nx11598, A=>nx11592);
   ix11601 : inv02 port map ( Y=>nx11602, A=>nx11600);
   ix11603 : inv02 port map ( Y=>nx11604, A=>nx11600);
   ix11605 : inv02 port map ( Y=>nx11606, A=>nx11600);
   ix11609 : inv02 port map ( Y=>nx11610, A=>nx11608);
   ix11611 : inv02 port map ( Y=>nx11612, A=>nx11608);
   ix11613 : inv02 port map ( Y=>nx11614, A=>nx11608);
   ix11615 : inv04 port map ( Y=>nx11616, A=>gen_18_cmp_pMux_1);
   ix11617 : inv04 port map ( Y=>nx11618, A=>gen_18_cmp_pMux_1);
   ix11619 : inv04 port map ( Y=>nx11620, A=>gen_18_cmp_pMux_1);
   ix11621 : inv04 port map ( Y=>nx11622, A=>gen_18_cmp_pMux_1);
   ix11625 : inv02 port map ( Y=>nx11626, A=>nx11624);
   ix11627 : inv02 port map ( Y=>nx11628, A=>nx11624);
   ix11629 : inv02 port map ( Y=>nx11630, A=>nx11624);
   ix11633 : inv02 port map ( Y=>nx11634, A=>nx11632);
   ix11635 : inv02 port map ( Y=>nx11636, A=>nx11632);
   ix11637 : inv02 port map ( Y=>nx11638, A=>nx11632);
   ix11641 : inv02 port map ( Y=>nx11642, A=>nx11640);
   ix11643 : inv02 port map ( Y=>nx11644, A=>nx11640);
   ix11645 : inv02 port map ( Y=>nx11646, A=>nx11640);
   ix11649 : inv02 port map ( Y=>nx11650, A=>nx11648);
   ix11651 : inv02 port map ( Y=>nx11652, A=>nx11648);
   ix11653 : inv02 port map ( Y=>nx11654, A=>nx11648);
   ix11655 : inv04 port map ( Y=>nx11656, A=>gen_19_cmp_pMux_1);
   ix11657 : inv04 port map ( Y=>nx11658, A=>gen_19_cmp_pMux_1);
   ix11659 : inv04 port map ( Y=>nx11660, A=>gen_19_cmp_pMux_1);
   ix11661 : inv04 port map ( Y=>nx11662, A=>gen_19_cmp_pMux_1);
   ix11665 : inv02 port map ( Y=>nx11666, A=>nx11664);
   ix11667 : inv02 port map ( Y=>nx11668, A=>nx11664);
   ix11669 : inv02 port map ( Y=>nx11670, A=>nx11664);
   ix11673 : inv02 port map ( Y=>nx11674, A=>nx11672);
   ix11675 : inv02 port map ( Y=>nx11676, A=>nx11672);
   ix11677 : inv02 port map ( Y=>nx11678, A=>nx11672);
   ix11681 : inv02 port map ( Y=>nx11682, A=>nx11680);
   ix11683 : inv02 port map ( Y=>nx11684, A=>nx11680);
   ix11685 : inv02 port map ( Y=>nx11686, A=>nx11680);
   ix11689 : inv02 port map ( Y=>nx11690, A=>nx11688);
   ix11691 : inv02 port map ( Y=>nx11692, A=>nx11688);
   ix11693 : inv02 port map ( Y=>nx11694, A=>nx11688);
   ix11695 : inv04 port map ( Y=>nx11696, A=>gen_20_cmp_pMux_1);
   ix11697 : inv04 port map ( Y=>nx11698, A=>gen_20_cmp_pMux_1);
   ix11699 : inv04 port map ( Y=>nx11700, A=>gen_20_cmp_pMux_1);
   ix11701 : inv04 port map ( Y=>nx11702, A=>gen_20_cmp_pMux_1);
   ix11705 : inv02 port map ( Y=>nx11706, A=>nx11704);
   ix11707 : inv02 port map ( Y=>nx11708, A=>nx11704);
   ix11709 : inv02 port map ( Y=>nx11710, A=>nx11704);
   ix11713 : inv02 port map ( Y=>nx11714, A=>nx11712);
   ix11715 : inv02 port map ( Y=>nx11716, A=>nx11712);
   ix11717 : inv02 port map ( Y=>nx11718, A=>nx11712);
   ix11721 : inv02 port map ( Y=>nx11722, A=>nx11720);
   ix11723 : inv02 port map ( Y=>nx11724, A=>nx11720);
   ix11725 : inv02 port map ( Y=>nx11726, A=>nx11720);
   ix11729 : inv02 port map ( Y=>nx11730, A=>nx11728);
   ix11731 : inv02 port map ( Y=>nx11732, A=>nx11728);
   ix11733 : inv02 port map ( Y=>nx11734, A=>nx11728);
   ix11735 : inv04 port map ( Y=>nx11736, A=>gen_21_cmp_pMux_1);
   ix11737 : inv04 port map ( Y=>nx11738, A=>gen_21_cmp_pMux_1);
   ix11739 : inv04 port map ( Y=>nx11740, A=>gen_21_cmp_pMux_1);
   ix11741 : inv04 port map ( Y=>nx11742, A=>gen_21_cmp_pMux_1);
   ix11745 : inv02 port map ( Y=>nx11746, A=>nx11744);
   ix11747 : inv02 port map ( Y=>nx11748, A=>nx11744);
   ix11749 : inv02 port map ( Y=>nx11750, A=>nx11744);
   ix11753 : inv02 port map ( Y=>nx11754, A=>nx11752);
   ix11755 : inv02 port map ( Y=>nx11756, A=>nx11752);
   ix11757 : inv02 port map ( Y=>nx11758, A=>nx11752);
   ix11761 : inv02 port map ( Y=>nx11762, A=>nx11760);
   ix11763 : inv02 port map ( Y=>nx11764, A=>nx11760);
   ix11765 : inv02 port map ( Y=>nx11766, A=>nx11760);
   ix11769 : inv02 port map ( Y=>nx11770, A=>nx11768);
   ix11771 : inv02 port map ( Y=>nx11772, A=>nx11768);
   ix11773 : inv02 port map ( Y=>nx11774, A=>nx11768);
   ix11775 : inv04 port map ( Y=>nx11776, A=>gen_22_cmp_pMux_1);
   ix11777 : inv04 port map ( Y=>nx11778, A=>gen_22_cmp_pMux_1);
   ix11779 : inv04 port map ( Y=>nx11780, A=>gen_22_cmp_pMux_1);
   ix11781 : inv04 port map ( Y=>nx11782, A=>gen_22_cmp_pMux_1);
   ix11785 : inv02 port map ( Y=>nx11786, A=>nx11784);
   ix11787 : inv02 port map ( Y=>nx11788, A=>nx11784);
   ix11789 : inv02 port map ( Y=>nx11790, A=>nx11784);
   ix11793 : inv02 port map ( Y=>nx11794, A=>nx11792);
   ix11795 : inv02 port map ( Y=>nx11796, A=>nx11792);
   ix11797 : inv02 port map ( Y=>nx11798, A=>nx11792);
   ix11801 : inv02 port map ( Y=>nx11802, A=>nx11800);
   ix11803 : inv02 port map ( Y=>nx11804, A=>nx11800);
   ix11805 : inv02 port map ( Y=>nx11806, A=>nx11800);
   ix11809 : inv02 port map ( Y=>nx11810, A=>nx11808);
   ix11811 : inv02 port map ( Y=>nx11812, A=>nx11808);
   ix11813 : inv02 port map ( Y=>nx11814, A=>nx11808);
   ix11815 : inv04 port map ( Y=>nx11816, A=>gen_23_cmp_pMux_1);
   ix11817 : inv04 port map ( Y=>nx11818, A=>gen_23_cmp_pMux_1);
   ix11819 : inv04 port map ( Y=>nx11820, A=>gen_23_cmp_pMux_1);
   ix11821 : inv04 port map ( Y=>nx11822, A=>gen_23_cmp_pMux_1);
   ix11825 : inv02 port map ( Y=>nx11826, A=>nx11824);
   ix11827 : inv02 port map ( Y=>nx11828, A=>nx11824);
   ix11829 : inv02 port map ( Y=>nx11830, A=>nx11824);
   ix11833 : inv02 port map ( Y=>nx11834, A=>nx11832);
   ix11835 : inv02 port map ( Y=>nx11836, A=>nx11832);
   ix11837 : inv02 port map ( Y=>nx11838, A=>nx11832);
   ix11841 : inv02 port map ( Y=>nx11842, A=>nx11840);
   ix11843 : inv02 port map ( Y=>nx11844, A=>nx11840);
   ix11845 : inv02 port map ( Y=>nx11846, A=>nx11840);
   ix11849 : inv02 port map ( Y=>nx11850, A=>nx11848);
   ix11851 : inv02 port map ( Y=>nx11852, A=>nx11848);
   ix11853 : inv02 port map ( Y=>nx11854, A=>nx11848);
   ix11855 : inv04 port map ( Y=>nx11856, A=>gen_24_cmp_pMux_1);
   ix11857 : inv04 port map ( Y=>nx11858, A=>gen_24_cmp_pMux_1);
   ix11859 : inv04 port map ( Y=>nx11860, A=>gen_24_cmp_pMux_1);
   ix11861 : inv04 port map ( Y=>nx11862, A=>gen_24_cmp_pMux_1);
   ix11865 : inv02 port map ( Y=>nx11866, A=>nx11864);
   ix11867 : inv02 port map ( Y=>nx11868, A=>nx11864);
   ix11869 : inv02 port map ( Y=>nx11870, A=>nx11864);
   ix11873 : inv02 port map ( Y=>nx11874, A=>nx11872);
   ix11875 : inv02 port map ( Y=>nx11876, A=>nx11872);
   ix11877 : inv02 port map ( Y=>nx11878, A=>nx11872);
   ix11881 : inv02 port map ( Y=>nx11882, A=>nx11880);
   ix11883 : inv02 port map ( Y=>nx11884, A=>nx11880);
   ix11885 : inv02 port map ( Y=>nx11886, A=>nx11880);
   ix3760 : nor02_2x port map ( Y=>nx10888, A0=>nx3769, A1=>gen_0_cmp_pMux_0
   );
   ix3768 : nor02_2x port map ( Y=>nx10904, A0=>gen_0_cmp_pMux_2, A1=>nx3761
   );
   ix3778 : xnor2 port map ( Y=>nx10912, A0=>gen_0_cmp_pMux_0, A1=>nx10900);
   ix3784 : aoi21 port map ( Y=>nx10920, A0=>gen_0_cmp_pMux_1, A1=>
      gen_0_cmp_pMux_0, B0=>nx3769);
   ix4004 : nor02_2x port map ( Y=>nx10928, A0=>nx4013, A1=>gen_1_cmp_pMux_0
   );
   ix4012 : nor02_2x port map ( Y=>nx10944, A0=>gen_1_cmp_pMux_2, A1=>nx4005
   );
   ix4022 : xnor2 port map ( Y=>nx10952, A0=>gen_1_cmp_pMux_0, A1=>nx10940);
   ix4028 : aoi21 port map ( Y=>nx10960, A0=>gen_1_cmp_pMux_1, A1=>
      gen_1_cmp_pMux_0, B0=>nx4013);
   ix4252 : nor02_2x port map ( Y=>nx10968, A0=>nx4260, A1=>gen_2_cmp_pMux_0
   );
   ix4259 : nor02_2x port map ( Y=>nx10984, A0=>gen_2_cmp_pMux_2, A1=>nx4253
   );
   ix4270 : xnor2 port map ( Y=>nx10992, A0=>gen_2_cmp_pMux_0, A1=>nx10980);
   ix4276 : aoi21 port map ( Y=>nx11000, A0=>gen_2_cmp_pMux_1, A1=>
      gen_2_cmp_pMux_0, B0=>nx4260);
   ix4500 : nor02_2x port map ( Y=>nx11008, A0=>nx4509, A1=>gen_3_cmp_pMux_0
   );
   ix4508 : nor02_2x port map ( Y=>nx11024, A0=>gen_3_cmp_pMux_2, A1=>nx4501
   );
   ix4518 : xnor2 port map ( Y=>nx11032, A0=>gen_3_cmp_pMux_0, A1=>nx11020);
   ix4524 : aoi21 port map ( Y=>nx11040, A0=>gen_3_cmp_pMux_1, A1=>
      gen_3_cmp_pMux_0, B0=>nx4509);
   ix4747 : nor02_2x port map ( Y=>nx11048, A0=>nx4757, A1=>gen_4_cmp_pMux_0
   );
   ix4756 : nor02_2x port map ( Y=>nx11064, A0=>gen_4_cmp_pMux_2, A1=>nx4748
   );
   ix4766 : xnor2 port map ( Y=>nx11072, A0=>gen_4_cmp_pMux_0, A1=>nx11060);
   ix4770 : aoi21 port map ( Y=>nx11080, A0=>gen_4_cmp_pMux_1, A1=>
      gen_4_cmp_pMux_0, B0=>nx4757);
   ix4994 : nor02_2x port map ( Y=>nx11088, A0=>nx5003, A1=>gen_5_cmp_pMux_0
   );
   ix5002 : nor02_2x port map ( Y=>nx11104, A0=>gen_5_cmp_pMux_2, A1=>nx4995
   );
   ix5012 : xnor2 port map ( Y=>nx11112, A0=>gen_5_cmp_pMux_0, A1=>nx11100);
   ix5018 : aoi21 port map ( Y=>nx11120, A0=>gen_5_cmp_pMux_1, A1=>
      gen_5_cmp_pMux_0, B0=>nx5003);
   ix5243 : nor02_2x port map ( Y=>nx11128, A0=>nx5253, A1=>gen_6_cmp_pMux_0
   );
   ix5252 : nor02_2x port map ( Y=>nx11144, A0=>gen_6_cmp_pMux_2, A1=>nx5244
   );
   ix5262 : xnor2 port map ( Y=>nx11152, A0=>gen_6_cmp_pMux_0, A1=>nx11140);
   ix5266 : aoi21 port map ( Y=>nx11160, A0=>gen_6_cmp_pMux_1, A1=>
      gen_6_cmp_pMux_0, B0=>nx5253);
   ix5490 : nor02_2x port map ( Y=>nx11168, A0=>nx5499, A1=>gen_7_cmp_pMux_0
   );
   ix5498 : nor02_2x port map ( Y=>nx11184, A0=>gen_7_cmp_pMux_2, A1=>nx5491
   );
   ix5508 : xnor2 port map ( Y=>nx11192, A0=>gen_7_cmp_pMux_0, A1=>nx11180);
   ix5512 : aoi21 port map ( Y=>nx11200, A0=>gen_7_cmp_pMux_1, A1=>
      gen_7_cmp_pMux_0, B0=>nx5499);
   ix5734 : nor02_2x port map ( Y=>nx11208, A0=>nx5743, A1=>gen_8_cmp_pMux_0
   );
   ix5742 : nor02_2x port map ( Y=>nx11224, A0=>gen_8_cmp_pMux_2, A1=>nx5735
   );
   ix5752 : xnor2 port map ( Y=>nx11232, A0=>gen_8_cmp_pMux_0, A1=>nx11220);
   ix5758 : aoi21 port map ( Y=>nx11240, A0=>gen_8_cmp_pMux_1, A1=>
      gen_8_cmp_pMux_0, B0=>nx5743);
   ix5978 : nor02_2x port map ( Y=>nx11248, A0=>nx5987, A1=>gen_9_cmp_pMux_0
   );
   ix5986 : nor02_2x port map ( Y=>nx11264, A0=>gen_9_cmp_pMux_2, A1=>nx5979
   );
   ix5996 : xnor2 port map ( Y=>nx11272, A0=>gen_9_cmp_pMux_0, A1=>nx11260);
   ix6002 : aoi21 port map ( Y=>nx11280, A0=>gen_9_cmp_pMux_1, A1=>
      gen_9_cmp_pMux_0, B0=>nx5987);
   ix6224 : nor02_2x port map ( Y=>nx11288, A0=>nx6233, A1=>
      gen_10_cmp_pMux_0);
   ix6232 : nor02_2x port map ( Y=>nx11304, A0=>gen_10_cmp_pMux_2, A1=>
      nx6225);
   ix6242 : xnor2 port map ( Y=>nx11312, A0=>gen_10_cmp_pMux_0, A1=>nx11300
   );
   ix6247 : aoi21 port map ( Y=>nx11320, A0=>gen_10_cmp_pMux_1, A1=>
      gen_10_cmp_pMux_0, B0=>nx6233);
   ix6467 : nor02_2x port map ( Y=>nx11328, A0=>nx6477, A1=>
      gen_11_cmp_pMux_0);
   ix6476 : nor02_2x port map ( Y=>nx11344, A0=>gen_11_cmp_pMux_2, A1=>
      nx6468);
   ix6486 : xnor2 port map ( Y=>nx11352, A0=>gen_11_cmp_pMux_0, A1=>nx11340
   );
   ix6490 : aoi21 port map ( Y=>nx11360, A0=>gen_11_cmp_pMux_1, A1=>
      gen_11_cmp_pMux_0, B0=>nx6477);
   ix6716 : nor02_2x port map ( Y=>nx11368, A0=>nx6725, A1=>
      gen_12_cmp_pMux_0);
   ix6724 : nor02_2x port map ( Y=>nx11384, A0=>gen_12_cmp_pMux_2, A1=>
      nx6717);
   ix6734 : xnor2 port map ( Y=>nx11392, A0=>gen_12_cmp_pMux_0, A1=>nx11380
   );
   ix6740 : aoi21 port map ( Y=>nx11400, A0=>gen_12_cmp_pMux_1, A1=>
      gen_12_cmp_pMux_0, B0=>nx6725);
   ix6963 : nor02_2x port map ( Y=>nx11408, A0=>nx6973, A1=>
      gen_13_cmp_pMux_0);
   ix6972 : nor02_2x port map ( Y=>nx11424, A0=>gen_13_cmp_pMux_2, A1=>
      nx6965);
   ix6982 : xnor2 port map ( Y=>nx11432, A0=>gen_13_cmp_pMux_0, A1=>nx11420
   );
   ix6988 : aoi21 port map ( Y=>nx11440, A0=>gen_13_cmp_pMux_1, A1=>
      gen_13_cmp_pMux_0, B0=>nx6973);
   ix7212 : nor02_2x port map ( Y=>nx11448, A0=>nx7221, A1=>
      gen_14_cmp_pMux_0);
   ix7220 : nor02_2x port map ( Y=>nx11464, A0=>gen_14_cmp_pMux_2, A1=>
      nx7213);
   ix7230 : xnor2 port map ( Y=>nx11472, A0=>gen_14_cmp_pMux_0, A1=>nx11460
   );
   ix7236 : aoi21 port map ( Y=>nx11480, A0=>gen_14_cmp_pMux_1, A1=>
      gen_14_cmp_pMux_0, B0=>nx7221);
   ix7461 : nor02_2x port map ( Y=>nx11488, A0=>nx7471, A1=>
      gen_15_cmp_pMux_0);
   ix7470 : nor02_2x port map ( Y=>nx11504, A0=>gen_15_cmp_pMux_2, A1=>
      nx7463);
   ix7480 : xnor2 port map ( Y=>nx11512, A0=>gen_15_cmp_pMux_0, A1=>nx11500
   );
   ix7486 : aoi21 port map ( Y=>nx11520, A0=>gen_15_cmp_pMux_1, A1=>
      gen_15_cmp_pMux_0, B0=>nx7471);
   ix7708 : nor02_2x port map ( Y=>nx11528, A0=>nx7717, A1=>
      gen_16_cmp_pMux_0);
   ix7716 : nor02_2x port map ( Y=>nx11544, A0=>gen_16_cmp_pMux_2, A1=>
      nx7709);
   ix7726 : xnor2 port map ( Y=>nx11552, A0=>gen_16_cmp_pMux_0, A1=>nx11540
   );
   ix7731 : aoi21 port map ( Y=>nx11560, A0=>gen_16_cmp_pMux_1, A1=>
      gen_16_cmp_pMux_0, B0=>nx7717);
   ix7952 : nor02_2x port map ( Y=>nx11568, A0=>nx7961, A1=>
      gen_17_cmp_pMux_0);
   ix7960 : nor02_2x port map ( Y=>nx11584, A0=>gen_17_cmp_pMux_2, A1=>
      nx7953);
   ix7970 : xnor2 port map ( Y=>nx11592, A0=>gen_17_cmp_pMux_0, A1=>nx11580
   );
   ix7976 : aoi21 port map ( Y=>nx11600, A0=>gen_17_cmp_pMux_1, A1=>
      gen_17_cmp_pMux_0, B0=>nx7961);
   ix8199 : nor02_2x port map ( Y=>nx11608, A0=>nx8209, A1=>
      gen_18_cmp_pMux_0);
   ix8208 : nor02_2x port map ( Y=>nx11624, A0=>gen_18_cmp_pMux_2, A1=>
      nx8200);
   ix8218 : xnor2 port map ( Y=>nx11632, A0=>gen_18_cmp_pMux_0, A1=>nx11620
   );
   ix8222 : aoi21 port map ( Y=>nx11640, A0=>gen_18_cmp_pMux_1, A1=>
      gen_18_cmp_pMux_0, B0=>nx8209);
   ix8446 : nor02_2x port map ( Y=>nx11648, A0=>nx8455, A1=>
      gen_19_cmp_pMux_0);
   ix8454 : nor02_2x port map ( Y=>nx11664, A0=>gen_19_cmp_pMux_2, A1=>
      nx8447);
   ix8464 : xnor2 port map ( Y=>nx11672, A0=>gen_19_cmp_pMux_0, A1=>nx11660
   );
   ix8470 : aoi21 port map ( Y=>nx11680, A0=>gen_19_cmp_pMux_1, A1=>
      gen_19_cmp_pMux_0, B0=>nx8455);
   ix8693 : nor02_2x port map ( Y=>nx11688, A0=>nx8701, A1=>
      gen_20_cmp_pMux_0);
   ix8700 : nor02_2x port map ( Y=>nx11704, A0=>gen_20_cmp_pMux_2, A1=>
      nx8694);
   ix8710 : xnor2 port map ( Y=>nx11712, A0=>gen_20_cmp_pMux_0, A1=>nx11700
   );
   ix8716 : aoi21 port map ( Y=>nx11720, A0=>gen_20_cmp_pMux_1, A1=>
      gen_20_cmp_pMux_0, B0=>nx8701);
   ix8936 : nor02_2x port map ( Y=>nx11728, A0=>nx8945, A1=>
      gen_21_cmp_pMux_0);
   ix8944 : nor02_2x port map ( Y=>nx11744, A0=>gen_21_cmp_pMux_2, A1=>
      nx8937);
   ix8954 : xnor2 port map ( Y=>nx11752, A0=>gen_21_cmp_pMux_0, A1=>nx11740
   );
   ix8960 : aoi21 port map ( Y=>nx11760, A0=>gen_21_cmp_pMux_1, A1=>
      gen_21_cmp_pMux_0, B0=>nx8945);
   ix9186 : nor02_2x port map ( Y=>nx11768, A0=>nx9195, A1=>
      gen_22_cmp_pMux_0);
   ix9194 : nor02_2x port map ( Y=>nx11784, A0=>gen_22_cmp_pMux_2, A1=>
      nx9187);
   ix9204 : xnor2 port map ( Y=>nx11792, A0=>gen_22_cmp_pMux_0, A1=>nx11780
   );
   ix9210 : aoi21 port map ( Y=>nx11800, A0=>gen_22_cmp_pMux_1, A1=>
      gen_22_cmp_pMux_0, B0=>nx9195);
   ix9435 : nor02_2x port map ( Y=>nx11808, A0=>nx9445, A1=>
      gen_23_cmp_pMux_0);
   ix9444 : nor02_2x port map ( Y=>nx11824, A0=>gen_23_cmp_pMux_2, A1=>
      nx9437);
   ix9454 : xnor2 port map ( Y=>nx11832, A0=>gen_23_cmp_pMux_0, A1=>nx11820
   );
   ix9460 : aoi21 port map ( Y=>nx11840, A0=>gen_23_cmp_pMux_1, A1=>
      gen_23_cmp_pMux_0, B0=>nx9445);
   ix9675 : nor02_2x port map ( Y=>nx11848, A0=>nx9683, A1=>
      gen_24_cmp_pMux_0);
   ix9682 : nor02_2x port map ( Y=>nx11864, A0=>gen_24_cmp_pMux_2, A1=>
      nx9676);
   ix9691 : xnor2 port map ( Y=>nx11872, A0=>gen_24_cmp_pMux_0, A1=>nx11860
   );
   ix9696 : aoi21 port map ( Y=>nx11880, A0=>gen_24_cmp_pMux_1, A1=>
      gen_24_cmp_pMux_0, B0=>nx9683);
   ix11895 : inv02 port map ( Y=>nx11896, A=>nx11938);
   ix11897 : inv02 port map ( Y=>nx11898, A=>nx11938);
   ix11899 : inv02 port map ( Y=>nx11900, A=>nx11938);
   ix11901 : inv02 port map ( Y=>nx11902, A=>nx11938);
   ix11903 : inv02 port map ( Y=>nx11904, A=>nx11938);
   ix11905 : inv02 port map ( Y=>nx11906, A=>nx11938);
   ix11907 : inv02 port map ( Y=>nx11908, A=>nx11940);
   ix11909 : inv02 port map ( Y=>nx11910, A=>nx11940);
   ix11911 : inv02 port map ( Y=>nx11912, A=>nx11940);
   ix11913 : inv01 port map ( Y=>nx11914, A=>nx11940);
   ix11915 : inv02 port map ( Y=>nx11916, A=>nx11934);
   ix11917 : inv02 port map ( Y=>nx11918, A=>nx11936);
   ix11919 : inv02 port map ( Y=>nx11920, A=>nx11936);
   ix11921 : inv02 port map ( Y=>nx11922, A=>nx11936);
   ix11923 : inv02 port map ( Y=>nx11924, A=>nx11936);
   ix11925 : inv02 port map ( Y=>nx11926, A=>nx11936);
   ix11927 : inv02 port map ( Y=>nx11928, A=>nx11936);
   ix11933 : inv02 port map ( Y=>nx11934, A=>nx10880);
   ix11935 : inv02 port map ( Y=>nx11936, A=>nx10880);
   ix11937 : inv02 port map ( Y=>nx11938, A=>nx10120);
   ix11939 : inv02 port map ( Y=>nx11940, A=>nx10120);
end CNNMulsArch ;

