
-- 
-- Definition of  CNNCores
-- 
--      Sun Apr 21 22:35:38 2019
--      
--      LeonardoSpectrum Level 3, 2018a.2
-- 

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity Reg_33 is
   port (
      D : IN std_logic_vector (32 DOWNTO 0) ;
      en : IN std_logic ;
      clk : IN std_logic ;
      rst : IN std_logic ;
      Q : OUT std_logic_vector (32 DOWNTO 0)) ;
end Reg_33 ;

architecture RegArch_unfold_1389 of Reg_33 is
   signal Q_30_EXMPLR, Q_29_EXMPLR, Q_28_EXMPLR, Q_27_EXMPLR, Q_26_EXMPLR, 
      Q_25_EXMPLR, Q_24_EXMPLR, Q_23_EXMPLR, Q_22_EXMPLR, Q_21_EXMPLR, 
      Q_20_EXMPLR, Q_19_EXMPLR, Q_18_EXMPLR, Q_17_EXMPLR, Q_16_EXMPLR, 
      Q_15_EXMPLR, Q_14_EXMPLR, Q_13_EXMPLR, Q_12_EXMPLR, Q_11_EXMPLR, 
      Q_10_EXMPLR, Q_9_EXMPLR, Q_8_EXMPLR, Q_7_EXMPLR, Q_6_EXMPLR, 
      Q_5_EXMPLR, Q_4_EXMPLR, Q_3_EXMPLR, Q_2_EXMPLR, Q_1_EXMPLR, Q_0_EXMPLR, 
      Q_32_EXMPLR, nx115, nx125, nx135, nx145, nx155, nx165, nx175, nx185, 
      nx195, nx205, nx215, nx225, nx235, nx245, nx255, nx265, nx275, nx285, 
      nx295, nx305, nx315, nx325, nx335, nx345, nx355, nx365, nx375, nx385, 
      nx395, nx405, nx415, nx427, nx431, nx436, nx438, nx443, nx445, nx450, 
      nx452, nx457, nx459, nx464, nx466, nx471, nx473, nx478, nx480, nx485, 
      nx487, nx492, nx494, nx499, nx501, nx506, nx508, nx513, nx515, nx520, 
      nx522, nx527, nx529, nx534, nx536, nx541, nx543, nx548, nx550, nx555, 
      nx557, nx562, nx564, nx569, nx571, nx576, nx578, nx583, nx585, nx590, 
      nx592, nx597, nx599, nx604, nx606, nx611, nx613, nx618, nx620, nx625, 
      nx627, nx632, nx634, nx639, nx641, nx649, nx651, nx653, nx655, nx657, 
      nx663, nx665, nx667, nx669, nx671, nx673, nx675, nx677, nx679, nx681, 
      nx683, nx685: std_logic ;

begin
   Q(32) <= Q_32_EXMPLR ;
   Q(31) <= Q_32_EXMPLR ;
   Q(30) <= Q_30_EXMPLR ;
   Q(29) <= Q_29_EXMPLR ;
   Q(28) <= Q_28_EXMPLR ;
   Q(27) <= Q_27_EXMPLR ;
   Q(26) <= Q_26_EXMPLR ;
   Q(25) <= Q_25_EXMPLR ;
   Q(24) <= Q_24_EXMPLR ;
   Q(23) <= Q_23_EXMPLR ;
   Q(22) <= Q_22_EXMPLR ;
   Q(21) <= Q_21_EXMPLR ;
   Q(20) <= Q_20_EXMPLR ;
   Q(19) <= Q_19_EXMPLR ;
   Q(18) <= Q_18_EXMPLR ;
   Q(17) <= Q_17_EXMPLR ;
   Q(16) <= Q_16_EXMPLR ;
   Q(15) <= Q_15_EXMPLR ;
   Q(14) <= Q_14_EXMPLR ;
   Q(13) <= Q_13_EXMPLR ;
   Q(12) <= Q_12_EXMPLR ;
   Q(11) <= Q_11_EXMPLR ;
   Q(10) <= Q_10_EXMPLR ;
   Q(9) <= Q_9_EXMPLR ;
   Q(8) <= Q_8_EXMPLR ;
   Q(7) <= Q_7_EXMPLR ;
   Q(6) <= Q_6_EXMPLR ;
   Q(5) <= Q_5_EXMPLR ;
   Q(4) <= Q_4_EXMPLR ;
   Q(3) <= Q_3_EXMPLR ;
   Q(2) <= Q_2_EXMPLR ;
   Q(1) <= Q_1_EXMPLR ;
   Q(0) <= Q_0_EXMPLR ;
   ix43 : fake_gnd port map ( Y=>Q_32_EXMPLR);
   reg_Q_0 : dffr port map ( Q=>Q_0_EXMPLR, QB=>OPEN, D=>nx115, CLK=>nx675, 
      R=>rst);
   ix116 : nand02 port map ( Y=>nx115, A0=>nx427, A1=>nx431);
   ix428 : nand02 port map ( Y=>nx427, A0=>Q_0_EXMPLR, A1=>nx685);
   ix432 : nand02 port map ( Y=>nx431, A0=>D(0), A1=>nx663);
   reg_Q_1 : dffr port map ( Q=>Q_1_EXMPLR, QB=>OPEN, D=>nx125, CLK=>nx675, 
      R=>rst);
   ix126 : nand02 port map ( Y=>nx125, A0=>nx436, A1=>nx438);
   ix437 : nand02 port map ( Y=>nx436, A0=>Q_1_EXMPLR, A1=>nx685);
   ix439 : nand02 port map ( Y=>nx438, A0=>D(1), A1=>nx663);
   reg_Q_2 : dffr port map ( Q=>Q_2_EXMPLR, QB=>OPEN, D=>nx135, CLK=>nx675, 
      R=>rst);
   ix136 : nand02 port map ( Y=>nx135, A0=>nx443, A1=>nx445);
   ix444 : nand02 port map ( Y=>nx443, A0=>Q_2_EXMPLR, A1=>nx685);
   ix446 : nand02 port map ( Y=>nx445, A0=>D(2), A1=>nx663);
   reg_Q_3 : dffr port map ( Q=>Q_3_EXMPLR, QB=>OPEN, D=>nx145, CLK=>nx675, 
      R=>rst);
   ix146 : nand02 port map ( Y=>nx145, A0=>nx450, A1=>nx452);
   ix451 : nand02 port map ( Y=>nx450, A0=>Q_3_EXMPLR, A1=>nx685);
   ix453 : nand02 port map ( Y=>nx452, A0=>D(3), A1=>nx663);
   reg_Q_4 : dffr port map ( Q=>Q_4_EXMPLR, QB=>OPEN, D=>nx155, CLK=>nx675, 
      R=>rst);
   ix156 : nand02 port map ( Y=>nx155, A0=>nx457, A1=>nx459);
   ix458 : nand02 port map ( Y=>nx457, A0=>Q_4_EXMPLR, A1=>nx685);
   ix460 : nand02 port map ( Y=>nx459, A0=>D(4), A1=>nx663);
   reg_Q_5 : dffr port map ( Q=>Q_5_EXMPLR, QB=>OPEN, D=>nx165, CLK=>nx675, 
      R=>rst);
   ix166 : nand02 port map ( Y=>nx165, A0=>nx464, A1=>nx466);
   ix465 : nand02 port map ( Y=>nx464, A0=>Q_5_EXMPLR, A1=>nx685);
   ix467 : nand02 port map ( Y=>nx466, A0=>D(5), A1=>nx663);
   reg_Q_6 : dffr port map ( Q=>Q_6_EXMPLR, QB=>OPEN, D=>nx175, CLK=>nx675, 
      R=>rst);
   ix176 : nand02 port map ( Y=>nx175, A0=>nx471, A1=>nx473);
   ix472 : nand02 port map ( Y=>nx471, A0=>Q_6_EXMPLR, A1=>nx685);
   ix474 : nand02 port map ( Y=>nx473, A0=>D(6), A1=>nx663);
   reg_Q_7 : dffr port map ( Q=>Q_7_EXMPLR, QB=>OPEN, D=>nx185, CLK=>nx677, 
      R=>rst);
   ix186 : nand02 port map ( Y=>nx185, A0=>nx478, A1=>nx480);
   ix479 : nand02 port map ( Y=>nx478, A0=>Q_7_EXMPLR, A1=>nx651);
   ix481 : nand02 port map ( Y=>nx480, A0=>D(7), A1=>nx665);
   reg_Q_8 : dffr port map ( Q=>Q_8_EXMPLR, QB=>OPEN, D=>nx195, CLK=>nx677, 
      R=>rst);
   ix196 : nand02 port map ( Y=>nx195, A0=>nx485, A1=>nx487);
   ix486 : nand02 port map ( Y=>nx485, A0=>Q_8_EXMPLR, A1=>nx651);
   ix488 : nand02 port map ( Y=>nx487, A0=>D(8), A1=>nx665);
   reg_Q_9 : dffr port map ( Q=>Q_9_EXMPLR, QB=>OPEN, D=>nx205, CLK=>nx677, 
      R=>rst);
   ix206 : nand02 port map ( Y=>nx205, A0=>nx492, A1=>nx494);
   ix493 : nand02 port map ( Y=>nx492, A0=>Q_9_EXMPLR, A1=>nx651);
   ix495 : nand02 port map ( Y=>nx494, A0=>D(9), A1=>nx665);
   reg_Q_10 : dffr port map ( Q=>Q_10_EXMPLR, QB=>OPEN, D=>nx215, CLK=>nx677, 
      R=>rst);
   ix216 : nand02 port map ( Y=>nx215, A0=>nx499, A1=>nx501);
   ix500 : nand02 port map ( Y=>nx499, A0=>Q_10_EXMPLR, A1=>nx651);
   ix502 : nand02 port map ( Y=>nx501, A0=>D(10), A1=>nx665);
   reg_Q_11 : dffr port map ( Q=>Q_11_EXMPLR, QB=>OPEN, D=>nx225, CLK=>nx677, 
      R=>rst);
   ix226 : nand02 port map ( Y=>nx225, A0=>nx506, A1=>nx508);
   ix507 : nand02 port map ( Y=>nx506, A0=>Q_11_EXMPLR, A1=>nx651);
   ix509 : nand02 port map ( Y=>nx508, A0=>D(11), A1=>nx665);
   reg_Q_12 : dffr port map ( Q=>Q_12_EXMPLR, QB=>OPEN, D=>nx235, CLK=>nx677, 
      R=>rst);
   ix236 : nand02 port map ( Y=>nx235, A0=>nx513, A1=>nx515);
   ix514 : nand02 port map ( Y=>nx513, A0=>Q_12_EXMPLR, A1=>nx651);
   ix516 : nand02 port map ( Y=>nx515, A0=>D(12), A1=>nx665);
   reg_Q_13 : dffr port map ( Q=>Q_13_EXMPLR, QB=>OPEN, D=>nx245, CLK=>nx677, 
      R=>rst);
   ix246 : nand02 port map ( Y=>nx245, A0=>nx520, A1=>nx522);
   ix521 : nand02 port map ( Y=>nx520, A0=>Q_13_EXMPLR, A1=>nx651);
   ix523 : nand02 port map ( Y=>nx522, A0=>D(13), A1=>nx665);
   reg_Q_14 : dffr port map ( Q=>Q_14_EXMPLR, QB=>OPEN, D=>nx255, CLK=>nx679, 
      R=>rst);
   ix256 : nand02 port map ( Y=>nx255, A0=>nx527, A1=>nx529);
   ix528 : nand02 port map ( Y=>nx527, A0=>Q_14_EXMPLR, A1=>nx653);
   ix530 : nand02 port map ( Y=>nx529, A0=>D(14), A1=>nx667);
   reg_Q_15 : dffr port map ( Q=>Q_15_EXMPLR, QB=>OPEN, D=>nx265, CLK=>nx679, 
      R=>rst);
   ix266 : nand02 port map ( Y=>nx265, A0=>nx534, A1=>nx536);
   ix535 : nand02 port map ( Y=>nx534, A0=>Q_15_EXMPLR, A1=>nx653);
   ix537 : nand02 port map ( Y=>nx536, A0=>D(15), A1=>nx667);
   reg_Q_16 : dffr port map ( Q=>Q_16_EXMPLR, QB=>OPEN, D=>nx275, CLK=>nx679, 
      R=>rst);
   ix276 : nand02 port map ( Y=>nx275, A0=>nx541, A1=>nx543);
   ix542 : nand02 port map ( Y=>nx541, A0=>Q_16_EXMPLR, A1=>nx653);
   ix544 : nand02 port map ( Y=>nx543, A0=>D(16), A1=>nx667);
   reg_Q_17 : dffr port map ( Q=>Q_17_EXMPLR, QB=>OPEN, D=>nx285, CLK=>nx679, 
      R=>rst);
   ix286 : nand02 port map ( Y=>nx285, A0=>nx548, A1=>nx550);
   ix549 : nand02 port map ( Y=>nx548, A0=>Q_17_EXMPLR, A1=>nx653);
   ix551 : nand02 port map ( Y=>nx550, A0=>D(17), A1=>nx667);
   reg_Q_18 : dffr port map ( Q=>Q_18_EXMPLR, QB=>OPEN, D=>nx295, CLK=>nx679, 
      R=>rst);
   ix296 : nand02 port map ( Y=>nx295, A0=>nx555, A1=>nx557);
   ix556 : nand02 port map ( Y=>nx555, A0=>Q_18_EXMPLR, A1=>nx653);
   ix558 : nand02 port map ( Y=>nx557, A0=>D(18), A1=>nx667);
   reg_Q_19 : dffr port map ( Q=>Q_19_EXMPLR, QB=>OPEN, D=>nx305, CLK=>nx679, 
      R=>rst);
   ix306 : nand02 port map ( Y=>nx305, A0=>nx562, A1=>nx564);
   ix563 : nand02 port map ( Y=>nx562, A0=>Q_19_EXMPLR, A1=>nx653);
   ix565 : nand02 port map ( Y=>nx564, A0=>D(19), A1=>nx667);
   reg_Q_20 : dffr port map ( Q=>Q_20_EXMPLR, QB=>OPEN, D=>nx315, CLK=>nx679, 
      R=>rst);
   ix316 : nand02 port map ( Y=>nx315, A0=>nx569, A1=>nx571);
   ix570 : nand02 port map ( Y=>nx569, A0=>Q_20_EXMPLR, A1=>nx653);
   ix572 : nand02 port map ( Y=>nx571, A0=>D(20), A1=>nx667);
   reg_Q_21 : dffr port map ( Q=>Q_21_EXMPLR, QB=>OPEN, D=>nx325, CLK=>nx681, 
      R=>rst);
   ix326 : nand02 port map ( Y=>nx325, A0=>nx576, A1=>nx578);
   ix577 : nand02 port map ( Y=>nx576, A0=>Q_21_EXMPLR, A1=>nx655);
   ix579 : nand02 port map ( Y=>nx578, A0=>D(21), A1=>nx669);
   reg_Q_22 : dffr port map ( Q=>Q_22_EXMPLR, QB=>OPEN, D=>nx335, CLK=>nx681, 
      R=>rst);
   ix336 : nand02 port map ( Y=>nx335, A0=>nx583, A1=>nx585);
   ix584 : nand02 port map ( Y=>nx583, A0=>Q_22_EXMPLR, A1=>nx655);
   ix586 : nand02 port map ( Y=>nx585, A0=>D(22), A1=>nx669);
   reg_Q_23 : dffr port map ( Q=>Q_23_EXMPLR, QB=>OPEN, D=>nx345, CLK=>nx681, 
      R=>rst);
   ix346 : nand02 port map ( Y=>nx345, A0=>nx590, A1=>nx592);
   ix591 : nand02 port map ( Y=>nx590, A0=>Q_23_EXMPLR, A1=>nx655);
   ix593 : nand02 port map ( Y=>nx592, A0=>D(23), A1=>nx669);
   reg_Q_24 : dffr port map ( Q=>Q_24_EXMPLR, QB=>OPEN, D=>nx355, CLK=>nx681, 
      R=>rst);
   ix356 : nand02 port map ( Y=>nx355, A0=>nx597, A1=>nx599);
   ix598 : nand02 port map ( Y=>nx597, A0=>Q_24_EXMPLR, A1=>nx655);
   ix600 : nand02 port map ( Y=>nx599, A0=>D(24), A1=>nx669);
   reg_Q_25 : dffr port map ( Q=>Q_25_EXMPLR, QB=>OPEN, D=>nx365, CLK=>nx681, 
      R=>rst);
   ix366 : nand02 port map ( Y=>nx365, A0=>nx604, A1=>nx606);
   ix605 : nand02 port map ( Y=>nx604, A0=>Q_25_EXMPLR, A1=>nx655);
   ix607 : nand02 port map ( Y=>nx606, A0=>D(25), A1=>nx669);
   reg_Q_26 : dffr port map ( Q=>Q_26_EXMPLR, QB=>OPEN, D=>nx375, CLK=>nx681, 
      R=>rst);
   ix376 : nand02 port map ( Y=>nx375, A0=>nx611, A1=>nx613);
   ix612 : nand02 port map ( Y=>nx611, A0=>Q_26_EXMPLR, A1=>nx655);
   ix614 : nand02 port map ( Y=>nx613, A0=>D(26), A1=>nx669);
   reg_Q_27 : dffr port map ( Q=>Q_27_EXMPLR, QB=>OPEN, D=>nx385, CLK=>nx681, 
      R=>rst);
   ix386 : nand02 port map ( Y=>nx385, A0=>nx618, A1=>nx620);
   ix619 : nand02 port map ( Y=>nx618, A0=>Q_27_EXMPLR, A1=>nx655);
   ix621 : nand02 port map ( Y=>nx620, A0=>D(27), A1=>nx669);
   reg_Q_28 : dffr port map ( Q=>Q_28_EXMPLR, QB=>OPEN, D=>nx395, CLK=>nx683, 
      R=>rst);
   ix396 : nand02 port map ( Y=>nx395, A0=>nx625, A1=>nx627);
   ix626 : nand02 port map ( Y=>nx625, A0=>Q_28_EXMPLR, A1=>nx657);
   ix628 : nand02 port map ( Y=>nx627, A0=>D(28), A1=>nx671);
   reg_Q_29 : dffr port map ( Q=>Q_29_EXMPLR, QB=>OPEN, D=>nx405, CLK=>nx683, 
      R=>rst);
   ix406 : nand02 port map ( Y=>nx405, A0=>nx632, A1=>nx634);
   ix633 : nand02 port map ( Y=>nx632, A0=>Q_29_EXMPLR, A1=>nx657);
   ix635 : nand02 port map ( Y=>nx634, A0=>D(29), A1=>nx671);
   reg_Q_30 : dffr port map ( Q=>Q_30_EXMPLR, QB=>OPEN, D=>nx415, CLK=>nx683, 
      R=>rst);
   ix416 : nand02 port map ( Y=>nx415, A0=>nx639, A1=>nx641);
   ix640 : nand02 port map ( Y=>nx639, A0=>Q_30_EXMPLR, A1=>nx657);
   ix642 : nand02 port map ( Y=>nx641, A0=>D(30), A1=>nx671);
   ix648 : inv02 port map ( Y=>nx649, A=>en);
   ix650 : inv02 port map ( Y=>nx651, A=>nx671);
   ix652 : inv02 port map ( Y=>nx653, A=>nx671);
   ix654 : inv02 port map ( Y=>nx655, A=>nx671);
   ix656 : inv02 port map ( Y=>nx657, A=>nx671);
   ix662 : inv02 port map ( Y=>nx663, A=>nx649);
   ix664 : inv02 port map ( Y=>nx665, A=>nx649);
   ix666 : inv02 port map ( Y=>nx667, A=>nx649);
   ix668 : inv02 port map ( Y=>nx669, A=>nx649);
   ix670 : inv02 port map ( Y=>nx671, A=>nx649);
   ix672 : inv01 port map ( Y=>nx673, A=>clk);
   ix674 : inv02 port map ( Y=>nx675, A=>nx673);
   ix676 : inv02 port map ( Y=>nx677, A=>nx673);
   ix678 : inv02 port map ( Y=>nx679, A=>nx673);
   ix680 : inv02 port map ( Y=>nx681, A=>nx673);
   ix682 : inv02 port map ( Y=>nx683, A=>nx673);
   ix684 : inv02 port map ( Y=>nx685, A=>en);
end RegArch_unfold_1389 ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity BinaryMux_33 is
   port (
      a : IN std_logic_vector (32 DOWNTO 0) ;
      b : IN std_logic_vector (32 DOWNTO 0) ;
      sel : IN std_logic ;
      f : OUT std_logic_vector (32 DOWNTO 0)) ;
end BinaryMux_33 ;

architecture BinaryMuxArch_unfold_1786 of BinaryMux_33 is
   signal f_32_EXMPLR, nx93, nx97, nx99, nx105, nx107, nx111, nx113, nx117, 
      nx119, nx123, nx125, nx129, nx131, nx135, nx137, nx141, nx143, nx147, 
      nx151, nx155, nx158, nx161, nx164, nx167, nx170, nx173, nx176, nx179, 
      nx182, nx185, nx188, nx191, nx194, nx197, nx200, nx203, nx206, nx209, 
      nx212, nx219, nx221, nx223, nx225, nx227, nx229, nx231: std_logic ;

begin
   f(32) <= f_32_EXMPLR ;
   f(31) <= f_32_EXMPLR ;
   ix44 : fake_gnd port map ( Y=>f_32_EXMPLR);
   ix3 : nor02_2x port map ( Y=>f(0), A0=>nx93, A1=>nx219);
   ix94 : inv01 port map ( Y=>nx93, A=>a(0));
   ix99 : nand02_2x port map ( Y=>f(1), A0=>nx97, A1=>nx99);
   ix98 : nand02 port map ( Y=>nx97, A0=>b(1), A1=>nx219);
   ix100 : nand02 port map ( Y=>nx99, A0=>a(1), A1=>nx229);
   ix107 : nand02 port map ( Y=>f(2), A0=>nx105, A1=>nx107);
   ix106 : nand02 port map ( Y=>nx105, A0=>b(2), A1=>nx219);
   ix108 : nand02 port map ( Y=>nx107, A0=>a(2), A1=>nx229);
   ix115 : nand02 port map ( Y=>f(3), A0=>nx111, A1=>nx113);
   ix112 : nand02 port map ( Y=>nx111, A0=>b(3), A1=>nx219);
   ix114 : nand02 port map ( Y=>nx113, A0=>a(3), A1=>nx229);
   ix123 : nand02 port map ( Y=>f(4), A0=>nx117, A1=>nx119);
   ix118 : nand02 port map ( Y=>nx117, A0=>b(4), A1=>nx219);
   ix120 : nand02 port map ( Y=>nx119, A0=>a(4), A1=>nx229);
   ix131 : nand02 port map ( Y=>f(5), A0=>nx123, A1=>nx125);
   ix124 : nand02 port map ( Y=>nx123, A0=>b(5), A1=>nx219);
   ix126 : nand02 port map ( Y=>nx125, A0=>a(5), A1=>nx229);
   ix139 : nand02 port map ( Y=>f(6), A0=>nx129, A1=>nx131);
   ix130 : nand02 port map ( Y=>nx129, A0=>b(6), A1=>nx219);
   ix132 : nand02 port map ( Y=>nx131, A0=>a(6), A1=>nx229);
   ix147 : nand02 port map ( Y=>f(7), A0=>nx135, A1=>nx137);
   ix136 : nand02 port map ( Y=>nx135, A0=>b(7), A1=>nx221);
   ix138 : nand02 port map ( Y=>nx137, A0=>a(7), A1=>nx229);
   ix155 : nand02 port map ( Y=>f(8), A0=>nx141, A1=>nx143);
   ix142 : nand02 port map ( Y=>nx141, A0=>nx221, A1=>b(8));
   ix144 : nand02 port map ( Y=>nx143, A0=>nx231, A1=>a(8));
   ix7 : nor02_2x port map ( Y=>f(9), A0=>nx147, A1=>nx221);
   ix148 : inv01 port map ( Y=>nx147, A=>a(9));
   ix11 : nor02_2x port map ( Y=>f(10), A0=>nx151, A1=>nx221);
   ix152 : inv01 port map ( Y=>nx151, A=>a(10));
   ix15 : nor02_2x port map ( Y=>f(11), A0=>nx155, A1=>nx221);
   ix156 : inv01 port map ( Y=>nx155, A=>a(11));
   ix19 : nor02_2x port map ( Y=>f(12), A0=>nx158, A1=>nx221);
   ix159 : inv01 port map ( Y=>nx158, A=>a(12));
   ix23 : nor02_2x port map ( Y=>f(13), A0=>nx161, A1=>nx221);
   ix162 : inv01 port map ( Y=>nx161, A=>a(13));
   ix27 : nor02_2x port map ( Y=>f(14), A0=>nx164, A1=>nx223);
   ix165 : inv01 port map ( Y=>nx164, A=>a(14));
   ix31 : nor02_2x port map ( Y=>f(15), A0=>nx167, A1=>nx223);
   ix168 : inv01 port map ( Y=>nx167, A=>a(15));
   ix35 : nor02_2x port map ( Y=>f(16), A0=>nx170, A1=>nx223);
   ix171 : inv01 port map ( Y=>nx170, A=>a(16));
   ix39 : nor02_2x port map ( Y=>f(17), A0=>nx173, A1=>nx223);
   ix174 : inv01 port map ( Y=>nx173, A=>a(17));
   ix43 : nor02_2x port map ( Y=>f(18), A0=>nx176, A1=>nx223);
   ix177 : inv01 port map ( Y=>nx176, A=>a(18));
   ix47 : nor02_2x port map ( Y=>f(19), A0=>nx179, A1=>nx223);
   ix180 : inv01 port map ( Y=>nx179, A=>a(19));
   ix51 : nor02_2x port map ( Y=>f(20), A0=>nx182, A1=>nx223);
   ix183 : inv01 port map ( Y=>nx182, A=>a(20));
   ix55 : nor02_2x port map ( Y=>f(21), A0=>nx185, A1=>nx225);
   ix186 : inv01 port map ( Y=>nx185, A=>a(21));
   ix59 : nor02_2x port map ( Y=>f(22), A0=>nx188, A1=>nx225);
   ix189 : inv01 port map ( Y=>nx188, A=>a(22));
   ix63 : nor02_2x port map ( Y=>f(23), A0=>nx191, A1=>nx225);
   ix192 : inv01 port map ( Y=>nx191, A=>a(23));
   ix67 : nor02_2x port map ( Y=>f(24), A0=>nx194, A1=>nx225);
   ix195 : inv01 port map ( Y=>nx194, A=>a(24));
   ix71 : nor02_2x port map ( Y=>f(25), A0=>nx197, A1=>nx225);
   ix198 : inv01 port map ( Y=>nx197, A=>a(25));
   ix75 : nor02_2x port map ( Y=>f(26), A0=>nx200, A1=>nx225);
   ix201 : inv01 port map ( Y=>nx200, A=>a(26));
   ix79 : nor02_2x port map ( Y=>f(27), A0=>nx203, A1=>nx225);
   ix204 : inv01 port map ( Y=>nx203, A=>a(27));
   ix83 : nor02_2x port map ( Y=>f(28), A0=>nx206, A1=>nx227);
   ix207 : inv01 port map ( Y=>nx206, A=>a(28));
   ix87 : nor02_2x port map ( Y=>f(29), A0=>nx209, A1=>nx227);
   ix210 : inv01 port map ( Y=>nx209, A=>a(29));
   ix91 : nor02_2x port map ( Y=>f(30), A0=>nx212, A1=>nx227);
   ix213 : inv01 port map ( Y=>nx212, A=>a(30));
   ix218 : inv02 port map ( Y=>nx219, A=>nx231);
   ix220 : inv02 port map ( Y=>nx221, A=>nx231);
   ix222 : inv02 port map ( Y=>nx223, A=>nx231);
   ix224 : inv02 port map ( Y=>nx225, A=>nx231);
   ix226 : inv02 port map ( Y=>nx227, A=>nx231);
   ix228 : inv02 port map ( Y=>nx229, A=>sel);
   ix230 : inv02 port map ( Y=>nx231, A=>sel);
end BinaryMuxArch_unfold_1786 ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity NBitAdder_24 is
   port (
      a : IN std_logic_vector (23 DOWNTO 0) ;
      b : IN std_logic_vector (23 DOWNTO 0) ;
      carryIn : IN std_logic ;
      sum : OUT std_logic_vector (23 DOWNTO 0) ;
      carryOut : OUT std_logic) ;
end NBitAdder_24 ;

architecture NBitAdderArch_unfold_2081 of NBitAdder_24 is
   signal nx6, nx8, nx16, nx18, nx22, nx24, nx30, nx32, nx38, nx40, nx46, 
      nx48, nx54, nx56, nx62, nx64, nx70, nx72, nx78, nx80, nx86, nx88, nx94, 
      nx96, nx102, nx104, nx110, nx112, nx118, nx120, nx126, nx128, nx134, 
      nx136, nx142, nx144, nx150, nx152, nx158, nx160, nx166, nx168, nx170, 
      nx172, nx103, nx109, nx111, nx113, nx115, nx119, nx123, nx127, nx133, 
      nx135, nx137, nx141, nx145, nx149, nx155, nx157, nx159, nx163, nx167, 
      nx171, nx177, nx179, nx181, nx185, nx189, nx193, nx199, nx201, nx203, 
      nx207, nx211, nx215, nx221, nx223, nx225, nx229, nx232, nx235, nx239, 
      nx241, nx243, nx246, nx249, nx252, nx256, nx258, nx260, nx263, nx266, 
      nx269, nx273, nx275, nx277, nx280, nx283, nx286, nx290, nx292, nx294, 
      nx297, nx300, nx303, nx307, nx309, nx311, nx314, nx317, nx320, nx323, 
      nx326, nx329, nx332, nx335, nx338, nx341, nx344, nx347, nx350, nx353, 
      nx356, nx358, nx360, nx362, nx364, nx366, nx368, nx370, nx372: 
   std_logic ;

begin
   ix44 : fake_gnd port map ( Y=>carryOut);
   ix229 : xnor2 port map ( Y=>sum(0), A0=>carryIn, A1=>nx103);
   ix104 : xnor2 port map ( Y=>nx103, A0=>a(0), A1=>b(0));
   ix227 : xnor2 port map ( Y=>sum(1), A0=>nx6, A1=>nx115);
   ix7 : oai22 port map ( Y=>nx6, A0=>nx109, A1=>nx103, B0=>nx111, B1=>nx113
   );
   ix110 : inv01 port map ( Y=>nx109, A=>carryIn);
   ix112 : inv01 port map ( Y=>nx111, A=>b(0));
   ix114 : inv01 port map ( Y=>nx113, A=>a(0));
   ix116 : xnor2 port map ( Y=>nx115, A0=>a(1), A1=>b(1));
   ix225 : xnor2 port map ( Y=>sum(2), A0=>nx119, A1=>nx16);
   ix120 : aoi22 port map ( Y=>nx119, A0=>b(1), A1=>a(1), B0=>nx6, B1=>nx8);
   ix9 : xnor2 port map ( Y=>nx8, A0=>a(1), A1=>nx123);
   ix124 : inv01 port map ( Y=>nx123, A=>b(1));
   ix17 : xnor2 port map ( Y=>nx16, A0=>a(2), A1=>nx127);
   ix128 : inv01 port map ( Y=>nx127, A=>b(2));
   ix223 : xnor2 port map ( Y=>sum(3), A0=>nx22, A1=>nx137);
   ix23 : oai21 port map ( Y=>nx22, A0=>nx119, A1=>nx133, B0=>nx135);
   ix134 : xnor2 port map ( Y=>nx133, A0=>a(2), A1=>b(2));
   ix136 : nand02 port map ( Y=>nx135, A0=>b(2), A1=>a(2));
   ix138 : xnor2 port map ( Y=>nx137, A0=>a(3), A1=>b(3));
   ix221 : xnor2 port map ( Y=>sum(4), A0=>nx141, A1=>nx32);
   ix142 : aoi22 port map ( Y=>nx141, A0=>b(3), A1=>a(3), B0=>nx22, B1=>nx24
   );
   ix25 : xnor2 port map ( Y=>nx24, A0=>a(3), A1=>nx145);
   ix146 : inv01 port map ( Y=>nx145, A=>b(3));
   ix33 : xnor2 port map ( Y=>nx32, A0=>a(4), A1=>nx149);
   ix150 : inv01 port map ( Y=>nx149, A=>b(4));
   ix219 : xnor2 port map ( Y=>sum(5), A0=>nx38, A1=>nx159);
   ix39 : oai21 port map ( Y=>nx38, A0=>nx141, A1=>nx155, B0=>nx157);
   ix156 : xnor2 port map ( Y=>nx155, A0=>a(4), A1=>b(4));
   ix158 : nand02 port map ( Y=>nx157, A0=>b(4), A1=>a(4));
   ix160 : xnor2 port map ( Y=>nx159, A0=>a(5), A1=>b(5));
   ix217 : xnor2 port map ( Y=>sum(6), A0=>nx163, A1=>nx48);
   ix164 : aoi22 port map ( Y=>nx163, A0=>b(5), A1=>a(5), B0=>nx38, B1=>nx40
   );
   ix41 : xnor2 port map ( Y=>nx40, A0=>a(5), A1=>nx167);
   ix168 : inv01 port map ( Y=>nx167, A=>b(5));
   ix49 : xnor2 port map ( Y=>nx48, A0=>a(6), A1=>nx171);
   ix172 : inv01 port map ( Y=>nx171, A=>b(6));
   ix215 : xnor2 port map ( Y=>sum(7), A0=>nx54, A1=>nx181);
   ix55 : oai21 port map ( Y=>nx54, A0=>nx163, A1=>nx177, B0=>nx179);
   ix178 : xnor2 port map ( Y=>nx177, A0=>a(6), A1=>b(6));
   ix180 : nand02 port map ( Y=>nx179, A0=>b(6), A1=>a(6));
   ix182 : xnor2 port map ( Y=>nx181, A0=>a(7), A1=>b(7));
   ix213 : xnor2 port map ( Y=>sum(8), A0=>nx185, A1=>nx64);
   ix186 : aoi22 port map ( Y=>nx185, A0=>b(7), A1=>a(7), B0=>nx54, B1=>nx56
   );
   ix57 : xnor2 port map ( Y=>nx56, A0=>a(7), A1=>nx189);
   ix190 : inv01 port map ( Y=>nx189, A=>b(7));
   ix65 : xnor2 port map ( Y=>nx64, A0=>a(8), A1=>nx193);
   ix194 : inv01 port map ( Y=>nx193, A=>b(8));
   ix211 : xnor2 port map ( Y=>sum(9), A0=>nx70, A1=>nx203);
   ix71 : oai21 port map ( Y=>nx70, A0=>nx185, A1=>nx199, B0=>nx201);
   ix200 : xnor2 port map ( Y=>nx199, A0=>a(8), A1=>b(8));
   ix202 : nand02 port map ( Y=>nx201, A0=>b(8), A1=>a(8));
   ix204 : xnor2 port map ( Y=>nx203, A0=>a(9), A1=>b(9));
   ix209 : xnor2 port map ( Y=>sum(10), A0=>nx207, A1=>nx80);
   ix208 : aoi22 port map ( Y=>nx207, A0=>b(9), A1=>a(9), B0=>nx70, B1=>nx72
   );
   ix73 : xnor2 port map ( Y=>nx72, A0=>a(9), A1=>nx211);
   ix212 : inv01 port map ( Y=>nx211, A=>b(9));
   ix81 : xnor2 port map ( Y=>nx80, A0=>a(10), A1=>nx215);
   ix216 : inv01 port map ( Y=>nx215, A=>b(10));
   ix207 : xnor2 port map ( Y=>sum(11), A0=>nx86, A1=>nx225);
   ix87 : oai21 port map ( Y=>nx86, A0=>nx207, A1=>nx221, B0=>nx223);
   ix222 : xnor2 port map ( Y=>nx221, A0=>a(10), A1=>b(10));
   ix224 : nand02 port map ( Y=>nx223, A0=>b(10), A1=>a(10));
   ix226 : xnor2 port map ( Y=>nx225, A0=>a(11), A1=>b(11));
   ix205 : xnor2 port map ( Y=>sum(12), A0=>nx229, A1=>nx96);
   ix230 : aoi22 port map ( Y=>nx229, A0=>b(11), A1=>a(11), B0=>nx86, B1=>
      nx88);
   ix89 : xnor2 port map ( Y=>nx88, A0=>a(11), A1=>nx232);
   ix233 : inv01 port map ( Y=>nx232, A=>b(11));
   ix97 : xnor2 port map ( Y=>nx96, A0=>a(12), A1=>nx235);
   ix236 : inv01 port map ( Y=>nx235, A=>b(12));
   ix203 : xnor2 port map ( Y=>sum(13), A0=>nx102, A1=>nx243);
   ix103 : oai21 port map ( Y=>nx102, A0=>nx229, A1=>nx239, B0=>nx241);
   ix240 : xnor2 port map ( Y=>nx239, A0=>a(12), A1=>b(12));
   ix242 : nand02 port map ( Y=>nx241, A0=>b(12), A1=>a(12));
   ix244 : xnor2 port map ( Y=>nx243, A0=>a(13), A1=>b(13));
   ix201 : xnor2 port map ( Y=>sum(14), A0=>nx246, A1=>nx112);
   ix247 : aoi22 port map ( Y=>nx246, A0=>b(13), A1=>a(13), B0=>nx102, B1=>
      nx104);
   ix105 : xnor2 port map ( Y=>nx104, A0=>a(13), A1=>nx249);
   ix250 : inv01 port map ( Y=>nx249, A=>b(13));
   ix113 : xnor2 port map ( Y=>nx112, A0=>a(14), A1=>nx252);
   ix253 : inv01 port map ( Y=>nx252, A=>b(14));
   ix199 : xnor2 port map ( Y=>sum(15), A0=>nx118, A1=>nx260);
   ix119 : oai21 port map ( Y=>nx118, A0=>nx246, A1=>nx256, B0=>nx258);
   ix257 : xnor2 port map ( Y=>nx256, A0=>a(14), A1=>b(14));
   ix259 : nand02 port map ( Y=>nx258, A0=>b(14), A1=>a(14));
   ix261 : xnor2 port map ( Y=>nx260, A0=>a(15), A1=>b(15));
   ix197 : xnor2 port map ( Y=>sum(16), A0=>nx263, A1=>nx128);
   ix264 : aoi22 port map ( Y=>nx263, A0=>b(15), A1=>a(15), B0=>nx118, B1=>
      nx120);
   ix121 : xnor2 port map ( Y=>nx120, A0=>a(15), A1=>nx266);
   ix267 : inv01 port map ( Y=>nx266, A=>b(15));
   ix129 : xnor2 port map ( Y=>nx128, A0=>a(16), A1=>nx269);
   ix270 : inv01 port map ( Y=>nx269, A=>b(16));
   ix195 : xnor2 port map ( Y=>sum(17), A0=>nx134, A1=>nx277);
   ix135 : oai21 port map ( Y=>nx134, A0=>nx263, A1=>nx273, B0=>nx275);
   ix274 : xnor2 port map ( Y=>nx273, A0=>a(16), A1=>b(16));
   ix276 : nand02 port map ( Y=>nx275, A0=>b(16), A1=>a(16));
   ix278 : xnor2 port map ( Y=>nx277, A0=>a(17), A1=>b(17));
   ix193 : xnor2 port map ( Y=>sum(18), A0=>nx280, A1=>nx144);
   ix281 : aoi22 port map ( Y=>nx280, A0=>b(17), A1=>a(17), B0=>nx134, B1=>
      nx136);
   ix137 : xnor2 port map ( Y=>nx136, A0=>a(17), A1=>nx283);
   ix284 : inv01 port map ( Y=>nx283, A=>b(17));
   ix145 : xnor2 port map ( Y=>nx144, A0=>a(18), A1=>nx286);
   ix287 : inv01 port map ( Y=>nx286, A=>b(18));
   ix191 : xnor2 port map ( Y=>sum(19), A0=>nx150, A1=>nx294);
   ix151 : oai21 port map ( Y=>nx150, A0=>nx280, A1=>nx290, B0=>nx292);
   ix291 : xnor2 port map ( Y=>nx290, A0=>a(18), A1=>b(18));
   ix293 : nand02 port map ( Y=>nx292, A0=>b(18), A1=>a(18));
   ix295 : xnor2 port map ( Y=>nx294, A0=>a(19), A1=>b(19));
   ix189 : xnor2 port map ( Y=>sum(20), A0=>nx297, A1=>nx160);
   ix298 : aoi22 port map ( Y=>nx297, A0=>b(19), A1=>a(19), B0=>nx150, B1=>
      nx152);
   ix153 : xnor2 port map ( Y=>nx152, A0=>a(19), A1=>nx300);
   ix301 : inv01 port map ( Y=>nx300, A=>b(19));
   ix161 : xnor2 port map ( Y=>nx160, A0=>a(20), A1=>nx303);
   ix304 : inv01 port map ( Y=>nx303, A=>b(20));
   ix187 : xnor2 port map ( Y=>sum(21), A0=>nx166, A1=>nx311);
   ix167 : oai21 port map ( Y=>nx166, A0=>nx297, A1=>nx307, B0=>nx309);
   ix308 : xnor2 port map ( Y=>nx307, A0=>a(20), A1=>b(20));
   ix310 : nand02 port map ( Y=>nx309, A0=>b(20), A1=>a(20));
   ix312 : xnor2 port map ( Y=>nx311, A0=>a(21), A1=>b(21));
   ix185 : xnor2 port map ( Y=>sum(22), A0=>b(22), A1=>nx314);
   ix315 : aoi22 port map ( Y=>nx314, A0=>b(21), A1=>a(21), B0=>nx166, B1=>
      nx168);
   ix169 : xnor2 port map ( Y=>nx168, A0=>a(21), A1=>nx317);
   ix318 : inv01 port map ( Y=>nx317, A=>b(21));
   ix179 : xnor2 port map ( Y=>sum(23), A0=>b(23), A1=>nx320);
   ix321 : oai21 port map ( Y=>nx320, A0=>nx172, A1=>nx170, B0=>b(22));
   ix173 : nor02_2x port map ( Y=>nx172, A0=>nx317, A1=>nx323);
   ix324 : inv01 port map ( Y=>nx323, A=>a(21));
   ix171 : nor02ii port map ( Y=>nx170, A0=>nx326, A1=>nx168);
   ix327 : aoi22 port map ( Y=>nx326, A0=>b(20), A1=>a(20), B0=>nx158, B1=>
      nx160);
   ix159 : oai21 port map ( Y=>nx158, A0=>nx329, A1=>nx294, B0=>nx372);
   ix330 : aoi22 port map ( Y=>nx329, A0=>b(18), A1=>a(18), B0=>nx142, B1=>
      nx144);
   ix143 : oai21 port map ( Y=>nx142, A0=>nx332, A1=>nx277, B0=>nx370);
   ix333 : aoi22 port map ( Y=>nx332, A0=>b(16), A1=>a(16), B0=>nx126, B1=>
      nx128);
   ix127 : oai21 port map ( Y=>nx126, A0=>nx335, A1=>nx260, B0=>nx368);
   ix336 : aoi22 port map ( Y=>nx335, A0=>b(14), A1=>a(14), B0=>nx110, B1=>
      nx112);
   ix111 : oai21 port map ( Y=>nx110, A0=>nx338, A1=>nx243, B0=>nx366);
   ix339 : aoi22 port map ( Y=>nx338, A0=>b(12), A1=>a(12), B0=>nx94, B1=>
      nx96);
   ix95 : oai21 port map ( Y=>nx94, A0=>nx341, A1=>nx225, B0=>nx364);
   ix342 : aoi22 port map ( Y=>nx341, A0=>b(10), A1=>a(10), B0=>nx78, B1=>
      nx80);
   ix79 : oai21 port map ( Y=>nx78, A0=>nx344, A1=>nx203, B0=>nx362);
   ix345 : aoi22 port map ( Y=>nx344, A0=>b(8), A1=>a(8), B0=>nx62, B1=>nx64
   );
   ix63 : oai21 port map ( Y=>nx62, A0=>nx347, A1=>nx181, B0=>nx360);
   ix348 : aoi22 port map ( Y=>nx347, A0=>b(6), A1=>a(6), B0=>nx46, B1=>nx48
   );
   ix47 : oai21 port map ( Y=>nx46, A0=>nx350, A1=>nx159, B0=>nx358);
   ix351 : aoi22 port map ( Y=>nx350, A0=>b(4), A1=>a(4), B0=>nx30, B1=>nx32
   );
   ix31 : oai21 port map ( Y=>nx30, A0=>nx353, A1=>nx137, B0=>nx356);
   ix354 : aoi21 port map ( Y=>nx353, A0=>b(2), A1=>a(2), B0=>nx18);
   ix19 : nor02ii port map ( Y=>nx18, A0=>nx119, A1=>nx16);
   ix357 : nand02 port map ( Y=>nx356, A0=>b(3), A1=>a(3));
   ix359 : nand02 port map ( Y=>nx358, A0=>b(5), A1=>a(5));
   ix361 : nand02 port map ( Y=>nx360, A0=>b(7), A1=>a(7));
   ix363 : nand02 port map ( Y=>nx362, A0=>b(9), A1=>a(9));
   ix365 : nand02 port map ( Y=>nx364, A0=>b(11), A1=>a(11));
   ix367 : nand02 port map ( Y=>nx366, A0=>b(13), A1=>a(13));
   ix369 : nand02 port map ( Y=>nx368, A0=>b(15), A1=>a(15));
   ix371 : nand02 port map ( Y=>nx370, A0=>b(17), A1=>a(17));
   ix373 : nand02 port map ( Y=>nx372, A0=>b(19), A1=>a(19));
end NBitAdderArch_unfold_2081 ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity CNNMuls_25 is
   port (
      filter_24_7 : IN std_logic ;
      filter_24_6 : IN std_logic ;
      filter_24_5 : IN std_logic ;
      filter_24_4 : IN std_logic ;
      filter_24_3 : IN std_logic ;
      filter_24_2 : IN std_logic ;
      filter_24_1 : IN std_logic ;
      filter_24_0 : IN std_logic ;
      filter_23_7 : IN std_logic ;
      filter_23_6 : IN std_logic ;
      filter_23_5 : IN std_logic ;
      filter_23_4 : IN std_logic ;
      filter_23_3 : IN std_logic ;
      filter_23_2 : IN std_logic ;
      filter_23_1 : IN std_logic ;
      filter_23_0 : IN std_logic ;
      filter_22_7 : IN std_logic ;
      filter_22_6 : IN std_logic ;
      filter_22_5 : IN std_logic ;
      filter_22_4 : IN std_logic ;
      filter_22_3 : IN std_logic ;
      filter_22_2 : IN std_logic ;
      filter_22_1 : IN std_logic ;
      filter_22_0 : IN std_logic ;
      filter_21_7 : IN std_logic ;
      filter_21_6 : IN std_logic ;
      filter_21_5 : IN std_logic ;
      filter_21_4 : IN std_logic ;
      filter_21_3 : IN std_logic ;
      filter_21_2 : IN std_logic ;
      filter_21_1 : IN std_logic ;
      filter_21_0 : IN std_logic ;
      filter_20_7 : IN std_logic ;
      filter_20_6 : IN std_logic ;
      filter_20_5 : IN std_logic ;
      filter_20_4 : IN std_logic ;
      filter_20_3 : IN std_logic ;
      filter_20_2 : IN std_logic ;
      filter_20_1 : IN std_logic ;
      filter_20_0 : IN std_logic ;
      filter_19_7 : IN std_logic ;
      filter_19_6 : IN std_logic ;
      filter_19_5 : IN std_logic ;
      filter_19_4 : IN std_logic ;
      filter_19_3 : IN std_logic ;
      filter_19_2 : IN std_logic ;
      filter_19_1 : IN std_logic ;
      filter_19_0 : IN std_logic ;
      filter_18_7 : IN std_logic ;
      filter_18_6 : IN std_logic ;
      filter_18_5 : IN std_logic ;
      filter_18_4 : IN std_logic ;
      filter_18_3 : IN std_logic ;
      filter_18_2 : IN std_logic ;
      filter_18_1 : IN std_logic ;
      filter_18_0 : IN std_logic ;
      filter_17_7 : IN std_logic ;
      filter_17_6 : IN std_logic ;
      filter_17_5 : IN std_logic ;
      filter_17_4 : IN std_logic ;
      filter_17_3 : IN std_logic ;
      filter_17_2 : IN std_logic ;
      filter_17_1 : IN std_logic ;
      filter_17_0 : IN std_logic ;
      filter_16_7 : IN std_logic ;
      filter_16_6 : IN std_logic ;
      filter_16_5 : IN std_logic ;
      filter_16_4 : IN std_logic ;
      filter_16_3 : IN std_logic ;
      filter_16_2 : IN std_logic ;
      filter_16_1 : IN std_logic ;
      filter_16_0 : IN std_logic ;
      filter_15_7 : IN std_logic ;
      filter_15_6 : IN std_logic ;
      filter_15_5 : IN std_logic ;
      filter_15_4 : IN std_logic ;
      filter_15_3 : IN std_logic ;
      filter_15_2 : IN std_logic ;
      filter_15_1 : IN std_logic ;
      filter_15_0 : IN std_logic ;
      filter_14_7 : IN std_logic ;
      filter_14_6 : IN std_logic ;
      filter_14_5 : IN std_logic ;
      filter_14_4 : IN std_logic ;
      filter_14_3 : IN std_logic ;
      filter_14_2 : IN std_logic ;
      filter_14_1 : IN std_logic ;
      filter_14_0 : IN std_logic ;
      filter_13_7 : IN std_logic ;
      filter_13_6 : IN std_logic ;
      filter_13_5 : IN std_logic ;
      filter_13_4 : IN std_logic ;
      filter_13_3 : IN std_logic ;
      filter_13_2 : IN std_logic ;
      filter_13_1 : IN std_logic ;
      filter_13_0 : IN std_logic ;
      filter_12_7 : IN std_logic ;
      filter_12_6 : IN std_logic ;
      filter_12_5 : IN std_logic ;
      filter_12_4 : IN std_logic ;
      filter_12_3 : IN std_logic ;
      filter_12_2 : IN std_logic ;
      filter_12_1 : IN std_logic ;
      filter_12_0 : IN std_logic ;
      filter_11_7 : IN std_logic ;
      filter_11_6 : IN std_logic ;
      filter_11_5 : IN std_logic ;
      filter_11_4 : IN std_logic ;
      filter_11_3 : IN std_logic ;
      filter_11_2 : IN std_logic ;
      filter_11_1 : IN std_logic ;
      filter_11_0 : IN std_logic ;
      filter_10_7 : IN std_logic ;
      filter_10_6 : IN std_logic ;
      filter_10_5 : IN std_logic ;
      filter_10_4 : IN std_logic ;
      filter_10_3 : IN std_logic ;
      filter_10_2 : IN std_logic ;
      filter_10_1 : IN std_logic ;
      filter_10_0 : IN std_logic ;
      filter_9_7 : IN std_logic ;
      filter_9_6 : IN std_logic ;
      filter_9_5 : IN std_logic ;
      filter_9_4 : IN std_logic ;
      filter_9_3 : IN std_logic ;
      filter_9_2 : IN std_logic ;
      filter_9_1 : IN std_logic ;
      filter_9_0 : IN std_logic ;
      filter_8_7 : IN std_logic ;
      filter_8_6 : IN std_logic ;
      filter_8_5 : IN std_logic ;
      filter_8_4 : IN std_logic ;
      filter_8_3 : IN std_logic ;
      filter_8_2 : IN std_logic ;
      filter_8_1 : IN std_logic ;
      filter_8_0 : IN std_logic ;
      filter_7_7 : IN std_logic ;
      filter_7_6 : IN std_logic ;
      filter_7_5 : IN std_logic ;
      filter_7_4 : IN std_logic ;
      filter_7_3 : IN std_logic ;
      filter_7_2 : IN std_logic ;
      filter_7_1 : IN std_logic ;
      filter_7_0 : IN std_logic ;
      filter_6_7 : IN std_logic ;
      filter_6_6 : IN std_logic ;
      filter_6_5 : IN std_logic ;
      filter_6_4 : IN std_logic ;
      filter_6_3 : IN std_logic ;
      filter_6_2 : IN std_logic ;
      filter_6_1 : IN std_logic ;
      filter_6_0 : IN std_logic ;
      filter_5_7 : IN std_logic ;
      filter_5_6 : IN std_logic ;
      filter_5_5 : IN std_logic ;
      filter_5_4 : IN std_logic ;
      filter_5_3 : IN std_logic ;
      filter_5_2 : IN std_logic ;
      filter_5_1 : IN std_logic ;
      filter_5_0 : IN std_logic ;
      filter_4_7 : IN std_logic ;
      filter_4_6 : IN std_logic ;
      filter_4_5 : IN std_logic ;
      filter_4_4 : IN std_logic ;
      filter_4_3 : IN std_logic ;
      filter_4_2 : IN std_logic ;
      filter_4_1 : IN std_logic ;
      filter_4_0 : IN std_logic ;
      filter_3_7 : IN std_logic ;
      filter_3_6 : IN std_logic ;
      filter_3_5 : IN std_logic ;
      filter_3_4 : IN std_logic ;
      filter_3_3 : IN std_logic ;
      filter_3_2 : IN std_logic ;
      filter_3_1 : IN std_logic ;
      filter_3_0 : IN std_logic ;
      filter_2_7 : IN std_logic ;
      filter_2_6 : IN std_logic ;
      filter_2_5 : IN std_logic ;
      filter_2_4 : IN std_logic ;
      filter_2_3 : IN std_logic ;
      filter_2_2 : IN std_logic ;
      filter_2_1 : IN std_logic ;
      filter_2_0 : IN std_logic ;
      filter_1_7 : IN std_logic ;
      filter_1_6 : IN std_logic ;
      filter_1_5 : IN std_logic ;
      filter_1_4 : IN std_logic ;
      filter_1_3 : IN std_logic ;
      filter_1_2 : IN std_logic ;
      filter_1_1 : IN std_logic ;
      filter_1_0 : IN std_logic ;
      filter_0_7 : IN std_logic ;
      filter_0_6 : IN std_logic ;
      filter_0_5 : IN std_logic ;
      filter_0_4 : IN std_logic ;
      filter_0_3 : IN std_logic ;
      filter_0_2 : IN std_logic ;
      filter_0_1 : IN std_logic ;
      filter_0_0 : IN std_logic ;
      window_24_15 : IN std_logic ;
      window_24_14 : IN std_logic ;
      window_24_13 : IN std_logic ;
      window_24_12 : IN std_logic ;
      window_24_11 : IN std_logic ;
      window_24_10 : IN std_logic ;
      window_24_9 : IN std_logic ;
      window_24_8 : IN std_logic ;
      window_24_7 : IN std_logic ;
      window_24_6 : IN std_logic ;
      window_24_5 : IN std_logic ;
      window_24_4 : IN std_logic ;
      window_24_3 : IN std_logic ;
      window_24_2 : IN std_logic ;
      window_24_1 : IN std_logic ;
      window_24_0 : IN std_logic ;
      window_23_15 : IN std_logic ;
      window_23_14 : IN std_logic ;
      window_23_13 : IN std_logic ;
      window_23_12 : IN std_logic ;
      window_23_11 : IN std_logic ;
      window_23_10 : IN std_logic ;
      window_23_9 : IN std_logic ;
      window_23_8 : IN std_logic ;
      window_23_7 : IN std_logic ;
      window_23_6 : IN std_logic ;
      window_23_5 : IN std_logic ;
      window_23_4 : IN std_logic ;
      window_23_3 : IN std_logic ;
      window_23_2 : IN std_logic ;
      window_23_1 : IN std_logic ;
      window_23_0 : IN std_logic ;
      window_22_15 : IN std_logic ;
      window_22_14 : IN std_logic ;
      window_22_13 : IN std_logic ;
      window_22_12 : IN std_logic ;
      window_22_11 : IN std_logic ;
      window_22_10 : IN std_logic ;
      window_22_9 : IN std_logic ;
      window_22_8 : IN std_logic ;
      window_22_7 : IN std_logic ;
      window_22_6 : IN std_logic ;
      window_22_5 : IN std_logic ;
      window_22_4 : IN std_logic ;
      window_22_3 : IN std_logic ;
      window_22_2 : IN std_logic ;
      window_22_1 : IN std_logic ;
      window_22_0 : IN std_logic ;
      window_21_15 : IN std_logic ;
      window_21_14 : IN std_logic ;
      window_21_13 : IN std_logic ;
      window_21_12 : IN std_logic ;
      window_21_11 : IN std_logic ;
      window_21_10 : IN std_logic ;
      window_21_9 : IN std_logic ;
      window_21_8 : IN std_logic ;
      window_21_7 : IN std_logic ;
      window_21_6 : IN std_logic ;
      window_21_5 : IN std_logic ;
      window_21_4 : IN std_logic ;
      window_21_3 : IN std_logic ;
      window_21_2 : IN std_logic ;
      window_21_1 : IN std_logic ;
      window_21_0 : IN std_logic ;
      window_20_15 : IN std_logic ;
      window_20_14 : IN std_logic ;
      window_20_13 : IN std_logic ;
      window_20_12 : IN std_logic ;
      window_20_11 : IN std_logic ;
      window_20_10 : IN std_logic ;
      window_20_9 : IN std_logic ;
      window_20_8 : IN std_logic ;
      window_20_7 : IN std_logic ;
      window_20_6 : IN std_logic ;
      window_20_5 : IN std_logic ;
      window_20_4 : IN std_logic ;
      window_20_3 : IN std_logic ;
      window_20_2 : IN std_logic ;
      window_20_1 : IN std_logic ;
      window_20_0 : IN std_logic ;
      window_19_15 : IN std_logic ;
      window_19_14 : IN std_logic ;
      window_19_13 : IN std_logic ;
      window_19_12 : IN std_logic ;
      window_19_11 : IN std_logic ;
      window_19_10 : IN std_logic ;
      window_19_9 : IN std_logic ;
      window_19_8 : IN std_logic ;
      window_19_7 : IN std_logic ;
      window_19_6 : IN std_logic ;
      window_19_5 : IN std_logic ;
      window_19_4 : IN std_logic ;
      window_19_3 : IN std_logic ;
      window_19_2 : IN std_logic ;
      window_19_1 : IN std_logic ;
      window_19_0 : IN std_logic ;
      window_18_15 : IN std_logic ;
      window_18_14 : IN std_logic ;
      window_18_13 : IN std_logic ;
      window_18_12 : IN std_logic ;
      window_18_11 : IN std_logic ;
      window_18_10 : IN std_logic ;
      window_18_9 : IN std_logic ;
      window_18_8 : IN std_logic ;
      window_18_7 : IN std_logic ;
      window_18_6 : IN std_logic ;
      window_18_5 : IN std_logic ;
      window_18_4 : IN std_logic ;
      window_18_3 : IN std_logic ;
      window_18_2 : IN std_logic ;
      window_18_1 : IN std_logic ;
      window_18_0 : IN std_logic ;
      window_17_15 : IN std_logic ;
      window_17_14 : IN std_logic ;
      window_17_13 : IN std_logic ;
      window_17_12 : IN std_logic ;
      window_17_11 : IN std_logic ;
      window_17_10 : IN std_logic ;
      window_17_9 : IN std_logic ;
      window_17_8 : IN std_logic ;
      window_17_7 : IN std_logic ;
      window_17_6 : IN std_logic ;
      window_17_5 : IN std_logic ;
      window_17_4 : IN std_logic ;
      window_17_3 : IN std_logic ;
      window_17_2 : IN std_logic ;
      window_17_1 : IN std_logic ;
      window_17_0 : IN std_logic ;
      window_16_15 : IN std_logic ;
      window_16_14 : IN std_logic ;
      window_16_13 : IN std_logic ;
      window_16_12 : IN std_logic ;
      window_16_11 : IN std_logic ;
      window_16_10 : IN std_logic ;
      window_16_9 : IN std_logic ;
      window_16_8 : IN std_logic ;
      window_16_7 : IN std_logic ;
      window_16_6 : IN std_logic ;
      window_16_5 : IN std_logic ;
      window_16_4 : IN std_logic ;
      window_16_3 : IN std_logic ;
      window_16_2 : IN std_logic ;
      window_16_1 : IN std_logic ;
      window_16_0 : IN std_logic ;
      window_15_15 : IN std_logic ;
      window_15_14 : IN std_logic ;
      window_15_13 : IN std_logic ;
      window_15_12 : IN std_logic ;
      window_15_11 : IN std_logic ;
      window_15_10 : IN std_logic ;
      window_15_9 : IN std_logic ;
      window_15_8 : IN std_logic ;
      window_15_7 : IN std_logic ;
      window_15_6 : IN std_logic ;
      window_15_5 : IN std_logic ;
      window_15_4 : IN std_logic ;
      window_15_3 : IN std_logic ;
      window_15_2 : IN std_logic ;
      window_15_1 : IN std_logic ;
      window_15_0 : IN std_logic ;
      window_14_15 : IN std_logic ;
      window_14_14 : IN std_logic ;
      window_14_13 : IN std_logic ;
      window_14_12 : IN std_logic ;
      window_14_11 : IN std_logic ;
      window_14_10 : IN std_logic ;
      window_14_9 : IN std_logic ;
      window_14_8 : IN std_logic ;
      window_14_7 : IN std_logic ;
      window_14_6 : IN std_logic ;
      window_14_5 : IN std_logic ;
      window_14_4 : IN std_logic ;
      window_14_3 : IN std_logic ;
      window_14_2 : IN std_logic ;
      window_14_1 : IN std_logic ;
      window_14_0 : IN std_logic ;
      window_13_15 : IN std_logic ;
      window_13_14 : IN std_logic ;
      window_13_13 : IN std_logic ;
      window_13_12 : IN std_logic ;
      window_13_11 : IN std_logic ;
      window_13_10 : IN std_logic ;
      window_13_9 : IN std_logic ;
      window_13_8 : IN std_logic ;
      window_13_7 : IN std_logic ;
      window_13_6 : IN std_logic ;
      window_13_5 : IN std_logic ;
      window_13_4 : IN std_logic ;
      window_13_3 : IN std_logic ;
      window_13_2 : IN std_logic ;
      window_13_1 : IN std_logic ;
      window_13_0 : IN std_logic ;
      window_12_15 : IN std_logic ;
      window_12_14 : IN std_logic ;
      window_12_13 : IN std_logic ;
      window_12_12 : IN std_logic ;
      window_12_11 : IN std_logic ;
      window_12_10 : IN std_logic ;
      window_12_9 : IN std_logic ;
      window_12_8 : IN std_logic ;
      window_12_7 : IN std_logic ;
      window_12_6 : IN std_logic ;
      window_12_5 : IN std_logic ;
      window_12_4 : IN std_logic ;
      window_12_3 : IN std_logic ;
      window_12_2 : IN std_logic ;
      window_12_1 : IN std_logic ;
      window_12_0 : IN std_logic ;
      window_11_15 : IN std_logic ;
      window_11_14 : IN std_logic ;
      window_11_13 : IN std_logic ;
      window_11_12 : IN std_logic ;
      window_11_11 : IN std_logic ;
      window_11_10 : IN std_logic ;
      window_11_9 : IN std_logic ;
      window_11_8 : IN std_logic ;
      window_11_7 : IN std_logic ;
      window_11_6 : IN std_logic ;
      window_11_5 : IN std_logic ;
      window_11_4 : IN std_logic ;
      window_11_3 : IN std_logic ;
      window_11_2 : IN std_logic ;
      window_11_1 : IN std_logic ;
      window_11_0 : IN std_logic ;
      window_10_15 : IN std_logic ;
      window_10_14 : IN std_logic ;
      window_10_13 : IN std_logic ;
      window_10_12 : IN std_logic ;
      window_10_11 : IN std_logic ;
      window_10_10 : IN std_logic ;
      window_10_9 : IN std_logic ;
      window_10_8 : IN std_logic ;
      window_10_7 : IN std_logic ;
      window_10_6 : IN std_logic ;
      window_10_5 : IN std_logic ;
      window_10_4 : IN std_logic ;
      window_10_3 : IN std_logic ;
      window_10_2 : IN std_logic ;
      window_10_1 : IN std_logic ;
      window_10_0 : IN std_logic ;
      window_9_15 : IN std_logic ;
      window_9_14 : IN std_logic ;
      window_9_13 : IN std_logic ;
      window_9_12 : IN std_logic ;
      window_9_11 : IN std_logic ;
      window_9_10 : IN std_logic ;
      window_9_9 : IN std_logic ;
      window_9_8 : IN std_logic ;
      window_9_7 : IN std_logic ;
      window_9_6 : IN std_logic ;
      window_9_5 : IN std_logic ;
      window_9_4 : IN std_logic ;
      window_9_3 : IN std_logic ;
      window_9_2 : IN std_logic ;
      window_9_1 : IN std_logic ;
      window_9_0 : IN std_logic ;
      window_8_15 : IN std_logic ;
      window_8_14 : IN std_logic ;
      window_8_13 : IN std_logic ;
      window_8_12 : IN std_logic ;
      window_8_11 : IN std_logic ;
      window_8_10 : IN std_logic ;
      window_8_9 : IN std_logic ;
      window_8_8 : IN std_logic ;
      window_8_7 : IN std_logic ;
      window_8_6 : IN std_logic ;
      window_8_5 : IN std_logic ;
      window_8_4 : IN std_logic ;
      window_8_3 : IN std_logic ;
      window_8_2 : IN std_logic ;
      window_8_1 : IN std_logic ;
      window_8_0 : IN std_logic ;
      window_7_15 : IN std_logic ;
      window_7_14 : IN std_logic ;
      window_7_13 : IN std_logic ;
      window_7_12 : IN std_logic ;
      window_7_11 : IN std_logic ;
      window_7_10 : IN std_logic ;
      window_7_9 : IN std_logic ;
      window_7_8 : IN std_logic ;
      window_7_7 : IN std_logic ;
      window_7_6 : IN std_logic ;
      window_7_5 : IN std_logic ;
      window_7_4 : IN std_logic ;
      window_7_3 : IN std_logic ;
      window_7_2 : IN std_logic ;
      window_7_1 : IN std_logic ;
      window_7_0 : IN std_logic ;
      window_6_15 : IN std_logic ;
      window_6_14 : IN std_logic ;
      window_6_13 : IN std_logic ;
      window_6_12 : IN std_logic ;
      window_6_11 : IN std_logic ;
      window_6_10 : IN std_logic ;
      window_6_9 : IN std_logic ;
      window_6_8 : IN std_logic ;
      window_6_7 : IN std_logic ;
      window_6_6 : IN std_logic ;
      window_6_5 : IN std_logic ;
      window_6_4 : IN std_logic ;
      window_6_3 : IN std_logic ;
      window_6_2 : IN std_logic ;
      window_6_1 : IN std_logic ;
      window_6_0 : IN std_logic ;
      window_5_15 : IN std_logic ;
      window_5_14 : IN std_logic ;
      window_5_13 : IN std_logic ;
      window_5_12 : IN std_logic ;
      window_5_11 : IN std_logic ;
      window_5_10 : IN std_logic ;
      window_5_9 : IN std_logic ;
      window_5_8 : IN std_logic ;
      window_5_7 : IN std_logic ;
      window_5_6 : IN std_logic ;
      window_5_5 : IN std_logic ;
      window_5_4 : IN std_logic ;
      window_5_3 : IN std_logic ;
      window_5_2 : IN std_logic ;
      window_5_1 : IN std_logic ;
      window_5_0 : IN std_logic ;
      window_4_15 : IN std_logic ;
      window_4_14 : IN std_logic ;
      window_4_13 : IN std_logic ;
      window_4_12 : IN std_logic ;
      window_4_11 : IN std_logic ;
      window_4_10 : IN std_logic ;
      window_4_9 : IN std_logic ;
      window_4_8 : IN std_logic ;
      window_4_7 : IN std_logic ;
      window_4_6 : IN std_logic ;
      window_4_5 : IN std_logic ;
      window_4_4 : IN std_logic ;
      window_4_3 : IN std_logic ;
      window_4_2 : IN std_logic ;
      window_4_1 : IN std_logic ;
      window_4_0 : IN std_logic ;
      window_3_15 : IN std_logic ;
      window_3_14 : IN std_logic ;
      window_3_13 : IN std_logic ;
      window_3_12 : IN std_logic ;
      window_3_11 : IN std_logic ;
      window_3_10 : IN std_logic ;
      window_3_9 : IN std_logic ;
      window_3_8 : IN std_logic ;
      window_3_7 : IN std_logic ;
      window_3_6 : IN std_logic ;
      window_3_5 : IN std_logic ;
      window_3_4 : IN std_logic ;
      window_3_3 : IN std_logic ;
      window_3_2 : IN std_logic ;
      window_3_1 : IN std_logic ;
      window_3_0 : IN std_logic ;
      window_2_15 : IN std_logic ;
      window_2_14 : IN std_logic ;
      window_2_13 : IN std_logic ;
      window_2_12 : IN std_logic ;
      window_2_11 : IN std_logic ;
      window_2_10 : IN std_logic ;
      window_2_9 : IN std_logic ;
      window_2_8 : IN std_logic ;
      window_2_7 : IN std_logic ;
      window_2_6 : IN std_logic ;
      window_2_5 : IN std_logic ;
      window_2_4 : IN std_logic ;
      window_2_3 : IN std_logic ;
      window_2_2 : IN std_logic ;
      window_2_1 : IN std_logic ;
      window_2_0 : IN std_logic ;
      window_1_15 : IN std_logic ;
      window_1_14 : IN std_logic ;
      window_1_13 : IN std_logic ;
      window_1_12 : IN std_logic ;
      window_1_11 : IN std_logic ;
      window_1_10 : IN std_logic ;
      window_1_9 : IN std_logic ;
      window_1_8 : IN std_logic ;
      window_1_7 : IN std_logic ;
      window_1_6 : IN std_logic ;
      window_1_5 : IN std_logic ;
      window_1_4 : IN std_logic ;
      window_1_3 : IN std_logic ;
      window_1_2 : IN std_logic ;
      window_1_1 : IN std_logic ;
      window_1_0 : IN std_logic ;
      window_0_15 : IN std_logic ;
      window_0_14 : IN std_logic ;
      window_0_13 : IN std_logic ;
      window_0_12 : IN std_logic ;
      window_0_11 : IN std_logic ;
      window_0_10 : IN std_logic ;
      window_0_9 : IN std_logic ;
      window_0_8 : IN std_logic ;
      window_0_7 : IN std_logic ;
      window_0_6 : IN std_logic ;
      window_0_5 : IN std_logic ;
      window_0_4 : IN std_logic ;
      window_0_3 : IN std_logic ;
      window_0_2 : IN std_logic ;
      window_0_1 : IN std_logic ;
      window_0_0 : IN std_logic ;
      outputs_24_15 : INOUT std_logic ;
      outputs_24_14 : INOUT std_logic ;
      outputs_24_13 : INOUT std_logic ;
      outputs_24_12 : INOUT std_logic ;
      outputs_24_11 : INOUT std_logic ;
      outputs_24_10 : INOUT std_logic ;
      outputs_24_9 : INOUT std_logic ;
      outputs_24_8 : INOUT std_logic ;
      outputs_24_7 : INOUT std_logic ;
      outputs_24_6 : INOUT std_logic ;
      outputs_24_5 : INOUT std_logic ;
      outputs_24_4 : INOUT std_logic ;
      outputs_24_3 : INOUT std_logic ;
      outputs_24_2 : INOUT std_logic ;
      outputs_24_1 : INOUT std_logic ;
      outputs_24_0 : INOUT std_logic ;
      outputs_23_15 : INOUT std_logic ;
      outputs_23_14 : INOUT std_logic ;
      outputs_23_13 : INOUT std_logic ;
      outputs_23_12 : INOUT std_logic ;
      outputs_23_11 : INOUT std_logic ;
      outputs_23_10 : INOUT std_logic ;
      outputs_23_9 : INOUT std_logic ;
      outputs_23_8 : INOUT std_logic ;
      outputs_23_7 : INOUT std_logic ;
      outputs_23_6 : INOUT std_logic ;
      outputs_23_5 : INOUT std_logic ;
      outputs_23_4 : INOUT std_logic ;
      outputs_23_3 : INOUT std_logic ;
      outputs_23_2 : INOUT std_logic ;
      outputs_23_1 : INOUT std_logic ;
      outputs_23_0 : INOUT std_logic ;
      outputs_22_15 : INOUT std_logic ;
      outputs_22_14 : INOUT std_logic ;
      outputs_22_13 : INOUT std_logic ;
      outputs_22_12 : INOUT std_logic ;
      outputs_22_11 : INOUT std_logic ;
      outputs_22_10 : INOUT std_logic ;
      outputs_22_9 : INOUT std_logic ;
      outputs_22_8 : INOUT std_logic ;
      outputs_22_7 : INOUT std_logic ;
      outputs_22_6 : INOUT std_logic ;
      outputs_22_5 : INOUT std_logic ;
      outputs_22_4 : INOUT std_logic ;
      outputs_22_3 : INOUT std_logic ;
      outputs_22_2 : INOUT std_logic ;
      outputs_22_1 : INOUT std_logic ;
      outputs_22_0 : INOUT std_logic ;
      outputs_21_15 : INOUT std_logic ;
      outputs_21_14 : INOUT std_logic ;
      outputs_21_13 : INOUT std_logic ;
      outputs_21_12 : INOUT std_logic ;
      outputs_21_11 : INOUT std_logic ;
      outputs_21_10 : INOUT std_logic ;
      outputs_21_9 : INOUT std_logic ;
      outputs_21_8 : INOUT std_logic ;
      outputs_21_7 : INOUT std_logic ;
      outputs_21_6 : INOUT std_logic ;
      outputs_21_5 : INOUT std_logic ;
      outputs_21_4 : INOUT std_logic ;
      outputs_21_3 : INOUT std_logic ;
      outputs_21_2 : INOUT std_logic ;
      outputs_21_1 : INOUT std_logic ;
      outputs_21_0 : INOUT std_logic ;
      outputs_20_15 : INOUT std_logic ;
      outputs_20_14 : INOUT std_logic ;
      outputs_20_13 : INOUT std_logic ;
      outputs_20_12 : INOUT std_logic ;
      outputs_20_11 : INOUT std_logic ;
      outputs_20_10 : INOUT std_logic ;
      outputs_20_9 : INOUT std_logic ;
      outputs_20_8 : INOUT std_logic ;
      outputs_20_7 : INOUT std_logic ;
      outputs_20_6 : INOUT std_logic ;
      outputs_20_5 : INOUT std_logic ;
      outputs_20_4 : INOUT std_logic ;
      outputs_20_3 : INOUT std_logic ;
      outputs_20_2 : INOUT std_logic ;
      outputs_20_1 : INOUT std_logic ;
      outputs_20_0 : INOUT std_logic ;
      outputs_19_15 : INOUT std_logic ;
      outputs_19_14 : INOUT std_logic ;
      outputs_19_13 : INOUT std_logic ;
      outputs_19_12 : INOUT std_logic ;
      outputs_19_11 : INOUT std_logic ;
      outputs_19_10 : INOUT std_logic ;
      outputs_19_9 : INOUT std_logic ;
      outputs_19_8 : INOUT std_logic ;
      outputs_19_7 : INOUT std_logic ;
      outputs_19_6 : INOUT std_logic ;
      outputs_19_5 : INOUT std_logic ;
      outputs_19_4 : INOUT std_logic ;
      outputs_19_3 : INOUT std_logic ;
      outputs_19_2 : INOUT std_logic ;
      outputs_19_1 : INOUT std_logic ;
      outputs_19_0 : INOUT std_logic ;
      outputs_18_15 : INOUT std_logic ;
      outputs_18_14 : INOUT std_logic ;
      outputs_18_13 : INOUT std_logic ;
      outputs_18_12 : INOUT std_logic ;
      outputs_18_11 : INOUT std_logic ;
      outputs_18_10 : INOUT std_logic ;
      outputs_18_9 : INOUT std_logic ;
      outputs_18_8 : INOUT std_logic ;
      outputs_18_7 : INOUT std_logic ;
      outputs_18_6 : INOUT std_logic ;
      outputs_18_5 : INOUT std_logic ;
      outputs_18_4 : INOUT std_logic ;
      outputs_18_3 : INOUT std_logic ;
      outputs_18_2 : INOUT std_logic ;
      outputs_18_1 : INOUT std_logic ;
      outputs_18_0 : INOUT std_logic ;
      outputs_17_15 : INOUT std_logic ;
      outputs_17_14 : INOUT std_logic ;
      outputs_17_13 : INOUT std_logic ;
      outputs_17_12 : INOUT std_logic ;
      outputs_17_11 : INOUT std_logic ;
      outputs_17_10 : INOUT std_logic ;
      outputs_17_9 : INOUT std_logic ;
      outputs_17_8 : INOUT std_logic ;
      outputs_17_7 : INOUT std_logic ;
      outputs_17_6 : INOUT std_logic ;
      outputs_17_5 : INOUT std_logic ;
      outputs_17_4 : INOUT std_logic ;
      outputs_17_3 : INOUT std_logic ;
      outputs_17_2 : INOUT std_logic ;
      outputs_17_1 : INOUT std_logic ;
      outputs_17_0 : INOUT std_logic ;
      outputs_16_15 : INOUT std_logic ;
      outputs_16_14 : INOUT std_logic ;
      outputs_16_13 : INOUT std_logic ;
      outputs_16_12 : INOUT std_logic ;
      outputs_16_11 : INOUT std_logic ;
      outputs_16_10 : INOUT std_logic ;
      outputs_16_9 : INOUT std_logic ;
      outputs_16_8 : INOUT std_logic ;
      outputs_16_7 : INOUT std_logic ;
      outputs_16_6 : INOUT std_logic ;
      outputs_16_5 : INOUT std_logic ;
      outputs_16_4 : INOUT std_logic ;
      outputs_16_3 : INOUT std_logic ;
      outputs_16_2 : INOUT std_logic ;
      outputs_16_1 : INOUT std_logic ;
      outputs_16_0 : INOUT std_logic ;
      outputs_15_15 : INOUT std_logic ;
      outputs_15_14 : INOUT std_logic ;
      outputs_15_13 : INOUT std_logic ;
      outputs_15_12 : INOUT std_logic ;
      outputs_15_11 : INOUT std_logic ;
      outputs_15_10 : INOUT std_logic ;
      outputs_15_9 : INOUT std_logic ;
      outputs_15_8 : INOUT std_logic ;
      outputs_15_7 : INOUT std_logic ;
      outputs_15_6 : INOUT std_logic ;
      outputs_15_5 : INOUT std_logic ;
      outputs_15_4 : INOUT std_logic ;
      outputs_15_3 : INOUT std_logic ;
      outputs_15_2 : INOUT std_logic ;
      outputs_15_1 : INOUT std_logic ;
      outputs_15_0 : INOUT std_logic ;
      outputs_14_15 : INOUT std_logic ;
      outputs_14_14 : INOUT std_logic ;
      outputs_14_13 : INOUT std_logic ;
      outputs_14_12 : INOUT std_logic ;
      outputs_14_11 : INOUT std_logic ;
      outputs_14_10 : INOUT std_logic ;
      outputs_14_9 : INOUT std_logic ;
      outputs_14_8 : INOUT std_logic ;
      outputs_14_7 : INOUT std_logic ;
      outputs_14_6 : INOUT std_logic ;
      outputs_14_5 : INOUT std_logic ;
      outputs_14_4 : INOUT std_logic ;
      outputs_14_3 : INOUT std_logic ;
      outputs_14_2 : INOUT std_logic ;
      outputs_14_1 : INOUT std_logic ;
      outputs_14_0 : INOUT std_logic ;
      outputs_13_15 : INOUT std_logic ;
      outputs_13_14 : INOUT std_logic ;
      outputs_13_13 : INOUT std_logic ;
      outputs_13_12 : INOUT std_logic ;
      outputs_13_11 : INOUT std_logic ;
      outputs_13_10 : INOUT std_logic ;
      outputs_13_9 : INOUT std_logic ;
      outputs_13_8 : INOUT std_logic ;
      outputs_13_7 : INOUT std_logic ;
      outputs_13_6 : INOUT std_logic ;
      outputs_13_5 : INOUT std_logic ;
      outputs_13_4 : INOUT std_logic ;
      outputs_13_3 : INOUT std_logic ;
      outputs_13_2 : INOUT std_logic ;
      outputs_13_1 : INOUT std_logic ;
      outputs_13_0 : INOUT std_logic ;
      outputs_12_15 : INOUT std_logic ;
      outputs_12_14 : INOUT std_logic ;
      outputs_12_13 : INOUT std_logic ;
      outputs_12_12 : INOUT std_logic ;
      outputs_12_11 : INOUT std_logic ;
      outputs_12_10 : INOUT std_logic ;
      outputs_12_9 : INOUT std_logic ;
      outputs_12_8 : INOUT std_logic ;
      outputs_12_7 : INOUT std_logic ;
      outputs_12_6 : INOUT std_logic ;
      outputs_12_5 : INOUT std_logic ;
      outputs_12_4 : INOUT std_logic ;
      outputs_12_3 : INOUT std_logic ;
      outputs_12_2 : INOUT std_logic ;
      outputs_12_1 : INOUT std_logic ;
      outputs_12_0 : INOUT std_logic ;
      outputs_11_15 : INOUT std_logic ;
      outputs_11_14 : INOUT std_logic ;
      outputs_11_13 : INOUT std_logic ;
      outputs_11_12 : INOUT std_logic ;
      outputs_11_11 : INOUT std_logic ;
      outputs_11_10 : INOUT std_logic ;
      outputs_11_9 : INOUT std_logic ;
      outputs_11_8 : INOUT std_logic ;
      outputs_11_7 : INOUT std_logic ;
      outputs_11_6 : INOUT std_logic ;
      outputs_11_5 : INOUT std_logic ;
      outputs_11_4 : INOUT std_logic ;
      outputs_11_3 : INOUT std_logic ;
      outputs_11_2 : INOUT std_logic ;
      outputs_11_1 : INOUT std_logic ;
      outputs_11_0 : INOUT std_logic ;
      outputs_10_15 : INOUT std_logic ;
      outputs_10_14 : INOUT std_logic ;
      outputs_10_13 : INOUT std_logic ;
      outputs_10_12 : INOUT std_logic ;
      outputs_10_11 : INOUT std_logic ;
      outputs_10_10 : INOUT std_logic ;
      outputs_10_9 : INOUT std_logic ;
      outputs_10_8 : INOUT std_logic ;
      outputs_10_7 : INOUT std_logic ;
      outputs_10_6 : INOUT std_logic ;
      outputs_10_5 : INOUT std_logic ;
      outputs_10_4 : INOUT std_logic ;
      outputs_10_3 : INOUT std_logic ;
      outputs_10_2 : INOUT std_logic ;
      outputs_10_1 : INOUT std_logic ;
      outputs_10_0 : INOUT std_logic ;
      outputs_9_15 : INOUT std_logic ;
      outputs_9_14 : INOUT std_logic ;
      outputs_9_13 : INOUT std_logic ;
      outputs_9_12 : INOUT std_logic ;
      outputs_9_11 : INOUT std_logic ;
      outputs_9_10 : INOUT std_logic ;
      outputs_9_9 : INOUT std_logic ;
      outputs_9_8 : INOUT std_logic ;
      outputs_9_7 : INOUT std_logic ;
      outputs_9_6 : INOUT std_logic ;
      outputs_9_5 : INOUT std_logic ;
      outputs_9_4 : INOUT std_logic ;
      outputs_9_3 : INOUT std_logic ;
      outputs_9_2 : INOUT std_logic ;
      outputs_9_1 : INOUT std_logic ;
      outputs_9_0 : INOUT std_logic ;
      outputs_8_15 : INOUT std_logic ;
      outputs_8_14 : INOUT std_logic ;
      outputs_8_13 : INOUT std_logic ;
      outputs_8_12 : INOUT std_logic ;
      outputs_8_11 : INOUT std_logic ;
      outputs_8_10 : INOUT std_logic ;
      outputs_8_9 : INOUT std_logic ;
      outputs_8_8 : INOUT std_logic ;
      outputs_8_7 : INOUT std_logic ;
      outputs_8_6 : INOUT std_logic ;
      outputs_8_5 : INOUT std_logic ;
      outputs_8_4 : INOUT std_logic ;
      outputs_8_3 : INOUT std_logic ;
      outputs_8_2 : INOUT std_logic ;
      outputs_8_1 : INOUT std_logic ;
      outputs_8_0 : INOUT std_logic ;
      outputs_7_15 : INOUT std_logic ;
      outputs_7_14 : INOUT std_logic ;
      outputs_7_13 : INOUT std_logic ;
      outputs_7_12 : INOUT std_logic ;
      outputs_7_11 : INOUT std_logic ;
      outputs_7_10 : INOUT std_logic ;
      outputs_7_9 : INOUT std_logic ;
      outputs_7_8 : INOUT std_logic ;
      outputs_7_7 : INOUT std_logic ;
      outputs_7_6 : INOUT std_logic ;
      outputs_7_5 : INOUT std_logic ;
      outputs_7_4 : INOUT std_logic ;
      outputs_7_3 : INOUT std_logic ;
      outputs_7_2 : INOUT std_logic ;
      outputs_7_1 : INOUT std_logic ;
      outputs_7_0 : INOUT std_logic ;
      outputs_6_15 : INOUT std_logic ;
      outputs_6_14 : INOUT std_logic ;
      outputs_6_13 : INOUT std_logic ;
      outputs_6_12 : INOUT std_logic ;
      outputs_6_11 : INOUT std_logic ;
      outputs_6_10 : INOUT std_logic ;
      outputs_6_9 : INOUT std_logic ;
      outputs_6_8 : INOUT std_logic ;
      outputs_6_7 : INOUT std_logic ;
      outputs_6_6 : INOUT std_logic ;
      outputs_6_5 : INOUT std_logic ;
      outputs_6_4 : INOUT std_logic ;
      outputs_6_3 : INOUT std_logic ;
      outputs_6_2 : INOUT std_logic ;
      outputs_6_1 : INOUT std_logic ;
      outputs_6_0 : INOUT std_logic ;
      outputs_5_15 : INOUT std_logic ;
      outputs_5_14 : INOUT std_logic ;
      outputs_5_13 : INOUT std_logic ;
      outputs_5_12 : INOUT std_logic ;
      outputs_5_11 : INOUT std_logic ;
      outputs_5_10 : INOUT std_logic ;
      outputs_5_9 : INOUT std_logic ;
      outputs_5_8 : INOUT std_logic ;
      outputs_5_7 : INOUT std_logic ;
      outputs_5_6 : INOUT std_logic ;
      outputs_5_5 : INOUT std_logic ;
      outputs_5_4 : INOUT std_logic ;
      outputs_5_3 : INOUT std_logic ;
      outputs_5_2 : INOUT std_logic ;
      outputs_5_1 : INOUT std_logic ;
      outputs_5_0 : INOUT std_logic ;
      outputs_4_15 : INOUT std_logic ;
      outputs_4_14 : INOUT std_logic ;
      outputs_4_13 : INOUT std_logic ;
      outputs_4_12 : INOUT std_logic ;
      outputs_4_11 : INOUT std_logic ;
      outputs_4_10 : INOUT std_logic ;
      outputs_4_9 : INOUT std_logic ;
      outputs_4_8 : INOUT std_logic ;
      outputs_4_7 : INOUT std_logic ;
      outputs_4_6 : INOUT std_logic ;
      outputs_4_5 : INOUT std_logic ;
      outputs_4_4 : INOUT std_logic ;
      outputs_4_3 : INOUT std_logic ;
      outputs_4_2 : INOUT std_logic ;
      outputs_4_1 : INOUT std_logic ;
      outputs_4_0 : INOUT std_logic ;
      outputs_3_15 : INOUT std_logic ;
      outputs_3_14 : INOUT std_logic ;
      outputs_3_13 : INOUT std_logic ;
      outputs_3_12 : INOUT std_logic ;
      outputs_3_11 : INOUT std_logic ;
      outputs_3_10 : INOUT std_logic ;
      outputs_3_9 : INOUT std_logic ;
      outputs_3_8 : INOUT std_logic ;
      outputs_3_7 : INOUT std_logic ;
      outputs_3_6 : INOUT std_logic ;
      outputs_3_5 : INOUT std_logic ;
      outputs_3_4 : INOUT std_logic ;
      outputs_3_3 : INOUT std_logic ;
      outputs_3_2 : INOUT std_logic ;
      outputs_3_1 : INOUT std_logic ;
      outputs_3_0 : INOUT std_logic ;
      outputs_2_15 : INOUT std_logic ;
      outputs_2_14 : INOUT std_logic ;
      outputs_2_13 : INOUT std_logic ;
      outputs_2_12 : INOUT std_logic ;
      outputs_2_11 : INOUT std_logic ;
      outputs_2_10 : INOUT std_logic ;
      outputs_2_9 : INOUT std_logic ;
      outputs_2_8 : INOUT std_logic ;
      outputs_2_7 : INOUT std_logic ;
      outputs_2_6 : INOUT std_logic ;
      outputs_2_5 : INOUT std_logic ;
      outputs_2_4 : INOUT std_logic ;
      outputs_2_3 : INOUT std_logic ;
      outputs_2_2 : INOUT std_logic ;
      outputs_2_1 : INOUT std_logic ;
      outputs_2_0 : INOUT std_logic ;
      outputs_1_15 : INOUT std_logic ;
      outputs_1_14 : INOUT std_logic ;
      outputs_1_13 : INOUT std_logic ;
      outputs_1_12 : INOUT std_logic ;
      outputs_1_11 : INOUT std_logic ;
      outputs_1_10 : INOUT std_logic ;
      outputs_1_9 : INOUT std_logic ;
      outputs_1_8 : INOUT std_logic ;
      outputs_1_7 : INOUT std_logic ;
      outputs_1_6 : INOUT std_logic ;
      outputs_1_5 : INOUT std_logic ;
      outputs_1_4 : INOUT std_logic ;
      outputs_1_3 : INOUT std_logic ;
      outputs_1_2 : INOUT std_logic ;
      outputs_1_1 : INOUT std_logic ;
      outputs_1_0 : INOUT std_logic ;
      outputs_0_15 : INOUT std_logic ;
      outputs_0_14 : INOUT std_logic ;
      outputs_0_13 : INOUT std_logic ;
      outputs_0_12 : INOUT std_logic ;
      outputs_0_11 : INOUT std_logic ;
      outputs_0_10 : INOUT std_logic ;
      outputs_0_9 : INOUT std_logic ;
      outputs_0_8 : INOUT std_logic ;
      outputs_0_7 : INOUT std_logic ;
      outputs_0_6 : INOUT std_logic ;
      outputs_0_5 : INOUT std_logic ;
      outputs_0_4 : INOUT std_logic ;
      outputs_0_3 : INOUT std_logic ;
      outputs_0_2 : INOUT std_logic ;
      outputs_0_1 : INOUT std_logic ;
      outputs_0_0 : INOUT std_logic ;
      clk : IN std_logic ;
      start : IN std_logic ;
      rst : IN std_logic ;
      done : INOUT std_logic ;
      working : INOUT std_logic) ;
end CNNMuls_25 ;

architecture CNNMulsArch_unfold_1782 of CNNMuls_25 is
   component Reg_33
      port (
         D : IN std_logic_vector (32 DOWNTO 0) ;
         en : IN std_logic ;
         clk : IN std_logic ;
         rst : IN std_logic ;
         Q : OUT std_logic_vector (32 DOWNTO 0)) ;
   end component ;
   component BinaryMux_33
      port (
         a : IN std_logic_vector (32 DOWNTO 0) ;
         b : IN std_logic_vector (32 DOWNTO 0) ;
         sel : IN std_logic ;
         f : OUT std_logic_vector (32 DOWNTO 0)) ;
   end component ;
   component NBitAdder_24
      port (
         a : IN std_logic_vector (23 DOWNTO 0) ;
         b : IN std_logic_vector (23 DOWNTO 0) ;
         carryIn : IN std_logic ;
         sum : OUT std_logic_vector (23 DOWNTO 0) ;
         carryOut : OUT std_logic) ;
   end component ;
   signal gen_24_cmp_pBs_30, gen_24_cmp_pBs_29, gen_24_cmp_pBs_28, 
      gen_24_cmp_pBs_27, gen_24_cmp_pBs_26, gen_24_cmp_pBs_25, 
      gen_24_cmp_pBs_24, gen_24_cmp_pBs_23, gen_24_cmp_pMux_30, 
      gen_24_cmp_pMux_29, gen_24_cmp_pMux_28, gen_24_cmp_pMux_27, 
      gen_24_cmp_pMux_26, gen_24_cmp_pMux_25, gen_24_cmp_pMux_24, 
      gen_24_cmp_pMux_23, gen_24_cmp_pMux_22, gen_24_cmp_pMux_21, 
      gen_24_cmp_pMux_20, gen_24_cmp_pMux_19, gen_24_cmp_pMux_18, 
      gen_24_cmp_pMux_17, gen_24_cmp_pMux_16, gen_24_cmp_pMux_15, 
      gen_24_cmp_pMux_14, gen_24_cmp_pMux_13, gen_24_cmp_pMux_12, 
      gen_24_cmp_pMux_11, gen_24_cmp_pMux_10, gen_24_cmp_pMux_9, 
      gen_24_cmp_pMux_8, gen_24_cmp_pMux_7, gen_24_cmp_pMux_6, 
      gen_24_cmp_pMux_5, gen_24_cmp_pMux_4, gen_24_cmp_pMux_3, 
      gen_24_cmp_pMux_2, gen_24_cmp_pMux_1, gen_24_cmp_pMux_0, 
      gen_24_cmp_pReg_30, gen_24_cmp_pReg_29, gen_24_cmp_pReg_28, 
      gen_24_cmp_pReg_27, gen_24_cmp_pReg_26, gen_24_cmp_pReg_25, 
      gen_24_cmp_pReg_24, gen_24_cmp_pReg_23, gen_24_cmp_pReg_22, 
      gen_24_cmp_pReg_21, gen_24_cmp_pReg_20, gen_24_cmp_pReg_19, 
      gen_24_cmp_pReg_18, gen_24_cmp_pReg_17, gen_24_cmp_pReg_16, 
      gen_24_cmp_pReg_15, gen_24_cmp_pReg_14, gen_24_cmp_pReg_13, 
      gen_24_cmp_pReg_12, gen_24_cmp_pReg_11, gen_24_cmp_pReg_10, 
      gen_24_cmp_pReg_9, gen_24_cmp_pReg_8, gen_24_cmp_pReg_7, 
      gen_24_cmp_pReg_6, gen_24_cmp_pReg_5, gen_24_cmp_pReg_4, 
      gen_24_cmp_pReg_3, gen_24_cmp_pReg_2, gen_24_cmp_pReg_1, 
      gen_24_cmp_pReg_0, gen_24_cmp_BSCmp_op2_0, gen_24_cmp_BSCmp_carryIn, 
      gen_23_cmp_pBs_30, gen_23_cmp_pBs_29, gen_23_cmp_pBs_28, 
      gen_23_cmp_pBs_27, gen_23_cmp_pBs_26, gen_23_cmp_pBs_25, 
      gen_23_cmp_pBs_24, gen_23_cmp_pBs_23, gen_23_cmp_pMux_30, 
      gen_23_cmp_pMux_29, gen_23_cmp_pMux_28, gen_23_cmp_pMux_27, 
      gen_23_cmp_pMux_26, gen_23_cmp_pMux_25, gen_23_cmp_pMux_24, 
      gen_23_cmp_pMux_23, gen_23_cmp_pMux_22, gen_23_cmp_pMux_21, 
      gen_23_cmp_pMux_20, gen_23_cmp_pMux_19, gen_23_cmp_pMux_18, 
      gen_23_cmp_pMux_17, gen_23_cmp_pMux_16, gen_23_cmp_pMux_15, 
      gen_23_cmp_pMux_14, gen_23_cmp_pMux_13, gen_23_cmp_pMux_12, 
      gen_23_cmp_pMux_11, gen_23_cmp_pMux_10, gen_23_cmp_pMux_9, 
      gen_23_cmp_pMux_8, gen_23_cmp_pMux_7, gen_23_cmp_pMux_6, 
      gen_23_cmp_pMux_5, gen_23_cmp_pMux_4, gen_23_cmp_pMux_3, 
      gen_23_cmp_pMux_2, gen_23_cmp_pMux_1, gen_23_cmp_pMux_0, 
      gen_23_cmp_pReg_30, gen_23_cmp_pReg_29, gen_23_cmp_pReg_28, 
      gen_23_cmp_pReg_27, gen_23_cmp_pReg_26, gen_23_cmp_pReg_25, 
      gen_23_cmp_pReg_24, gen_23_cmp_pReg_23, gen_23_cmp_pReg_22, 
      gen_23_cmp_pReg_21, gen_23_cmp_pReg_20, gen_23_cmp_pReg_19, 
      gen_23_cmp_pReg_18, gen_23_cmp_pReg_17, gen_23_cmp_pReg_16, 
      gen_23_cmp_pReg_15, gen_23_cmp_pReg_14, gen_23_cmp_pReg_13, 
      gen_23_cmp_pReg_12, gen_23_cmp_pReg_11, gen_23_cmp_pReg_10, 
      gen_23_cmp_pReg_9, gen_23_cmp_pReg_8, gen_23_cmp_pReg_7, 
      gen_23_cmp_pReg_6, gen_23_cmp_pReg_5, gen_23_cmp_pReg_4, 
      gen_23_cmp_pReg_3, gen_23_cmp_pReg_2, gen_23_cmp_pReg_1, 
      gen_23_cmp_pReg_0, gen_23_cmp_BSCmp_op2_0, gen_23_cmp_BSCmp_carryIn, 
      gen_22_cmp_pBs_30, gen_22_cmp_pBs_29, gen_22_cmp_pBs_28, 
      gen_22_cmp_pBs_27, gen_22_cmp_pBs_26, gen_22_cmp_pBs_25, 
      gen_22_cmp_pBs_24, gen_22_cmp_pBs_23, gen_22_cmp_pMux_30, 
      gen_22_cmp_pMux_29, gen_22_cmp_pMux_28, gen_22_cmp_pMux_27, 
      gen_22_cmp_pMux_26, gen_22_cmp_pMux_25, gen_22_cmp_pMux_24, 
      gen_22_cmp_pMux_23, gen_22_cmp_pMux_22, gen_22_cmp_pMux_21, 
      gen_22_cmp_pMux_20, gen_22_cmp_pMux_19, gen_22_cmp_pMux_18, 
      gen_22_cmp_pMux_17, gen_22_cmp_pMux_16, gen_22_cmp_pMux_15, 
      gen_22_cmp_pMux_14, gen_22_cmp_pMux_13, gen_22_cmp_pMux_12, 
      gen_22_cmp_pMux_11, gen_22_cmp_pMux_10, gen_22_cmp_pMux_9, 
      gen_22_cmp_pMux_8, gen_22_cmp_pMux_7, gen_22_cmp_pMux_6, 
      gen_22_cmp_pMux_5, gen_22_cmp_pMux_4, gen_22_cmp_pMux_3, 
      gen_22_cmp_pMux_2, gen_22_cmp_pMux_1, gen_22_cmp_pMux_0, 
      gen_22_cmp_pReg_30, gen_22_cmp_pReg_29, gen_22_cmp_pReg_28, 
      gen_22_cmp_pReg_27, gen_22_cmp_pReg_26, gen_22_cmp_pReg_25, 
      gen_22_cmp_pReg_24, gen_22_cmp_pReg_23, gen_22_cmp_pReg_22, 
      gen_22_cmp_pReg_21, gen_22_cmp_pReg_20, gen_22_cmp_pReg_19, 
      gen_22_cmp_pReg_18, gen_22_cmp_pReg_17, gen_22_cmp_pReg_16, 
      gen_22_cmp_pReg_15, gen_22_cmp_pReg_14, gen_22_cmp_pReg_13, 
      gen_22_cmp_pReg_12, gen_22_cmp_pReg_11, gen_22_cmp_pReg_10, 
      gen_22_cmp_pReg_9, gen_22_cmp_pReg_8, gen_22_cmp_pReg_7, 
      gen_22_cmp_pReg_6, gen_22_cmp_pReg_5, gen_22_cmp_pReg_4, 
      gen_22_cmp_pReg_3, gen_22_cmp_pReg_2, gen_22_cmp_pReg_1, 
      gen_22_cmp_pReg_0, gen_22_cmp_BSCmp_op2_0, gen_22_cmp_BSCmp_carryIn, 
      gen_21_cmp_pBs_30, gen_21_cmp_pBs_29, gen_21_cmp_pBs_28, 
      gen_21_cmp_pBs_27, gen_21_cmp_pBs_26, gen_21_cmp_pBs_25, 
      gen_21_cmp_pBs_24, gen_21_cmp_pBs_23, gen_21_cmp_pMux_30, 
      gen_21_cmp_pMux_29, gen_21_cmp_pMux_28, gen_21_cmp_pMux_27, 
      gen_21_cmp_pMux_26, gen_21_cmp_pMux_25, gen_21_cmp_pMux_24, 
      gen_21_cmp_pMux_23, gen_21_cmp_pMux_22, gen_21_cmp_pMux_21, 
      gen_21_cmp_pMux_20, gen_21_cmp_pMux_19, gen_21_cmp_pMux_18, 
      gen_21_cmp_pMux_17, gen_21_cmp_pMux_16, gen_21_cmp_pMux_15, 
      gen_21_cmp_pMux_14, gen_21_cmp_pMux_13, gen_21_cmp_pMux_12, 
      gen_21_cmp_pMux_11, gen_21_cmp_pMux_10, gen_21_cmp_pMux_9, 
      gen_21_cmp_pMux_8, gen_21_cmp_pMux_7, gen_21_cmp_pMux_6, 
      gen_21_cmp_pMux_5, gen_21_cmp_pMux_4, gen_21_cmp_pMux_3, 
      gen_21_cmp_pMux_2, gen_21_cmp_pMux_1, gen_21_cmp_pMux_0, 
      gen_21_cmp_pReg_30, gen_21_cmp_pReg_29, gen_21_cmp_pReg_28, 
      gen_21_cmp_pReg_27, gen_21_cmp_pReg_26, gen_21_cmp_pReg_25, 
      gen_21_cmp_pReg_24, gen_21_cmp_pReg_23, gen_21_cmp_pReg_22, 
      gen_21_cmp_pReg_21, gen_21_cmp_pReg_20, gen_21_cmp_pReg_19, 
      gen_21_cmp_pReg_18, gen_21_cmp_pReg_17, gen_21_cmp_pReg_16, 
      gen_21_cmp_pReg_15, gen_21_cmp_pReg_14, gen_21_cmp_pReg_13, 
      gen_21_cmp_pReg_12, gen_21_cmp_pReg_11, gen_21_cmp_pReg_10, 
      gen_21_cmp_pReg_9, gen_21_cmp_pReg_8, gen_21_cmp_pReg_7, 
      gen_21_cmp_pReg_6, gen_21_cmp_pReg_5, gen_21_cmp_pReg_4, 
      gen_21_cmp_pReg_3, gen_21_cmp_pReg_2, gen_21_cmp_pReg_1, 
      gen_21_cmp_pReg_0, gen_21_cmp_BSCmp_op2_0, gen_21_cmp_BSCmp_carryIn, 
      gen_20_cmp_pBs_30, gen_20_cmp_pBs_29, gen_20_cmp_pBs_28, 
      gen_20_cmp_pBs_27, gen_20_cmp_pBs_26, gen_20_cmp_pBs_25, 
      gen_20_cmp_pBs_24, gen_20_cmp_pBs_23, gen_20_cmp_pMux_30, 
      gen_20_cmp_pMux_29, gen_20_cmp_pMux_28, gen_20_cmp_pMux_27, 
      gen_20_cmp_pMux_26, gen_20_cmp_pMux_25, gen_20_cmp_pMux_24, 
      gen_20_cmp_pMux_23, gen_20_cmp_pMux_22, gen_20_cmp_pMux_21, 
      gen_20_cmp_pMux_20, gen_20_cmp_pMux_19, gen_20_cmp_pMux_18, 
      gen_20_cmp_pMux_17, gen_20_cmp_pMux_16, gen_20_cmp_pMux_15, 
      gen_20_cmp_pMux_14, gen_20_cmp_pMux_13, gen_20_cmp_pMux_12, 
      gen_20_cmp_pMux_11, gen_20_cmp_pMux_10, gen_20_cmp_pMux_9, 
      gen_20_cmp_pMux_8, gen_20_cmp_pMux_7, gen_20_cmp_pMux_6, 
      gen_20_cmp_pMux_5, gen_20_cmp_pMux_4, gen_20_cmp_pMux_3, 
      gen_20_cmp_pMux_2, gen_20_cmp_pMux_1, gen_20_cmp_pMux_0, 
      gen_20_cmp_pReg_30, gen_20_cmp_pReg_29, gen_20_cmp_pReg_28, 
      gen_20_cmp_pReg_27, gen_20_cmp_pReg_26, gen_20_cmp_pReg_25, 
      gen_20_cmp_pReg_24, gen_20_cmp_pReg_23, gen_20_cmp_pReg_22, 
      gen_20_cmp_pReg_21, gen_20_cmp_pReg_20, gen_20_cmp_pReg_19, 
      gen_20_cmp_pReg_18, gen_20_cmp_pReg_17, gen_20_cmp_pReg_16, 
      gen_20_cmp_pReg_15, gen_20_cmp_pReg_14, gen_20_cmp_pReg_13, 
      gen_20_cmp_pReg_12, gen_20_cmp_pReg_11, gen_20_cmp_pReg_10, 
      gen_20_cmp_pReg_9, gen_20_cmp_pReg_8, gen_20_cmp_pReg_7, 
      gen_20_cmp_pReg_6, gen_20_cmp_pReg_5, gen_20_cmp_pReg_4, 
      gen_20_cmp_pReg_3, gen_20_cmp_pReg_2, gen_20_cmp_pReg_1, 
      gen_20_cmp_pReg_0, gen_20_cmp_BSCmp_op2_0, gen_20_cmp_BSCmp_carryIn, 
      gen_19_cmp_pBs_30, gen_19_cmp_pBs_29, gen_19_cmp_pBs_28, 
      gen_19_cmp_pBs_27, gen_19_cmp_pBs_26, gen_19_cmp_pBs_25, 
      gen_19_cmp_pBs_24, gen_19_cmp_pBs_23, gen_19_cmp_pMux_30, 
      gen_19_cmp_pMux_29, gen_19_cmp_pMux_28, gen_19_cmp_pMux_27, 
      gen_19_cmp_pMux_26, gen_19_cmp_pMux_25, gen_19_cmp_pMux_24, 
      gen_19_cmp_pMux_23, gen_19_cmp_pMux_22, gen_19_cmp_pMux_21, 
      gen_19_cmp_pMux_20, gen_19_cmp_pMux_19, gen_19_cmp_pMux_18, 
      gen_19_cmp_pMux_17, gen_19_cmp_pMux_16, gen_19_cmp_pMux_15, 
      gen_19_cmp_pMux_14, gen_19_cmp_pMux_13, gen_19_cmp_pMux_12, 
      gen_19_cmp_pMux_11, gen_19_cmp_pMux_10, gen_19_cmp_pMux_9, 
      gen_19_cmp_pMux_8, gen_19_cmp_pMux_7, gen_19_cmp_pMux_6, 
      gen_19_cmp_pMux_5, gen_19_cmp_pMux_4, gen_19_cmp_pMux_3, 
      gen_19_cmp_pMux_2, gen_19_cmp_pMux_1, gen_19_cmp_pMux_0, 
      gen_19_cmp_pReg_30, gen_19_cmp_pReg_29, gen_19_cmp_pReg_28, 
      gen_19_cmp_pReg_27, gen_19_cmp_pReg_26, gen_19_cmp_pReg_25, 
      gen_19_cmp_pReg_24, gen_19_cmp_pReg_23, gen_19_cmp_pReg_22, 
      gen_19_cmp_pReg_21, gen_19_cmp_pReg_20, gen_19_cmp_pReg_19, 
      gen_19_cmp_pReg_18, gen_19_cmp_pReg_17, gen_19_cmp_pReg_16, 
      gen_19_cmp_pReg_15, gen_19_cmp_pReg_14, gen_19_cmp_pReg_13, 
      gen_19_cmp_pReg_12, gen_19_cmp_pReg_11, gen_19_cmp_pReg_10, 
      gen_19_cmp_pReg_9, gen_19_cmp_pReg_8, gen_19_cmp_pReg_7, 
      gen_19_cmp_pReg_6, gen_19_cmp_pReg_5, gen_19_cmp_pReg_4, 
      gen_19_cmp_pReg_3, gen_19_cmp_pReg_2, gen_19_cmp_pReg_1, 
      gen_19_cmp_pReg_0, gen_19_cmp_BSCmp_op2_0, gen_19_cmp_BSCmp_carryIn, 
      gen_18_cmp_pBs_30, gen_18_cmp_pBs_29, gen_18_cmp_pBs_28, 
      gen_18_cmp_pBs_27, gen_18_cmp_pBs_26, gen_18_cmp_pBs_25, 
      gen_18_cmp_pBs_24, gen_18_cmp_pBs_23, gen_18_cmp_pMux_30, 
      gen_18_cmp_pMux_29, gen_18_cmp_pMux_28, gen_18_cmp_pMux_27, 
      gen_18_cmp_pMux_26, gen_18_cmp_pMux_25, gen_18_cmp_pMux_24, 
      gen_18_cmp_pMux_23, gen_18_cmp_pMux_22, gen_18_cmp_pMux_21, 
      gen_18_cmp_pMux_20, gen_18_cmp_pMux_19, gen_18_cmp_pMux_18, 
      gen_18_cmp_pMux_17, gen_18_cmp_pMux_16, gen_18_cmp_pMux_15, 
      gen_18_cmp_pMux_14, gen_18_cmp_pMux_13, gen_18_cmp_pMux_12, 
      gen_18_cmp_pMux_11, gen_18_cmp_pMux_10, gen_18_cmp_pMux_9, 
      gen_18_cmp_pMux_8, gen_18_cmp_pMux_7, gen_18_cmp_pMux_6, 
      gen_18_cmp_pMux_5, gen_18_cmp_pMux_4, gen_18_cmp_pMux_3, 
      gen_18_cmp_pMux_2, gen_18_cmp_pMux_1, gen_18_cmp_pMux_0, 
      gen_18_cmp_pReg_30, gen_18_cmp_pReg_29, gen_18_cmp_pReg_28, 
      gen_18_cmp_pReg_27, gen_18_cmp_pReg_26, gen_18_cmp_pReg_25, 
      gen_18_cmp_pReg_24, gen_18_cmp_pReg_23, gen_18_cmp_pReg_22, 
      gen_18_cmp_pReg_21, gen_18_cmp_pReg_20, gen_18_cmp_pReg_19, 
      gen_18_cmp_pReg_18, gen_18_cmp_pReg_17, gen_18_cmp_pReg_16, 
      gen_18_cmp_pReg_15, gen_18_cmp_pReg_14, gen_18_cmp_pReg_13, 
      gen_18_cmp_pReg_12, gen_18_cmp_pReg_11, gen_18_cmp_pReg_10, 
      gen_18_cmp_pReg_9, gen_18_cmp_pReg_8, gen_18_cmp_pReg_7, 
      gen_18_cmp_pReg_6, gen_18_cmp_pReg_5, gen_18_cmp_pReg_4, 
      gen_18_cmp_pReg_3, gen_18_cmp_pReg_2, gen_18_cmp_pReg_1, 
      gen_18_cmp_pReg_0, gen_18_cmp_BSCmp_op2_0, gen_18_cmp_BSCmp_carryIn, 
      gen_17_cmp_pBs_30, gen_17_cmp_pBs_29, gen_17_cmp_pBs_28, 
      gen_17_cmp_pBs_27, gen_17_cmp_pBs_26, gen_17_cmp_pBs_25, 
      gen_17_cmp_pBs_24, gen_17_cmp_pBs_23, gen_17_cmp_pMux_30, 
      gen_17_cmp_pMux_29, gen_17_cmp_pMux_28, gen_17_cmp_pMux_27, 
      gen_17_cmp_pMux_26, gen_17_cmp_pMux_25, gen_17_cmp_pMux_24, 
      gen_17_cmp_pMux_23, gen_17_cmp_pMux_22, gen_17_cmp_pMux_21, 
      gen_17_cmp_pMux_20, gen_17_cmp_pMux_19, gen_17_cmp_pMux_18, 
      gen_17_cmp_pMux_17, gen_17_cmp_pMux_16, gen_17_cmp_pMux_15, 
      gen_17_cmp_pMux_14, gen_17_cmp_pMux_13, gen_17_cmp_pMux_12, 
      gen_17_cmp_pMux_11, gen_17_cmp_pMux_10, gen_17_cmp_pMux_9, 
      gen_17_cmp_pMux_8, gen_17_cmp_pMux_7, gen_17_cmp_pMux_6, 
      gen_17_cmp_pMux_5, gen_17_cmp_pMux_4, gen_17_cmp_pMux_3, 
      gen_17_cmp_pMux_2, gen_17_cmp_pMux_1, gen_17_cmp_pMux_0, 
      gen_17_cmp_pReg_30, gen_17_cmp_pReg_29, gen_17_cmp_pReg_28, 
      gen_17_cmp_pReg_27, gen_17_cmp_pReg_26, gen_17_cmp_pReg_25, 
      gen_17_cmp_pReg_24, gen_17_cmp_pReg_23, gen_17_cmp_pReg_22, 
      gen_17_cmp_pReg_21, gen_17_cmp_pReg_20, gen_17_cmp_pReg_19, 
      gen_17_cmp_pReg_18, gen_17_cmp_pReg_17, gen_17_cmp_pReg_16, 
      gen_17_cmp_pReg_15, gen_17_cmp_pReg_14, gen_17_cmp_pReg_13, 
      gen_17_cmp_pReg_12, gen_17_cmp_pReg_11, gen_17_cmp_pReg_10, 
      gen_17_cmp_pReg_9, gen_17_cmp_pReg_8, gen_17_cmp_pReg_7, 
      gen_17_cmp_pReg_6, gen_17_cmp_pReg_5, gen_17_cmp_pReg_4, 
      gen_17_cmp_pReg_3, gen_17_cmp_pReg_2, gen_17_cmp_pReg_1, 
      gen_17_cmp_pReg_0, gen_17_cmp_BSCmp_op2_0, gen_17_cmp_BSCmp_carryIn, 
      gen_16_cmp_pBs_30, gen_16_cmp_pBs_29, gen_16_cmp_pBs_28, 
      gen_16_cmp_pBs_27, gen_16_cmp_pBs_26, gen_16_cmp_pBs_25, 
      gen_16_cmp_pBs_24, gen_16_cmp_pBs_23, gen_16_cmp_pMux_30, 
      gen_16_cmp_pMux_29, gen_16_cmp_pMux_28, gen_16_cmp_pMux_27, 
      gen_16_cmp_pMux_26, gen_16_cmp_pMux_25, gen_16_cmp_pMux_24, 
      gen_16_cmp_pMux_23, gen_16_cmp_pMux_22, gen_16_cmp_pMux_21, 
      gen_16_cmp_pMux_20, gen_16_cmp_pMux_19, gen_16_cmp_pMux_18, 
      gen_16_cmp_pMux_17, gen_16_cmp_pMux_16, gen_16_cmp_pMux_15, 
      gen_16_cmp_pMux_14, gen_16_cmp_pMux_13, gen_16_cmp_pMux_12, 
      gen_16_cmp_pMux_11, gen_16_cmp_pMux_10, gen_16_cmp_pMux_9, 
      gen_16_cmp_pMux_8, gen_16_cmp_pMux_7, gen_16_cmp_pMux_6, 
      gen_16_cmp_pMux_5, gen_16_cmp_pMux_4, gen_16_cmp_pMux_3, 
      gen_16_cmp_pMux_2, gen_16_cmp_pMux_1, gen_16_cmp_pMux_0, 
      gen_16_cmp_pReg_30, gen_16_cmp_pReg_29, gen_16_cmp_pReg_28, 
      gen_16_cmp_pReg_27, gen_16_cmp_pReg_26, gen_16_cmp_pReg_25, 
      gen_16_cmp_pReg_24, gen_16_cmp_pReg_23, gen_16_cmp_pReg_22, 
      gen_16_cmp_pReg_21, gen_16_cmp_pReg_20, gen_16_cmp_pReg_19, 
      gen_16_cmp_pReg_18, gen_16_cmp_pReg_17, gen_16_cmp_pReg_16, 
      gen_16_cmp_pReg_15, gen_16_cmp_pReg_14, gen_16_cmp_pReg_13, 
      gen_16_cmp_pReg_12, gen_16_cmp_pReg_11, gen_16_cmp_pReg_10, 
      gen_16_cmp_pReg_9, gen_16_cmp_pReg_8, gen_16_cmp_pReg_7, 
      gen_16_cmp_pReg_6, gen_16_cmp_pReg_5, gen_16_cmp_pReg_4, 
      gen_16_cmp_pReg_3, gen_16_cmp_pReg_2, gen_16_cmp_pReg_1, 
      gen_16_cmp_pReg_0, gen_16_cmp_BSCmp_op2_0, gen_16_cmp_BSCmp_carryIn, 
      gen_15_cmp_pBs_30, gen_15_cmp_pBs_29, gen_15_cmp_pBs_28, 
      gen_15_cmp_pBs_27, gen_15_cmp_pBs_26, gen_15_cmp_pBs_25, 
      gen_15_cmp_pBs_24, gen_15_cmp_pBs_23, gen_15_cmp_pMux_30, 
      gen_15_cmp_pMux_29, gen_15_cmp_pMux_28, gen_15_cmp_pMux_27, 
      gen_15_cmp_pMux_26, gen_15_cmp_pMux_25, gen_15_cmp_pMux_24, 
      gen_15_cmp_pMux_23, gen_15_cmp_pMux_22, gen_15_cmp_pMux_21, 
      gen_15_cmp_pMux_20, gen_15_cmp_pMux_19, gen_15_cmp_pMux_18, 
      gen_15_cmp_pMux_17, gen_15_cmp_pMux_16, gen_15_cmp_pMux_15, 
      gen_15_cmp_pMux_14, gen_15_cmp_pMux_13, gen_15_cmp_pMux_12, 
      gen_15_cmp_pMux_11, gen_15_cmp_pMux_10, gen_15_cmp_pMux_9, 
      gen_15_cmp_pMux_8, gen_15_cmp_pMux_7, gen_15_cmp_pMux_6, 
      gen_15_cmp_pMux_5, gen_15_cmp_pMux_4, gen_15_cmp_pMux_3, 
      gen_15_cmp_pMux_2, gen_15_cmp_pMux_1, gen_15_cmp_pMux_0, 
      gen_15_cmp_pReg_30, gen_15_cmp_pReg_29, gen_15_cmp_pReg_28, 
      gen_15_cmp_pReg_27, gen_15_cmp_pReg_26, gen_15_cmp_pReg_25, 
      gen_15_cmp_pReg_24, gen_15_cmp_pReg_23, gen_15_cmp_pReg_22, 
      gen_15_cmp_pReg_21, gen_15_cmp_pReg_20, gen_15_cmp_pReg_19, 
      gen_15_cmp_pReg_18, gen_15_cmp_pReg_17, gen_15_cmp_pReg_16, 
      gen_15_cmp_pReg_15, gen_15_cmp_pReg_14, gen_15_cmp_pReg_13, 
      gen_15_cmp_pReg_12, gen_15_cmp_pReg_11, gen_15_cmp_pReg_10, 
      gen_15_cmp_pReg_9, gen_15_cmp_pReg_8, gen_15_cmp_pReg_7, 
      gen_15_cmp_pReg_6, gen_15_cmp_pReg_5, gen_15_cmp_pReg_4, 
      gen_15_cmp_pReg_3, gen_15_cmp_pReg_2, gen_15_cmp_pReg_1, 
      gen_15_cmp_pReg_0, gen_15_cmp_BSCmp_op2_0, gen_15_cmp_BSCmp_carryIn, 
      gen_14_cmp_pBs_30, gen_14_cmp_pBs_29, gen_14_cmp_pBs_28, 
      gen_14_cmp_pBs_27, gen_14_cmp_pBs_26, gen_14_cmp_pBs_25, 
      gen_14_cmp_pBs_24, gen_14_cmp_pBs_23, gen_14_cmp_pMux_30, 
      gen_14_cmp_pMux_29, gen_14_cmp_pMux_28, gen_14_cmp_pMux_27, 
      gen_14_cmp_pMux_26, gen_14_cmp_pMux_25, gen_14_cmp_pMux_24, 
      gen_14_cmp_pMux_23, gen_14_cmp_pMux_22, gen_14_cmp_pMux_21, 
      gen_14_cmp_pMux_20, gen_14_cmp_pMux_19, gen_14_cmp_pMux_18, 
      gen_14_cmp_pMux_17, gen_14_cmp_pMux_16, gen_14_cmp_pMux_15, 
      gen_14_cmp_pMux_14, gen_14_cmp_pMux_13, gen_14_cmp_pMux_12, 
      gen_14_cmp_pMux_11, gen_14_cmp_pMux_10, gen_14_cmp_pMux_9, 
      gen_14_cmp_pMux_8, gen_14_cmp_pMux_7, gen_14_cmp_pMux_6, 
      gen_14_cmp_pMux_5, gen_14_cmp_pMux_4, gen_14_cmp_pMux_3, 
      gen_14_cmp_pMux_2, gen_14_cmp_pMux_1, gen_14_cmp_pMux_0, 
      gen_14_cmp_pReg_30, gen_14_cmp_pReg_29, gen_14_cmp_pReg_28, 
      gen_14_cmp_pReg_27, gen_14_cmp_pReg_26, gen_14_cmp_pReg_25, 
      gen_14_cmp_pReg_24, gen_14_cmp_pReg_23, gen_14_cmp_pReg_22, 
      gen_14_cmp_pReg_21, gen_14_cmp_pReg_20, gen_14_cmp_pReg_19, 
      gen_14_cmp_pReg_18, gen_14_cmp_pReg_17, gen_14_cmp_pReg_16, 
      gen_14_cmp_pReg_15, gen_14_cmp_pReg_14, gen_14_cmp_pReg_13, 
      gen_14_cmp_pReg_12, gen_14_cmp_pReg_11, gen_14_cmp_pReg_10, 
      gen_14_cmp_pReg_9, gen_14_cmp_pReg_8, gen_14_cmp_pReg_7, 
      gen_14_cmp_pReg_6, gen_14_cmp_pReg_5, gen_14_cmp_pReg_4, 
      gen_14_cmp_pReg_3, gen_14_cmp_pReg_2, gen_14_cmp_pReg_1, 
      gen_14_cmp_pReg_0, gen_14_cmp_BSCmp_op2_0, gen_14_cmp_BSCmp_carryIn, 
      gen_13_cmp_pBs_30, gen_13_cmp_pBs_29, gen_13_cmp_pBs_28, 
      gen_13_cmp_pBs_27, gen_13_cmp_pBs_26, gen_13_cmp_pBs_25, 
      gen_13_cmp_pBs_24, gen_13_cmp_pBs_23, gen_13_cmp_pMux_30, 
      gen_13_cmp_pMux_29, gen_13_cmp_pMux_28, gen_13_cmp_pMux_27, 
      gen_13_cmp_pMux_26, gen_13_cmp_pMux_25, gen_13_cmp_pMux_24, 
      gen_13_cmp_pMux_23, gen_13_cmp_pMux_22, gen_13_cmp_pMux_21, 
      gen_13_cmp_pMux_20, gen_13_cmp_pMux_19, gen_13_cmp_pMux_18, 
      gen_13_cmp_pMux_17, gen_13_cmp_pMux_16, gen_13_cmp_pMux_15, 
      gen_13_cmp_pMux_14, gen_13_cmp_pMux_13, gen_13_cmp_pMux_12, 
      gen_13_cmp_pMux_11, gen_13_cmp_pMux_10, gen_13_cmp_pMux_9, 
      gen_13_cmp_pMux_8, gen_13_cmp_pMux_7, gen_13_cmp_pMux_6, 
      gen_13_cmp_pMux_5, gen_13_cmp_pMux_4, gen_13_cmp_pMux_3, 
      gen_13_cmp_pMux_2, gen_13_cmp_pMux_1, gen_13_cmp_pMux_0, 
      gen_13_cmp_pReg_30, gen_13_cmp_pReg_29, gen_13_cmp_pReg_28, 
      gen_13_cmp_pReg_27, gen_13_cmp_pReg_26, gen_13_cmp_pReg_25, 
      gen_13_cmp_pReg_24, gen_13_cmp_pReg_23, gen_13_cmp_pReg_22, 
      gen_13_cmp_pReg_21, gen_13_cmp_pReg_20, gen_13_cmp_pReg_19, 
      gen_13_cmp_pReg_18, gen_13_cmp_pReg_17, gen_13_cmp_pReg_16, 
      gen_13_cmp_pReg_15, gen_13_cmp_pReg_14, gen_13_cmp_pReg_13, 
      gen_13_cmp_pReg_12, gen_13_cmp_pReg_11, gen_13_cmp_pReg_10, 
      gen_13_cmp_pReg_9, gen_13_cmp_pReg_8, gen_13_cmp_pReg_7, 
      gen_13_cmp_pReg_6, gen_13_cmp_pReg_5, gen_13_cmp_pReg_4, 
      gen_13_cmp_pReg_3, gen_13_cmp_pReg_2, gen_13_cmp_pReg_1, 
      gen_13_cmp_pReg_0, gen_13_cmp_BSCmp_op2_0, gen_13_cmp_BSCmp_carryIn, 
      gen_12_cmp_pBs_30, gen_12_cmp_pBs_29, gen_12_cmp_pBs_28, 
      gen_12_cmp_pBs_27, gen_12_cmp_pBs_26, gen_12_cmp_pBs_25, 
      gen_12_cmp_pBs_24, gen_12_cmp_pBs_23, gen_12_cmp_pMux_30, 
      gen_12_cmp_pMux_29, gen_12_cmp_pMux_28, gen_12_cmp_pMux_27, 
      gen_12_cmp_pMux_26, gen_12_cmp_pMux_25, gen_12_cmp_pMux_24, 
      gen_12_cmp_pMux_23, gen_12_cmp_pMux_22, gen_12_cmp_pMux_21, 
      gen_12_cmp_pMux_20, gen_12_cmp_pMux_19, gen_12_cmp_pMux_18, 
      gen_12_cmp_pMux_17, gen_12_cmp_pMux_16, gen_12_cmp_pMux_15, 
      gen_12_cmp_pMux_14, gen_12_cmp_pMux_13, gen_12_cmp_pMux_12, 
      gen_12_cmp_pMux_11, gen_12_cmp_pMux_10, gen_12_cmp_pMux_9, 
      gen_12_cmp_pMux_8, gen_12_cmp_pMux_7, gen_12_cmp_pMux_6, 
      gen_12_cmp_pMux_5, gen_12_cmp_pMux_4, gen_12_cmp_pMux_3, 
      gen_12_cmp_pMux_2, gen_12_cmp_pMux_1, gen_12_cmp_pMux_0, 
      gen_12_cmp_pReg_30, gen_12_cmp_pReg_29, gen_12_cmp_pReg_28, 
      gen_12_cmp_pReg_27, gen_12_cmp_pReg_26, gen_12_cmp_pReg_25, 
      gen_12_cmp_pReg_24, gen_12_cmp_pReg_23, gen_12_cmp_pReg_22, 
      gen_12_cmp_pReg_21, gen_12_cmp_pReg_20, gen_12_cmp_pReg_19, 
      gen_12_cmp_pReg_18, gen_12_cmp_pReg_17, gen_12_cmp_pReg_16, 
      gen_12_cmp_pReg_15, gen_12_cmp_pReg_14, gen_12_cmp_pReg_13, 
      gen_12_cmp_pReg_12, gen_12_cmp_pReg_11, gen_12_cmp_pReg_10, 
      gen_12_cmp_pReg_9, gen_12_cmp_pReg_8, gen_12_cmp_pReg_7, 
      gen_12_cmp_pReg_6, gen_12_cmp_pReg_5, gen_12_cmp_pReg_4, 
      gen_12_cmp_pReg_3, gen_12_cmp_pReg_2, gen_12_cmp_pReg_1, 
      gen_12_cmp_pReg_0, gen_12_cmp_BSCmp_op2_0, gen_12_cmp_BSCmp_carryIn, 
      gen_11_cmp_pBs_30, gen_11_cmp_pBs_29, gen_11_cmp_pBs_28, 
      gen_11_cmp_pBs_27, gen_11_cmp_pBs_26, gen_11_cmp_pBs_25, 
      gen_11_cmp_pBs_24, gen_11_cmp_pBs_23, gen_11_cmp_pMux_30, 
      gen_11_cmp_pMux_29, gen_11_cmp_pMux_28, gen_11_cmp_pMux_27, 
      gen_11_cmp_pMux_26, gen_11_cmp_pMux_25, gen_11_cmp_pMux_24, 
      gen_11_cmp_pMux_23, gen_11_cmp_pMux_22, gen_11_cmp_pMux_21, 
      gen_11_cmp_pMux_20, gen_11_cmp_pMux_19, gen_11_cmp_pMux_18, 
      gen_11_cmp_pMux_17, gen_11_cmp_pMux_16, gen_11_cmp_pMux_15, 
      gen_11_cmp_pMux_14, gen_11_cmp_pMux_13, gen_11_cmp_pMux_12, 
      gen_11_cmp_pMux_11, gen_11_cmp_pMux_10, gen_11_cmp_pMux_9, 
      gen_11_cmp_pMux_8, gen_11_cmp_pMux_7, gen_11_cmp_pMux_6, 
      gen_11_cmp_pMux_5, gen_11_cmp_pMux_4, gen_11_cmp_pMux_3, 
      gen_11_cmp_pMux_2, gen_11_cmp_pMux_1, gen_11_cmp_pMux_0, 
      gen_11_cmp_pReg_30, gen_11_cmp_pReg_29, gen_11_cmp_pReg_28, 
      gen_11_cmp_pReg_27, gen_11_cmp_pReg_26, gen_11_cmp_pReg_25, 
      gen_11_cmp_pReg_24, gen_11_cmp_pReg_23, gen_11_cmp_pReg_22, 
      gen_11_cmp_pReg_21, gen_11_cmp_pReg_20, gen_11_cmp_pReg_19, 
      gen_11_cmp_pReg_18, gen_11_cmp_pReg_17, gen_11_cmp_pReg_16, 
      gen_11_cmp_pReg_15, gen_11_cmp_pReg_14, gen_11_cmp_pReg_13, 
      gen_11_cmp_pReg_12, gen_11_cmp_pReg_11, gen_11_cmp_pReg_10, 
      gen_11_cmp_pReg_9, gen_11_cmp_pReg_8, gen_11_cmp_pReg_7, 
      gen_11_cmp_pReg_6, gen_11_cmp_pReg_5, gen_11_cmp_pReg_4, 
      gen_11_cmp_pReg_3, gen_11_cmp_pReg_2, gen_11_cmp_pReg_1, 
      gen_11_cmp_pReg_0, gen_11_cmp_BSCmp_op2_0, gen_11_cmp_BSCmp_carryIn, 
      gen_10_cmp_pBs_30, gen_10_cmp_pBs_29, gen_10_cmp_pBs_28, 
      gen_10_cmp_pBs_27, gen_10_cmp_pBs_26, gen_10_cmp_pBs_25, 
      gen_10_cmp_pBs_24, gen_10_cmp_pBs_23, gen_10_cmp_pMux_30, 
      gen_10_cmp_pMux_29, gen_10_cmp_pMux_28, gen_10_cmp_pMux_27, 
      gen_10_cmp_pMux_26, gen_10_cmp_pMux_25, gen_10_cmp_pMux_24, 
      gen_10_cmp_pMux_23, gen_10_cmp_pMux_22, gen_10_cmp_pMux_21, 
      gen_10_cmp_pMux_20, gen_10_cmp_pMux_19, gen_10_cmp_pMux_18, 
      gen_10_cmp_pMux_17, gen_10_cmp_pMux_16, gen_10_cmp_pMux_15, 
      gen_10_cmp_pMux_14, gen_10_cmp_pMux_13, gen_10_cmp_pMux_12, 
      gen_10_cmp_pMux_11, gen_10_cmp_pMux_10, gen_10_cmp_pMux_9, 
      gen_10_cmp_pMux_8, gen_10_cmp_pMux_7, gen_10_cmp_pMux_6, 
      gen_10_cmp_pMux_5, gen_10_cmp_pMux_4, gen_10_cmp_pMux_3, 
      gen_10_cmp_pMux_2, gen_10_cmp_pMux_1, gen_10_cmp_pMux_0, 
      gen_10_cmp_pReg_30, gen_10_cmp_pReg_29, gen_10_cmp_pReg_28, 
      gen_10_cmp_pReg_27, gen_10_cmp_pReg_26, gen_10_cmp_pReg_25, 
      gen_10_cmp_pReg_24, gen_10_cmp_pReg_23, gen_10_cmp_pReg_22, 
      gen_10_cmp_pReg_21, gen_10_cmp_pReg_20, gen_10_cmp_pReg_19, 
      gen_10_cmp_pReg_18, gen_10_cmp_pReg_17, gen_10_cmp_pReg_16, 
      gen_10_cmp_pReg_15, gen_10_cmp_pReg_14, gen_10_cmp_pReg_13, 
      gen_10_cmp_pReg_12, gen_10_cmp_pReg_11, gen_10_cmp_pReg_10, 
      gen_10_cmp_pReg_9, gen_10_cmp_pReg_8, gen_10_cmp_pReg_7, 
      gen_10_cmp_pReg_6, gen_10_cmp_pReg_5, gen_10_cmp_pReg_4, 
      gen_10_cmp_pReg_3, gen_10_cmp_pReg_2, gen_10_cmp_pReg_1, 
      gen_10_cmp_pReg_0, gen_10_cmp_BSCmp_op2_0, gen_10_cmp_BSCmp_carryIn, 
      gen_9_cmp_pBs_30, gen_9_cmp_pBs_29, gen_9_cmp_pBs_28, gen_9_cmp_pBs_27, 
      gen_9_cmp_pBs_26, gen_9_cmp_pBs_25, gen_9_cmp_pBs_24, gen_9_cmp_pBs_23, 
      gen_9_cmp_pMux_30, gen_9_cmp_pMux_29, gen_9_cmp_pMux_28, 
      gen_9_cmp_pMux_27, gen_9_cmp_pMux_26, gen_9_cmp_pMux_25, 
      gen_9_cmp_pMux_24, gen_9_cmp_pMux_23, gen_9_cmp_pMux_22, 
      gen_9_cmp_pMux_21, gen_9_cmp_pMux_20, gen_9_cmp_pMux_19, 
      gen_9_cmp_pMux_18, gen_9_cmp_pMux_17, gen_9_cmp_pMux_16, 
      gen_9_cmp_pMux_15, gen_9_cmp_pMux_14, gen_9_cmp_pMux_13, 
      gen_9_cmp_pMux_12, gen_9_cmp_pMux_11, gen_9_cmp_pMux_10, 
      gen_9_cmp_pMux_9, gen_9_cmp_pMux_8, gen_9_cmp_pMux_7, gen_9_cmp_pMux_6, 
      gen_9_cmp_pMux_5, gen_9_cmp_pMux_4, gen_9_cmp_pMux_3, gen_9_cmp_pMux_2, 
      gen_9_cmp_pMux_1, gen_9_cmp_pMux_0, gen_9_cmp_pReg_30, 
      gen_9_cmp_pReg_29, gen_9_cmp_pReg_28, gen_9_cmp_pReg_27, 
      gen_9_cmp_pReg_26, gen_9_cmp_pReg_25, gen_9_cmp_pReg_24, 
      gen_9_cmp_pReg_23, gen_9_cmp_pReg_22, gen_9_cmp_pReg_21, 
      gen_9_cmp_pReg_20, gen_9_cmp_pReg_19, gen_9_cmp_pReg_18, 
      gen_9_cmp_pReg_17, gen_9_cmp_pReg_16, gen_9_cmp_pReg_15, 
      gen_9_cmp_pReg_14, gen_9_cmp_pReg_13, gen_9_cmp_pReg_12, 
      gen_9_cmp_pReg_11, gen_9_cmp_pReg_10, gen_9_cmp_pReg_9, 
      gen_9_cmp_pReg_8, gen_9_cmp_pReg_7, gen_9_cmp_pReg_6, gen_9_cmp_pReg_5, 
      gen_9_cmp_pReg_4, gen_9_cmp_pReg_3, gen_9_cmp_pReg_2, gen_9_cmp_pReg_1, 
      gen_9_cmp_pReg_0, gen_9_cmp_BSCmp_op2_0, gen_9_cmp_BSCmp_carryIn, 
      gen_8_cmp_pBs_30, gen_8_cmp_pBs_29, gen_8_cmp_pBs_28, gen_8_cmp_pBs_27, 
      gen_8_cmp_pBs_26, gen_8_cmp_pBs_25, gen_8_cmp_pBs_24, gen_8_cmp_pBs_23, 
      gen_8_cmp_pMux_30, gen_8_cmp_pMux_29, gen_8_cmp_pMux_28, 
      gen_8_cmp_pMux_27, gen_8_cmp_pMux_26, gen_8_cmp_pMux_25, 
      gen_8_cmp_pMux_24, gen_8_cmp_pMux_23, gen_8_cmp_pMux_22, 
      gen_8_cmp_pMux_21, gen_8_cmp_pMux_20, gen_8_cmp_pMux_19, 
      gen_8_cmp_pMux_18, gen_8_cmp_pMux_17, gen_8_cmp_pMux_16, 
      gen_8_cmp_pMux_15, gen_8_cmp_pMux_14, gen_8_cmp_pMux_13, 
      gen_8_cmp_pMux_12, gen_8_cmp_pMux_11, gen_8_cmp_pMux_10, 
      gen_8_cmp_pMux_9, gen_8_cmp_pMux_8, gen_8_cmp_pMux_7, gen_8_cmp_pMux_6, 
      gen_8_cmp_pMux_5, gen_8_cmp_pMux_4, gen_8_cmp_pMux_3, gen_8_cmp_pMux_2, 
      gen_8_cmp_pMux_1, gen_8_cmp_pMux_0, gen_8_cmp_pReg_30, 
      gen_8_cmp_pReg_29, gen_8_cmp_pReg_28, gen_8_cmp_pReg_27, 
      gen_8_cmp_pReg_26, gen_8_cmp_pReg_25, gen_8_cmp_pReg_24, 
      gen_8_cmp_pReg_23, gen_8_cmp_pReg_22, gen_8_cmp_pReg_21, 
      gen_8_cmp_pReg_20, gen_8_cmp_pReg_19, gen_8_cmp_pReg_18, 
      gen_8_cmp_pReg_17, gen_8_cmp_pReg_16, gen_8_cmp_pReg_15, 
      gen_8_cmp_pReg_14, gen_8_cmp_pReg_13, gen_8_cmp_pReg_12, 
      gen_8_cmp_pReg_11, gen_8_cmp_pReg_10, gen_8_cmp_pReg_9, 
      gen_8_cmp_pReg_8, gen_8_cmp_pReg_7, gen_8_cmp_pReg_6, gen_8_cmp_pReg_5, 
      gen_8_cmp_pReg_4, gen_8_cmp_pReg_3, gen_8_cmp_pReg_2, gen_8_cmp_pReg_1, 
      gen_8_cmp_pReg_0, gen_8_cmp_BSCmp_op2_0, gen_8_cmp_BSCmp_carryIn, 
      gen_7_cmp_pBs_30, gen_7_cmp_pBs_29, gen_7_cmp_pBs_28, gen_7_cmp_pBs_27, 
      gen_7_cmp_pBs_26, gen_7_cmp_pBs_25, gen_7_cmp_pBs_24, gen_7_cmp_pBs_23, 
      gen_7_cmp_pMux_30, gen_7_cmp_pMux_29, gen_7_cmp_pMux_28, 
      gen_7_cmp_pMux_27, gen_7_cmp_pMux_26, gen_7_cmp_pMux_25, 
      gen_7_cmp_pMux_24, gen_7_cmp_pMux_23, gen_7_cmp_pMux_22, 
      gen_7_cmp_pMux_21, gen_7_cmp_pMux_20, gen_7_cmp_pMux_19, 
      gen_7_cmp_pMux_18, gen_7_cmp_pMux_17, gen_7_cmp_pMux_16, 
      gen_7_cmp_pMux_15, gen_7_cmp_pMux_14, gen_7_cmp_pMux_13, 
      gen_7_cmp_pMux_12, gen_7_cmp_pMux_11, gen_7_cmp_pMux_10, 
      gen_7_cmp_pMux_9, gen_7_cmp_pMux_8, gen_7_cmp_pMux_7, gen_7_cmp_pMux_6, 
      gen_7_cmp_pMux_5, gen_7_cmp_pMux_4, gen_7_cmp_pMux_3, gen_7_cmp_pMux_2, 
      gen_7_cmp_pMux_1, gen_7_cmp_pMux_0, gen_7_cmp_pReg_30, 
      gen_7_cmp_pReg_29, gen_7_cmp_pReg_28, gen_7_cmp_pReg_27, 
      gen_7_cmp_pReg_26, gen_7_cmp_pReg_25, gen_7_cmp_pReg_24, 
      gen_7_cmp_pReg_23, gen_7_cmp_pReg_22, gen_7_cmp_pReg_21, 
      gen_7_cmp_pReg_20, gen_7_cmp_pReg_19, gen_7_cmp_pReg_18, 
      gen_7_cmp_pReg_17, gen_7_cmp_pReg_16, gen_7_cmp_pReg_15, 
      gen_7_cmp_pReg_14, gen_7_cmp_pReg_13, gen_7_cmp_pReg_12, 
      gen_7_cmp_pReg_11, gen_7_cmp_pReg_10, gen_7_cmp_pReg_9, 
      gen_7_cmp_pReg_8, gen_7_cmp_pReg_7, gen_7_cmp_pReg_6, gen_7_cmp_pReg_5, 
      gen_7_cmp_pReg_4, gen_7_cmp_pReg_3, gen_7_cmp_pReg_2, gen_7_cmp_pReg_1, 
      gen_7_cmp_pReg_0, gen_7_cmp_BSCmp_op2_0, gen_7_cmp_BSCmp_carryIn, 
      gen_6_cmp_pBs_30, gen_6_cmp_pBs_29, gen_6_cmp_pBs_28, gen_6_cmp_pBs_27, 
      gen_6_cmp_pBs_26, gen_6_cmp_pBs_25, gen_6_cmp_pBs_24, gen_6_cmp_pBs_23, 
      gen_6_cmp_pMux_30, gen_6_cmp_pMux_29, gen_6_cmp_pMux_28, 
      gen_6_cmp_pMux_27, gen_6_cmp_pMux_26, gen_6_cmp_pMux_25, 
      gen_6_cmp_pMux_24, gen_6_cmp_pMux_23, gen_6_cmp_pMux_22, 
      gen_6_cmp_pMux_21, gen_6_cmp_pMux_20, gen_6_cmp_pMux_19, 
      gen_6_cmp_pMux_18, gen_6_cmp_pMux_17, gen_6_cmp_pMux_16, 
      gen_6_cmp_pMux_15, gen_6_cmp_pMux_14, gen_6_cmp_pMux_13, 
      gen_6_cmp_pMux_12, gen_6_cmp_pMux_11, gen_6_cmp_pMux_10, 
      gen_6_cmp_pMux_9, gen_6_cmp_pMux_8, gen_6_cmp_pMux_7, gen_6_cmp_pMux_6, 
      gen_6_cmp_pMux_5, gen_6_cmp_pMux_4, gen_6_cmp_pMux_3, gen_6_cmp_pMux_2, 
      gen_6_cmp_pMux_1, gen_6_cmp_pMux_0, gen_6_cmp_pReg_30, 
      gen_6_cmp_pReg_29, gen_6_cmp_pReg_28, gen_6_cmp_pReg_27, 
      gen_6_cmp_pReg_26, gen_6_cmp_pReg_25, gen_6_cmp_pReg_24, 
      gen_6_cmp_pReg_23, gen_6_cmp_pReg_22, gen_6_cmp_pReg_21, 
      gen_6_cmp_pReg_20, gen_6_cmp_pReg_19, gen_6_cmp_pReg_18, 
      gen_6_cmp_pReg_17, gen_6_cmp_pReg_16, gen_6_cmp_pReg_15, 
      gen_6_cmp_pReg_14, gen_6_cmp_pReg_13, gen_6_cmp_pReg_12, 
      gen_6_cmp_pReg_11, gen_6_cmp_pReg_10, gen_6_cmp_pReg_9, 
      gen_6_cmp_pReg_8, gen_6_cmp_pReg_7, gen_6_cmp_pReg_6, gen_6_cmp_pReg_5, 
      gen_6_cmp_pReg_4, gen_6_cmp_pReg_3, gen_6_cmp_pReg_2, gen_6_cmp_pReg_1, 
      gen_6_cmp_pReg_0, gen_6_cmp_BSCmp_op2_0, gen_6_cmp_BSCmp_carryIn, 
      gen_5_cmp_pBs_30, gen_5_cmp_pBs_29, gen_5_cmp_pBs_28, gen_5_cmp_pBs_27, 
      gen_5_cmp_pBs_26, gen_5_cmp_pBs_25, gen_5_cmp_pBs_24, gen_5_cmp_pBs_23, 
      gen_5_cmp_pMux_30, gen_5_cmp_pMux_29, gen_5_cmp_pMux_28, 
      gen_5_cmp_pMux_27, gen_5_cmp_pMux_26, gen_5_cmp_pMux_25, 
      gen_5_cmp_pMux_24, gen_5_cmp_pMux_23, gen_5_cmp_pMux_22, 
      gen_5_cmp_pMux_21, gen_5_cmp_pMux_20, gen_5_cmp_pMux_19, 
      gen_5_cmp_pMux_18, gen_5_cmp_pMux_17, gen_5_cmp_pMux_16, 
      gen_5_cmp_pMux_15, gen_5_cmp_pMux_14, gen_5_cmp_pMux_13, 
      gen_5_cmp_pMux_12, gen_5_cmp_pMux_11, gen_5_cmp_pMux_10, 
      gen_5_cmp_pMux_9, gen_5_cmp_pMux_8, gen_5_cmp_pMux_7, gen_5_cmp_pMux_6, 
      gen_5_cmp_pMux_5, gen_5_cmp_pMux_4, gen_5_cmp_pMux_3, gen_5_cmp_pMux_2, 
      gen_5_cmp_pMux_1, gen_5_cmp_pMux_0, gen_5_cmp_pReg_30, 
      gen_5_cmp_pReg_29, gen_5_cmp_pReg_28, gen_5_cmp_pReg_27, 
      gen_5_cmp_pReg_26, gen_5_cmp_pReg_25, gen_5_cmp_pReg_24, 
      gen_5_cmp_pReg_23, gen_5_cmp_pReg_22, gen_5_cmp_pReg_21, 
      gen_5_cmp_pReg_20, gen_5_cmp_pReg_19, gen_5_cmp_pReg_18, 
      gen_5_cmp_pReg_17, gen_5_cmp_pReg_16, gen_5_cmp_pReg_15, 
      gen_5_cmp_pReg_14, gen_5_cmp_pReg_13, gen_5_cmp_pReg_12, 
      gen_5_cmp_pReg_11, gen_5_cmp_pReg_10, gen_5_cmp_pReg_9, 
      gen_5_cmp_pReg_8, gen_5_cmp_pReg_7, gen_5_cmp_pReg_6, gen_5_cmp_pReg_5, 
      gen_5_cmp_pReg_4, gen_5_cmp_pReg_3, gen_5_cmp_pReg_2, gen_5_cmp_pReg_1, 
      gen_5_cmp_pReg_0, gen_5_cmp_BSCmp_op2_0, gen_5_cmp_BSCmp_carryIn, 
      gen_4_cmp_pBs_30, gen_4_cmp_pBs_29, gen_4_cmp_pBs_28, gen_4_cmp_pBs_27, 
      gen_4_cmp_pBs_26, gen_4_cmp_pBs_25, gen_4_cmp_pBs_24, gen_4_cmp_pBs_23, 
      gen_4_cmp_pMux_30, gen_4_cmp_pMux_29, gen_4_cmp_pMux_28, 
      gen_4_cmp_pMux_27, gen_4_cmp_pMux_26, gen_4_cmp_pMux_25, 
      gen_4_cmp_pMux_24, gen_4_cmp_pMux_23, gen_4_cmp_pMux_22, 
      gen_4_cmp_pMux_21, gen_4_cmp_pMux_20, gen_4_cmp_pMux_19, 
      gen_4_cmp_pMux_18, gen_4_cmp_pMux_17, gen_4_cmp_pMux_16, 
      gen_4_cmp_pMux_15, gen_4_cmp_pMux_14, gen_4_cmp_pMux_13, 
      gen_4_cmp_pMux_12, gen_4_cmp_pMux_11, gen_4_cmp_pMux_10, 
      gen_4_cmp_pMux_9, gen_4_cmp_pMux_8, gen_4_cmp_pMux_7, gen_4_cmp_pMux_6, 
      gen_4_cmp_pMux_5, gen_4_cmp_pMux_4, gen_4_cmp_pMux_3, gen_4_cmp_pMux_2, 
      gen_4_cmp_pMux_1, gen_4_cmp_pMux_0, gen_4_cmp_pReg_30, 
      gen_4_cmp_pReg_29, gen_4_cmp_pReg_28, gen_4_cmp_pReg_27, 
      gen_4_cmp_pReg_26, gen_4_cmp_pReg_25, gen_4_cmp_pReg_24, 
      gen_4_cmp_pReg_23, gen_4_cmp_pReg_22, gen_4_cmp_pReg_21, 
      gen_4_cmp_pReg_20, gen_4_cmp_pReg_19, gen_4_cmp_pReg_18, 
      gen_4_cmp_pReg_17, gen_4_cmp_pReg_16, gen_4_cmp_pReg_15, 
      gen_4_cmp_pReg_14, gen_4_cmp_pReg_13, gen_4_cmp_pReg_12, 
      gen_4_cmp_pReg_11, gen_4_cmp_pReg_10, gen_4_cmp_pReg_9, 
      gen_4_cmp_pReg_8, gen_4_cmp_pReg_7, gen_4_cmp_pReg_6, gen_4_cmp_pReg_5, 
      gen_4_cmp_pReg_4, gen_4_cmp_pReg_3, gen_4_cmp_pReg_2, gen_4_cmp_pReg_1, 
      gen_4_cmp_pReg_0, gen_4_cmp_BSCmp_op2_0, gen_4_cmp_BSCmp_carryIn, 
      gen_3_cmp_pBs_30, gen_3_cmp_pBs_29, gen_3_cmp_pBs_28, gen_3_cmp_pBs_27, 
      gen_3_cmp_pBs_26, gen_3_cmp_pBs_25, gen_3_cmp_pBs_24, gen_3_cmp_pBs_23, 
      gen_3_cmp_pMux_30, gen_3_cmp_pMux_29, gen_3_cmp_pMux_28, 
      gen_3_cmp_pMux_27, gen_3_cmp_pMux_26, gen_3_cmp_pMux_25, 
      gen_3_cmp_pMux_24, gen_3_cmp_pMux_23, gen_3_cmp_pMux_22, 
      gen_3_cmp_pMux_21, gen_3_cmp_pMux_20, gen_3_cmp_pMux_19, 
      gen_3_cmp_pMux_18, gen_3_cmp_pMux_17, gen_3_cmp_pMux_16, 
      gen_3_cmp_pMux_15, gen_3_cmp_pMux_14, gen_3_cmp_pMux_13, 
      gen_3_cmp_pMux_12, gen_3_cmp_pMux_11, gen_3_cmp_pMux_10, 
      gen_3_cmp_pMux_9, gen_3_cmp_pMux_8, gen_3_cmp_pMux_7, gen_3_cmp_pMux_6, 
      gen_3_cmp_pMux_5, gen_3_cmp_pMux_4, gen_3_cmp_pMux_3, gen_3_cmp_pMux_2, 
      gen_3_cmp_pMux_1, gen_3_cmp_pMux_0, gen_3_cmp_pReg_30, 
      gen_3_cmp_pReg_29, gen_3_cmp_pReg_28, gen_3_cmp_pReg_27, 
      gen_3_cmp_pReg_26, gen_3_cmp_pReg_25, gen_3_cmp_pReg_24, 
      gen_3_cmp_pReg_23, gen_3_cmp_pReg_22, gen_3_cmp_pReg_21, 
      gen_3_cmp_pReg_20, gen_3_cmp_pReg_19, gen_3_cmp_pReg_18, 
      gen_3_cmp_pReg_17, gen_3_cmp_pReg_16, gen_3_cmp_pReg_15, 
      gen_3_cmp_pReg_14, gen_3_cmp_pReg_13, gen_3_cmp_pReg_12, 
      gen_3_cmp_pReg_11, gen_3_cmp_pReg_10, gen_3_cmp_pReg_9, 
      gen_3_cmp_pReg_8, gen_3_cmp_pReg_7, gen_3_cmp_pReg_6, gen_3_cmp_pReg_5, 
      gen_3_cmp_pReg_4, gen_3_cmp_pReg_3, gen_3_cmp_pReg_2, gen_3_cmp_pReg_1, 
      gen_3_cmp_pReg_0, gen_3_cmp_BSCmp_op2_0, gen_3_cmp_BSCmp_carryIn, 
      gen_2_cmp_pBs_30, gen_2_cmp_pBs_29, gen_2_cmp_pBs_28, gen_2_cmp_pBs_27, 
      gen_2_cmp_pBs_26, gen_2_cmp_pBs_25, gen_2_cmp_pBs_24, gen_2_cmp_pBs_23, 
      gen_2_cmp_pMux_30, gen_2_cmp_pMux_29, gen_2_cmp_pMux_28, 
      gen_2_cmp_pMux_27, gen_2_cmp_pMux_26, gen_2_cmp_pMux_25, 
      gen_2_cmp_pMux_24, gen_2_cmp_pMux_23, gen_2_cmp_pMux_22, 
      gen_2_cmp_pMux_21, gen_2_cmp_pMux_20, gen_2_cmp_pMux_19, 
      gen_2_cmp_pMux_18, gen_2_cmp_pMux_17, gen_2_cmp_pMux_16, 
      gen_2_cmp_pMux_15, gen_2_cmp_pMux_14, gen_2_cmp_pMux_13, 
      gen_2_cmp_pMux_12, gen_2_cmp_pMux_11, gen_2_cmp_pMux_10, 
      gen_2_cmp_pMux_9, gen_2_cmp_pMux_8, gen_2_cmp_pMux_7, gen_2_cmp_pMux_6, 
      gen_2_cmp_pMux_5, gen_2_cmp_pMux_4, gen_2_cmp_pMux_3, gen_2_cmp_pMux_2, 
      gen_2_cmp_pMux_1, gen_2_cmp_pMux_0, gen_2_cmp_pReg_30, 
      gen_2_cmp_pReg_29, gen_2_cmp_pReg_28, gen_2_cmp_pReg_27, 
      gen_2_cmp_pReg_26, gen_2_cmp_pReg_25, gen_2_cmp_pReg_24, 
      gen_2_cmp_pReg_23, gen_2_cmp_pReg_22, gen_2_cmp_pReg_21, 
      gen_2_cmp_pReg_20, gen_2_cmp_pReg_19, gen_2_cmp_pReg_18, 
      gen_2_cmp_pReg_17, gen_2_cmp_pReg_16, gen_2_cmp_pReg_15, 
      gen_2_cmp_pReg_14, gen_2_cmp_pReg_13, gen_2_cmp_pReg_12, 
      gen_2_cmp_pReg_11, gen_2_cmp_pReg_10, gen_2_cmp_pReg_9, 
      gen_2_cmp_pReg_8, gen_2_cmp_pReg_7, gen_2_cmp_pReg_6, gen_2_cmp_pReg_5, 
      gen_2_cmp_pReg_4, gen_2_cmp_pReg_3, gen_2_cmp_pReg_2, gen_2_cmp_pReg_1, 
      gen_2_cmp_pReg_0, gen_2_cmp_BSCmp_op2_0, gen_2_cmp_BSCmp_carryIn, 
      gen_1_cmp_pBs_30, gen_1_cmp_pBs_29, gen_1_cmp_pBs_28, gen_1_cmp_pBs_27, 
      gen_1_cmp_pBs_26, gen_1_cmp_pBs_25, gen_1_cmp_pBs_24, gen_1_cmp_pBs_23, 
      gen_1_cmp_pMux_30, gen_1_cmp_pMux_29, gen_1_cmp_pMux_28, 
      gen_1_cmp_pMux_27, gen_1_cmp_pMux_26, gen_1_cmp_pMux_25, 
      gen_1_cmp_pMux_24, gen_1_cmp_pMux_23, gen_1_cmp_pMux_22, 
      gen_1_cmp_pMux_21, gen_1_cmp_pMux_20, gen_1_cmp_pMux_19, 
      gen_1_cmp_pMux_18, gen_1_cmp_pMux_17, gen_1_cmp_pMux_16, 
      gen_1_cmp_pMux_15, gen_1_cmp_pMux_14, gen_1_cmp_pMux_13, 
      gen_1_cmp_pMux_12, gen_1_cmp_pMux_11, gen_1_cmp_pMux_10, 
      gen_1_cmp_pMux_9, gen_1_cmp_pMux_8, gen_1_cmp_pMux_7, gen_1_cmp_pMux_6, 
      gen_1_cmp_pMux_5, gen_1_cmp_pMux_4, gen_1_cmp_pMux_3, gen_1_cmp_pMux_2, 
      gen_1_cmp_pMux_1, gen_1_cmp_pMux_0, gen_1_cmp_pReg_30, 
      gen_1_cmp_pReg_29, gen_1_cmp_pReg_28, gen_1_cmp_pReg_27, 
      gen_1_cmp_pReg_26, gen_1_cmp_pReg_25, gen_1_cmp_pReg_24, 
      gen_1_cmp_pReg_23, gen_1_cmp_pReg_22, gen_1_cmp_pReg_21, 
      gen_1_cmp_pReg_20, gen_1_cmp_pReg_19, gen_1_cmp_pReg_18, 
      gen_1_cmp_pReg_17, gen_1_cmp_pReg_16, gen_1_cmp_pReg_15, 
      gen_1_cmp_pReg_14, gen_1_cmp_pReg_13, gen_1_cmp_pReg_12, 
      gen_1_cmp_pReg_11, gen_1_cmp_pReg_10, gen_1_cmp_pReg_9, 
      gen_1_cmp_pReg_8, gen_1_cmp_pReg_7, gen_1_cmp_pReg_6, gen_1_cmp_pReg_5, 
      gen_1_cmp_pReg_4, gen_1_cmp_pReg_3, gen_1_cmp_pReg_2, gen_1_cmp_pReg_1, 
      gen_1_cmp_pReg_0, gen_1_cmp_BSCmp_op2_0, gen_1_cmp_BSCmp_carryIn, 
      gen_0_cmp_pBs_30, gen_0_cmp_pBs_29, gen_0_cmp_pBs_28, gen_0_cmp_pBs_27, 
      gen_0_cmp_pBs_26, gen_0_cmp_pBs_25, gen_0_cmp_pBs_24, gen_0_cmp_pBs_23, 
      gen_0_cmp_pMux_30, gen_0_cmp_pMux_29, gen_0_cmp_pMux_28, 
      gen_0_cmp_pMux_27, gen_0_cmp_pMux_26, gen_0_cmp_pMux_25, 
      gen_0_cmp_pMux_24, gen_0_cmp_pMux_23, gen_0_cmp_pMux_22, 
      gen_0_cmp_pMux_21, gen_0_cmp_pMux_20, gen_0_cmp_pMux_19, 
      gen_0_cmp_pMux_18, gen_0_cmp_pMux_17, gen_0_cmp_pMux_16, 
      gen_0_cmp_pMux_15, gen_0_cmp_pMux_14, gen_0_cmp_pMux_13, 
      gen_0_cmp_pMux_12, gen_0_cmp_pMux_11, gen_0_cmp_pMux_10, 
      gen_0_cmp_pMux_9, gen_0_cmp_pMux_8, gen_0_cmp_pMux_7, gen_0_cmp_pMux_6, 
      gen_0_cmp_pMux_5, gen_0_cmp_pMux_4, gen_0_cmp_pMux_3, gen_0_cmp_pMux_2, 
      gen_0_cmp_pMux_1, gen_0_cmp_pMux_0, gen_0_cmp_pReg_30, 
      gen_0_cmp_pReg_29, gen_0_cmp_pReg_28, gen_0_cmp_pReg_27, 
      gen_0_cmp_pReg_26, gen_0_cmp_pReg_25, gen_0_cmp_pReg_24, 
      gen_0_cmp_pReg_23, gen_0_cmp_pReg_22, gen_0_cmp_pReg_21, 
      gen_0_cmp_pReg_20, gen_0_cmp_pReg_19, gen_0_cmp_pReg_18, 
      gen_0_cmp_pReg_17, gen_0_cmp_pReg_16, gen_0_cmp_pReg_15, 
      gen_0_cmp_pReg_14, gen_0_cmp_pReg_13, gen_0_cmp_pReg_12, 
      gen_0_cmp_pReg_11, gen_0_cmp_pReg_10, gen_0_cmp_pReg_9, 
      gen_0_cmp_pReg_8, gen_0_cmp_pReg_7, gen_0_cmp_pReg_6, gen_0_cmp_pReg_5, 
      gen_0_cmp_pReg_4, gen_0_cmp_pReg_3, gen_0_cmp_pReg_2, gen_0_cmp_pReg_1, 
      gen_0_cmp_pReg_0, gen_0_cmp_BSCmp_op2_0, gen_0_cmp_BSCmp_carryIn, 
      gen_24_cmp_BSCmp_op2_16, gen_24_cmp_BSCmp_op2_15, 
      gen_24_cmp_BSCmp_op2_14, gen_24_cmp_BSCmp_op2_13, 
      gen_24_cmp_BSCmp_op2_12, gen_24_cmp_BSCmp_op2_11, 
      gen_24_cmp_BSCmp_op2_10, gen_24_cmp_BSCmp_op2_9, 
      gen_24_cmp_BSCmp_op2_8, gen_24_cmp_BSCmp_op2_7, gen_24_cmp_BSCmp_op2_6, 
      gen_24_cmp_BSCmp_op2_5, gen_24_cmp_BSCmp_op2_4, gen_24_cmp_BSCmp_op2_3, 
      gen_24_cmp_BSCmp_op2_2, gen_24_cmp_BSCmp_op2_1, 
      gen_23_cmp_BSCmp_op2_16, gen_23_cmp_BSCmp_op2_15, 
      gen_23_cmp_BSCmp_op2_14, gen_23_cmp_BSCmp_op2_13, 
      gen_23_cmp_BSCmp_op2_12, gen_23_cmp_BSCmp_op2_11, 
      gen_23_cmp_BSCmp_op2_10, gen_23_cmp_BSCmp_op2_9, 
      gen_23_cmp_BSCmp_op2_8, gen_23_cmp_BSCmp_op2_7, gen_23_cmp_BSCmp_op2_6, 
      gen_23_cmp_BSCmp_op2_5, gen_23_cmp_BSCmp_op2_4, gen_23_cmp_BSCmp_op2_3, 
      gen_23_cmp_BSCmp_op2_2, gen_23_cmp_BSCmp_op2_1, 
      gen_22_cmp_BSCmp_op2_16, gen_22_cmp_BSCmp_op2_15, 
      gen_22_cmp_BSCmp_op2_14, gen_22_cmp_BSCmp_op2_13, 
      gen_22_cmp_BSCmp_op2_12, gen_22_cmp_BSCmp_op2_11, 
      gen_22_cmp_BSCmp_op2_10, gen_22_cmp_BSCmp_op2_9, 
      gen_22_cmp_BSCmp_op2_8, gen_22_cmp_BSCmp_op2_7, gen_22_cmp_BSCmp_op2_6, 
      gen_22_cmp_BSCmp_op2_5, gen_22_cmp_BSCmp_op2_4, gen_22_cmp_BSCmp_op2_3, 
      gen_22_cmp_BSCmp_op2_2, gen_22_cmp_BSCmp_op2_1, 
      gen_21_cmp_BSCmp_op2_16, gen_21_cmp_BSCmp_op2_15, 
      gen_21_cmp_BSCmp_op2_14, gen_21_cmp_BSCmp_op2_13, 
      gen_21_cmp_BSCmp_op2_12, gen_21_cmp_BSCmp_op2_11, 
      gen_21_cmp_BSCmp_op2_10, gen_21_cmp_BSCmp_op2_9, 
      gen_21_cmp_BSCmp_op2_8, gen_21_cmp_BSCmp_op2_7, gen_21_cmp_BSCmp_op2_6, 
      gen_21_cmp_BSCmp_op2_5, gen_21_cmp_BSCmp_op2_4, gen_21_cmp_BSCmp_op2_3, 
      gen_21_cmp_BSCmp_op2_2, gen_21_cmp_BSCmp_op2_1, 
      gen_20_cmp_BSCmp_op2_16, gen_20_cmp_BSCmp_op2_15, 
      gen_20_cmp_BSCmp_op2_14, gen_20_cmp_BSCmp_op2_13, 
      gen_20_cmp_BSCmp_op2_12, gen_20_cmp_BSCmp_op2_11, 
      gen_20_cmp_BSCmp_op2_10, gen_20_cmp_BSCmp_op2_9, 
      gen_20_cmp_BSCmp_op2_8, gen_20_cmp_BSCmp_op2_7, gen_20_cmp_BSCmp_op2_6, 
      gen_20_cmp_BSCmp_op2_5, gen_20_cmp_BSCmp_op2_4, gen_20_cmp_BSCmp_op2_3, 
      gen_20_cmp_BSCmp_op2_2, gen_20_cmp_BSCmp_op2_1, 
      gen_19_cmp_BSCmp_op2_16, gen_19_cmp_BSCmp_op2_15, 
      gen_19_cmp_BSCmp_op2_14, gen_19_cmp_BSCmp_op2_13, 
      gen_19_cmp_BSCmp_op2_12, gen_19_cmp_BSCmp_op2_11, 
      gen_19_cmp_BSCmp_op2_10, gen_19_cmp_BSCmp_op2_9, 
      gen_19_cmp_BSCmp_op2_8, gen_19_cmp_BSCmp_op2_7, gen_19_cmp_BSCmp_op2_6, 
      gen_19_cmp_BSCmp_op2_5, gen_19_cmp_BSCmp_op2_4, gen_19_cmp_BSCmp_op2_3, 
      gen_19_cmp_BSCmp_op2_2, gen_19_cmp_BSCmp_op2_1, 
      gen_18_cmp_BSCmp_op2_16, gen_18_cmp_BSCmp_op2_15, 
      gen_18_cmp_BSCmp_op2_14, gen_18_cmp_BSCmp_op2_13, 
      gen_18_cmp_BSCmp_op2_12, gen_18_cmp_BSCmp_op2_11, 
      gen_18_cmp_BSCmp_op2_10, gen_18_cmp_BSCmp_op2_9, 
      gen_18_cmp_BSCmp_op2_8, gen_18_cmp_BSCmp_op2_7, gen_18_cmp_BSCmp_op2_6, 
      gen_18_cmp_BSCmp_op2_5, gen_18_cmp_BSCmp_op2_4, gen_18_cmp_BSCmp_op2_3, 
      gen_18_cmp_BSCmp_op2_2, gen_18_cmp_BSCmp_op2_1, 
      gen_17_cmp_BSCmp_op2_16, gen_17_cmp_BSCmp_op2_15, 
      gen_17_cmp_BSCmp_op2_14, gen_17_cmp_BSCmp_op2_13, 
      gen_17_cmp_BSCmp_op2_12, gen_17_cmp_BSCmp_op2_11, 
      gen_17_cmp_BSCmp_op2_10, gen_17_cmp_BSCmp_op2_9, 
      gen_17_cmp_BSCmp_op2_8, gen_17_cmp_BSCmp_op2_7, gen_17_cmp_BSCmp_op2_6, 
      gen_17_cmp_BSCmp_op2_5, gen_17_cmp_BSCmp_op2_4, gen_17_cmp_BSCmp_op2_3, 
      gen_17_cmp_BSCmp_op2_2, gen_17_cmp_BSCmp_op2_1, 
      gen_16_cmp_BSCmp_op2_16, gen_16_cmp_BSCmp_op2_15, 
      gen_16_cmp_BSCmp_op2_14, gen_16_cmp_BSCmp_op2_13, 
      gen_16_cmp_BSCmp_op2_12, gen_16_cmp_BSCmp_op2_11, 
      gen_16_cmp_BSCmp_op2_10, gen_16_cmp_BSCmp_op2_9, 
      gen_16_cmp_BSCmp_op2_8, gen_16_cmp_BSCmp_op2_7, gen_16_cmp_BSCmp_op2_6, 
      gen_16_cmp_BSCmp_op2_5, gen_16_cmp_BSCmp_op2_4, gen_16_cmp_BSCmp_op2_3, 
      gen_16_cmp_BSCmp_op2_2, gen_16_cmp_BSCmp_op2_1, 
      gen_15_cmp_BSCmp_op2_16, gen_15_cmp_BSCmp_op2_15, 
      gen_15_cmp_BSCmp_op2_14, gen_15_cmp_BSCmp_op2_13, 
      gen_15_cmp_BSCmp_op2_12, gen_15_cmp_BSCmp_op2_11, 
      gen_15_cmp_BSCmp_op2_10, gen_15_cmp_BSCmp_op2_9, 
      gen_15_cmp_BSCmp_op2_8, gen_15_cmp_BSCmp_op2_7, gen_15_cmp_BSCmp_op2_6, 
      gen_15_cmp_BSCmp_op2_5, gen_15_cmp_BSCmp_op2_4, gen_15_cmp_BSCmp_op2_3, 
      gen_15_cmp_BSCmp_op2_2, gen_15_cmp_BSCmp_op2_1, 
      gen_14_cmp_BSCmp_op2_16, gen_14_cmp_BSCmp_op2_15, 
      gen_14_cmp_BSCmp_op2_14, gen_14_cmp_BSCmp_op2_13, 
      gen_14_cmp_BSCmp_op2_12, gen_14_cmp_BSCmp_op2_11, 
      gen_14_cmp_BSCmp_op2_10, gen_14_cmp_BSCmp_op2_9, 
      gen_14_cmp_BSCmp_op2_8, gen_14_cmp_BSCmp_op2_7, gen_14_cmp_BSCmp_op2_6, 
      gen_14_cmp_BSCmp_op2_5, gen_14_cmp_BSCmp_op2_4, gen_14_cmp_BSCmp_op2_3, 
      gen_14_cmp_BSCmp_op2_2, gen_14_cmp_BSCmp_op2_1, 
      gen_13_cmp_BSCmp_op2_16, gen_13_cmp_BSCmp_op2_15, 
      gen_13_cmp_BSCmp_op2_14, gen_13_cmp_BSCmp_op2_13, 
      gen_13_cmp_BSCmp_op2_12, gen_13_cmp_BSCmp_op2_11, 
      gen_13_cmp_BSCmp_op2_10, gen_13_cmp_BSCmp_op2_9, 
      gen_13_cmp_BSCmp_op2_8, gen_13_cmp_BSCmp_op2_7, gen_13_cmp_BSCmp_op2_6, 
      gen_13_cmp_BSCmp_op2_5, gen_13_cmp_BSCmp_op2_4, gen_13_cmp_BSCmp_op2_3, 
      gen_13_cmp_BSCmp_op2_2, gen_13_cmp_BSCmp_op2_1, 
      gen_12_cmp_BSCmp_op2_16, gen_12_cmp_BSCmp_op2_15, 
      gen_12_cmp_BSCmp_op2_14, gen_12_cmp_BSCmp_op2_13, 
      gen_12_cmp_BSCmp_op2_12, gen_12_cmp_BSCmp_op2_11, 
      gen_12_cmp_BSCmp_op2_10, gen_12_cmp_BSCmp_op2_9, 
      gen_12_cmp_BSCmp_op2_8, gen_12_cmp_BSCmp_op2_7, gen_12_cmp_BSCmp_op2_6, 
      gen_12_cmp_BSCmp_op2_5, gen_12_cmp_BSCmp_op2_4, gen_12_cmp_BSCmp_op2_3, 
      gen_12_cmp_BSCmp_op2_2, gen_12_cmp_BSCmp_op2_1, 
      gen_11_cmp_BSCmp_op2_16, gen_11_cmp_BSCmp_op2_15, 
      gen_11_cmp_BSCmp_op2_14, gen_11_cmp_BSCmp_op2_13, 
      gen_11_cmp_BSCmp_op2_12, gen_11_cmp_BSCmp_op2_11, 
      gen_11_cmp_BSCmp_op2_10, gen_11_cmp_BSCmp_op2_9, 
      gen_11_cmp_BSCmp_op2_8, gen_11_cmp_BSCmp_op2_7, gen_11_cmp_BSCmp_op2_6, 
      gen_11_cmp_BSCmp_op2_5, gen_11_cmp_BSCmp_op2_4, gen_11_cmp_BSCmp_op2_3, 
      gen_11_cmp_BSCmp_op2_2, gen_11_cmp_BSCmp_op2_1, 
      gen_10_cmp_BSCmp_op2_16, gen_10_cmp_BSCmp_op2_15, 
      gen_10_cmp_BSCmp_op2_14, gen_10_cmp_BSCmp_op2_13, 
      gen_10_cmp_BSCmp_op2_12, gen_10_cmp_BSCmp_op2_11, 
      gen_10_cmp_BSCmp_op2_10, gen_10_cmp_BSCmp_op2_9, 
      gen_10_cmp_BSCmp_op2_8, gen_10_cmp_BSCmp_op2_7, gen_10_cmp_BSCmp_op2_6, 
      gen_10_cmp_BSCmp_op2_5, gen_10_cmp_BSCmp_op2_4, gen_10_cmp_BSCmp_op2_3, 
      gen_10_cmp_BSCmp_op2_2, gen_10_cmp_BSCmp_op2_1, gen_9_cmp_BSCmp_op2_16, 
      gen_9_cmp_BSCmp_op2_15, gen_9_cmp_BSCmp_op2_14, gen_9_cmp_BSCmp_op2_13, 
      gen_9_cmp_BSCmp_op2_12, gen_9_cmp_BSCmp_op2_11, gen_9_cmp_BSCmp_op2_10, 
      gen_9_cmp_BSCmp_op2_9, gen_9_cmp_BSCmp_op2_8, gen_9_cmp_BSCmp_op2_7, 
      gen_9_cmp_BSCmp_op2_6, gen_9_cmp_BSCmp_op2_5, gen_9_cmp_BSCmp_op2_4, 
      gen_9_cmp_BSCmp_op2_3, gen_9_cmp_BSCmp_op2_2, gen_9_cmp_BSCmp_op2_1, 
      gen_8_cmp_BSCmp_op2_16, gen_8_cmp_BSCmp_op2_15, gen_8_cmp_BSCmp_op2_14, 
      gen_8_cmp_BSCmp_op2_13, gen_8_cmp_BSCmp_op2_12, gen_8_cmp_BSCmp_op2_11, 
      gen_8_cmp_BSCmp_op2_10, gen_8_cmp_BSCmp_op2_9, gen_8_cmp_BSCmp_op2_8, 
      gen_8_cmp_BSCmp_op2_7, gen_8_cmp_BSCmp_op2_6, gen_8_cmp_BSCmp_op2_5, 
      gen_8_cmp_BSCmp_op2_4, gen_8_cmp_BSCmp_op2_3, gen_8_cmp_BSCmp_op2_2, 
      gen_8_cmp_BSCmp_op2_1, gen_7_cmp_BSCmp_op2_16, gen_7_cmp_BSCmp_op2_15, 
      gen_7_cmp_BSCmp_op2_14, gen_7_cmp_BSCmp_op2_13, gen_7_cmp_BSCmp_op2_12, 
      gen_7_cmp_BSCmp_op2_11, gen_7_cmp_BSCmp_op2_10, gen_7_cmp_BSCmp_op2_9, 
      gen_7_cmp_BSCmp_op2_8, gen_7_cmp_BSCmp_op2_7, gen_7_cmp_BSCmp_op2_6, 
      gen_7_cmp_BSCmp_op2_5, gen_7_cmp_BSCmp_op2_4, gen_7_cmp_BSCmp_op2_3, 
      gen_7_cmp_BSCmp_op2_2, gen_7_cmp_BSCmp_op2_1, gen_6_cmp_BSCmp_op2_16, 
      gen_6_cmp_BSCmp_op2_15, gen_6_cmp_BSCmp_op2_14, gen_6_cmp_BSCmp_op2_13, 
      gen_6_cmp_BSCmp_op2_12, gen_6_cmp_BSCmp_op2_11, gen_6_cmp_BSCmp_op2_10, 
      gen_6_cmp_BSCmp_op2_9, gen_6_cmp_BSCmp_op2_8, gen_6_cmp_BSCmp_op2_7, 
      gen_6_cmp_BSCmp_op2_6, gen_6_cmp_BSCmp_op2_5, gen_6_cmp_BSCmp_op2_4, 
      gen_6_cmp_BSCmp_op2_3, gen_6_cmp_BSCmp_op2_2, gen_6_cmp_BSCmp_op2_1, 
      gen_5_cmp_BSCmp_op2_16, gen_5_cmp_BSCmp_op2_15, gen_5_cmp_BSCmp_op2_14, 
      gen_5_cmp_BSCmp_op2_13, gen_5_cmp_BSCmp_op2_12, gen_5_cmp_BSCmp_op2_11, 
      gen_5_cmp_BSCmp_op2_10, gen_5_cmp_BSCmp_op2_9, gen_5_cmp_BSCmp_op2_8, 
      gen_5_cmp_BSCmp_op2_7, gen_5_cmp_BSCmp_op2_6, gen_5_cmp_BSCmp_op2_5, 
      gen_5_cmp_BSCmp_op2_4, gen_5_cmp_BSCmp_op2_3, gen_5_cmp_BSCmp_op2_2, 
      gen_5_cmp_BSCmp_op2_1, gen_4_cmp_BSCmp_op2_16, gen_4_cmp_BSCmp_op2_15, 
      gen_4_cmp_BSCmp_op2_14, gen_4_cmp_BSCmp_op2_13, gen_4_cmp_BSCmp_op2_12, 
      gen_4_cmp_BSCmp_op2_11, gen_4_cmp_BSCmp_op2_10, gen_4_cmp_BSCmp_op2_9, 
      gen_4_cmp_BSCmp_op2_8, gen_4_cmp_BSCmp_op2_7, gen_4_cmp_BSCmp_op2_6, 
      gen_4_cmp_BSCmp_op2_5, gen_4_cmp_BSCmp_op2_4, gen_4_cmp_BSCmp_op2_3, 
      gen_4_cmp_BSCmp_op2_2, gen_4_cmp_BSCmp_op2_1, gen_3_cmp_BSCmp_op2_16, 
      gen_3_cmp_BSCmp_op2_15, gen_3_cmp_BSCmp_op2_14, gen_3_cmp_BSCmp_op2_13, 
      gen_3_cmp_BSCmp_op2_12, gen_3_cmp_BSCmp_op2_11, gen_3_cmp_BSCmp_op2_10, 
      gen_3_cmp_BSCmp_op2_9, gen_3_cmp_BSCmp_op2_8, gen_3_cmp_BSCmp_op2_7, 
      gen_3_cmp_BSCmp_op2_6, gen_3_cmp_BSCmp_op2_5, gen_3_cmp_BSCmp_op2_4, 
      gen_3_cmp_BSCmp_op2_3, gen_3_cmp_BSCmp_op2_2, gen_3_cmp_BSCmp_op2_1, 
      gen_2_cmp_BSCmp_op2_16, gen_2_cmp_BSCmp_op2_15, gen_2_cmp_BSCmp_op2_14, 
      gen_2_cmp_BSCmp_op2_13, gen_2_cmp_BSCmp_op2_12, gen_2_cmp_BSCmp_op2_11, 
      gen_2_cmp_BSCmp_op2_10, gen_2_cmp_BSCmp_op2_9, gen_2_cmp_BSCmp_op2_8, 
      gen_2_cmp_BSCmp_op2_7, gen_2_cmp_BSCmp_op2_6, gen_2_cmp_BSCmp_op2_5, 
      gen_2_cmp_BSCmp_op2_4, gen_2_cmp_BSCmp_op2_3, gen_2_cmp_BSCmp_op2_2, 
      gen_2_cmp_BSCmp_op2_1, gen_1_cmp_BSCmp_op2_16, gen_1_cmp_BSCmp_op2_15, 
      gen_1_cmp_BSCmp_op2_14, gen_1_cmp_BSCmp_op2_13, gen_1_cmp_BSCmp_op2_12, 
      gen_1_cmp_BSCmp_op2_11, gen_1_cmp_BSCmp_op2_10, gen_1_cmp_BSCmp_op2_9, 
      gen_1_cmp_BSCmp_op2_8, gen_1_cmp_BSCmp_op2_7, gen_1_cmp_BSCmp_op2_6, 
      gen_1_cmp_BSCmp_op2_5, gen_1_cmp_BSCmp_op2_4, gen_1_cmp_BSCmp_op2_3, 
      gen_1_cmp_BSCmp_op2_2, gen_1_cmp_BSCmp_op2_1, gen_0_cmp_BSCmp_op2_16, 
      gen_0_cmp_BSCmp_op2_15, gen_0_cmp_BSCmp_op2_14, gen_0_cmp_BSCmp_op2_13, 
      gen_0_cmp_BSCmp_op2_12, gen_0_cmp_BSCmp_op2_11, gen_0_cmp_BSCmp_op2_10, 
      gen_0_cmp_BSCmp_op2_9, gen_0_cmp_BSCmp_op2_8, gen_0_cmp_BSCmp_op2_7, 
      gen_0_cmp_BSCmp_op2_6, gen_0_cmp_BSCmp_op2_5, gen_0_cmp_BSCmp_op2_4, 
      gen_0_cmp_BSCmp_op2_3, gen_0_cmp_BSCmp_op2_2, gen_0_cmp_BSCmp_op2_1, 
      nx6, gen_0_cmp_mReg_0, nx26, nx34, gen_0_cmp_mReg_1, nx46, nx48, nx58, 
      nx62, gen_0_cmp_mReg_2, nx74, nx76, nx80, nx84, gen_0_cmp_mReg_3, nx96, 
      nx98, nx102, nx106, gen_0_cmp_mReg_4, nx118, nx120, nx124, nx128, 
      gen_0_cmp_mReg_5, nx140, nx142, nx146, nx150, gen_0_cmp_mReg_6, nx162, 
      nx164, nx168, nx172, gen_0_cmp_mReg_7, nx184, nx186, nx190, nx194, 
      gen_0_cmp_mReg_8, nx206, nx208, nx212, nx216, gen_0_cmp_mReg_9, nx228, 
      nx230, nx234, nx238, gen_0_cmp_mReg_10, nx250, nx252, nx256, nx260, 
      gen_0_cmp_mReg_11, nx272, nx274, nx278, nx282, gen_0_cmp_mReg_12, 
      nx294, nx296, nx300, nx304, gen_0_cmp_mReg_13, nx316, nx318, nx322, 
      nx326, gen_0_cmp_mReg_14, nx338, nx340, nx344, nx348, 
      gen_0_cmp_mReg_15, nx360, nx362, nx366, nx370, nx376, nx380, nx392, 
      gen_1_cmp_mReg_0, nx412, nx420, gen_1_cmp_mReg_1, nx432, nx434, nx444, 
      nx448, gen_1_cmp_mReg_2, nx460, nx462, nx466, nx470, gen_1_cmp_mReg_3, 
      nx482, nx484, nx488, nx492, gen_1_cmp_mReg_4, nx504, nx506, nx510, 
      nx514, gen_1_cmp_mReg_5, nx526, nx528, nx532, nx536, gen_1_cmp_mReg_6, 
      nx548, nx550, nx554, nx558, gen_1_cmp_mReg_7, nx570, nx572, nx576, 
      nx580, gen_1_cmp_mReg_8, nx592, nx594, nx598, nx602, gen_1_cmp_mReg_9, 
      nx614, nx616, nx620, nx624, gen_1_cmp_mReg_10, nx636, nx638, nx642, 
      nx646, gen_1_cmp_mReg_11, nx658, nx660, nx664, nx668, 
      gen_1_cmp_mReg_12, nx680, nx682, nx686, nx690, gen_1_cmp_mReg_13, 
      nx702, nx704, nx708, nx712, gen_1_cmp_mReg_14, nx724, nx726, nx730, 
      nx734, gen_1_cmp_mReg_15, nx746, nx748, nx752, nx756, nx762, nx766, 
      nx778, gen_2_cmp_mReg_0, nx798, nx806, gen_2_cmp_mReg_1, nx818, nx820, 
      nx830, nx834, gen_2_cmp_mReg_2, nx846, nx848, nx852, nx856, 
      gen_2_cmp_mReg_3, nx868, nx870, nx874, nx878, gen_2_cmp_mReg_4, nx890, 
      nx892, nx896, nx900, gen_2_cmp_mReg_5, nx912, nx914, nx918, nx922, 
      gen_2_cmp_mReg_6, nx934, nx936, nx940, nx944, gen_2_cmp_mReg_7, nx956, 
      nx958, nx962, nx966, gen_2_cmp_mReg_8, nx978, nx980, nx984, nx988, 
      gen_2_cmp_mReg_9, nx1000, nx1002, nx1006, nx1010, gen_2_cmp_mReg_10, 
      nx1022, nx1024, nx1028, nx1032, gen_2_cmp_mReg_11, nx1044, nx1046, 
      nx1050, nx1054, gen_2_cmp_mReg_12, nx1066, nx1068, nx1072, nx1076, 
      gen_2_cmp_mReg_13, nx1088, nx1090, nx1094, nx1098, gen_2_cmp_mReg_14, 
      nx1110, nx1112, nx1116, nx1120, gen_2_cmp_mReg_15, nx1132, nx1134, 
      nx1138, nx1142, nx1148, nx1152, nx1164, gen_3_cmp_mReg_0, nx1184, 
      nx1192, gen_3_cmp_mReg_1, nx1204, nx1206, nx1216, nx1220, 
      gen_3_cmp_mReg_2, nx1232, nx1234, nx1238, nx1242, gen_3_cmp_mReg_3, 
      nx1254, nx1256, nx1260, nx1264, gen_3_cmp_mReg_4, nx1276, nx1278, 
      nx1282, nx1286, gen_3_cmp_mReg_5, nx1298, nx1300, nx1304, nx1308, 
      gen_3_cmp_mReg_6, nx1320, nx1322, nx1326, nx1330, gen_3_cmp_mReg_7, 
      nx1342, nx1344, nx1348, nx1352, gen_3_cmp_mReg_8, nx1364, nx1366, 
      nx1370, nx1374, gen_3_cmp_mReg_9, nx1386, nx1388, nx1392, nx1396, 
      gen_3_cmp_mReg_10, nx1408, nx1410, nx1414, nx1418, gen_3_cmp_mReg_11, 
      nx1430, nx1432, nx1436, nx1440, gen_3_cmp_mReg_12, nx1452, nx1454, 
      nx1458, nx1462, gen_3_cmp_mReg_13, nx1474, nx1476, nx1480, nx1484, 
      gen_3_cmp_mReg_14, nx1496, nx1498, nx1502, nx1506, gen_3_cmp_mReg_15, 
      nx1518, nx1520, nx1524, nx1528, nx1534, nx1538, nx1550, 
      gen_4_cmp_mReg_0, nx1570, nx1578, gen_4_cmp_mReg_1, nx1590, nx1592, 
      nx1602, nx1606, gen_4_cmp_mReg_2, nx1618, nx1620, nx1624, nx1628, 
      gen_4_cmp_mReg_3, nx1640, nx1642, nx1646, nx1650, gen_4_cmp_mReg_4, 
      nx1662, nx1664, nx1668, nx1672, gen_4_cmp_mReg_5, nx1684, nx1686, 
      nx1690, nx1694, gen_4_cmp_mReg_6, nx1706, nx1708, nx1712, nx1716, 
      gen_4_cmp_mReg_7, nx1728, nx1730, nx1734, nx1738, gen_4_cmp_mReg_8, 
      nx1750, nx1752, nx1756, nx1760, gen_4_cmp_mReg_9, nx1772, nx1774, 
      nx1778, nx1782, gen_4_cmp_mReg_10, nx1794, nx1796, nx1800, nx1804, 
      gen_4_cmp_mReg_11, nx1816, nx1818, nx1822, nx1826, gen_4_cmp_mReg_12, 
      nx1838, nx1840, nx1844, nx1848, gen_4_cmp_mReg_13, nx1860, nx1862, 
      nx1866, nx1870, gen_4_cmp_mReg_14, nx1882, nx1884, nx1888, nx1892, 
      gen_4_cmp_mReg_15, nx1904, nx1906, nx1910, nx1914, nx1920, nx1924, 
      nx1936, gen_5_cmp_mReg_0, nx1956, nx1964, gen_5_cmp_mReg_1, nx1976, 
      nx1978, nx1988, nx1992, gen_5_cmp_mReg_2, nx2004, nx2006, nx2010, 
      nx2014, gen_5_cmp_mReg_3, nx2026, nx2028, nx2032, nx2036, 
      gen_5_cmp_mReg_4, nx2048, nx2050, nx2054, nx2058, gen_5_cmp_mReg_5, 
      nx2070, nx2072, nx2076, nx2080, gen_5_cmp_mReg_6, nx2092, nx2094, 
      nx2098, nx2102, gen_5_cmp_mReg_7, nx2114, nx2116, nx2120, nx2124, 
      gen_5_cmp_mReg_8, nx2136, nx2138, nx2142, nx2146, gen_5_cmp_mReg_9, 
      nx2158, nx2160, nx2164, nx2168, gen_5_cmp_mReg_10, nx2180, nx2182, 
      nx2186, nx2190, gen_5_cmp_mReg_11, nx2202, nx2204, nx2208, nx2212, 
      gen_5_cmp_mReg_12, nx2224, nx2226, nx2230, nx2234, gen_5_cmp_mReg_13, 
      nx2246, nx2248, nx2252, nx2256, gen_5_cmp_mReg_14, nx2268, nx2270, 
      nx2274, nx2278, gen_5_cmp_mReg_15, nx2290, nx2292, nx2296, nx2300, 
      nx2306, nx2310, nx2322, gen_6_cmp_mReg_0, nx2342, nx2350, 
      gen_6_cmp_mReg_1, nx2362, nx2364, nx2374, nx2378, gen_6_cmp_mReg_2, 
      nx2390, nx2392, nx2396, nx2400, gen_6_cmp_mReg_3, nx2412, nx2414, 
      nx2418, nx2422, gen_6_cmp_mReg_4, nx2434, nx2436, nx2440, nx2444, 
      gen_6_cmp_mReg_5, nx2456, nx2458, nx2462, nx2466, gen_6_cmp_mReg_6, 
      nx2478, nx2480, nx2484, nx2488, gen_6_cmp_mReg_7, nx2500, nx2502, 
      nx2506, nx2510, gen_6_cmp_mReg_8, nx2522, nx2524, nx2528, nx2532, 
      gen_6_cmp_mReg_9, nx2544, nx2546, nx2550, nx2554, gen_6_cmp_mReg_10, 
      nx2566, nx2568, nx2572, nx2576, gen_6_cmp_mReg_11, nx2588, nx2590, 
      nx2594, nx2598, gen_6_cmp_mReg_12, nx2610, nx2612, nx2616, nx2620, 
      gen_6_cmp_mReg_13, nx2632, nx2634, nx2638, nx2642, gen_6_cmp_mReg_14, 
      nx2654, nx2656, nx2660, nx2664, gen_6_cmp_mReg_15, nx2676, nx2678, 
      nx2682, nx2686, nx2692, nx2696, nx2708, gen_7_cmp_mReg_0, nx2728, 
      nx2736, gen_7_cmp_mReg_1, nx2748, nx2750, nx2760, nx2764, 
      gen_7_cmp_mReg_2, nx2776, nx2778, nx2782, nx2786, gen_7_cmp_mReg_3, 
      nx2798, nx2800, nx2804, nx2808, gen_7_cmp_mReg_4, nx2820, nx2822, 
      nx2826, nx2830, gen_7_cmp_mReg_5, nx2842, nx2844, nx2848, nx2852, 
      gen_7_cmp_mReg_6, nx2864, nx2866, nx2870, nx2874, gen_7_cmp_mReg_7, 
      nx2886, nx2888, nx2892, nx2896, gen_7_cmp_mReg_8, nx2908, nx2910, 
      nx2914, nx2918, gen_7_cmp_mReg_9, nx2930, nx2932, nx2936, nx2940, 
      gen_7_cmp_mReg_10, nx2952, nx2954, nx2958, nx2962, gen_7_cmp_mReg_11, 
      nx2974, nx2976, nx2980, nx2984, gen_7_cmp_mReg_12, nx2996, nx2998, 
      nx3002, nx3006, gen_7_cmp_mReg_13, nx3018, nx3020, nx3024, nx3028, 
      gen_7_cmp_mReg_14, nx3040, nx3042, nx3046, nx3050, gen_7_cmp_mReg_15, 
      nx3062, nx3064, nx3068, nx3072, nx3078, nx3082, nx3094, 
      gen_8_cmp_mReg_0, nx3114, nx3122, gen_8_cmp_mReg_1, nx3134, nx3136, 
      nx3146, nx3150, gen_8_cmp_mReg_2, nx3162, nx3164, nx3168, nx3172, 
      gen_8_cmp_mReg_3, nx3184, nx3186, nx3190, nx3194, gen_8_cmp_mReg_4, 
      nx3206, nx3208, nx3212, nx3216, gen_8_cmp_mReg_5, nx3228, nx3230, 
      nx3234, nx3238, gen_8_cmp_mReg_6, nx3250, nx3252, nx3256, nx3260, 
      gen_8_cmp_mReg_7, nx3272, nx3274, nx3278, nx3282, gen_8_cmp_mReg_8, 
      nx3294, nx3296, nx3300, nx3304, gen_8_cmp_mReg_9, nx3316, nx3318, 
      nx3322, nx3326, gen_8_cmp_mReg_10, nx3338, nx3340, nx3344, nx3348, 
      gen_8_cmp_mReg_11, nx3360, nx3362, nx3366, nx3370, gen_8_cmp_mReg_12, 
      nx3382, nx3384, nx3388, nx3392, gen_8_cmp_mReg_13, nx3404, nx3406, 
      nx3410, nx3414, gen_8_cmp_mReg_14, nx3426, nx3428, nx3432, nx3436, 
      gen_8_cmp_mReg_15, nx3448, nx3450, nx3454, nx3458, nx3464, nx3468, 
      nx3480, gen_9_cmp_mReg_0, nx3500, nx3508, gen_9_cmp_mReg_1, nx3520, 
      nx3522, nx3532, nx3536, gen_9_cmp_mReg_2, nx3548, nx3550, nx3554, 
      nx3558, gen_9_cmp_mReg_3, nx3570, nx3572, nx3576, nx3580, 
      gen_9_cmp_mReg_4, nx3592, nx3594, nx3598, nx3602, gen_9_cmp_mReg_5, 
      nx3614, nx3616, nx3620, nx3624, gen_9_cmp_mReg_6, nx3636, nx3638, 
      nx3642, nx3646, gen_9_cmp_mReg_7, nx3658, nx3660, nx3664, nx3668, 
      gen_9_cmp_mReg_8, nx3680, nx3682, nx3686, nx3690, gen_9_cmp_mReg_9, 
      nx3702, nx3704, nx3708, nx3712, gen_9_cmp_mReg_10, nx3724, nx3726, 
      nx3730, nx3734, gen_9_cmp_mReg_11, nx3746, nx3748, nx3752, nx3756, 
      gen_9_cmp_mReg_12, nx3768, nx3770, nx3774, nx3778, gen_9_cmp_mReg_13, 
      nx3790, nx3792, nx3796, nx3800, gen_9_cmp_mReg_14, nx3812, nx3814, 
      nx3818, nx3822, gen_9_cmp_mReg_15, nx3834, nx3836, nx3840, nx3844, 
      nx3850, nx3854, nx3866, gen_10_cmp_mReg_0, nx3886, nx3894, 
      gen_10_cmp_mReg_1, nx3906, nx3908, nx3918, nx3922, gen_10_cmp_mReg_2, 
      nx3934, nx3936, nx3940, nx3944, gen_10_cmp_mReg_3, nx3956, nx3958, 
      nx3962, nx3966, gen_10_cmp_mReg_4, nx3978, nx3980, nx3984, nx3988, 
      gen_10_cmp_mReg_5, nx4000, nx4002, nx4006, nx4010, gen_10_cmp_mReg_6, 
      nx4022, nx4024, nx4028, nx4032, gen_10_cmp_mReg_7, nx4044, nx4046, 
      nx4050, nx4054, gen_10_cmp_mReg_8, nx4066, nx4068, nx4072, nx4076, 
      gen_10_cmp_mReg_9, nx4088, nx4090, nx4094, nx4098, gen_10_cmp_mReg_10, 
      nx4110, nx4112, nx4116, nx4120, gen_10_cmp_mReg_11, nx4132, nx4134, 
      nx4138, nx4142, gen_10_cmp_mReg_12, nx4154, nx4156, nx4160, nx4164, 
      gen_10_cmp_mReg_13, nx4176, nx4178, nx4182, nx4186, gen_10_cmp_mReg_14, 
      nx4198, nx4200, nx4204, nx4208, gen_10_cmp_mReg_15, nx4220, nx4222, 
      nx4226, nx4230, nx4236, nx4240, nx4252, gen_11_cmp_mReg_0, nx4272, 
      nx4280, gen_11_cmp_mReg_1, nx4292, nx4294, nx4304, nx4308, 
      gen_11_cmp_mReg_2, nx4320, nx4322, nx4326, nx4330, gen_11_cmp_mReg_3, 
      nx4342, nx4344, nx4348, nx4352, gen_11_cmp_mReg_4, nx4364, nx4366, 
      nx4370, nx4374, gen_11_cmp_mReg_5, nx4386, nx4388, nx4392, nx4396, 
      gen_11_cmp_mReg_6, nx4408, nx4410, nx4414, nx4418, gen_11_cmp_mReg_7, 
      nx4430, nx4432, nx4436, nx4440, gen_11_cmp_mReg_8, nx4452, nx4454, 
      nx4458, nx4462, gen_11_cmp_mReg_9, nx4474, nx4476, nx4480, nx4484, 
      gen_11_cmp_mReg_10, nx4496, nx4498, nx4502, nx4506, gen_11_cmp_mReg_11, 
      nx4518, nx4520, nx4524, nx4528, gen_11_cmp_mReg_12, nx4540, nx4542, 
      nx4546, nx4550, gen_11_cmp_mReg_13, nx4562, nx4564, nx4568, nx4572, 
      gen_11_cmp_mReg_14, nx4584, nx4586, nx4590, nx4594, gen_11_cmp_mReg_15, 
      nx4606, nx4608, nx4612, nx4616, nx4622, nx4626, nx4638, 
      gen_12_cmp_mReg_0, nx4658, nx4666, gen_12_cmp_mReg_1, nx4678, nx4680, 
      nx4690, nx4694, gen_12_cmp_mReg_2, nx4706, nx4708, nx4712, nx4716, 
      gen_12_cmp_mReg_3, nx4728, nx4730, nx4734, nx4738, gen_12_cmp_mReg_4, 
      nx4750, nx4752, nx4756, nx4760, gen_12_cmp_mReg_5, nx4772, nx4774, 
      nx4778, nx4782, gen_12_cmp_mReg_6, nx4794, nx4796, nx4800, nx4804, 
      gen_12_cmp_mReg_7, nx4816, nx4818, nx4822, nx4826, gen_12_cmp_mReg_8, 
      nx4838, nx4840, nx4844, nx4848, gen_12_cmp_mReg_9, nx4860, nx4862, 
      nx4866, nx4870, gen_12_cmp_mReg_10, nx4882, nx4884, nx4888, nx4892, 
      gen_12_cmp_mReg_11, nx4904, nx4906, nx4910, nx4914, gen_12_cmp_mReg_12, 
      nx4926, nx4928, nx4932, nx4936, gen_12_cmp_mReg_13, nx4948, nx4950, 
      nx4954, nx4958, gen_12_cmp_mReg_14, nx4970, nx4972, nx4976, nx4980, 
      gen_12_cmp_mReg_15, nx4992, nx4994, nx4998, nx5002, nx5008, nx5012, 
      nx5024, gen_13_cmp_mReg_0, nx5044, nx5052, gen_13_cmp_mReg_1, nx5064, 
      nx5066, nx5076, nx5080, gen_13_cmp_mReg_2, nx5092, nx5094, nx5098, 
      nx5102, gen_13_cmp_mReg_3, nx5114, nx5116, nx5120, nx5124, 
      gen_13_cmp_mReg_4, nx5136, nx5138, nx5142, nx5146, gen_13_cmp_mReg_5, 
      nx5158, nx5160, nx5164, nx5168, gen_13_cmp_mReg_6, nx5180, nx5182, 
      nx5186, nx5190, gen_13_cmp_mReg_7, nx5202, nx5204, nx5208, nx5212, 
      gen_13_cmp_mReg_8, nx5224, nx5226, nx5230, nx5234, gen_13_cmp_mReg_9, 
      nx5246, nx5248, nx5252, nx5256, gen_13_cmp_mReg_10, nx5268, nx5270, 
      nx5274, nx5278, gen_13_cmp_mReg_11, nx5290, nx5292, nx5296, nx5300, 
      gen_13_cmp_mReg_12, nx5312, nx5314, nx5318, nx5322, gen_13_cmp_mReg_13, 
      nx5334, nx5336, nx5340, nx5344, gen_13_cmp_mReg_14, nx5356, nx5358, 
      nx5362, nx5366, gen_13_cmp_mReg_15, nx5378, nx5380, nx5384, nx5388, 
      nx5394, nx5398, nx5410, gen_14_cmp_mReg_0, nx5430, nx5438, 
      gen_14_cmp_mReg_1, nx5450, nx5452, nx5462, nx5466, gen_14_cmp_mReg_2, 
      nx5478, nx5480, nx5484, nx5488, gen_14_cmp_mReg_3, nx5500, nx5502, 
      nx5506, nx5510, gen_14_cmp_mReg_4, nx5522, nx5524, nx5528, nx5532, 
      gen_14_cmp_mReg_5, nx5544, nx5546, nx5550, nx5554, gen_14_cmp_mReg_6, 
      nx5566, nx5568, nx5572, nx5576, gen_14_cmp_mReg_7, nx5588, nx5590, 
      nx5594, nx5598, gen_14_cmp_mReg_8, nx5610, nx5612, nx5616, nx5620, 
      gen_14_cmp_mReg_9, nx5632, nx5634, nx5638, nx5642, gen_14_cmp_mReg_10, 
      nx5654, nx5656, nx5660, nx5664, gen_14_cmp_mReg_11, nx5676, nx5678, 
      nx5682, nx5686, gen_14_cmp_mReg_12, nx5698, nx5700, nx5704, nx5708, 
      gen_14_cmp_mReg_13, nx5720, nx5722, nx5726, nx5730, gen_14_cmp_mReg_14, 
      nx5742, nx5744, nx5748, nx5752, gen_14_cmp_mReg_15, nx5764, nx5766, 
      nx5770, nx5774, nx5780, nx5784, nx5796, gen_15_cmp_mReg_0, nx5816, 
      nx5824, gen_15_cmp_mReg_1, nx5836, nx5838, nx5848, nx5852, 
      gen_15_cmp_mReg_2, nx5864, nx5866, nx5870, nx5874, gen_15_cmp_mReg_3, 
      nx5886, nx5888, nx5892, nx5896, gen_15_cmp_mReg_4, nx5908, nx5910, 
      nx5914, nx5918, gen_15_cmp_mReg_5, nx5930, nx5932, nx5936, nx5940, 
      gen_15_cmp_mReg_6, nx5952, nx5954, nx5958, nx5962, gen_15_cmp_mReg_7, 
      nx5974, nx5976, nx5980, nx5984, gen_15_cmp_mReg_8, nx5996, nx5998, 
      nx6002, nx6006, gen_15_cmp_mReg_9, nx6018, nx6020, nx6024, nx6028, 
      gen_15_cmp_mReg_10, nx6040, nx6042, nx6046, nx6050, gen_15_cmp_mReg_11, 
      nx6062, nx6064, nx6068, nx6072, gen_15_cmp_mReg_12, nx6084, nx6086, 
      nx6090, nx6094, gen_15_cmp_mReg_13, nx6106, nx6108, nx6112, nx6116, 
      gen_15_cmp_mReg_14, nx6128, nx6130, nx6134, nx6138, gen_15_cmp_mReg_15, 
      nx6150, nx6152, nx6156, nx6160, nx6166, nx6170, nx6182, 
      gen_16_cmp_mReg_0, nx6202, nx6210, gen_16_cmp_mReg_1, nx6222, nx6224, 
      nx6234, nx6238, gen_16_cmp_mReg_2, nx6250, nx6252, nx6256, nx6260, 
      gen_16_cmp_mReg_3, nx6272, nx6274, nx6278, nx6282, gen_16_cmp_mReg_4, 
      nx6294, nx6296, nx6300, nx6304, gen_16_cmp_mReg_5, nx6316, nx6318, 
      nx6322, nx6326, gen_16_cmp_mReg_6, nx6338, nx6340, nx6344, nx6348, 
      gen_16_cmp_mReg_7, nx6360, nx6362, nx6366, nx6370, gen_16_cmp_mReg_8, 
      nx6382, nx6384, nx6388, nx6392, gen_16_cmp_mReg_9, nx6404, nx6406, 
      nx6410, nx6414, gen_16_cmp_mReg_10, nx6426, nx6428, nx6432, nx6436, 
      gen_16_cmp_mReg_11, nx6448, nx6450, nx6454, nx6458, gen_16_cmp_mReg_12, 
      nx6470, nx6472, nx6476, nx6480, gen_16_cmp_mReg_13, nx6492, nx6494, 
      nx6498, nx6502, gen_16_cmp_mReg_14, nx6514, nx6516, nx6520, nx6524, 
      gen_16_cmp_mReg_15, nx6536, nx6538, nx6542, nx6546, nx6552, nx6556, 
      nx6568, gen_17_cmp_mReg_0, nx6588, nx6596, gen_17_cmp_mReg_1, nx6608, 
      nx6610, nx6620, nx6624, gen_17_cmp_mReg_2, nx6636, nx6638, nx6642, 
      nx6646, gen_17_cmp_mReg_3, nx6658, nx6660, nx6664, nx6668, 
      gen_17_cmp_mReg_4, nx6680, nx6682, nx6686, nx6690, gen_17_cmp_mReg_5, 
      nx6702, nx6704, nx6708, nx6712, gen_17_cmp_mReg_6, nx6724, nx6726, 
      nx6730, nx6734, gen_17_cmp_mReg_7, nx6746, nx6748, nx6752, nx6756, 
      gen_17_cmp_mReg_8, nx6768, nx6770, nx6774, nx6778, gen_17_cmp_mReg_9, 
      nx6790, nx6792, nx6796, nx6800, gen_17_cmp_mReg_10, nx6812, nx6814, 
      nx6818, nx6822, gen_17_cmp_mReg_11, nx6834, nx6836, nx6840, nx6844, 
      gen_17_cmp_mReg_12, nx6856, nx6858, nx6862, nx6866, gen_17_cmp_mReg_13, 
      nx6878, nx6880, nx6884, nx6888, gen_17_cmp_mReg_14, nx6900, nx6902, 
      nx6906, nx6910, gen_17_cmp_mReg_15, nx6922, nx6924, nx6928, nx6932, 
      nx6938, nx6942, nx6954, gen_18_cmp_mReg_0, nx6974, nx6982, 
      gen_18_cmp_mReg_1, nx6994, nx6996, nx7006, nx7010, gen_18_cmp_mReg_2, 
      nx7022, nx7024, nx7028, nx7032, gen_18_cmp_mReg_3, nx7044, nx7046, 
      nx7050, nx7054, gen_18_cmp_mReg_4, nx7066, nx7068, nx7072, nx7076, 
      gen_18_cmp_mReg_5, nx7088, nx7090, nx7094, nx7098, gen_18_cmp_mReg_6, 
      nx7110, nx7112, nx7116, nx7120, gen_18_cmp_mReg_7, nx7132, nx7134, 
      nx7138, nx7142, gen_18_cmp_mReg_8, nx7154, nx7156, nx7160, nx7164, 
      gen_18_cmp_mReg_9, nx7176, nx7178, nx7182, nx7186, gen_18_cmp_mReg_10, 
      nx7198, nx7200, nx7204, nx7208, gen_18_cmp_mReg_11, nx7220, nx7222, 
      nx7226, nx7230, gen_18_cmp_mReg_12, nx7242, nx7244, nx7248, nx7252, 
      gen_18_cmp_mReg_13, nx7264, nx7266, nx7270, nx7274, gen_18_cmp_mReg_14, 
      nx7286, nx7288, nx7292, nx7296, gen_18_cmp_mReg_15, nx7308, nx7310, 
      nx7314, nx7318, nx7324, nx7328, nx7340, gen_19_cmp_mReg_0, nx7360, 
      nx7368, gen_19_cmp_mReg_1, nx7380, nx7382, nx7392, nx7396, 
      gen_19_cmp_mReg_2, nx7408, nx7410, nx7414, nx7418, gen_19_cmp_mReg_3, 
      nx7430, nx7432, nx7436, nx7440, gen_19_cmp_mReg_4, nx7452, nx7454, 
      nx7458, nx7462, gen_19_cmp_mReg_5, nx7474, nx7476, nx7480, nx7484, 
      gen_19_cmp_mReg_6, nx7496, nx7498, nx7502, nx7506, gen_19_cmp_mReg_7, 
      nx7518, nx7520, nx7524, nx7528, gen_19_cmp_mReg_8, nx7540, nx7542, 
      nx7546, nx7550, gen_19_cmp_mReg_9, nx7562, nx7564, nx7568, nx7572, 
      gen_19_cmp_mReg_10, nx7584, nx7586, nx7590, nx7594, gen_19_cmp_mReg_11, 
      nx7606, nx7608, nx7612, nx7616, gen_19_cmp_mReg_12, nx7628, nx7630, 
      nx7634, nx7638, gen_19_cmp_mReg_13, nx7650, nx7652, nx7656, nx7660, 
      gen_19_cmp_mReg_14, nx7672, nx7674, nx7678, nx7682, gen_19_cmp_mReg_15, 
      nx7694, nx7696, nx7700, nx7704, nx7710, nx7714, nx7726, 
      gen_20_cmp_mReg_0, nx7746, nx7754, gen_20_cmp_mReg_1, nx7766, nx7768, 
      nx7778, nx7782, gen_20_cmp_mReg_2, nx7794, nx7796, nx7800, nx7804, 
      gen_20_cmp_mReg_3, nx7816, nx7818, nx7822, nx7826, gen_20_cmp_mReg_4, 
      nx7838, nx7840, nx7844, nx7848, gen_20_cmp_mReg_5, nx7860, nx7862, 
      nx7866, nx7870, gen_20_cmp_mReg_6, nx7882, nx7884, nx7888, nx7892, 
      gen_20_cmp_mReg_7, nx7904, nx7906, nx7910, nx7914, gen_20_cmp_mReg_8, 
      nx7926, nx7928, nx7932, nx7936, gen_20_cmp_mReg_9, nx7948, nx7950, 
      nx7954, nx7958, gen_20_cmp_mReg_10, nx7970, nx7972, nx7976, nx7980, 
      gen_20_cmp_mReg_11, nx7992, nx7994, nx7998, nx8002, gen_20_cmp_mReg_12, 
      nx8014, nx8016, nx8020, nx8024, gen_20_cmp_mReg_13, nx8036, nx8038, 
      nx8042, nx8046, gen_20_cmp_mReg_14, nx8058, nx8060, nx8064, nx8068, 
      gen_20_cmp_mReg_15, nx8080, nx8082, nx8086, nx8090, nx8096, nx8100, 
      nx8112, gen_21_cmp_mReg_0, nx8132, nx8140, gen_21_cmp_mReg_1, nx8152, 
      nx8154, nx8164, nx8168, gen_21_cmp_mReg_2, nx8180, nx8182, nx8186, 
      nx8190, gen_21_cmp_mReg_3, nx8202, nx8204, nx8208, nx8212, 
      gen_21_cmp_mReg_4, nx8224, nx8226, nx8230, nx8234, gen_21_cmp_mReg_5, 
      nx8246, nx8248, nx8252, nx8256, gen_21_cmp_mReg_6, nx8268, nx8270, 
      nx8274, nx8278, gen_21_cmp_mReg_7, nx8290, nx8292, nx8296, nx8300, 
      gen_21_cmp_mReg_8, nx8312, nx8314, nx8318, nx8322, gen_21_cmp_mReg_9, 
      nx8334, nx8336, nx8340, nx8344, gen_21_cmp_mReg_10, nx8356, nx8358, 
      nx8362, nx8366, gen_21_cmp_mReg_11, nx8378, nx8380, nx8384, nx8388, 
      gen_21_cmp_mReg_12, nx8400, nx8402, nx8406, nx8410, gen_21_cmp_mReg_13, 
      nx8422, nx8424, nx8428, nx8432, gen_21_cmp_mReg_14, nx8444, nx8446, 
      nx8450, nx8454, gen_21_cmp_mReg_15, nx8466, nx8468, nx8472, nx8476, 
      nx8482, nx8486, nx8498, gen_22_cmp_mReg_0, nx8518, nx8526, 
      gen_22_cmp_mReg_1, nx8538, nx8540, nx8550, nx8554, gen_22_cmp_mReg_2, 
      nx8566, nx8568, nx8572, nx8576, gen_22_cmp_mReg_3, nx8588, nx8590, 
      nx8594, nx8598, gen_22_cmp_mReg_4, nx8610, nx8612, nx8616, nx8620, 
      gen_22_cmp_mReg_5, nx8632, nx8634, nx8638, nx8642, gen_22_cmp_mReg_6, 
      nx8654, nx8656, nx8660, nx8664, gen_22_cmp_mReg_7, nx8676, nx8678, 
      nx8682, nx8686, gen_22_cmp_mReg_8, nx8698, nx8700, nx8704, nx8708, 
      gen_22_cmp_mReg_9, nx8720, nx8722, nx8726, nx8730, gen_22_cmp_mReg_10, 
      nx8742, nx8744, nx8748, nx8752, gen_22_cmp_mReg_11, nx8764, nx8766, 
      nx8770, nx8774, gen_22_cmp_mReg_12, nx8786, nx8788, nx8792, nx8796, 
      gen_22_cmp_mReg_13, nx8808, nx8810, nx8814, nx8818, gen_22_cmp_mReg_14, 
      nx8830, nx8832, nx8836, nx8840, gen_22_cmp_mReg_15, nx8852, nx8854, 
      nx8858, nx8862, nx8868, nx8872, nx8884, gen_23_cmp_mReg_0, nx8904, 
      nx8912, gen_23_cmp_mReg_1, nx8924, nx8926, nx8936, nx8940, 
      gen_23_cmp_mReg_2, nx8952, nx8954, nx8958, nx8962, gen_23_cmp_mReg_3, 
      nx8974, nx8976, nx8980, nx8984, gen_23_cmp_mReg_4, nx8996, nx8998, 
      nx9002, nx9006, gen_23_cmp_mReg_5, nx9018, nx9020, nx9024, nx9028, 
      gen_23_cmp_mReg_6, nx9040, nx9042, nx9046, nx9050, gen_23_cmp_mReg_7, 
      nx9062, nx9064, nx9068, nx9072, gen_23_cmp_mReg_8, nx9084, nx9086, 
      nx9090, nx9094, gen_23_cmp_mReg_9, nx9106, nx9108, nx9112, nx9116, 
      gen_23_cmp_mReg_10, nx9128, nx9130, nx9134, nx9138, gen_23_cmp_mReg_11, 
      nx9150, nx9152, nx9156, nx9160, gen_23_cmp_mReg_12, nx9172, nx9174, 
      nx9178, nx9182, gen_23_cmp_mReg_13, nx9194, nx9196, nx9200, nx9204, 
      gen_23_cmp_mReg_14, nx9216, nx9218, nx9222, nx9226, gen_23_cmp_mReg_15, 
      nx9238, nx9240, nx9244, nx9248, nx9254, nx9258, nx9270, 
      gen_24_cmp_mReg_0, nx9290, nx9298, gen_24_cmp_mReg_1, nx9310, nx9312, 
      nx9322, nx9326, gen_24_cmp_mReg_2, nx9338, nx9340, nx9344, nx9348, 
      gen_24_cmp_mReg_3, nx9360, nx9362, nx9366, nx9370, gen_24_cmp_mReg_4, 
      nx9382, nx9384, nx9388, nx9392, gen_24_cmp_mReg_5, nx9404, nx9406, 
      nx9410, nx9414, gen_24_cmp_mReg_6, nx9426, nx9428, nx9432, nx9436, 
      gen_24_cmp_mReg_7, nx9448, nx9450, nx9454, nx9458, gen_24_cmp_mReg_8, 
      nx9470, nx9472, nx9476, nx9480, gen_24_cmp_mReg_9, nx9492, nx9494, 
      nx9498, nx9502, gen_24_cmp_mReg_10, nx9514, nx9516, nx9520, nx9524, 
      gen_24_cmp_mReg_11, nx9536, nx9538, nx9542, nx9546, gen_24_cmp_mReg_12, 
      nx9558, nx9560, nx9564, nx9568, gen_24_cmp_mReg_13, nx9580, nx9582, 
      nx9586, nx9590, gen_24_cmp_mReg_14, nx9602, nx9604, nx9608, nx9612, 
      gen_24_cmp_mReg_15, nx9624, nx9626, nx9630, nx9634, nx9640, nx9644, 
      nx9650, restartDetection, StartCaptuerCmp_d, nx9664, nx9670, nx2813, 
      nx2823, nx2833, nx2839, nx2853, nx2859, nx2862, nx2871, nx2873, nx2877, 
      nx2887, nx2893, nx2897, nx2903, nx2907, nx2911, nx2917, nx2923, nx2926, 
      nx2931, nx2937, nx2941, nx2947, nx2951, nx2955, nx2961, nx2967, nx2970, 
      nx2975, nx2981, nx2985, nx2991, nx2995, nx2999, nx3005, nx3011, nx3014, 
      nx3019, nx3025, nx3029, nx3035, nx3039, nx3043, nx3049, nx3055, nx3058, 
      nx3063, nx3069, nx3073, nx3079, nx3083, nx3087, nx3093, nx3099, nx3103, 
      nx3107, nx3115, nx3117, nx3121, nx3132, nx3139, nx3143, nx3149, nx3155, 
      nx3158, nx3163, nx3169, nx3173, nx3179, nx3183, nx3187, nx3193, nx3199, 
      nx3202, nx3207, nx3213, nx3217, nx3223, nx3227, nx3231, nx3237, nx3243, 
      nx3246, nx3251, nx3257, nx3261, nx3267, nx3271, nx3275, nx3281, nx3287, 
      nx3290, nx3295, nx3301, nx3305, nx3311, nx3315, nx3319, nx3325, nx3331, 
      nx3334, nx3339, nx3347, nx3353, nx3356, nx3363, nx3365, nx3369, nx3380, 
      nx3387, nx3391, nx3397, nx3401, nx3405, nx3411, nx3415, nx3419, nx3423, 
      nx3429, nx3433, nx3437, nx3443, nx3446, nx3453, nx3459, nx3463, nx3469, 
      nx3475, nx3479, nx3484, nx3488, nx3491, nx3497, nx3503, nx3507, nx3513, 
      nx3517, nx3521, nx3527, nx3533, nx3537, nx3543, nx3547, nx3551, nx3557, 
      nx3563, nx3566, nx3571, nx3577, nx3581, nx3587, nx3593, nx3599, nx3603, 
      nx3611, nx3613, nx3617, nx3629, nx3633, nx3637, nx3643, nx3647, nx3651, 
      nx3655, nx3661, nx3665, nx3669, nx3675, nx3678, nx3685, nx3691, nx3695, 
      nx3699, nx3705, nx3709, nx3713, nx3719, nx3722, nx3729, nx3735, nx3739, 
      nx3743, nx3749, nx3753, nx3757, nx3763, nx3766, nx3773, nx3779, nx3783, 
      nx3787, nx3793, nx3797, nx3801, nx3807, nx3810, nx3817, nx3823, nx3827, 
      nx3831, nx3839, nx3845, nx3849, nx3857, nx3859, nx3863, nx3873, nx3877, 
      nx3881, nx3887, nx3893, nx3897, nx3902, nx3907, nx3911, nx3915, nx3921, 
      nx3925, nx3930, nx3935, nx3939, nx3945, nx3951, nx3954, nx3961, nx3967, 
      nx3971, nx3975, nx3981, nx3985, nx3989, nx3995, nx3998, nx4005, nx4011, 
      nx4015, nx4019, nx4025, nx4029, nx4033, nx4039, nx4042, nx4049, nx4055, 
      nx4059, nx4063, nx4069, nx4073, nx4077, nx4084, nx4089, nx4093, nx4101, 
      nx4103, nx4106, nx4119, nx4125, nx4128, nx4133, nx4139, nx4143, nx4149, 
      nx4153, nx4157, nx4163, nx4169, nx4172, nx4177, nx4183, nx4187, nx4193, 
      nx4197, nx4201, nx4207, nx4213, nx4216, nx4221, nx4227, nx4231, nx4237, 
      nx4241, nx4245, nx4251, nx4256, nx4259, nx4263, nx4269, nx4273, nx4279, 
      nx4285, nx4288, nx4293, nx4299, nx4303, nx4309, nx4315, nx4318, nx4325, 
      nx4331, nx4337, nx4340, nx4349, nx4351, nx4355, nx4365, nx4371, nx4375, 
      nx4381, nx4385, nx4389, nx4395, nx4401, nx4404, nx4409, nx4415, nx4419, 
      nx4425, nx4429, nx4433, nx4439, nx4445, nx4448, nx4453, nx4459, nx4463, 
      nx4469, nx4473, nx4477, nx4483, nx4489, nx4492, nx4497, nx4503, nx4507, 
      nx4513, nx4517, nx4521, nx4527, nx4533, nx4536, nx4541, nx4547, nx4551, 
      nx4557, nx4561, nx4565, nx4571, nx4579, nx4583, nx4587, nx4595, nx4597, 
      nx4601, nx4613, nx4617, nx4621, nx4627, nx4633, nx4637, nx4642, nx4646, 
      nx4649, nx4655, nx4661, nx4665, nx4671, nx4675, nx4679, nx4685, nx4691, 
      nx4695, nx4701, nx4705, nx4709, nx4715, nx4721, nx4724, nx4729, nx4735, 
      nx4739, nx4745, nx4749, nx4753, nx4759, nx4765, nx4768, nx4773, nx4779, 
      nx4783, nx4789, nx4793, nx4797, nx4803, nx4809, nx4812, nx4817, nx4825, 
      nx4831, nx4834, nx4841, nx4843, nx4847, nx4858, nx4865, nx4869, nx4875, 
      nx4879, nx4883, nx4889, nx4893, nx4897, nx4901, nx4907, nx4911, nx4915, 
      nx4921, nx4924, nx4931, nx4937, nx4941, nx4945, nx4951, nx4955, nx4959, 
      nx4965, nx4968, nx4975, nx4981, nx4985, nx4989, nx4995, nx4999, nx5003, 
      nx5009, nx5013, nx5019, nx5025, nx5028, nx5032, nx5037, nx5041, nx5047, 
      nx5053, nx5057, nx5061, nx5069, nx5073, nx5077, nx5085, nx5087, nx5090, 
      nx5103, nx5109, nx5112, nx5119, nx5125, nx5129, nx5133, nx5139, nx5143, 
      nx5147, nx5153, nx5156, nx5163, nx5169, nx5173, nx5177, nx5183, nx5187, 
      nx5191, nx5197, nx5200, nx5207, nx5213, nx5217, nx5221, nx5227, nx5231, 
      nx5235, nx5241, nx5244, nx5251, nx5257, nx5261, nx5265, nx5271, nx5275, 
      nx5279, nx5285, nx5288, nx5295, nx5301, nx5305, nx5309, nx5317, nx5323, 
      nx5327, nx5335, nx5337, nx5341, nx5352, nx5357, nx5361, nx5367, nx5373, 
      nx5376, nx5383, nx5389, nx5393, nx5399, nx5405, nx5409, nx5414, nx5418, 
      nx5421, nx5427, nx5433, nx5437, nx5443, nx5447, nx5451, nx5457, nx5463, 
      nx5467, nx5473, nx5477, nx5481, nx5487, nx5493, nx5496, nx5501, nx5507, 
      nx5511, nx5517, nx5521, nx5525, nx5531, nx5537, nx5540, nx5545, nx5551, 
      nx5555, nx5561, nx5567, nx5573, nx5577, nx5585, nx5587, nx5591, nx5603, 
      nx5607, nx5611, nx5617, nx5621, nx5625, nx5629, nx5635, nx5639, nx5643, 
      nx5649, nx5652, nx5659, nx5665, nx5669, nx5673, nx5679, nx5683, nx5687, 
      nx5693, nx5696, nx5703, nx5709, nx5713, nx5717, nx5723, nx5727, nx5731, 
      nx5737, nx5740, nx5747, nx5753, nx5757, nx5761, nx5767, nx5771, nx5775, 
      nx5781, nx5785, nx5791, nx5797, nx5800, nx5804, nx5811, nx5817, nx5821, 
      nx5829, nx5831, nx5834, nx5847, nx5853, nx5857, nx5861, nx5867, nx5871, 
      nx5875, nx5881, nx5884, nx5891, nx5897, nx5901, nx5905, nx5911, nx5915, 
      nx5919, nx5925, nx5928, nx5935, nx5941, nx5945, nx5949, nx5955, nx5959, 
      nx5963, nx5969, nx5972, nx5979, nx5985, nx5989, nx5993, nx5999, nx6003, 
      nx6007, nx6013, nx6016, nx6023, nx6029, nx6033, nx6037, nx6043, nx6047, 
      nx6051, nx6058, nx6063, nx6067, nx6075, nx6077, nx6080, nx6093, nx6099, 
      nx6102, nx6107, nx6113, nx6117, nx6123, nx6127, nx6131, nx6137, nx6143, 
      nx6146, nx6151, nx6157, nx6161, nx6167, nx6171, nx6175, nx6181, nx6186, 
      nx6189, nx6193, nx6199, nx6203, nx6209, nx6215, nx6218, nx6223, nx6229, 
      nx6233, nx6239, nx6245, nx6248, nx6255, nx6261, nx6265, nx6269, nx6275, 
      nx6279, nx6283, nx6289, nx6292, nx6299, nx6305, nx6311, nx6314, nx6323, 
      nx6325, nx6329, nx6339, nx6345, nx6349, nx6355, nx6359, nx6363, nx6369, 
      nx6375, nx6378, nx6383, nx6389, nx6393, nx6399, nx6403, nx6407, nx6413, 
      nx6419, nx6422, nx6427, nx6433, nx6437, nx6443, nx6447, nx6451, nx6457, 
      nx6463, nx6466, nx6471, nx6477, nx6481, nx6487, nx6491, nx6495, nx6501, 
      nx6507, nx6510, nx6515, nx6521, nx6525, nx6531, nx6535, nx6539, nx6545, 
      nx6553, nx6557, nx6561, nx6569, nx6571, nx6574, nx6585, nx6591, nx6595, 
      nx6601, nx6605, nx6609, nx6615, nx6621, nx6625, nx6631, nx6635, nx6639, 
      nx6645, nx6651, nx6654, nx6659, nx6665, nx6669, nx6675, nx6679, nx6683, 
      nx6689, nx6695, nx6698, nx6703, nx6709, nx6713, nx6719, nx6723, nx6727, 
      nx6733, nx6739, nx6742, nx6747, nx6753, nx6757, nx6763, nx6767, nx6771, 
      nx6777, nx6783, nx6786, nx6791, nx6799, nx6805, nx6808, nx6815, nx6817, 
      nx6821, nx6832, nx6839, nx6843, nx6849, nx6853, nx6857, nx6863, nx6867, 
      nx6871, nx6875, nx6881, nx6885, nx6889, nx6895, nx6898, nx6905, nx6911, 
      nx6915, nx6919, nx6925, nx6929, nx6933, nx6939, nx6943, nx6949, nx6955, 
      nx6958, nx6962, nx6967, nx6971, nx6977, nx6983, nx6987, nx6991, nx6997, 
      nx7001, nx7007, nx7011, nx7015, nx7019, nx7025, nx7029, nx7033, nx7040, 
      nx7045, nx7049, nx7057, nx7059, nx7062, nx7075, nx7081, nx7084, nx7089, 
      nx7095, nx7099, nx7105, nx7109, nx7113, nx7119, nx7125, nx7128, nx7133, 
      nx7139, nx7143, nx7149, nx7153, nx7157, nx7163, nx7169, nx7172, nx7177, 
      nx7183, nx7187, nx7193, nx7197, nx7201, nx7207, nx7213, nx7216, nx7221, 
      nx7227, nx7231, nx7237, nx7241, nx7245, nx7251, nx7257, nx7260, nx7265, 
      nx7271, nx7275, nx7281, nx7287, nx7293, nx7297, nx7305, nx7307, nx7311, 
      nx7323, nx7329, nx7333, nx7339, nx7344, nx7347, nx7351, nx7357, nx7361, 
      nx7367, nx7373, nx7376, nx7381, nx7387, nx7391, nx7397, nx7403, nx7406, 
      nx7413, nx7419, nx7423, nx7427, nx7433, nx7437, nx7441, nx7447, nx7450, 
      nx7457, nx7463, nx7467, nx7471, nx7477, nx7481, nx7485, nx7491, nx7494, 
      nx7501, nx7507, nx7511, nx7515, nx7521, nx7525, nx7529, nx7536, nx7541, 
      nx7545, nx7553, nx7555, nx7558, nx7571, nx7577, nx7580, nx7585, nx7591, 
      nx7595, nx7601, nx7605, nx7609, nx7615, nx7621, nx7624, nx7629, nx7635, 
      nx7639, nx7645, nx7649, nx7653, nx7659, nx7665, nx7668, nx7673, nx7679, 
      nx7683, nx7689, nx7693, nx7697, nx7703, nx7709, nx7713, nx7719, nx7725, 
      nx7729, nx7733, nx7737, nx7741, nx7747, nx7753, nx7757, nx7762, nx7767, 
      nx7771, nx7775, nx7783, nx7789, nx7792, nx7801, nx7803, nx7807, nx7817, 
      nx7823, nx7827, nx7833, nx7837, nx7841, nx7847, nx7853, nx7856, nx7861, 
      nx7867, nx7871, nx7877, nx7881, nx7885, nx7891, nx7897, nx7900, nx7905, 
      nx7911, nx7915, nx7921, nx7925, nx7929, nx7935, nx7941, nx7944, nx7949, 
      nx7955, nx7959, nx7965, nx7969, nx7973, nx7979, nx7985, nx7988, nx7993, 
      nx7999, nx8003, nx8009, nx8013, nx8017, nx8023, nx8031, nx8035, nx8039, 
      nx8047, nx8049, nx8053, nx8065, nx8069, nx8073, nx8077, nx8083, nx8087, 
      nx8091, nx8097, nx8101, nx8107, nx8113, nx8116, nx8120, nx8125, nx8129, 
      nx8135, nx8141, nx8145, nx8149, nx8155, nx8159, nx8165, nx8169, nx8173, 
      nx8177, nx8183, nx8187, nx8191, nx8197, nx8200, nx8207, nx8213, nx8217, 
      nx8221, nx8227, nx8231, nx8235, nx8241, nx8244, nx8251, nx8257, nx8261, 
      nx8265, nx8273, nx8279, nx8283, nx8291, nx8293, nx8297, nx8308, nx8313, 
      nx8317, nx8323, nx8329, nx8332, nx8339, nx8345, nx8349, nx8353, nx8359, 
      nx8363, nx8367, nx8373, nx8376, nx8383, nx8389, nx8393, nx8397, nx8403, 
      nx8407, nx8411, nx8417, nx8420, nx8427, nx8433, nx8437, nx8441, nx8447, 
      nx8451, nx8455, nx8461, nx8464, nx8471, nx8477, nx8481, nx8487, nx8493, 
      nx8497, nx8502, nx8506, nx8509, nx8515, nx8523, nx8529, nx8533, nx8541, 
      nx8543, nx8547, nx8559, nx8563, nx8567, nx8573, nx8577, nx8581, nx8585, 
      nx8591, nx8595, nx8599, nx8605, nx8608, nx8615, nx8621, nx8625, nx8629, 
      nx8635, nx8639, nx8643, nx8649, nx8652, nx8659, nx8665, nx8669, nx8673, 
      nx8679, nx8683, nx8687, nx8693, nx8696, nx8703, nx8709, nx8713, nx8717, 
      nx8723, nx8727, nx8731, nx8737, nx8740, nx8747, nx8753, nx8757, nx8761, 
      nx8769, nx8775, nx8779, nx8787, nx8789, nx8793, nx8804, nx8809, nx8813, 
      nx8819, nx8825, nx8828, nx8835, nx8841, nx8845, nx8849, nx8855, nx8859, 
      nx8863, nx8869, nx8873, nx8879, nx8885, nx8888, nx8892, nx8897, nx8901, 
      nx8907, nx8913, nx8917, nx8921, nx8927, nx8931, nx8937, nx8941, nx8945, 
      nx8949, nx8955, nx8959, nx8963, nx8969, nx8972, nx8979, nx8985, nx8989, 
      nx8993, nx8999, nx9003, nx9007, nx9014, nx9017, nx9023, nx9027, nx9031, 
      nx9036, nx9039, nx9043, nx9049, nx9053, nx9057, nx9061, nx9065, nx9069, 
      nx9073, nx9077, nx9080, nx9085, nx9089, nx9093, nx9099, nx9102, nx9105, 
      nx9111, nx9115, nx9119, nx9124, nx9127, nx9131, nx9137, nx9141, nx9145, 
      nx9149, nx9153, nx9157, nx9161, nx9165, nx9168, nx9173, nx9177, nx9181, 
      nx9187, nx9190, nx9193, nx9199, nx9203, nx9207, nx9212, nx9215, nx9219, 
      nx9225, nx9229, nx9233, nx9237, nx9241, nx9245, nx9249, nx9253, nx9257, 
      nx9263, nx9267, nx9271, nx9275, nx9278, nx9281, nx9287, nx9291, nx9295, 
      nx9301, nx9305, nx9308, nx9315, nx9319, nx9323, nx9327, nx9333, nx9336, 
      nx9343, nx9353, nx9357, nx9361, nx9365, nx9373, nx9375, nx9377, nx9379, 
      nx9381, nx9389, nx9391, nx9393, nx9395, nx9397, nx9399, nx9401, nx9403, 
      nx9405, nx9407, nx9409, nx9411, nx9413, nx9415, nx9417, nx9419, nx9421, 
      nx9423, nx9425, nx9427, nx9429, nx9431, nx9433, nx9435, nx9437, nx9439, 
      nx9441, nx9443, nx9445, nx9447, nx9449, nx9451, nx9453, nx9455, nx9457, 
      nx9459, nx9461, nx9463, nx9465, nx9467, nx9469, nx9471, nx9473, nx9475, 
      nx9477, nx9479, nx9481, nx9483, nx9485, nx9487, nx9489, nx9491, nx9493, 
      nx9495, nx9497, nx9499, nx9501, nx9503, nx9505, nx9507, nx9509, nx9511, 
      nx9513, nx9515, nx9517, nx9519, nx9521, nx9523, nx9525, nx9527, nx9529, 
      nx9531, nx9533, nx9535, nx9537, nx9539, nx9541, nx9543, nx9545, nx9547, 
      nx9549, nx9551, nx9553, nx9555, nx9557, nx9559, nx9561, nx9563, nx9565, 
      nx9567, nx9569, nx9571, nx9573, nx9575, nx9577, nx9579, nx9581, nx9583, 
      nx9585, nx9587, nx9589, nx9591, nx9593, nx9595, nx9597, nx9599, nx9601, 
      nx9603, nx9605, nx9607, nx9609, nx9611, nx9613, nx9615, nx9617, nx9619, 
      nx9621, nx9623, nx9625, nx9627, nx9629, nx9631, nx9633, nx9635, nx9637, 
      nx9639, nx9641, nx9643, nx9645, nx9647, nx9649, nx9651, nx9653, nx9655, 
      nx9657, nx9659, nx9661, nx9663, nx9665, nx9667, nx9669, nx9671, nx9673, 
      nx9675, nx9677, nx9679, nx9681, nx9683, nx9685, nx9687, nx9689, nx9691, 
      nx9693, nx9695, nx9697, nx9699, nx9701, nx9703, nx9705, nx9707, nx9709, 
      nx9711, nx9713, nx9715, nx9717, nx9719, nx9721, nx9723, nx9725, nx9727, 
      nx9729, nx9731, nx9733, nx9735, nx9737, nx9739, nx9741, nx9743, nx9745, 
      nx9747, nx9749, nx9751, nx9753, nx9755, nx9757, nx9759, nx9761, nx9763, 
      nx9765, nx9767, nx9769, nx9771, nx9773, nx9775, nx9777, nx9779, nx9781, 
      nx9783, nx9785, nx9787, nx9789, nx9791, nx9793, nx9795, nx9797, nx9799, 
      nx9801, nx9803, nx9805, nx9807, nx9809, nx9811, nx9813, nx9815, nx9817, 
      nx9819, nx9821, nx9823, nx9825, nx9827, nx9829, nx9831, nx9833, nx9835, 
      nx9837, nx9839, nx9841, nx9843, nx9845, nx9847, nx9849, nx9851, nx9853, 
      nx9855, nx9857, nx9859, nx9861, nx9863, nx9865, nx9867, nx9869, nx9871, 
      nx9873, nx9875, nx9877, nx9879, nx9881, nx9883, nx9885, nx9887, nx9889, 
      nx9891, nx9893, nx9895, nx9897, nx9899, nx9901, nx9903, nx9905, nx9907, 
      nx9909, nx9911, nx9913, nx9915, nx9917, nx9919, nx9921, nx9923, nx9925, 
      nx9927, nx9929, nx9931, nx9933, nx9935, nx9937, nx9939, nx9941, nx9943, 
      nx9945, nx9947, nx9949, nx9951, nx9953, nx9955, nx9957, nx9959, nx9961, 
      nx9963, nx9965, nx9967, nx9969, nx9971, nx9973, nx9975, nx9977, nx9979, 
      nx9981, nx9983, nx9985, nx9987, nx9989, nx9991, nx9993, nx9995, nx9997, 
      nx9999, nx10001, nx10003, nx10005, nx10007, nx10009, nx10011, nx10013, 
      nx10015, nx10017, nx10019, nx10021, nx10023, nx10025, nx10027, nx10029, 
      nx10031, nx10033, nx10035, nx10037, nx10039, nx10041, nx10043, nx10045, 
      nx10047, nx10049, nx10051, nx10053, nx10055, nx10057, nx10059, nx10061, 
      nx10063, nx10065, nx10067, nx10069, nx10071, nx10073, nx10075, nx10077, 
      nx10079, nx10081, nx10083, nx10085, nx10087, nx10089, nx10091, nx10093, 
      nx10095, nx10097, nx10099, nx10101, nx10103, nx10105, nx10107, nx10109, 
      nx10111, nx10113, nx10115, nx10117, nx10119, nx10121, nx10123, nx10125, 
      nx10127, nx10129, nx10131, nx10133, nx10135, nx10137, nx10139, nx10141, 
      nx10143, nx10145, nx10147, nx10149, nx10151, nx10153, nx10155, nx10157, 
      nx10159, nx10161, nx10163, nx10165, nx10167, nx10169, nx10171, nx10173, 
      nx10175, nx10177, nx10179, nx10181, nx10183, nx10185, nx10187, nx10189, 
      nx10191, nx10193, nx10195, nx10197, nx10199, nx10201, nx10203, nx10205, 
      nx10207, nx10209, nx10211, nx10213, nx10215, nx10217, nx10219, nx10221, 
      nx10223, nx10225, nx10227, nx10229, nx10231, nx10233, nx10235, nx10237, 
      nx10239, nx10241, nx10243, nx10245, nx10247, nx10249, nx10251, nx10253, 
      nx10255, nx10257, nx10259, nx10261, nx10263, nx10265, nx10267, nx10269, 
      nx10271, nx10273, nx10275, nx10277, nx10279, nx10281, nx10283, nx10285, 
      nx10287, nx10289, nx10291, nx10293, nx10295, nx10297, nx10299, nx10301, 
      nx10303, nx10305, nx10307, nx10309, nx10311, nx10313, nx10315, nx10317, 
      nx10319, nx10321, nx10323, nx10325, nx10327, nx10329, nx10331, nx10333, 
      nx10335, nx10337, nx10339, nx10341, nx10343, nx10345, nx10347, nx10349, 
      nx10351, nx10353, nx10355, nx10357, nx10359, nx10361, nx10363, nx10365, 
      nx10367, nx10369, nx10371, nx10373, nx10375, nx10377, nx10379, nx10381, 
      nx10383, nx10385, nx10387, nx10389, nx10391, nx10393, nx10395, nx10397, 
      nx10399, nx10401, nx10403, nx10405, nx10407, nx10409, nx10411, nx10413, 
      nx10415, nx10417, nx10419, nx10421, nx10423, nx10425, nx10427, nx10429, 
      nx10431, nx10433, nx10435, nx10437, nx10439, nx10441, nx10443, nx10445, 
      nx10447, nx10449, nx10451, nx10453, nx10455, nx10457, nx10459, nx10461, 
      nx10463, nx10465, nx10467, nx10469, nx10471, nx10473, nx10475, nx10477, 
      nx10479, nx10481, nx10483, nx10485, nx10487, nx10489, nx10491, nx10493, 
      nx10495, nx10497, nx10499, nx10501, nx10503, nx10505, nx10507, nx10509, 
      nx10511, nx10513, nx10515, nx10517, nx10519, nx10521, nx10523, nx10525, 
      nx10527, nx10529, nx10531, nx10533, nx10535, nx10537, nx10539, nx10541, 
      nx10543, nx10545, nx10547, nx10549, nx10551, nx10553, nx10555, nx10557, 
      nx10559, nx10561, nx10563, nx10565, nx10567, nx10569, nx10571, nx10573, 
      nx10575, nx10577, nx10579, nx10581, nx10583, nx10585, nx10587, nx10589, 
      nx10591, nx10593, nx10595, nx10597, nx10599, nx10601, nx10603, nx10605, 
      nx10607, nx10609, nx10611, nx10613, nx10615, nx10617, nx10619, nx10621, 
      nx10623, nx10625, nx10627, nx10629, nx10631, nx10633, nx10635, nx10637, 
      nx10639, nx10641, nx10643, nx10645, nx10647, nx10649, nx10651, nx10653, 
      nx10655, nx10657, nx10659, nx10661, nx10663, nx10665, nx10667, nx10669, 
      nx10671, nx10673, nx10675, nx10677, nx10679, nx10681, nx10683, nx10685, 
      nx10687, nx10689, nx10691, nx10693, nx10695, nx10697, nx10699, nx10701, 
      nx10703, nx10705, nx10707, nx10709, nx10711, nx10713, nx10715, nx10717, 
      nx10719, nx10721, nx10723, nx10725, nx10727, nx10729, nx10731, nx10733, 
      nx10735, nx10737, nx10739, nx10741, nx10743, nx10745, nx10747, nx10749, 
      nx10751, nx10753, nx10755, nx10757, nx10759, nx10761, nx10763, nx10765, 
      nx10767, nx10769, nx10771, nx10773, nx10775, nx10777, nx10779, nx10781, 
      nx10783, nx10785, nx10787, nx10789, nx10791, nx10793, nx10795, nx10797, 
      nx10799, nx10801, nx10803, nx10805, nx10807, nx10809, nx10811, nx10813, 
      nx10815, nx10817, nx10819, nx10821, nx10823, nx10825, nx10827, nx10829, 
      nx10831, nx10833, nx10835, nx10837, nx10839, nx10841, nx10843, nx10845, 
      nx10847, nx10849, nx10851, nx10853, nx10855, nx10857, nx10859, nx10861, 
      nx10863, nx10865, nx10867, nx10869, nx10871, nx10873, nx10875, nx10877, 
      nx10879, nx10881, nx10883, nx10885, nx10887, nx10889, nx10891, nx10893, 
      nx10895, nx10897, nx10899, nx10901, nx10903, nx10905, nx10907, nx10909, 
      nx10911, nx10913, nx10915, nx10917, nx10919, nx10921, nx10923, nx10925, 
      nx10927, nx10929, nx10931, nx10933, nx10935, nx10937, nx10939, nx10941, 
      nx10943, nx10945, nx10947, nx10949, nx10951, nx10953, nx10955, nx10957, 
      nx10959, nx10961, nx10963, nx10965, nx10967, nx10969, nx10971, nx10973, 
      nx10975, nx10977, nx10979, nx10981, nx10983, nx10985, nx10987, nx10989, 
      nx10991, nx10993, nx10995, nx10997, nx10999, nx11001, nx11003, nx11005, 
      nx11007, nx11009, nx11011, nx11013, nx11015, nx11017, nx11019, nx11021, 
      nx11023, nx11025, nx11027, nx11029, nx11031, nx11033, nx11035, nx11037, 
      nx11039, nx11041, nx11043, nx11045, nx11047, nx11049, nx11051, nx11053, 
      nx11055, nx11057, nx11059, nx11061, nx11063, nx11065, nx11067, nx11069, 
      nx11071, nx11073, nx11075, nx11077, nx11079, nx11081, nx11083, nx11085, 
      nx11087, nx11089, nx11091, nx11093, nx11095, nx11097, nx11099, nx11101, 
      nx11103, nx11105, nx11107, nx11109, nx11111, nx11113, nx11115, nx11117, 
      nx11119, nx11121, nx11123, nx11125, nx11127, nx11129, nx11131, nx11133, 
      nx11135, nx11137, nx11139, nx11141, nx11143, nx11145, nx11147, nx11157, 
      nx11159, nx11161, nx11163, nx11165, nx11167, nx11169, nx11171, nx11173, 
      nx11175, nx11177, nx11179, nx11181, nx11183, nx11185, nx11187, nx11189, 
      nx11191, nx11197, nx11199, nx11201, nx11203: std_logic ;
   
   signal DANGLING : std_logic_vector (124 downto 0 );

begin
   gen_24_cmp_pRegCmp : Reg_33 port map ( D(32)=>working, D(31)=>working, 
      D(30)=>gen_24_cmp_pBs_30, D(29)=>gen_24_cmp_pBs_29, D(28)=>
      gen_24_cmp_pBs_28, D(27)=>gen_24_cmp_pBs_27, D(26)=>gen_24_cmp_pBs_26, 
      D(25)=>gen_24_cmp_pBs_25, D(24)=>gen_24_cmp_pBs_24, D(23)=>
      gen_24_cmp_pBs_23, D(22)=>outputs_24_15, D(21)=>outputs_24_14, D(20)=>
      outputs_24_13, D(19)=>outputs_24_12, D(18)=>outputs_24_11, D(17)=>
      outputs_24_10, D(16)=>outputs_24_9, D(15)=>outputs_24_8, D(14)=>
      outputs_24_7, D(13)=>outputs_24_6, D(12)=>outputs_24_5, D(11)=>
      outputs_24_4, D(10)=>outputs_24_3, D(9)=>outputs_24_2, D(8)=>
      outputs_24_1, D(7)=>outputs_24_0, D(6)=>gen_24_cmp_pMux_8, D(5)=>
      gen_24_cmp_pMux_7, D(4)=>gen_24_cmp_pMux_6, D(3)=>gen_24_cmp_pMux_5, 
      D(2)=>gen_24_cmp_pMux_4, D(1)=>gen_24_cmp_pMux_3, D(0)=>nx9399, en=>
      nx11159, clk=>nx9391, rst=>rst, Q(32)=>DANGLING(0), Q(31)=>DANGLING(1), 
      Q(30)=>gen_24_cmp_pReg_30, Q(29)=>gen_24_cmp_pReg_29, Q(28)=>
      gen_24_cmp_pReg_28, Q(27)=>gen_24_cmp_pReg_27, Q(26)=>
      gen_24_cmp_pReg_26, Q(25)=>gen_24_cmp_pReg_25, Q(24)=>
      gen_24_cmp_pReg_24, Q(23)=>gen_24_cmp_pReg_23, Q(22)=>
      gen_24_cmp_pReg_22, Q(21)=>gen_24_cmp_pReg_21, Q(20)=>
      gen_24_cmp_pReg_20, Q(19)=>gen_24_cmp_pReg_19, Q(18)=>
      gen_24_cmp_pReg_18, Q(17)=>gen_24_cmp_pReg_17, Q(16)=>
      gen_24_cmp_pReg_16, Q(15)=>gen_24_cmp_pReg_15, Q(14)=>
      gen_24_cmp_pReg_14, Q(13)=>gen_24_cmp_pReg_13, Q(12)=>
      gen_24_cmp_pReg_12, Q(11)=>gen_24_cmp_pReg_11, Q(10)=>
      gen_24_cmp_pReg_10, Q(9)=>gen_24_cmp_pReg_9, Q(8)=>gen_24_cmp_pReg_8, 
      Q(7)=>gen_24_cmp_pReg_7, Q(6)=>gen_24_cmp_pReg_6, Q(5)=>
      gen_24_cmp_pReg_5, Q(4)=>gen_24_cmp_pReg_4, Q(3)=>gen_24_cmp_pReg_3, 
      Q(2)=>gen_24_cmp_pReg_2, Q(1)=>gen_24_cmp_pReg_1, Q(0)=>
      gen_24_cmp_pReg_0);
   gen_24_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>working, a(31)=>
      working, a(30)=>gen_24_cmp_pReg_30, a(29)=>gen_24_cmp_pReg_29, a(28)=>
      gen_24_cmp_pReg_28, a(27)=>gen_24_cmp_pReg_27, a(26)=>
      gen_24_cmp_pReg_26, a(25)=>gen_24_cmp_pReg_25, a(24)=>
      gen_24_cmp_pReg_24, a(23)=>gen_24_cmp_pReg_23, a(22)=>
      gen_24_cmp_pReg_22, a(21)=>gen_24_cmp_pReg_21, a(20)=>
      gen_24_cmp_pReg_20, a(19)=>gen_24_cmp_pReg_19, a(18)=>
      gen_24_cmp_pReg_18, a(17)=>gen_24_cmp_pReg_17, a(16)=>
      gen_24_cmp_pReg_16, a(15)=>gen_24_cmp_pReg_15, a(14)=>
      gen_24_cmp_pReg_14, a(13)=>gen_24_cmp_pReg_13, a(12)=>
      gen_24_cmp_pReg_12, a(11)=>gen_24_cmp_pReg_11, a(10)=>
      gen_24_cmp_pReg_10, a(9)=>gen_24_cmp_pReg_9, a(8)=>gen_24_cmp_pReg_8, 
      a(7)=>gen_24_cmp_pReg_7, a(6)=>gen_24_cmp_pReg_6, a(5)=>
      gen_24_cmp_pReg_5, a(4)=>gen_24_cmp_pReg_4, a(3)=>gen_24_cmp_pReg_3, 
      a(2)=>gen_24_cmp_pReg_2, a(1)=>gen_24_cmp_pReg_1, a(0)=>
      gen_24_cmp_pReg_0, b(32)=>working, b(31)=>working, b(30)=>working, 
      b(29)=>working, b(28)=>working, b(27)=>working, b(26)=>working, b(25)
      =>working, b(24)=>working, b(23)=>working, b(22)=>working, b(21)=>
      working, b(20)=>working, b(19)=>working, b(18)=>working, b(17)=>
      working, b(16)=>working, b(15)=>working, b(14)=>working, b(13)=>
      working, b(12)=>working, b(11)=>working, b(10)=>working, b(9)=>working, 
      b(8)=>filter_24_7, b(7)=>filter_24_6, b(6)=>filter_24_5, b(5)=>
      filter_24_4, b(4)=>filter_24_3, b(3)=>filter_24_2, b(2)=>filter_24_1, 
      b(1)=>filter_24_0, b(0)=>working, sel=>nx11173, f(32)=>DANGLING(2), 
      f(31)=>DANGLING(3), f(30)=>gen_24_cmp_pMux_30, f(29)=>
      gen_24_cmp_pMux_29, f(28)=>gen_24_cmp_pMux_28, f(27)=>
      gen_24_cmp_pMux_27, f(26)=>gen_24_cmp_pMux_26, f(25)=>
      gen_24_cmp_pMux_25, f(24)=>gen_24_cmp_pMux_24, f(23)=>
      gen_24_cmp_pMux_23, f(22)=>gen_24_cmp_pMux_22, f(21)=>
      gen_24_cmp_pMux_21, f(20)=>gen_24_cmp_pMux_20, f(19)=>
      gen_24_cmp_pMux_19, f(18)=>gen_24_cmp_pMux_18, f(17)=>
      gen_24_cmp_pMux_17, f(16)=>gen_24_cmp_pMux_16, f(15)=>
      gen_24_cmp_pMux_15, f(14)=>gen_24_cmp_pMux_14, f(13)=>
      gen_24_cmp_pMux_13, f(12)=>gen_24_cmp_pMux_12, f(11)=>
      gen_24_cmp_pMux_11, f(10)=>gen_24_cmp_pMux_10, f(9)=>gen_24_cmp_pMux_9, 
      f(8)=>gen_24_cmp_pMux_8, f(7)=>gen_24_cmp_pMux_7, f(6)=>
      gen_24_cmp_pMux_6, f(5)=>gen_24_cmp_pMux_5, f(4)=>gen_24_cmp_pMux_4, 
      f(3)=>gen_24_cmp_pMux_3, f(2)=>gen_24_cmp_pMux_2, f(1)=>
      gen_24_cmp_pMux_1, f(0)=>gen_24_cmp_pMux_0);
   gen_24_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>working, a(22)
      =>working, a(21)=>gen_24_cmp_pMux_30, a(20)=>gen_24_cmp_pMux_29, a(19)
      =>gen_24_cmp_pMux_28, a(18)=>gen_24_cmp_pMux_27, a(17)=>
      gen_24_cmp_pMux_26, a(16)=>gen_24_cmp_pMux_25, a(15)=>
      gen_24_cmp_pMux_24, a(14)=>gen_24_cmp_pMux_23, a(13)=>
      gen_24_cmp_pMux_22, a(12)=>gen_24_cmp_pMux_21, a(11)=>
      gen_24_cmp_pMux_20, a(10)=>gen_24_cmp_pMux_19, a(9)=>
      gen_24_cmp_pMux_18, a(8)=>gen_24_cmp_pMux_17, a(7)=>gen_24_cmp_pMux_16, 
      a(6)=>gen_24_cmp_pMux_15, a(5)=>gen_24_cmp_pMux_14, a(4)=>
      gen_24_cmp_pMux_13, a(3)=>gen_24_cmp_pMux_12, a(2)=>gen_24_cmp_pMux_11, 
      a(1)=>gen_24_cmp_pMux_10, a(0)=>gen_24_cmp_pMux_9, b(23)=>nx9703, 
      b(22)=>nx9703, b(21)=>nx9701, b(20)=>nx9709, b(19)=>nx9707, b(18)=>
      nx9705, b(17)=>nx9703, b(16)=>nx9701, b(15)=>gen_24_cmp_BSCmp_op2_15, 
      b(14)=>gen_24_cmp_BSCmp_op2_14, b(13)=>gen_24_cmp_BSCmp_op2_13, b(12)
      =>gen_24_cmp_BSCmp_op2_12, b(11)=>gen_24_cmp_BSCmp_op2_11, b(10)=>
      gen_24_cmp_BSCmp_op2_10, b(9)=>gen_24_cmp_BSCmp_op2_9, b(8)=>
      gen_24_cmp_BSCmp_op2_8, b(7)=>gen_24_cmp_BSCmp_op2_7, b(6)=>
      gen_24_cmp_BSCmp_op2_6, b(5)=>gen_24_cmp_BSCmp_op2_5, b(4)=>
      gen_24_cmp_BSCmp_op2_4, b(3)=>gen_24_cmp_BSCmp_op2_3, b(2)=>
      gen_24_cmp_BSCmp_op2_2, b(1)=>gen_24_cmp_BSCmp_op2_1, b(0)=>
      gen_24_cmp_BSCmp_op2_0, carryIn=>gen_24_cmp_BSCmp_carryIn, sum(23)=>
      gen_24_cmp_pBs_30, sum(22)=>gen_24_cmp_pBs_29, sum(21)=>
      gen_24_cmp_pBs_28, sum(20)=>gen_24_cmp_pBs_27, sum(19)=>
      gen_24_cmp_pBs_26, sum(18)=>gen_24_cmp_pBs_25, sum(17)=>
      gen_24_cmp_pBs_24, sum(16)=>gen_24_cmp_pBs_23, sum(15)=>outputs_24_15, 
      sum(14)=>outputs_24_14, sum(13)=>outputs_24_13, sum(12)=>outputs_24_12, 
      sum(11)=>outputs_24_11, sum(10)=>outputs_24_10, sum(9)=>outputs_24_9, 
      sum(8)=>outputs_24_8, sum(7)=>outputs_24_7, sum(6)=>outputs_24_6, 
      sum(5)=>outputs_24_5, sum(4)=>outputs_24_4, sum(3)=>outputs_24_3, 
      sum(2)=>outputs_24_2, sum(1)=>outputs_24_1, sum(0)=>outputs_24_0, 
      carryOut=>DANGLING(4));
   gen_23_cmp_pRegCmp : Reg_33 port map ( D(32)=>working, D(31)=>working, 
      D(30)=>gen_23_cmp_pBs_30, D(29)=>gen_23_cmp_pBs_29, D(28)=>
      gen_23_cmp_pBs_28, D(27)=>gen_23_cmp_pBs_27, D(26)=>gen_23_cmp_pBs_26, 
      D(25)=>gen_23_cmp_pBs_25, D(24)=>gen_23_cmp_pBs_24, D(23)=>
      gen_23_cmp_pBs_23, D(22)=>outputs_23_15, D(21)=>outputs_23_14, D(20)=>
      outputs_23_13, D(19)=>outputs_23_12, D(18)=>outputs_23_11, D(17)=>
      outputs_23_10, D(16)=>outputs_23_9, D(15)=>outputs_23_8, D(14)=>
      outputs_23_7, D(13)=>outputs_23_6, D(12)=>outputs_23_5, D(11)=>
      outputs_23_4, D(10)=>outputs_23_3, D(9)=>outputs_23_2, D(8)=>
      outputs_23_1, D(7)=>outputs_23_0, D(6)=>gen_23_cmp_pMux_8, D(5)=>
      gen_23_cmp_pMux_7, D(4)=>gen_23_cmp_pMux_6, D(3)=>gen_23_cmp_pMux_5, 
      D(2)=>gen_23_cmp_pMux_4, D(1)=>gen_23_cmp_pMux_3, D(0)=>nx9411, en=>
      nx11159, clk=>nx9391, rst=>rst, Q(32)=>DANGLING(5), Q(31)=>DANGLING(6), 
      Q(30)=>gen_23_cmp_pReg_30, Q(29)=>gen_23_cmp_pReg_29, Q(28)=>
      gen_23_cmp_pReg_28, Q(27)=>gen_23_cmp_pReg_27, Q(26)=>
      gen_23_cmp_pReg_26, Q(25)=>gen_23_cmp_pReg_25, Q(24)=>
      gen_23_cmp_pReg_24, Q(23)=>gen_23_cmp_pReg_23, Q(22)=>
      gen_23_cmp_pReg_22, Q(21)=>gen_23_cmp_pReg_21, Q(20)=>
      gen_23_cmp_pReg_20, Q(19)=>gen_23_cmp_pReg_19, Q(18)=>
      gen_23_cmp_pReg_18, Q(17)=>gen_23_cmp_pReg_17, Q(16)=>
      gen_23_cmp_pReg_16, Q(15)=>gen_23_cmp_pReg_15, Q(14)=>
      gen_23_cmp_pReg_14, Q(13)=>gen_23_cmp_pReg_13, Q(12)=>
      gen_23_cmp_pReg_12, Q(11)=>gen_23_cmp_pReg_11, Q(10)=>
      gen_23_cmp_pReg_10, Q(9)=>gen_23_cmp_pReg_9, Q(8)=>gen_23_cmp_pReg_8, 
      Q(7)=>gen_23_cmp_pReg_7, Q(6)=>gen_23_cmp_pReg_6, Q(5)=>
      gen_23_cmp_pReg_5, Q(4)=>gen_23_cmp_pReg_4, Q(3)=>gen_23_cmp_pReg_3, 
      Q(2)=>gen_23_cmp_pReg_2, Q(1)=>gen_23_cmp_pReg_1, Q(0)=>
      gen_23_cmp_pReg_0);
   gen_23_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>working, a(31)=>
      working, a(30)=>gen_23_cmp_pReg_30, a(29)=>gen_23_cmp_pReg_29, a(28)=>
      gen_23_cmp_pReg_28, a(27)=>gen_23_cmp_pReg_27, a(26)=>
      gen_23_cmp_pReg_26, a(25)=>gen_23_cmp_pReg_25, a(24)=>
      gen_23_cmp_pReg_24, a(23)=>gen_23_cmp_pReg_23, a(22)=>
      gen_23_cmp_pReg_22, a(21)=>gen_23_cmp_pReg_21, a(20)=>
      gen_23_cmp_pReg_20, a(19)=>gen_23_cmp_pReg_19, a(18)=>
      gen_23_cmp_pReg_18, a(17)=>gen_23_cmp_pReg_17, a(16)=>
      gen_23_cmp_pReg_16, a(15)=>gen_23_cmp_pReg_15, a(14)=>
      gen_23_cmp_pReg_14, a(13)=>gen_23_cmp_pReg_13, a(12)=>
      gen_23_cmp_pReg_12, a(11)=>gen_23_cmp_pReg_11, a(10)=>
      gen_23_cmp_pReg_10, a(9)=>gen_23_cmp_pReg_9, a(8)=>gen_23_cmp_pReg_8, 
      a(7)=>gen_23_cmp_pReg_7, a(6)=>gen_23_cmp_pReg_6, a(5)=>
      gen_23_cmp_pReg_5, a(4)=>gen_23_cmp_pReg_4, a(3)=>gen_23_cmp_pReg_3, 
      a(2)=>gen_23_cmp_pReg_2, a(1)=>gen_23_cmp_pReg_1, a(0)=>
      gen_23_cmp_pReg_0, b(32)=>working, b(31)=>working, b(30)=>working, 
      b(29)=>working, b(28)=>working, b(27)=>working, b(26)=>working, b(25)
      =>working, b(24)=>working, b(23)=>working, b(22)=>working, b(21)=>
      working, b(20)=>working, b(19)=>working, b(18)=>working, b(17)=>
      working, b(16)=>working, b(15)=>working, b(14)=>working, b(13)=>
      working, b(12)=>working, b(11)=>working, b(10)=>working, b(9)=>working, 
      b(8)=>filter_23_7, b(7)=>filter_23_6, b(6)=>filter_23_5, b(5)=>
      filter_23_4, b(4)=>filter_23_3, b(3)=>filter_23_2, b(2)=>filter_23_1, 
      b(1)=>filter_23_0, b(0)=>working, sel=>nx11173, f(32)=>DANGLING(7), 
      f(31)=>DANGLING(8), f(30)=>gen_23_cmp_pMux_30, f(29)=>
      gen_23_cmp_pMux_29, f(28)=>gen_23_cmp_pMux_28, f(27)=>
      gen_23_cmp_pMux_27, f(26)=>gen_23_cmp_pMux_26, f(25)=>
      gen_23_cmp_pMux_25, f(24)=>gen_23_cmp_pMux_24, f(23)=>
      gen_23_cmp_pMux_23, f(22)=>gen_23_cmp_pMux_22, f(21)=>
      gen_23_cmp_pMux_21, f(20)=>gen_23_cmp_pMux_20, f(19)=>
      gen_23_cmp_pMux_19, f(18)=>gen_23_cmp_pMux_18, f(17)=>
      gen_23_cmp_pMux_17, f(16)=>gen_23_cmp_pMux_16, f(15)=>
      gen_23_cmp_pMux_15, f(14)=>gen_23_cmp_pMux_14, f(13)=>
      gen_23_cmp_pMux_13, f(12)=>gen_23_cmp_pMux_12, f(11)=>
      gen_23_cmp_pMux_11, f(10)=>gen_23_cmp_pMux_10, f(9)=>gen_23_cmp_pMux_9, 
      f(8)=>gen_23_cmp_pMux_8, f(7)=>gen_23_cmp_pMux_7, f(6)=>
      gen_23_cmp_pMux_6, f(5)=>gen_23_cmp_pMux_5, f(4)=>gen_23_cmp_pMux_4, 
      f(3)=>gen_23_cmp_pMux_3, f(2)=>gen_23_cmp_pMux_2, f(1)=>
      gen_23_cmp_pMux_1, f(0)=>gen_23_cmp_pMux_0);
   gen_23_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>working, a(22)
      =>working, a(21)=>gen_23_cmp_pMux_30, a(20)=>gen_23_cmp_pMux_29, a(19)
      =>gen_23_cmp_pMux_28, a(18)=>gen_23_cmp_pMux_27, a(17)=>
      gen_23_cmp_pMux_26, a(16)=>gen_23_cmp_pMux_25, a(15)=>
      gen_23_cmp_pMux_24, a(14)=>gen_23_cmp_pMux_23, a(13)=>
      gen_23_cmp_pMux_22, a(12)=>gen_23_cmp_pMux_21, a(11)=>
      gen_23_cmp_pMux_20, a(10)=>gen_23_cmp_pMux_19, a(9)=>
      gen_23_cmp_pMux_18, a(8)=>gen_23_cmp_pMux_17, a(7)=>gen_23_cmp_pMux_16, 
      a(6)=>gen_23_cmp_pMux_15, a(5)=>gen_23_cmp_pMux_14, a(4)=>
      gen_23_cmp_pMux_13, a(3)=>gen_23_cmp_pMux_12, a(2)=>gen_23_cmp_pMux_11, 
      a(1)=>gen_23_cmp_pMux_10, a(0)=>gen_23_cmp_pMux_9, b(23)=>nx9715, 
      b(22)=>nx9715, b(21)=>nx9713, b(20)=>nx9721, b(19)=>nx9719, b(18)=>
      nx9717, b(17)=>nx9715, b(16)=>nx9713, b(15)=>gen_23_cmp_BSCmp_op2_15, 
      b(14)=>gen_23_cmp_BSCmp_op2_14, b(13)=>gen_23_cmp_BSCmp_op2_13, b(12)
      =>gen_23_cmp_BSCmp_op2_12, b(11)=>gen_23_cmp_BSCmp_op2_11, b(10)=>
      gen_23_cmp_BSCmp_op2_10, b(9)=>gen_23_cmp_BSCmp_op2_9, b(8)=>
      gen_23_cmp_BSCmp_op2_8, b(7)=>gen_23_cmp_BSCmp_op2_7, b(6)=>
      gen_23_cmp_BSCmp_op2_6, b(5)=>gen_23_cmp_BSCmp_op2_5, b(4)=>
      gen_23_cmp_BSCmp_op2_4, b(3)=>gen_23_cmp_BSCmp_op2_3, b(2)=>
      gen_23_cmp_BSCmp_op2_2, b(1)=>gen_23_cmp_BSCmp_op2_1, b(0)=>
      gen_23_cmp_BSCmp_op2_0, carryIn=>gen_23_cmp_BSCmp_carryIn, sum(23)=>
      gen_23_cmp_pBs_30, sum(22)=>gen_23_cmp_pBs_29, sum(21)=>
      gen_23_cmp_pBs_28, sum(20)=>gen_23_cmp_pBs_27, sum(19)=>
      gen_23_cmp_pBs_26, sum(18)=>gen_23_cmp_pBs_25, sum(17)=>
      gen_23_cmp_pBs_24, sum(16)=>gen_23_cmp_pBs_23, sum(15)=>outputs_23_15, 
      sum(14)=>outputs_23_14, sum(13)=>outputs_23_13, sum(12)=>outputs_23_12, 
      sum(11)=>outputs_23_11, sum(10)=>outputs_23_10, sum(9)=>outputs_23_9, 
      sum(8)=>outputs_23_8, sum(7)=>outputs_23_7, sum(6)=>outputs_23_6, 
      sum(5)=>outputs_23_5, sum(4)=>outputs_23_4, sum(3)=>outputs_23_3, 
      sum(2)=>outputs_23_2, sum(1)=>outputs_23_1, sum(0)=>outputs_23_0, 
      carryOut=>DANGLING(9));
   gen_22_cmp_pRegCmp : Reg_33 port map ( D(32)=>working, D(31)=>working, 
      D(30)=>gen_22_cmp_pBs_30, D(29)=>gen_22_cmp_pBs_29, D(28)=>
      gen_22_cmp_pBs_28, D(27)=>gen_22_cmp_pBs_27, D(26)=>gen_22_cmp_pBs_26, 
      D(25)=>gen_22_cmp_pBs_25, D(24)=>gen_22_cmp_pBs_24, D(23)=>
      gen_22_cmp_pBs_23, D(22)=>outputs_22_15, D(21)=>outputs_22_14, D(20)=>
      outputs_22_13, D(19)=>outputs_22_12, D(18)=>outputs_22_11, D(17)=>
      outputs_22_10, D(16)=>outputs_22_9, D(15)=>outputs_22_8, D(14)=>
      outputs_22_7, D(13)=>outputs_22_6, D(12)=>outputs_22_5, D(11)=>
      outputs_22_4, D(10)=>outputs_22_3, D(9)=>outputs_22_2, D(8)=>
      outputs_22_1, D(7)=>outputs_22_0, D(6)=>gen_22_cmp_pMux_8, D(5)=>
      gen_22_cmp_pMux_7, D(4)=>gen_22_cmp_pMux_6, D(3)=>gen_22_cmp_pMux_5, 
      D(2)=>gen_22_cmp_pMux_4, D(1)=>gen_22_cmp_pMux_3, D(0)=>nx9423, en=>
      nx11159, clk=>nx9391, rst=>rst, Q(32)=>DANGLING(10), Q(31)=>DANGLING(
      11), Q(30)=>gen_22_cmp_pReg_30, Q(29)=>gen_22_cmp_pReg_29, Q(28)=>
      gen_22_cmp_pReg_28, Q(27)=>gen_22_cmp_pReg_27, Q(26)=>
      gen_22_cmp_pReg_26, Q(25)=>gen_22_cmp_pReg_25, Q(24)=>
      gen_22_cmp_pReg_24, Q(23)=>gen_22_cmp_pReg_23, Q(22)=>
      gen_22_cmp_pReg_22, Q(21)=>gen_22_cmp_pReg_21, Q(20)=>
      gen_22_cmp_pReg_20, Q(19)=>gen_22_cmp_pReg_19, Q(18)=>
      gen_22_cmp_pReg_18, Q(17)=>gen_22_cmp_pReg_17, Q(16)=>
      gen_22_cmp_pReg_16, Q(15)=>gen_22_cmp_pReg_15, Q(14)=>
      gen_22_cmp_pReg_14, Q(13)=>gen_22_cmp_pReg_13, Q(12)=>
      gen_22_cmp_pReg_12, Q(11)=>gen_22_cmp_pReg_11, Q(10)=>
      gen_22_cmp_pReg_10, Q(9)=>gen_22_cmp_pReg_9, Q(8)=>gen_22_cmp_pReg_8, 
      Q(7)=>gen_22_cmp_pReg_7, Q(6)=>gen_22_cmp_pReg_6, Q(5)=>
      gen_22_cmp_pReg_5, Q(4)=>gen_22_cmp_pReg_4, Q(3)=>gen_22_cmp_pReg_3, 
      Q(2)=>gen_22_cmp_pReg_2, Q(1)=>gen_22_cmp_pReg_1, Q(0)=>
      gen_22_cmp_pReg_0);
   gen_22_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>working, a(31)=>
      working, a(30)=>gen_22_cmp_pReg_30, a(29)=>gen_22_cmp_pReg_29, a(28)=>
      gen_22_cmp_pReg_28, a(27)=>gen_22_cmp_pReg_27, a(26)=>
      gen_22_cmp_pReg_26, a(25)=>gen_22_cmp_pReg_25, a(24)=>
      gen_22_cmp_pReg_24, a(23)=>gen_22_cmp_pReg_23, a(22)=>
      gen_22_cmp_pReg_22, a(21)=>gen_22_cmp_pReg_21, a(20)=>
      gen_22_cmp_pReg_20, a(19)=>gen_22_cmp_pReg_19, a(18)=>
      gen_22_cmp_pReg_18, a(17)=>gen_22_cmp_pReg_17, a(16)=>
      gen_22_cmp_pReg_16, a(15)=>gen_22_cmp_pReg_15, a(14)=>
      gen_22_cmp_pReg_14, a(13)=>gen_22_cmp_pReg_13, a(12)=>
      gen_22_cmp_pReg_12, a(11)=>gen_22_cmp_pReg_11, a(10)=>
      gen_22_cmp_pReg_10, a(9)=>gen_22_cmp_pReg_9, a(8)=>gen_22_cmp_pReg_8, 
      a(7)=>gen_22_cmp_pReg_7, a(6)=>gen_22_cmp_pReg_6, a(5)=>
      gen_22_cmp_pReg_5, a(4)=>gen_22_cmp_pReg_4, a(3)=>gen_22_cmp_pReg_3, 
      a(2)=>gen_22_cmp_pReg_2, a(1)=>gen_22_cmp_pReg_1, a(0)=>
      gen_22_cmp_pReg_0, b(32)=>working, b(31)=>working, b(30)=>working, 
      b(29)=>working, b(28)=>working, b(27)=>working, b(26)=>working, b(25)
      =>working, b(24)=>working, b(23)=>working, b(22)=>working, b(21)=>
      working, b(20)=>working, b(19)=>working, b(18)=>working, b(17)=>
      working, b(16)=>working, b(15)=>working, b(14)=>working, b(13)=>
      working, b(12)=>working, b(11)=>working, b(10)=>working, b(9)=>working, 
      b(8)=>filter_22_7, b(7)=>filter_22_6, b(6)=>filter_22_5, b(5)=>
      filter_22_4, b(4)=>filter_22_3, b(3)=>filter_22_2, b(2)=>filter_22_1, 
      b(1)=>filter_22_0, b(0)=>working, sel=>nx11173, f(32)=>DANGLING(12), 
      f(31)=>DANGLING(13), f(30)=>gen_22_cmp_pMux_30, f(29)=>
      gen_22_cmp_pMux_29, f(28)=>gen_22_cmp_pMux_28, f(27)=>
      gen_22_cmp_pMux_27, f(26)=>gen_22_cmp_pMux_26, f(25)=>
      gen_22_cmp_pMux_25, f(24)=>gen_22_cmp_pMux_24, f(23)=>
      gen_22_cmp_pMux_23, f(22)=>gen_22_cmp_pMux_22, f(21)=>
      gen_22_cmp_pMux_21, f(20)=>gen_22_cmp_pMux_20, f(19)=>
      gen_22_cmp_pMux_19, f(18)=>gen_22_cmp_pMux_18, f(17)=>
      gen_22_cmp_pMux_17, f(16)=>gen_22_cmp_pMux_16, f(15)=>
      gen_22_cmp_pMux_15, f(14)=>gen_22_cmp_pMux_14, f(13)=>
      gen_22_cmp_pMux_13, f(12)=>gen_22_cmp_pMux_12, f(11)=>
      gen_22_cmp_pMux_11, f(10)=>gen_22_cmp_pMux_10, f(9)=>gen_22_cmp_pMux_9, 
      f(8)=>gen_22_cmp_pMux_8, f(7)=>gen_22_cmp_pMux_7, f(6)=>
      gen_22_cmp_pMux_6, f(5)=>gen_22_cmp_pMux_5, f(4)=>gen_22_cmp_pMux_4, 
      f(3)=>gen_22_cmp_pMux_3, f(2)=>gen_22_cmp_pMux_2, f(1)=>
      gen_22_cmp_pMux_1, f(0)=>gen_22_cmp_pMux_0);
   gen_22_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>working, a(22)
      =>working, a(21)=>gen_22_cmp_pMux_30, a(20)=>gen_22_cmp_pMux_29, a(19)
      =>gen_22_cmp_pMux_28, a(18)=>gen_22_cmp_pMux_27, a(17)=>
      gen_22_cmp_pMux_26, a(16)=>gen_22_cmp_pMux_25, a(15)=>
      gen_22_cmp_pMux_24, a(14)=>gen_22_cmp_pMux_23, a(13)=>
      gen_22_cmp_pMux_22, a(12)=>gen_22_cmp_pMux_21, a(11)=>
      gen_22_cmp_pMux_20, a(10)=>gen_22_cmp_pMux_19, a(9)=>
      gen_22_cmp_pMux_18, a(8)=>gen_22_cmp_pMux_17, a(7)=>gen_22_cmp_pMux_16, 
      a(6)=>gen_22_cmp_pMux_15, a(5)=>gen_22_cmp_pMux_14, a(4)=>
      gen_22_cmp_pMux_13, a(3)=>gen_22_cmp_pMux_12, a(2)=>gen_22_cmp_pMux_11, 
      a(1)=>gen_22_cmp_pMux_10, a(0)=>gen_22_cmp_pMux_9, b(23)=>nx9727, 
      b(22)=>nx9727, b(21)=>nx9725, b(20)=>nx9733, b(19)=>nx9731, b(18)=>
      nx9729, b(17)=>nx9727, b(16)=>nx9725, b(15)=>gen_22_cmp_BSCmp_op2_15, 
      b(14)=>gen_22_cmp_BSCmp_op2_14, b(13)=>gen_22_cmp_BSCmp_op2_13, b(12)
      =>gen_22_cmp_BSCmp_op2_12, b(11)=>gen_22_cmp_BSCmp_op2_11, b(10)=>
      gen_22_cmp_BSCmp_op2_10, b(9)=>gen_22_cmp_BSCmp_op2_9, b(8)=>
      gen_22_cmp_BSCmp_op2_8, b(7)=>gen_22_cmp_BSCmp_op2_7, b(6)=>
      gen_22_cmp_BSCmp_op2_6, b(5)=>gen_22_cmp_BSCmp_op2_5, b(4)=>
      gen_22_cmp_BSCmp_op2_4, b(3)=>gen_22_cmp_BSCmp_op2_3, b(2)=>
      gen_22_cmp_BSCmp_op2_2, b(1)=>gen_22_cmp_BSCmp_op2_1, b(0)=>
      gen_22_cmp_BSCmp_op2_0, carryIn=>gen_22_cmp_BSCmp_carryIn, sum(23)=>
      gen_22_cmp_pBs_30, sum(22)=>gen_22_cmp_pBs_29, sum(21)=>
      gen_22_cmp_pBs_28, sum(20)=>gen_22_cmp_pBs_27, sum(19)=>
      gen_22_cmp_pBs_26, sum(18)=>gen_22_cmp_pBs_25, sum(17)=>
      gen_22_cmp_pBs_24, sum(16)=>gen_22_cmp_pBs_23, sum(15)=>outputs_22_15, 
      sum(14)=>outputs_22_14, sum(13)=>outputs_22_13, sum(12)=>outputs_22_12, 
      sum(11)=>outputs_22_11, sum(10)=>outputs_22_10, sum(9)=>outputs_22_9, 
      sum(8)=>outputs_22_8, sum(7)=>outputs_22_7, sum(6)=>outputs_22_6, 
      sum(5)=>outputs_22_5, sum(4)=>outputs_22_4, sum(3)=>outputs_22_3, 
      sum(2)=>outputs_22_2, sum(1)=>outputs_22_1, sum(0)=>outputs_22_0, 
      carryOut=>DANGLING(14));
   gen_21_cmp_pRegCmp : Reg_33 port map ( D(32)=>working, D(31)=>working, 
      D(30)=>gen_21_cmp_pBs_30, D(29)=>gen_21_cmp_pBs_29, D(28)=>
      gen_21_cmp_pBs_28, D(27)=>gen_21_cmp_pBs_27, D(26)=>gen_21_cmp_pBs_26, 
      D(25)=>gen_21_cmp_pBs_25, D(24)=>gen_21_cmp_pBs_24, D(23)=>
      gen_21_cmp_pBs_23, D(22)=>outputs_21_15, D(21)=>outputs_21_14, D(20)=>
      outputs_21_13, D(19)=>outputs_21_12, D(18)=>outputs_21_11, D(17)=>
      outputs_21_10, D(16)=>outputs_21_9, D(15)=>outputs_21_8, D(14)=>
      outputs_21_7, D(13)=>outputs_21_6, D(12)=>outputs_21_5, D(11)=>
      outputs_21_4, D(10)=>outputs_21_3, D(9)=>outputs_21_2, D(8)=>
      outputs_21_1, D(7)=>outputs_21_0, D(6)=>gen_21_cmp_pMux_8, D(5)=>
      gen_21_cmp_pMux_7, D(4)=>gen_21_cmp_pMux_6, D(3)=>gen_21_cmp_pMux_5, 
      D(2)=>gen_21_cmp_pMux_4, D(1)=>gen_21_cmp_pMux_3, D(0)=>nx9435, en=>
      nx11161, clk=>nx9391, rst=>rst, Q(32)=>DANGLING(15), Q(31)=>DANGLING(
      16), Q(30)=>gen_21_cmp_pReg_30, Q(29)=>gen_21_cmp_pReg_29, Q(28)=>
      gen_21_cmp_pReg_28, Q(27)=>gen_21_cmp_pReg_27, Q(26)=>
      gen_21_cmp_pReg_26, Q(25)=>gen_21_cmp_pReg_25, Q(24)=>
      gen_21_cmp_pReg_24, Q(23)=>gen_21_cmp_pReg_23, Q(22)=>
      gen_21_cmp_pReg_22, Q(21)=>gen_21_cmp_pReg_21, Q(20)=>
      gen_21_cmp_pReg_20, Q(19)=>gen_21_cmp_pReg_19, Q(18)=>
      gen_21_cmp_pReg_18, Q(17)=>gen_21_cmp_pReg_17, Q(16)=>
      gen_21_cmp_pReg_16, Q(15)=>gen_21_cmp_pReg_15, Q(14)=>
      gen_21_cmp_pReg_14, Q(13)=>gen_21_cmp_pReg_13, Q(12)=>
      gen_21_cmp_pReg_12, Q(11)=>gen_21_cmp_pReg_11, Q(10)=>
      gen_21_cmp_pReg_10, Q(9)=>gen_21_cmp_pReg_9, Q(8)=>gen_21_cmp_pReg_8, 
      Q(7)=>gen_21_cmp_pReg_7, Q(6)=>gen_21_cmp_pReg_6, Q(5)=>
      gen_21_cmp_pReg_5, Q(4)=>gen_21_cmp_pReg_4, Q(3)=>gen_21_cmp_pReg_3, 
      Q(2)=>gen_21_cmp_pReg_2, Q(1)=>gen_21_cmp_pReg_1, Q(0)=>
      gen_21_cmp_pReg_0);
   gen_21_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>working, a(31)=>
      working, a(30)=>gen_21_cmp_pReg_30, a(29)=>gen_21_cmp_pReg_29, a(28)=>
      gen_21_cmp_pReg_28, a(27)=>gen_21_cmp_pReg_27, a(26)=>
      gen_21_cmp_pReg_26, a(25)=>gen_21_cmp_pReg_25, a(24)=>
      gen_21_cmp_pReg_24, a(23)=>gen_21_cmp_pReg_23, a(22)=>
      gen_21_cmp_pReg_22, a(21)=>gen_21_cmp_pReg_21, a(20)=>
      gen_21_cmp_pReg_20, a(19)=>gen_21_cmp_pReg_19, a(18)=>
      gen_21_cmp_pReg_18, a(17)=>gen_21_cmp_pReg_17, a(16)=>
      gen_21_cmp_pReg_16, a(15)=>gen_21_cmp_pReg_15, a(14)=>
      gen_21_cmp_pReg_14, a(13)=>gen_21_cmp_pReg_13, a(12)=>
      gen_21_cmp_pReg_12, a(11)=>gen_21_cmp_pReg_11, a(10)=>
      gen_21_cmp_pReg_10, a(9)=>gen_21_cmp_pReg_9, a(8)=>gen_21_cmp_pReg_8, 
      a(7)=>gen_21_cmp_pReg_7, a(6)=>gen_21_cmp_pReg_6, a(5)=>
      gen_21_cmp_pReg_5, a(4)=>gen_21_cmp_pReg_4, a(3)=>gen_21_cmp_pReg_3, 
      a(2)=>gen_21_cmp_pReg_2, a(1)=>gen_21_cmp_pReg_1, a(0)=>
      gen_21_cmp_pReg_0, b(32)=>working, b(31)=>working, b(30)=>working, 
      b(29)=>working, b(28)=>working, b(27)=>working, b(26)=>working, b(25)
      =>working, b(24)=>working, b(23)=>working, b(22)=>working, b(21)=>
      working, b(20)=>working, b(19)=>working, b(18)=>working, b(17)=>
      working, b(16)=>working, b(15)=>working, b(14)=>working, b(13)=>
      working, b(12)=>working, b(11)=>working, b(10)=>working, b(9)=>working, 
      b(8)=>filter_21_7, b(7)=>filter_21_6, b(6)=>filter_21_5, b(5)=>
      filter_21_4, b(4)=>filter_21_3, b(3)=>filter_21_2, b(2)=>filter_21_1, 
      b(1)=>filter_21_0, b(0)=>working, sel=>nx11175, f(32)=>DANGLING(17), 
      f(31)=>DANGLING(18), f(30)=>gen_21_cmp_pMux_30, f(29)=>
      gen_21_cmp_pMux_29, f(28)=>gen_21_cmp_pMux_28, f(27)=>
      gen_21_cmp_pMux_27, f(26)=>gen_21_cmp_pMux_26, f(25)=>
      gen_21_cmp_pMux_25, f(24)=>gen_21_cmp_pMux_24, f(23)=>
      gen_21_cmp_pMux_23, f(22)=>gen_21_cmp_pMux_22, f(21)=>
      gen_21_cmp_pMux_21, f(20)=>gen_21_cmp_pMux_20, f(19)=>
      gen_21_cmp_pMux_19, f(18)=>gen_21_cmp_pMux_18, f(17)=>
      gen_21_cmp_pMux_17, f(16)=>gen_21_cmp_pMux_16, f(15)=>
      gen_21_cmp_pMux_15, f(14)=>gen_21_cmp_pMux_14, f(13)=>
      gen_21_cmp_pMux_13, f(12)=>gen_21_cmp_pMux_12, f(11)=>
      gen_21_cmp_pMux_11, f(10)=>gen_21_cmp_pMux_10, f(9)=>gen_21_cmp_pMux_9, 
      f(8)=>gen_21_cmp_pMux_8, f(7)=>gen_21_cmp_pMux_7, f(6)=>
      gen_21_cmp_pMux_6, f(5)=>gen_21_cmp_pMux_5, f(4)=>gen_21_cmp_pMux_4, 
      f(3)=>gen_21_cmp_pMux_3, f(2)=>gen_21_cmp_pMux_2, f(1)=>
      gen_21_cmp_pMux_1, f(0)=>gen_21_cmp_pMux_0);
   gen_21_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>working, a(22)
      =>working, a(21)=>gen_21_cmp_pMux_30, a(20)=>gen_21_cmp_pMux_29, a(19)
      =>gen_21_cmp_pMux_28, a(18)=>gen_21_cmp_pMux_27, a(17)=>
      gen_21_cmp_pMux_26, a(16)=>gen_21_cmp_pMux_25, a(15)=>
      gen_21_cmp_pMux_24, a(14)=>gen_21_cmp_pMux_23, a(13)=>
      gen_21_cmp_pMux_22, a(12)=>gen_21_cmp_pMux_21, a(11)=>
      gen_21_cmp_pMux_20, a(10)=>gen_21_cmp_pMux_19, a(9)=>
      gen_21_cmp_pMux_18, a(8)=>gen_21_cmp_pMux_17, a(7)=>gen_21_cmp_pMux_16, 
      a(6)=>gen_21_cmp_pMux_15, a(5)=>gen_21_cmp_pMux_14, a(4)=>
      gen_21_cmp_pMux_13, a(3)=>gen_21_cmp_pMux_12, a(2)=>gen_21_cmp_pMux_11, 
      a(1)=>gen_21_cmp_pMux_10, a(0)=>gen_21_cmp_pMux_9, b(23)=>nx9739, 
      b(22)=>nx9739, b(21)=>nx9737, b(20)=>nx9745, b(19)=>nx9743, b(18)=>
      nx9741, b(17)=>nx9739, b(16)=>nx9737, b(15)=>gen_21_cmp_BSCmp_op2_15, 
      b(14)=>gen_21_cmp_BSCmp_op2_14, b(13)=>gen_21_cmp_BSCmp_op2_13, b(12)
      =>gen_21_cmp_BSCmp_op2_12, b(11)=>gen_21_cmp_BSCmp_op2_11, b(10)=>
      gen_21_cmp_BSCmp_op2_10, b(9)=>gen_21_cmp_BSCmp_op2_9, b(8)=>
      gen_21_cmp_BSCmp_op2_8, b(7)=>gen_21_cmp_BSCmp_op2_7, b(6)=>
      gen_21_cmp_BSCmp_op2_6, b(5)=>gen_21_cmp_BSCmp_op2_5, b(4)=>
      gen_21_cmp_BSCmp_op2_4, b(3)=>gen_21_cmp_BSCmp_op2_3, b(2)=>
      gen_21_cmp_BSCmp_op2_2, b(1)=>gen_21_cmp_BSCmp_op2_1, b(0)=>
      gen_21_cmp_BSCmp_op2_0, carryIn=>gen_21_cmp_BSCmp_carryIn, sum(23)=>
      gen_21_cmp_pBs_30, sum(22)=>gen_21_cmp_pBs_29, sum(21)=>
      gen_21_cmp_pBs_28, sum(20)=>gen_21_cmp_pBs_27, sum(19)=>
      gen_21_cmp_pBs_26, sum(18)=>gen_21_cmp_pBs_25, sum(17)=>
      gen_21_cmp_pBs_24, sum(16)=>gen_21_cmp_pBs_23, sum(15)=>outputs_21_15, 
      sum(14)=>outputs_21_14, sum(13)=>outputs_21_13, sum(12)=>outputs_21_12, 
      sum(11)=>outputs_21_11, sum(10)=>outputs_21_10, sum(9)=>outputs_21_9, 
      sum(8)=>outputs_21_8, sum(7)=>outputs_21_7, sum(6)=>outputs_21_6, 
      sum(5)=>outputs_21_5, sum(4)=>outputs_21_4, sum(3)=>outputs_21_3, 
      sum(2)=>outputs_21_2, sum(1)=>outputs_21_1, sum(0)=>outputs_21_0, 
      carryOut=>DANGLING(19));
   gen_20_cmp_pRegCmp : Reg_33 port map ( D(32)=>working, D(31)=>working, 
      D(30)=>gen_20_cmp_pBs_30, D(29)=>gen_20_cmp_pBs_29, D(28)=>
      gen_20_cmp_pBs_28, D(27)=>gen_20_cmp_pBs_27, D(26)=>gen_20_cmp_pBs_26, 
      D(25)=>gen_20_cmp_pBs_25, D(24)=>gen_20_cmp_pBs_24, D(23)=>
      gen_20_cmp_pBs_23, D(22)=>outputs_20_15, D(21)=>outputs_20_14, D(20)=>
      outputs_20_13, D(19)=>outputs_20_12, D(18)=>outputs_20_11, D(17)=>
      outputs_20_10, D(16)=>outputs_20_9, D(15)=>outputs_20_8, D(14)=>
      outputs_20_7, D(13)=>outputs_20_6, D(12)=>outputs_20_5, D(11)=>
      outputs_20_4, D(10)=>outputs_20_3, D(9)=>outputs_20_2, D(8)=>
      outputs_20_1, D(7)=>outputs_20_0, D(6)=>gen_20_cmp_pMux_8, D(5)=>
      gen_20_cmp_pMux_7, D(4)=>gen_20_cmp_pMux_6, D(3)=>gen_20_cmp_pMux_5, 
      D(2)=>gen_20_cmp_pMux_4, D(1)=>gen_20_cmp_pMux_3, D(0)=>nx9447, en=>
      nx11161, clk=>nx9391, rst=>rst, Q(32)=>DANGLING(20), Q(31)=>DANGLING(
      21), Q(30)=>gen_20_cmp_pReg_30, Q(29)=>gen_20_cmp_pReg_29, Q(28)=>
      gen_20_cmp_pReg_28, Q(27)=>gen_20_cmp_pReg_27, Q(26)=>
      gen_20_cmp_pReg_26, Q(25)=>gen_20_cmp_pReg_25, Q(24)=>
      gen_20_cmp_pReg_24, Q(23)=>gen_20_cmp_pReg_23, Q(22)=>
      gen_20_cmp_pReg_22, Q(21)=>gen_20_cmp_pReg_21, Q(20)=>
      gen_20_cmp_pReg_20, Q(19)=>gen_20_cmp_pReg_19, Q(18)=>
      gen_20_cmp_pReg_18, Q(17)=>gen_20_cmp_pReg_17, Q(16)=>
      gen_20_cmp_pReg_16, Q(15)=>gen_20_cmp_pReg_15, Q(14)=>
      gen_20_cmp_pReg_14, Q(13)=>gen_20_cmp_pReg_13, Q(12)=>
      gen_20_cmp_pReg_12, Q(11)=>gen_20_cmp_pReg_11, Q(10)=>
      gen_20_cmp_pReg_10, Q(9)=>gen_20_cmp_pReg_9, Q(8)=>gen_20_cmp_pReg_8, 
      Q(7)=>gen_20_cmp_pReg_7, Q(6)=>gen_20_cmp_pReg_6, Q(5)=>
      gen_20_cmp_pReg_5, Q(4)=>gen_20_cmp_pReg_4, Q(3)=>gen_20_cmp_pReg_3, 
      Q(2)=>gen_20_cmp_pReg_2, Q(1)=>gen_20_cmp_pReg_1, Q(0)=>
      gen_20_cmp_pReg_0);
   gen_20_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>working, a(31)=>
      working, a(30)=>gen_20_cmp_pReg_30, a(29)=>gen_20_cmp_pReg_29, a(28)=>
      gen_20_cmp_pReg_28, a(27)=>gen_20_cmp_pReg_27, a(26)=>
      gen_20_cmp_pReg_26, a(25)=>gen_20_cmp_pReg_25, a(24)=>
      gen_20_cmp_pReg_24, a(23)=>gen_20_cmp_pReg_23, a(22)=>
      gen_20_cmp_pReg_22, a(21)=>gen_20_cmp_pReg_21, a(20)=>
      gen_20_cmp_pReg_20, a(19)=>gen_20_cmp_pReg_19, a(18)=>
      gen_20_cmp_pReg_18, a(17)=>gen_20_cmp_pReg_17, a(16)=>
      gen_20_cmp_pReg_16, a(15)=>gen_20_cmp_pReg_15, a(14)=>
      gen_20_cmp_pReg_14, a(13)=>gen_20_cmp_pReg_13, a(12)=>
      gen_20_cmp_pReg_12, a(11)=>gen_20_cmp_pReg_11, a(10)=>
      gen_20_cmp_pReg_10, a(9)=>gen_20_cmp_pReg_9, a(8)=>gen_20_cmp_pReg_8, 
      a(7)=>gen_20_cmp_pReg_7, a(6)=>gen_20_cmp_pReg_6, a(5)=>
      gen_20_cmp_pReg_5, a(4)=>gen_20_cmp_pReg_4, a(3)=>gen_20_cmp_pReg_3, 
      a(2)=>gen_20_cmp_pReg_2, a(1)=>gen_20_cmp_pReg_1, a(0)=>
      gen_20_cmp_pReg_0, b(32)=>working, b(31)=>working, b(30)=>working, 
      b(29)=>working, b(28)=>working, b(27)=>working, b(26)=>working, b(25)
      =>working, b(24)=>working, b(23)=>working, b(22)=>working, b(21)=>
      working, b(20)=>working, b(19)=>working, b(18)=>working, b(17)=>
      working, b(16)=>working, b(15)=>working, b(14)=>working, b(13)=>
      working, b(12)=>working, b(11)=>working, b(10)=>working, b(9)=>working, 
      b(8)=>filter_20_7, b(7)=>filter_20_6, b(6)=>filter_20_5, b(5)=>
      filter_20_4, b(4)=>filter_20_3, b(3)=>filter_20_2, b(2)=>filter_20_1, 
      b(1)=>filter_20_0, b(0)=>working, sel=>nx11175, f(32)=>DANGLING(22), 
      f(31)=>DANGLING(23), f(30)=>gen_20_cmp_pMux_30, f(29)=>
      gen_20_cmp_pMux_29, f(28)=>gen_20_cmp_pMux_28, f(27)=>
      gen_20_cmp_pMux_27, f(26)=>gen_20_cmp_pMux_26, f(25)=>
      gen_20_cmp_pMux_25, f(24)=>gen_20_cmp_pMux_24, f(23)=>
      gen_20_cmp_pMux_23, f(22)=>gen_20_cmp_pMux_22, f(21)=>
      gen_20_cmp_pMux_21, f(20)=>gen_20_cmp_pMux_20, f(19)=>
      gen_20_cmp_pMux_19, f(18)=>gen_20_cmp_pMux_18, f(17)=>
      gen_20_cmp_pMux_17, f(16)=>gen_20_cmp_pMux_16, f(15)=>
      gen_20_cmp_pMux_15, f(14)=>gen_20_cmp_pMux_14, f(13)=>
      gen_20_cmp_pMux_13, f(12)=>gen_20_cmp_pMux_12, f(11)=>
      gen_20_cmp_pMux_11, f(10)=>gen_20_cmp_pMux_10, f(9)=>gen_20_cmp_pMux_9, 
      f(8)=>gen_20_cmp_pMux_8, f(7)=>gen_20_cmp_pMux_7, f(6)=>
      gen_20_cmp_pMux_6, f(5)=>gen_20_cmp_pMux_5, f(4)=>gen_20_cmp_pMux_4, 
      f(3)=>gen_20_cmp_pMux_3, f(2)=>gen_20_cmp_pMux_2, f(1)=>
      gen_20_cmp_pMux_1, f(0)=>gen_20_cmp_pMux_0);
   gen_20_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>working, a(22)
      =>working, a(21)=>gen_20_cmp_pMux_30, a(20)=>gen_20_cmp_pMux_29, a(19)
      =>gen_20_cmp_pMux_28, a(18)=>gen_20_cmp_pMux_27, a(17)=>
      gen_20_cmp_pMux_26, a(16)=>gen_20_cmp_pMux_25, a(15)=>
      gen_20_cmp_pMux_24, a(14)=>gen_20_cmp_pMux_23, a(13)=>
      gen_20_cmp_pMux_22, a(12)=>gen_20_cmp_pMux_21, a(11)=>
      gen_20_cmp_pMux_20, a(10)=>gen_20_cmp_pMux_19, a(9)=>
      gen_20_cmp_pMux_18, a(8)=>gen_20_cmp_pMux_17, a(7)=>gen_20_cmp_pMux_16, 
      a(6)=>gen_20_cmp_pMux_15, a(5)=>gen_20_cmp_pMux_14, a(4)=>
      gen_20_cmp_pMux_13, a(3)=>gen_20_cmp_pMux_12, a(2)=>gen_20_cmp_pMux_11, 
      a(1)=>gen_20_cmp_pMux_10, a(0)=>gen_20_cmp_pMux_9, b(23)=>nx9751, 
      b(22)=>nx9751, b(21)=>nx9749, b(20)=>nx9757, b(19)=>nx9755, b(18)=>
      nx9753, b(17)=>nx9751, b(16)=>nx9749, b(15)=>gen_20_cmp_BSCmp_op2_15, 
      b(14)=>gen_20_cmp_BSCmp_op2_14, b(13)=>gen_20_cmp_BSCmp_op2_13, b(12)
      =>gen_20_cmp_BSCmp_op2_12, b(11)=>gen_20_cmp_BSCmp_op2_11, b(10)=>
      gen_20_cmp_BSCmp_op2_10, b(9)=>gen_20_cmp_BSCmp_op2_9, b(8)=>
      gen_20_cmp_BSCmp_op2_8, b(7)=>gen_20_cmp_BSCmp_op2_7, b(6)=>
      gen_20_cmp_BSCmp_op2_6, b(5)=>gen_20_cmp_BSCmp_op2_5, b(4)=>
      gen_20_cmp_BSCmp_op2_4, b(3)=>gen_20_cmp_BSCmp_op2_3, b(2)=>
      gen_20_cmp_BSCmp_op2_2, b(1)=>gen_20_cmp_BSCmp_op2_1, b(0)=>
      gen_20_cmp_BSCmp_op2_0, carryIn=>gen_20_cmp_BSCmp_carryIn, sum(23)=>
      gen_20_cmp_pBs_30, sum(22)=>gen_20_cmp_pBs_29, sum(21)=>
      gen_20_cmp_pBs_28, sum(20)=>gen_20_cmp_pBs_27, sum(19)=>
      gen_20_cmp_pBs_26, sum(18)=>gen_20_cmp_pBs_25, sum(17)=>
      gen_20_cmp_pBs_24, sum(16)=>gen_20_cmp_pBs_23, sum(15)=>outputs_20_15, 
      sum(14)=>outputs_20_14, sum(13)=>outputs_20_13, sum(12)=>outputs_20_12, 
      sum(11)=>outputs_20_11, sum(10)=>outputs_20_10, sum(9)=>outputs_20_9, 
      sum(8)=>outputs_20_8, sum(7)=>outputs_20_7, sum(6)=>outputs_20_6, 
      sum(5)=>outputs_20_5, sum(4)=>outputs_20_4, sum(3)=>outputs_20_3, 
      sum(2)=>outputs_20_2, sum(1)=>outputs_20_1, sum(0)=>outputs_20_0, 
      carryOut=>DANGLING(24));
   gen_19_cmp_pRegCmp : Reg_33 port map ( D(32)=>working, D(31)=>working, 
      D(30)=>gen_19_cmp_pBs_30, D(29)=>gen_19_cmp_pBs_29, D(28)=>
      gen_19_cmp_pBs_28, D(27)=>gen_19_cmp_pBs_27, D(26)=>gen_19_cmp_pBs_26, 
      D(25)=>gen_19_cmp_pBs_25, D(24)=>gen_19_cmp_pBs_24, D(23)=>
      gen_19_cmp_pBs_23, D(22)=>outputs_19_15, D(21)=>outputs_19_14, D(20)=>
      outputs_19_13, D(19)=>outputs_19_12, D(18)=>outputs_19_11, D(17)=>
      outputs_19_10, D(16)=>outputs_19_9, D(15)=>outputs_19_8, D(14)=>
      outputs_19_7, D(13)=>outputs_19_6, D(12)=>outputs_19_5, D(11)=>
      outputs_19_4, D(10)=>outputs_19_3, D(9)=>outputs_19_2, D(8)=>
      outputs_19_1, D(7)=>outputs_19_0, D(6)=>gen_19_cmp_pMux_8, D(5)=>
      gen_19_cmp_pMux_7, D(4)=>gen_19_cmp_pMux_6, D(3)=>gen_19_cmp_pMux_5, 
      D(2)=>gen_19_cmp_pMux_4, D(1)=>gen_19_cmp_pMux_3, D(0)=>nx9459, en=>
      nx11161, clk=>nx9391, rst=>rst, Q(32)=>DANGLING(25), Q(31)=>DANGLING(
      26), Q(30)=>gen_19_cmp_pReg_30, Q(29)=>gen_19_cmp_pReg_29, Q(28)=>
      gen_19_cmp_pReg_28, Q(27)=>gen_19_cmp_pReg_27, Q(26)=>
      gen_19_cmp_pReg_26, Q(25)=>gen_19_cmp_pReg_25, Q(24)=>
      gen_19_cmp_pReg_24, Q(23)=>gen_19_cmp_pReg_23, Q(22)=>
      gen_19_cmp_pReg_22, Q(21)=>gen_19_cmp_pReg_21, Q(20)=>
      gen_19_cmp_pReg_20, Q(19)=>gen_19_cmp_pReg_19, Q(18)=>
      gen_19_cmp_pReg_18, Q(17)=>gen_19_cmp_pReg_17, Q(16)=>
      gen_19_cmp_pReg_16, Q(15)=>gen_19_cmp_pReg_15, Q(14)=>
      gen_19_cmp_pReg_14, Q(13)=>gen_19_cmp_pReg_13, Q(12)=>
      gen_19_cmp_pReg_12, Q(11)=>gen_19_cmp_pReg_11, Q(10)=>
      gen_19_cmp_pReg_10, Q(9)=>gen_19_cmp_pReg_9, Q(8)=>gen_19_cmp_pReg_8, 
      Q(7)=>gen_19_cmp_pReg_7, Q(6)=>gen_19_cmp_pReg_6, Q(5)=>
      gen_19_cmp_pReg_5, Q(4)=>gen_19_cmp_pReg_4, Q(3)=>gen_19_cmp_pReg_3, 
      Q(2)=>gen_19_cmp_pReg_2, Q(1)=>gen_19_cmp_pReg_1, Q(0)=>
      gen_19_cmp_pReg_0);
   gen_19_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>working, a(31)=>
      working, a(30)=>gen_19_cmp_pReg_30, a(29)=>gen_19_cmp_pReg_29, a(28)=>
      gen_19_cmp_pReg_28, a(27)=>gen_19_cmp_pReg_27, a(26)=>
      gen_19_cmp_pReg_26, a(25)=>gen_19_cmp_pReg_25, a(24)=>
      gen_19_cmp_pReg_24, a(23)=>gen_19_cmp_pReg_23, a(22)=>
      gen_19_cmp_pReg_22, a(21)=>gen_19_cmp_pReg_21, a(20)=>
      gen_19_cmp_pReg_20, a(19)=>gen_19_cmp_pReg_19, a(18)=>
      gen_19_cmp_pReg_18, a(17)=>gen_19_cmp_pReg_17, a(16)=>
      gen_19_cmp_pReg_16, a(15)=>gen_19_cmp_pReg_15, a(14)=>
      gen_19_cmp_pReg_14, a(13)=>gen_19_cmp_pReg_13, a(12)=>
      gen_19_cmp_pReg_12, a(11)=>gen_19_cmp_pReg_11, a(10)=>
      gen_19_cmp_pReg_10, a(9)=>gen_19_cmp_pReg_9, a(8)=>gen_19_cmp_pReg_8, 
      a(7)=>gen_19_cmp_pReg_7, a(6)=>gen_19_cmp_pReg_6, a(5)=>
      gen_19_cmp_pReg_5, a(4)=>gen_19_cmp_pReg_4, a(3)=>gen_19_cmp_pReg_3, 
      a(2)=>gen_19_cmp_pReg_2, a(1)=>gen_19_cmp_pReg_1, a(0)=>
      gen_19_cmp_pReg_0, b(32)=>working, b(31)=>working, b(30)=>working, 
      b(29)=>working, b(28)=>working, b(27)=>working, b(26)=>working, b(25)
      =>working, b(24)=>working, b(23)=>working, b(22)=>working, b(21)=>
      working, b(20)=>working, b(19)=>working, b(18)=>working, b(17)=>
      working, b(16)=>working, b(15)=>working, b(14)=>working, b(13)=>
      working, b(12)=>working, b(11)=>working, b(10)=>working, b(9)=>working, 
      b(8)=>filter_19_7, b(7)=>filter_19_6, b(6)=>filter_19_5, b(5)=>
      filter_19_4, b(4)=>filter_19_3, b(3)=>filter_19_2, b(2)=>filter_19_1, 
      b(1)=>filter_19_0, b(0)=>working, sel=>nx11175, f(32)=>DANGLING(27), 
      f(31)=>DANGLING(28), f(30)=>gen_19_cmp_pMux_30, f(29)=>
      gen_19_cmp_pMux_29, f(28)=>gen_19_cmp_pMux_28, f(27)=>
      gen_19_cmp_pMux_27, f(26)=>gen_19_cmp_pMux_26, f(25)=>
      gen_19_cmp_pMux_25, f(24)=>gen_19_cmp_pMux_24, f(23)=>
      gen_19_cmp_pMux_23, f(22)=>gen_19_cmp_pMux_22, f(21)=>
      gen_19_cmp_pMux_21, f(20)=>gen_19_cmp_pMux_20, f(19)=>
      gen_19_cmp_pMux_19, f(18)=>gen_19_cmp_pMux_18, f(17)=>
      gen_19_cmp_pMux_17, f(16)=>gen_19_cmp_pMux_16, f(15)=>
      gen_19_cmp_pMux_15, f(14)=>gen_19_cmp_pMux_14, f(13)=>
      gen_19_cmp_pMux_13, f(12)=>gen_19_cmp_pMux_12, f(11)=>
      gen_19_cmp_pMux_11, f(10)=>gen_19_cmp_pMux_10, f(9)=>gen_19_cmp_pMux_9, 
      f(8)=>gen_19_cmp_pMux_8, f(7)=>gen_19_cmp_pMux_7, f(6)=>
      gen_19_cmp_pMux_6, f(5)=>gen_19_cmp_pMux_5, f(4)=>gen_19_cmp_pMux_4, 
      f(3)=>gen_19_cmp_pMux_3, f(2)=>gen_19_cmp_pMux_2, f(1)=>
      gen_19_cmp_pMux_1, f(0)=>gen_19_cmp_pMux_0);
   gen_19_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>working, a(22)
      =>working, a(21)=>gen_19_cmp_pMux_30, a(20)=>gen_19_cmp_pMux_29, a(19)
      =>gen_19_cmp_pMux_28, a(18)=>gen_19_cmp_pMux_27, a(17)=>
      gen_19_cmp_pMux_26, a(16)=>gen_19_cmp_pMux_25, a(15)=>
      gen_19_cmp_pMux_24, a(14)=>gen_19_cmp_pMux_23, a(13)=>
      gen_19_cmp_pMux_22, a(12)=>gen_19_cmp_pMux_21, a(11)=>
      gen_19_cmp_pMux_20, a(10)=>gen_19_cmp_pMux_19, a(9)=>
      gen_19_cmp_pMux_18, a(8)=>gen_19_cmp_pMux_17, a(7)=>gen_19_cmp_pMux_16, 
      a(6)=>gen_19_cmp_pMux_15, a(5)=>gen_19_cmp_pMux_14, a(4)=>
      gen_19_cmp_pMux_13, a(3)=>gen_19_cmp_pMux_12, a(2)=>gen_19_cmp_pMux_11, 
      a(1)=>gen_19_cmp_pMux_10, a(0)=>gen_19_cmp_pMux_9, b(23)=>nx9763, 
      b(22)=>nx9763, b(21)=>nx9761, b(20)=>nx9769, b(19)=>nx9767, b(18)=>
      nx9765, b(17)=>nx9763, b(16)=>nx9761, b(15)=>gen_19_cmp_BSCmp_op2_15, 
      b(14)=>gen_19_cmp_BSCmp_op2_14, b(13)=>gen_19_cmp_BSCmp_op2_13, b(12)
      =>gen_19_cmp_BSCmp_op2_12, b(11)=>gen_19_cmp_BSCmp_op2_11, b(10)=>
      gen_19_cmp_BSCmp_op2_10, b(9)=>gen_19_cmp_BSCmp_op2_9, b(8)=>
      gen_19_cmp_BSCmp_op2_8, b(7)=>gen_19_cmp_BSCmp_op2_7, b(6)=>
      gen_19_cmp_BSCmp_op2_6, b(5)=>gen_19_cmp_BSCmp_op2_5, b(4)=>
      gen_19_cmp_BSCmp_op2_4, b(3)=>gen_19_cmp_BSCmp_op2_3, b(2)=>
      gen_19_cmp_BSCmp_op2_2, b(1)=>gen_19_cmp_BSCmp_op2_1, b(0)=>
      gen_19_cmp_BSCmp_op2_0, carryIn=>gen_19_cmp_BSCmp_carryIn, sum(23)=>
      gen_19_cmp_pBs_30, sum(22)=>gen_19_cmp_pBs_29, sum(21)=>
      gen_19_cmp_pBs_28, sum(20)=>gen_19_cmp_pBs_27, sum(19)=>
      gen_19_cmp_pBs_26, sum(18)=>gen_19_cmp_pBs_25, sum(17)=>
      gen_19_cmp_pBs_24, sum(16)=>gen_19_cmp_pBs_23, sum(15)=>outputs_19_15, 
      sum(14)=>outputs_19_14, sum(13)=>outputs_19_13, sum(12)=>outputs_19_12, 
      sum(11)=>outputs_19_11, sum(10)=>outputs_19_10, sum(9)=>outputs_19_9, 
      sum(8)=>outputs_19_8, sum(7)=>outputs_19_7, sum(6)=>outputs_19_6, 
      sum(5)=>outputs_19_5, sum(4)=>outputs_19_4, sum(3)=>outputs_19_3, 
      sum(2)=>outputs_19_2, sum(1)=>outputs_19_1, sum(0)=>outputs_19_0, 
      carryOut=>DANGLING(29));
   gen_18_cmp_pRegCmp : Reg_33 port map ( D(32)=>working, D(31)=>working, 
      D(30)=>gen_18_cmp_pBs_30, D(29)=>gen_18_cmp_pBs_29, D(28)=>
      gen_18_cmp_pBs_28, D(27)=>gen_18_cmp_pBs_27, D(26)=>gen_18_cmp_pBs_26, 
      D(25)=>gen_18_cmp_pBs_25, D(24)=>gen_18_cmp_pBs_24, D(23)=>
      gen_18_cmp_pBs_23, D(22)=>outputs_18_15, D(21)=>outputs_18_14, D(20)=>
      outputs_18_13, D(19)=>outputs_18_12, D(18)=>outputs_18_11, D(17)=>
      outputs_18_10, D(16)=>outputs_18_9, D(15)=>outputs_18_8, D(14)=>
      outputs_18_7, D(13)=>outputs_18_6, D(12)=>outputs_18_5, D(11)=>
      outputs_18_4, D(10)=>outputs_18_3, D(9)=>outputs_18_2, D(8)=>
      outputs_18_1, D(7)=>outputs_18_0, D(6)=>gen_18_cmp_pMux_8, D(5)=>
      gen_18_cmp_pMux_7, D(4)=>gen_18_cmp_pMux_6, D(3)=>gen_18_cmp_pMux_5, 
      D(2)=>gen_18_cmp_pMux_4, D(1)=>gen_18_cmp_pMux_3, D(0)=>nx9471, en=>
      nx9375, clk=>nx9391, rst=>rst, Q(32)=>DANGLING(30), Q(31)=>DANGLING(31
      ), Q(30)=>gen_18_cmp_pReg_30, Q(29)=>gen_18_cmp_pReg_29, Q(28)=>
      gen_18_cmp_pReg_28, Q(27)=>gen_18_cmp_pReg_27, Q(26)=>
      gen_18_cmp_pReg_26, Q(25)=>gen_18_cmp_pReg_25, Q(24)=>
      gen_18_cmp_pReg_24, Q(23)=>gen_18_cmp_pReg_23, Q(22)=>
      gen_18_cmp_pReg_22, Q(21)=>gen_18_cmp_pReg_21, Q(20)=>
      gen_18_cmp_pReg_20, Q(19)=>gen_18_cmp_pReg_19, Q(18)=>
      gen_18_cmp_pReg_18, Q(17)=>gen_18_cmp_pReg_17, Q(16)=>
      gen_18_cmp_pReg_16, Q(15)=>gen_18_cmp_pReg_15, Q(14)=>
      gen_18_cmp_pReg_14, Q(13)=>gen_18_cmp_pReg_13, Q(12)=>
      gen_18_cmp_pReg_12, Q(11)=>gen_18_cmp_pReg_11, Q(10)=>
      gen_18_cmp_pReg_10, Q(9)=>gen_18_cmp_pReg_9, Q(8)=>gen_18_cmp_pReg_8, 
      Q(7)=>gen_18_cmp_pReg_7, Q(6)=>gen_18_cmp_pReg_6, Q(5)=>
      gen_18_cmp_pReg_5, Q(4)=>gen_18_cmp_pReg_4, Q(3)=>gen_18_cmp_pReg_3, 
      Q(2)=>gen_18_cmp_pReg_2, Q(1)=>gen_18_cmp_pReg_1, Q(0)=>
      gen_18_cmp_pReg_0);
   gen_18_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>working, a(31)=>
      working, a(30)=>gen_18_cmp_pReg_30, a(29)=>gen_18_cmp_pReg_29, a(28)=>
      gen_18_cmp_pReg_28, a(27)=>gen_18_cmp_pReg_27, a(26)=>
      gen_18_cmp_pReg_26, a(25)=>gen_18_cmp_pReg_25, a(24)=>
      gen_18_cmp_pReg_24, a(23)=>gen_18_cmp_pReg_23, a(22)=>
      gen_18_cmp_pReg_22, a(21)=>gen_18_cmp_pReg_21, a(20)=>
      gen_18_cmp_pReg_20, a(19)=>gen_18_cmp_pReg_19, a(18)=>
      gen_18_cmp_pReg_18, a(17)=>gen_18_cmp_pReg_17, a(16)=>
      gen_18_cmp_pReg_16, a(15)=>gen_18_cmp_pReg_15, a(14)=>
      gen_18_cmp_pReg_14, a(13)=>gen_18_cmp_pReg_13, a(12)=>
      gen_18_cmp_pReg_12, a(11)=>gen_18_cmp_pReg_11, a(10)=>
      gen_18_cmp_pReg_10, a(9)=>gen_18_cmp_pReg_9, a(8)=>gen_18_cmp_pReg_8, 
      a(7)=>gen_18_cmp_pReg_7, a(6)=>gen_18_cmp_pReg_6, a(5)=>
      gen_18_cmp_pReg_5, a(4)=>gen_18_cmp_pReg_4, a(3)=>gen_18_cmp_pReg_3, 
      a(2)=>gen_18_cmp_pReg_2, a(1)=>gen_18_cmp_pReg_1, a(0)=>
      gen_18_cmp_pReg_0, b(32)=>working, b(31)=>working, b(30)=>working, 
      b(29)=>working, b(28)=>working, b(27)=>working, b(26)=>working, b(25)
      =>working, b(24)=>working, b(23)=>working, b(22)=>working, b(21)=>
      working, b(20)=>working, b(19)=>working, b(18)=>working, b(17)=>
      working, b(16)=>working, b(15)=>working, b(14)=>working, b(13)=>
      working, b(12)=>working, b(11)=>working, b(10)=>working, b(9)=>working, 
      b(8)=>filter_18_7, b(7)=>filter_18_6, b(6)=>filter_18_5, b(5)=>
      filter_18_4, b(4)=>filter_18_3, b(3)=>filter_18_2, b(2)=>filter_18_1, 
      b(1)=>filter_18_0, b(0)=>working, sel=>nx11177, f(32)=>DANGLING(32), 
      f(31)=>DANGLING(33), f(30)=>gen_18_cmp_pMux_30, f(29)=>
      gen_18_cmp_pMux_29, f(28)=>gen_18_cmp_pMux_28, f(27)=>
      gen_18_cmp_pMux_27, f(26)=>gen_18_cmp_pMux_26, f(25)=>
      gen_18_cmp_pMux_25, f(24)=>gen_18_cmp_pMux_24, f(23)=>
      gen_18_cmp_pMux_23, f(22)=>gen_18_cmp_pMux_22, f(21)=>
      gen_18_cmp_pMux_21, f(20)=>gen_18_cmp_pMux_20, f(19)=>
      gen_18_cmp_pMux_19, f(18)=>gen_18_cmp_pMux_18, f(17)=>
      gen_18_cmp_pMux_17, f(16)=>gen_18_cmp_pMux_16, f(15)=>
      gen_18_cmp_pMux_15, f(14)=>gen_18_cmp_pMux_14, f(13)=>
      gen_18_cmp_pMux_13, f(12)=>gen_18_cmp_pMux_12, f(11)=>
      gen_18_cmp_pMux_11, f(10)=>gen_18_cmp_pMux_10, f(9)=>gen_18_cmp_pMux_9, 
      f(8)=>gen_18_cmp_pMux_8, f(7)=>gen_18_cmp_pMux_7, f(6)=>
      gen_18_cmp_pMux_6, f(5)=>gen_18_cmp_pMux_5, f(4)=>gen_18_cmp_pMux_4, 
      f(3)=>gen_18_cmp_pMux_3, f(2)=>gen_18_cmp_pMux_2, f(1)=>
      gen_18_cmp_pMux_1, f(0)=>gen_18_cmp_pMux_0);
   gen_18_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>working, a(22)
      =>working, a(21)=>gen_18_cmp_pMux_30, a(20)=>gen_18_cmp_pMux_29, a(19)
      =>gen_18_cmp_pMux_28, a(18)=>gen_18_cmp_pMux_27, a(17)=>
      gen_18_cmp_pMux_26, a(16)=>gen_18_cmp_pMux_25, a(15)=>
      gen_18_cmp_pMux_24, a(14)=>gen_18_cmp_pMux_23, a(13)=>
      gen_18_cmp_pMux_22, a(12)=>gen_18_cmp_pMux_21, a(11)=>
      gen_18_cmp_pMux_20, a(10)=>gen_18_cmp_pMux_19, a(9)=>
      gen_18_cmp_pMux_18, a(8)=>gen_18_cmp_pMux_17, a(7)=>gen_18_cmp_pMux_16, 
      a(6)=>gen_18_cmp_pMux_15, a(5)=>gen_18_cmp_pMux_14, a(4)=>
      gen_18_cmp_pMux_13, a(3)=>gen_18_cmp_pMux_12, a(2)=>gen_18_cmp_pMux_11, 
      a(1)=>gen_18_cmp_pMux_10, a(0)=>gen_18_cmp_pMux_9, b(23)=>nx9775, 
      b(22)=>nx9775, b(21)=>nx9773, b(20)=>nx9781, b(19)=>nx9779, b(18)=>
      nx9777, b(17)=>nx9775, b(16)=>nx9773, b(15)=>gen_18_cmp_BSCmp_op2_15, 
      b(14)=>gen_18_cmp_BSCmp_op2_14, b(13)=>gen_18_cmp_BSCmp_op2_13, b(12)
      =>gen_18_cmp_BSCmp_op2_12, b(11)=>gen_18_cmp_BSCmp_op2_11, b(10)=>
      gen_18_cmp_BSCmp_op2_10, b(9)=>gen_18_cmp_BSCmp_op2_9, b(8)=>
      gen_18_cmp_BSCmp_op2_8, b(7)=>gen_18_cmp_BSCmp_op2_7, b(6)=>
      gen_18_cmp_BSCmp_op2_6, b(5)=>gen_18_cmp_BSCmp_op2_5, b(4)=>
      gen_18_cmp_BSCmp_op2_4, b(3)=>gen_18_cmp_BSCmp_op2_3, b(2)=>
      gen_18_cmp_BSCmp_op2_2, b(1)=>gen_18_cmp_BSCmp_op2_1, b(0)=>
      gen_18_cmp_BSCmp_op2_0, carryIn=>gen_18_cmp_BSCmp_carryIn, sum(23)=>
      gen_18_cmp_pBs_30, sum(22)=>gen_18_cmp_pBs_29, sum(21)=>
      gen_18_cmp_pBs_28, sum(20)=>gen_18_cmp_pBs_27, sum(19)=>
      gen_18_cmp_pBs_26, sum(18)=>gen_18_cmp_pBs_25, sum(17)=>
      gen_18_cmp_pBs_24, sum(16)=>gen_18_cmp_pBs_23, sum(15)=>outputs_18_15, 
      sum(14)=>outputs_18_14, sum(13)=>outputs_18_13, sum(12)=>outputs_18_12, 
      sum(11)=>outputs_18_11, sum(10)=>outputs_18_10, sum(9)=>outputs_18_9, 
      sum(8)=>outputs_18_8, sum(7)=>outputs_18_7, sum(6)=>outputs_18_6, 
      sum(5)=>outputs_18_5, sum(4)=>outputs_18_4, sum(3)=>outputs_18_3, 
      sum(2)=>outputs_18_2, sum(1)=>outputs_18_1, sum(0)=>outputs_18_0, 
      carryOut=>DANGLING(34));
   gen_17_cmp_pRegCmp : Reg_33 port map ( D(32)=>working, D(31)=>working, 
      D(30)=>gen_17_cmp_pBs_30, D(29)=>gen_17_cmp_pBs_29, D(28)=>
      gen_17_cmp_pBs_28, D(27)=>gen_17_cmp_pBs_27, D(26)=>gen_17_cmp_pBs_26, 
      D(25)=>gen_17_cmp_pBs_25, D(24)=>gen_17_cmp_pBs_24, D(23)=>
      gen_17_cmp_pBs_23, D(22)=>outputs_17_15, D(21)=>outputs_17_14, D(20)=>
      outputs_17_13, D(19)=>outputs_17_12, D(18)=>outputs_17_11, D(17)=>
      outputs_17_10, D(16)=>outputs_17_9, D(15)=>outputs_17_8, D(14)=>
      outputs_17_7, D(13)=>outputs_17_6, D(12)=>outputs_17_5, D(11)=>
      outputs_17_4, D(10)=>outputs_17_3, D(9)=>outputs_17_2, D(8)=>
      outputs_17_1, D(7)=>outputs_17_0, D(6)=>gen_17_cmp_pMux_8, D(5)=>
      gen_17_cmp_pMux_7, D(4)=>gen_17_cmp_pMux_6, D(3)=>gen_17_cmp_pMux_5, 
      D(2)=>gen_17_cmp_pMux_4, D(1)=>gen_17_cmp_pMux_3, D(0)=>nx9483, en=>
      nx11163, clk=>nx9393, rst=>rst, Q(32)=>DANGLING(35), Q(31)=>DANGLING(
      36), Q(30)=>gen_17_cmp_pReg_30, Q(29)=>gen_17_cmp_pReg_29, Q(28)=>
      gen_17_cmp_pReg_28, Q(27)=>gen_17_cmp_pReg_27, Q(26)=>
      gen_17_cmp_pReg_26, Q(25)=>gen_17_cmp_pReg_25, Q(24)=>
      gen_17_cmp_pReg_24, Q(23)=>gen_17_cmp_pReg_23, Q(22)=>
      gen_17_cmp_pReg_22, Q(21)=>gen_17_cmp_pReg_21, Q(20)=>
      gen_17_cmp_pReg_20, Q(19)=>gen_17_cmp_pReg_19, Q(18)=>
      gen_17_cmp_pReg_18, Q(17)=>gen_17_cmp_pReg_17, Q(16)=>
      gen_17_cmp_pReg_16, Q(15)=>gen_17_cmp_pReg_15, Q(14)=>
      gen_17_cmp_pReg_14, Q(13)=>gen_17_cmp_pReg_13, Q(12)=>
      gen_17_cmp_pReg_12, Q(11)=>gen_17_cmp_pReg_11, Q(10)=>
      gen_17_cmp_pReg_10, Q(9)=>gen_17_cmp_pReg_9, Q(8)=>gen_17_cmp_pReg_8, 
      Q(7)=>gen_17_cmp_pReg_7, Q(6)=>gen_17_cmp_pReg_6, Q(5)=>
      gen_17_cmp_pReg_5, Q(4)=>gen_17_cmp_pReg_4, Q(3)=>gen_17_cmp_pReg_3, 
      Q(2)=>gen_17_cmp_pReg_2, Q(1)=>gen_17_cmp_pReg_1, Q(0)=>
      gen_17_cmp_pReg_0);
   gen_17_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>working, a(31)=>
      working, a(30)=>gen_17_cmp_pReg_30, a(29)=>gen_17_cmp_pReg_29, a(28)=>
      gen_17_cmp_pReg_28, a(27)=>gen_17_cmp_pReg_27, a(26)=>
      gen_17_cmp_pReg_26, a(25)=>gen_17_cmp_pReg_25, a(24)=>
      gen_17_cmp_pReg_24, a(23)=>gen_17_cmp_pReg_23, a(22)=>
      gen_17_cmp_pReg_22, a(21)=>gen_17_cmp_pReg_21, a(20)=>
      gen_17_cmp_pReg_20, a(19)=>gen_17_cmp_pReg_19, a(18)=>
      gen_17_cmp_pReg_18, a(17)=>gen_17_cmp_pReg_17, a(16)=>
      gen_17_cmp_pReg_16, a(15)=>gen_17_cmp_pReg_15, a(14)=>
      gen_17_cmp_pReg_14, a(13)=>gen_17_cmp_pReg_13, a(12)=>
      gen_17_cmp_pReg_12, a(11)=>gen_17_cmp_pReg_11, a(10)=>
      gen_17_cmp_pReg_10, a(9)=>gen_17_cmp_pReg_9, a(8)=>gen_17_cmp_pReg_8, 
      a(7)=>gen_17_cmp_pReg_7, a(6)=>gen_17_cmp_pReg_6, a(5)=>
      gen_17_cmp_pReg_5, a(4)=>gen_17_cmp_pReg_4, a(3)=>gen_17_cmp_pReg_3, 
      a(2)=>gen_17_cmp_pReg_2, a(1)=>gen_17_cmp_pReg_1, a(0)=>
      gen_17_cmp_pReg_0, b(32)=>working, b(31)=>working, b(30)=>working, 
      b(29)=>working, b(28)=>working, b(27)=>working, b(26)=>working, b(25)
      =>working, b(24)=>working, b(23)=>working, b(22)=>working, b(21)=>
      working, b(20)=>working, b(19)=>working, b(18)=>working, b(17)=>
      working, b(16)=>working, b(15)=>working, b(14)=>working, b(13)=>
      working, b(12)=>working, b(11)=>working, b(10)=>working, b(9)=>working, 
      b(8)=>filter_17_7, b(7)=>filter_17_6, b(6)=>filter_17_5, b(5)=>
      filter_17_4, b(4)=>filter_17_3, b(3)=>filter_17_2, b(2)=>filter_17_1, 
      b(1)=>filter_17_0, b(0)=>working, sel=>nx11179, f(32)=>DANGLING(37), 
      f(31)=>DANGLING(38), f(30)=>gen_17_cmp_pMux_30, f(29)=>
      gen_17_cmp_pMux_29, f(28)=>gen_17_cmp_pMux_28, f(27)=>
      gen_17_cmp_pMux_27, f(26)=>gen_17_cmp_pMux_26, f(25)=>
      gen_17_cmp_pMux_25, f(24)=>gen_17_cmp_pMux_24, f(23)=>
      gen_17_cmp_pMux_23, f(22)=>gen_17_cmp_pMux_22, f(21)=>
      gen_17_cmp_pMux_21, f(20)=>gen_17_cmp_pMux_20, f(19)=>
      gen_17_cmp_pMux_19, f(18)=>gen_17_cmp_pMux_18, f(17)=>
      gen_17_cmp_pMux_17, f(16)=>gen_17_cmp_pMux_16, f(15)=>
      gen_17_cmp_pMux_15, f(14)=>gen_17_cmp_pMux_14, f(13)=>
      gen_17_cmp_pMux_13, f(12)=>gen_17_cmp_pMux_12, f(11)=>
      gen_17_cmp_pMux_11, f(10)=>gen_17_cmp_pMux_10, f(9)=>gen_17_cmp_pMux_9, 
      f(8)=>gen_17_cmp_pMux_8, f(7)=>gen_17_cmp_pMux_7, f(6)=>
      gen_17_cmp_pMux_6, f(5)=>gen_17_cmp_pMux_5, f(4)=>gen_17_cmp_pMux_4, 
      f(3)=>gen_17_cmp_pMux_3, f(2)=>gen_17_cmp_pMux_2, f(1)=>
      gen_17_cmp_pMux_1, f(0)=>gen_17_cmp_pMux_0);
   gen_17_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>working, a(22)
      =>working, a(21)=>gen_17_cmp_pMux_30, a(20)=>gen_17_cmp_pMux_29, a(19)
      =>gen_17_cmp_pMux_28, a(18)=>gen_17_cmp_pMux_27, a(17)=>
      gen_17_cmp_pMux_26, a(16)=>gen_17_cmp_pMux_25, a(15)=>
      gen_17_cmp_pMux_24, a(14)=>gen_17_cmp_pMux_23, a(13)=>
      gen_17_cmp_pMux_22, a(12)=>gen_17_cmp_pMux_21, a(11)=>
      gen_17_cmp_pMux_20, a(10)=>gen_17_cmp_pMux_19, a(9)=>
      gen_17_cmp_pMux_18, a(8)=>gen_17_cmp_pMux_17, a(7)=>gen_17_cmp_pMux_16, 
      a(6)=>gen_17_cmp_pMux_15, a(5)=>gen_17_cmp_pMux_14, a(4)=>
      gen_17_cmp_pMux_13, a(3)=>gen_17_cmp_pMux_12, a(2)=>gen_17_cmp_pMux_11, 
      a(1)=>gen_17_cmp_pMux_10, a(0)=>gen_17_cmp_pMux_9, b(23)=>nx9787, 
      b(22)=>nx9787, b(21)=>nx9785, b(20)=>nx9793, b(19)=>nx9791, b(18)=>
      nx9789, b(17)=>nx9787, b(16)=>nx9785, b(15)=>gen_17_cmp_BSCmp_op2_15, 
      b(14)=>gen_17_cmp_BSCmp_op2_14, b(13)=>gen_17_cmp_BSCmp_op2_13, b(12)
      =>gen_17_cmp_BSCmp_op2_12, b(11)=>gen_17_cmp_BSCmp_op2_11, b(10)=>
      gen_17_cmp_BSCmp_op2_10, b(9)=>gen_17_cmp_BSCmp_op2_9, b(8)=>
      gen_17_cmp_BSCmp_op2_8, b(7)=>gen_17_cmp_BSCmp_op2_7, b(6)=>
      gen_17_cmp_BSCmp_op2_6, b(5)=>gen_17_cmp_BSCmp_op2_5, b(4)=>
      gen_17_cmp_BSCmp_op2_4, b(3)=>gen_17_cmp_BSCmp_op2_3, b(2)=>
      gen_17_cmp_BSCmp_op2_2, b(1)=>gen_17_cmp_BSCmp_op2_1, b(0)=>
      gen_17_cmp_BSCmp_op2_0, carryIn=>gen_17_cmp_BSCmp_carryIn, sum(23)=>
      gen_17_cmp_pBs_30, sum(22)=>gen_17_cmp_pBs_29, sum(21)=>
      gen_17_cmp_pBs_28, sum(20)=>gen_17_cmp_pBs_27, sum(19)=>
      gen_17_cmp_pBs_26, sum(18)=>gen_17_cmp_pBs_25, sum(17)=>
      gen_17_cmp_pBs_24, sum(16)=>gen_17_cmp_pBs_23, sum(15)=>outputs_17_15, 
      sum(14)=>outputs_17_14, sum(13)=>outputs_17_13, sum(12)=>outputs_17_12, 
      sum(11)=>outputs_17_11, sum(10)=>outputs_17_10, sum(9)=>outputs_17_9, 
      sum(8)=>outputs_17_8, sum(7)=>outputs_17_7, sum(6)=>outputs_17_6, 
      sum(5)=>outputs_17_5, sum(4)=>outputs_17_4, sum(3)=>outputs_17_3, 
      sum(2)=>outputs_17_2, sum(1)=>outputs_17_1, sum(0)=>outputs_17_0, 
      carryOut=>DANGLING(39));
   gen_16_cmp_pRegCmp : Reg_33 port map ( D(32)=>working, D(31)=>working, 
      D(30)=>gen_16_cmp_pBs_30, D(29)=>gen_16_cmp_pBs_29, D(28)=>
      gen_16_cmp_pBs_28, D(27)=>gen_16_cmp_pBs_27, D(26)=>gen_16_cmp_pBs_26, 
      D(25)=>gen_16_cmp_pBs_25, D(24)=>gen_16_cmp_pBs_24, D(23)=>
      gen_16_cmp_pBs_23, D(22)=>outputs_16_15, D(21)=>outputs_16_14, D(20)=>
      outputs_16_13, D(19)=>outputs_16_12, D(18)=>outputs_16_11, D(17)=>
      outputs_16_10, D(16)=>outputs_16_9, D(15)=>outputs_16_8, D(14)=>
      outputs_16_7, D(13)=>outputs_16_6, D(12)=>outputs_16_5, D(11)=>
      outputs_16_4, D(10)=>outputs_16_3, D(9)=>outputs_16_2, D(8)=>
      outputs_16_1, D(7)=>outputs_16_0, D(6)=>gen_16_cmp_pMux_8, D(5)=>
      gen_16_cmp_pMux_7, D(4)=>gen_16_cmp_pMux_6, D(3)=>gen_16_cmp_pMux_5, 
      D(2)=>gen_16_cmp_pMux_4, D(1)=>gen_16_cmp_pMux_3, D(0)=>nx9495, en=>
      nx11163, clk=>nx9393, rst=>rst, Q(32)=>DANGLING(40), Q(31)=>DANGLING(
      41), Q(30)=>gen_16_cmp_pReg_30, Q(29)=>gen_16_cmp_pReg_29, Q(28)=>
      gen_16_cmp_pReg_28, Q(27)=>gen_16_cmp_pReg_27, Q(26)=>
      gen_16_cmp_pReg_26, Q(25)=>gen_16_cmp_pReg_25, Q(24)=>
      gen_16_cmp_pReg_24, Q(23)=>gen_16_cmp_pReg_23, Q(22)=>
      gen_16_cmp_pReg_22, Q(21)=>gen_16_cmp_pReg_21, Q(20)=>
      gen_16_cmp_pReg_20, Q(19)=>gen_16_cmp_pReg_19, Q(18)=>
      gen_16_cmp_pReg_18, Q(17)=>gen_16_cmp_pReg_17, Q(16)=>
      gen_16_cmp_pReg_16, Q(15)=>gen_16_cmp_pReg_15, Q(14)=>
      gen_16_cmp_pReg_14, Q(13)=>gen_16_cmp_pReg_13, Q(12)=>
      gen_16_cmp_pReg_12, Q(11)=>gen_16_cmp_pReg_11, Q(10)=>
      gen_16_cmp_pReg_10, Q(9)=>gen_16_cmp_pReg_9, Q(8)=>gen_16_cmp_pReg_8, 
      Q(7)=>gen_16_cmp_pReg_7, Q(6)=>gen_16_cmp_pReg_6, Q(5)=>
      gen_16_cmp_pReg_5, Q(4)=>gen_16_cmp_pReg_4, Q(3)=>gen_16_cmp_pReg_3, 
      Q(2)=>gen_16_cmp_pReg_2, Q(1)=>gen_16_cmp_pReg_1, Q(0)=>
      gen_16_cmp_pReg_0);
   gen_16_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>working, a(31)=>
      working, a(30)=>gen_16_cmp_pReg_30, a(29)=>gen_16_cmp_pReg_29, a(28)=>
      gen_16_cmp_pReg_28, a(27)=>gen_16_cmp_pReg_27, a(26)=>
      gen_16_cmp_pReg_26, a(25)=>gen_16_cmp_pReg_25, a(24)=>
      gen_16_cmp_pReg_24, a(23)=>gen_16_cmp_pReg_23, a(22)=>
      gen_16_cmp_pReg_22, a(21)=>gen_16_cmp_pReg_21, a(20)=>
      gen_16_cmp_pReg_20, a(19)=>gen_16_cmp_pReg_19, a(18)=>
      gen_16_cmp_pReg_18, a(17)=>gen_16_cmp_pReg_17, a(16)=>
      gen_16_cmp_pReg_16, a(15)=>gen_16_cmp_pReg_15, a(14)=>
      gen_16_cmp_pReg_14, a(13)=>gen_16_cmp_pReg_13, a(12)=>
      gen_16_cmp_pReg_12, a(11)=>gen_16_cmp_pReg_11, a(10)=>
      gen_16_cmp_pReg_10, a(9)=>gen_16_cmp_pReg_9, a(8)=>gen_16_cmp_pReg_8, 
      a(7)=>gen_16_cmp_pReg_7, a(6)=>gen_16_cmp_pReg_6, a(5)=>
      gen_16_cmp_pReg_5, a(4)=>gen_16_cmp_pReg_4, a(3)=>gen_16_cmp_pReg_3, 
      a(2)=>gen_16_cmp_pReg_2, a(1)=>gen_16_cmp_pReg_1, a(0)=>
      gen_16_cmp_pReg_0, b(32)=>working, b(31)=>working, b(30)=>working, 
      b(29)=>working, b(28)=>working, b(27)=>working, b(26)=>working, b(25)
      =>working, b(24)=>working, b(23)=>working, b(22)=>working, b(21)=>
      working, b(20)=>working, b(19)=>working, b(18)=>working, b(17)=>
      working, b(16)=>working, b(15)=>working, b(14)=>working, b(13)=>
      working, b(12)=>working, b(11)=>working, b(10)=>working, b(9)=>working, 
      b(8)=>filter_16_7, b(7)=>filter_16_6, b(6)=>filter_16_5, b(5)=>
      filter_16_4, b(4)=>filter_16_3, b(3)=>filter_16_2, b(2)=>filter_16_1, 
      b(1)=>filter_16_0, b(0)=>working, sel=>nx11179, f(32)=>DANGLING(42), 
      f(31)=>DANGLING(43), f(30)=>gen_16_cmp_pMux_30, f(29)=>
      gen_16_cmp_pMux_29, f(28)=>gen_16_cmp_pMux_28, f(27)=>
      gen_16_cmp_pMux_27, f(26)=>gen_16_cmp_pMux_26, f(25)=>
      gen_16_cmp_pMux_25, f(24)=>gen_16_cmp_pMux_24, f(23)=>
      gen_16_cmp_pMux_23, f(22)=>gen_16_cmp_pMux_22, f(21)=>
      gen_16_cmp_pMux_21, f(20)=>gen_16_cmp_pMux_20, f(19)=>
      gen_16_cmp_pMux_19, f(18)=>gen_16_cmp_pMux_18, f(17)=>
      gen_16_cmp_pMux_17, f(16)=>gen_16_cmp_pMux_16, f(15)=>
      gen_16_cmp_pMux_15, f(14)=>gen_16_cmp_pMux_14, f(13)=>
      gen_16_cmp_pMux_13, f(12)=>gen_16_cmp_pMux_12, f(11)=>
      gen_16_cmp_pMux_11, f(10)=>gen_16_cmp_pMux_10, f(9)=>gen_16_cmp_pMux_9, 
      f(8)=>gen_16_cmp_pMux_8, f(7)=>gen_16_cmp_pMux_7, f(6)=>
      gen_16_cmp_pMux_6, f(5)=>gen_16_cmp_pMux_5, f(4)=>gen_16_cmp_pMux_4, 
      f(3)=>gen_16_cmp_pMux_3, f(2)=>gen_16_cmp_pMux_2, f(1)=>
      gen_16_cmp_pMux_1, f(0)=>gen_16_cmp_pMux_0);
   gen_16_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>working, a(22)
      =>working, a(21)=>gen_16_cmp_pMux_30, a(20)=>gen_16_cmp_pMux_29, a(19)
      =>gen_16_cmp_pMux_28, a(18)=>gen_16_cmp_pMux_27, a(17)=>
      gen_16_cmp_pMux_26, a(16)=>gen_16_cmp_pMux_25, a(15)=>
      gen_16_cmp_pMux_24, a(14)=>gen_16_cmp_pMux_23, a(13)=>
      gen_16_cmp_pMux_22, a(12)=>gen_16_cmp_pMux_21, a(11)=>
      gen_16_cmp_pMux_20, a(10)=>gen_16_cmp_pMux_19, a(9)=>
      gen_16_cmp_pMux_18, a(8)=>gen_16_cmp_pMux_17, a(7)=>gen_16_cmp_pMux_16, 
      a(6)=>gen_16_cmp_pMux_15, a(5)=>gen_16_cmp_pMux_14, a(4)=>
      gen_16_cmp_pMux_13, a(3)=>gen_16_cmp_pMux_12, a(2)=>gen_16_cmp_pMux_11, 
      a(1)=>gen_16_cmp_pMux_10, a(0)=>gen_16_cmp_pMux_9, b(23)=>nx9799, 
      b(22)=>nx9799, b(21)=>nx9797, b(20)=>nx9805, b(19)=>nx9803, b(18)=>
      nx9801, b(17)=>nx9799, b(16)=>nx9797, b(15)=>gen_16_cmp_BSCmp_op2_15, 
      b(14)=>gen_16_cmp_BSCmp_op2_14, b(13)=>gen_16_cmp_BSCmp_op2_13, b(12)
      =>gen_16_cmp_BSCmp_op2_12, b(11)=>gen_16_cmp_BSCmp_op2_11, b(10)=>
      gen_16_cmp_BSCmp_op2_10, b(9)=>gen_16_cmp_BSCmp_op2_9, b(8)=>
      gen_16_cmp_BSCmp_op2_8, b(7)=>gen_16_cmp_BSCmp_op2_7, b(6)=>
      gen_16_cmp_BSCmp_op2_6, b(5)=>gen_16_cmp_BSCmp_op2_5, b(4)=>
      gen_16_cmp_BSCmp_op2_4, b(3)=>gen_16_cmp_BSCmp_op2_3, b(2)=>
      gen_16_cmp_BSCmp_op2_2, b(1)=>gen_16_cmp_BSCmp_op2_1, b(0)=>
      gen_16_cmp_BSCmp_op2_0, carryIn=>gen_16_cmp_BSCmp_carryIn, sum(23)=>
      gen_16_cmp_pBs_30, sum(22)=>gen_16_cmp_pBs_29, sum(21)=>
      gen_16_cmp_pBs_28, sum(20)=>gen_16_cmp_pBs_27, sum(19)=>
      gen_16_cmp_pBs_26, sum(18)=>gen_16_cmp_pBs_25, sum(17)=>
      gen_16_cmp_pBs_24, sum(16)=>gen_16_cmp_pBs_23, sum(15)=>outputs_16_15, 
      sum(14)=>outputs_16_14, sum(13)=>outputs_16_13, sum(12)=>outputs_16_12, 
      sum(11)=>outputs_16_11, sum(10)=>outputs_16_10, sum(9)=>outputs_16_9, 
      sum(8)=>outputs_16_8, sum(7)=>outputs_16_7, sum(6)=>outputs_16_6, 
      sum(5)=>outputs_16_5, sum(4)=>outputs_16_4, sum(3)=>outputs_16_3, 
      sum(2)=>outputs_16_2, sum(1)=>outputs_16_1, sum(0)=>outputs_16_0, 
      carryOut=>DANGLING(44));
   gen_15_cmp_pRegCmp : Reg_33 port map ( D(32)=>working, D(31)=>working, 
      D(30)=>gen_15_cmp_pBs_30, D(29)=>gen_15_cmp_pBs_29, D(28)=>
      gen_15_cmp_pBs_28, D(27)=>gen_15_cmp_pBs_27, D(26)=>gen_15_cmp_pBs_26, 
      D(25)=>gen_15_cmp_pBs_25, D(24)=>gen_15_cmp_pBs_24, D(23)=>
      gen_15_cmp_pBs_23, D(22)=>outputs_15_15, D(21)=>outputs_15_14, D(20)=>
      outputs_15_13, D(19)=>outputs_15_12, D(18)=>outputs_15_11, D(17)=>
      outputs_15_10, D(16)=>outputs_15_9, D(15)=>outputs_15_8, D(14)=>
      outputs_15_7, D(13)=>outputs_15_6, D(12)=>outputs_15_5, D(11)=>
      outputs_15_4, D(10)=>outputs_15_3, D(9)=>outputs_15_2, D(8)=>
      outputs_15_1, D(7)=>outputs_15_0, D(6)=>gen_15_cmp_pMux_8, D(5)=>
      gen_15_cmp_pMux_7, D(4)=>gen_15_cmp_pMux_6, D(3)=>gen_15_cmp_pMux_5, 
      D(2)=>gen_15_cmp_pMux_4, D(1)=>gen_15_cmp_pMux_3, D(0)=>nx9507, en=>
      nx11163, clk=>nx9393, rst=>rst, Q(32)=>DANGLING(45), Q(31)=>DANGLING(
      46), Q(30)=>gen_15_cmp_pReg_30, Q(29)=>gen_15_cmp_pReg_29, Q(28)=>
      gen_15_cmp_pReg_28, Q(27)=>gen_15_cmp_pReg_27, Q(26)=>
      gen_15_cmp_pReg_26, Q(25)=>gen_15_cmp_pReg_25, Q(24)=>
      gen_15_cmp_pReg_24, Q(23)=>gen_15_cmp_pReg_23, Q(22)=>
      gen_15_cmp_pReg_22, Q(21)=>gen_15_cmp_pReg_21, Q(20)=>
      gen_15_cmp_pReg_20, Q(19)=>gen_15_cmp_pReg_19, Q(18)=>
      gen_15_cmp_pReg_18, Q(17)=>gen_15_cmp_pReg_17, Q(16)=>
      gen_15_cmp_pReg_16, Q(15)=>gen_15_cmp_pReg_15, Q(14)=>
      gen_15_cmp_pReg_14, Q(13)=>gen_15_cmp_pReg_13, Q(12)=>
      gen_15_cmp_pReg_12, Q(11)=>gen_15_cmp_pReg_11, Q(10)=>
      gen_15_cmp_pReg_10, Q(9)=>gen_15_cmp_pReg_9, Q(8)=>gen_15_cmp_pReg_8, 
      Q(7)=>gen_15_cmp_pReg_7, Q(6)=>gen_15_cmp_pReg_6, Q(5)=>
      gen_15_cmp_pReg_5, Q(4)=>gen_15_cmp_pReg_4, Q(3)=>gen_15_cmp_pReg_3, 
      Q(2)=>gen_15_cmp_pReg_2, Q(1)=>gen_15_cmp_pReg_1, Q(0)=>
      gen_15_cmp_pReg_0);
   gen_15_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>working, a(31)=>
      working, a(30)=>gen_15_cmp_pReg_30, a(29)=>gen_15_cmp_pReg_29, a(28)=>
      gen_15_cmp_pReg_28, a(27)=>gen_15_cmp_pReg_27, a(26)=>
      gen_15_cmp_pReg_26, a(25)=>gen_15_cmp_pReg_25, a(24)=>
      gen_15_cmp_pReg_24, a(23)=>gen_15_cmp_pReg_23, a(22)=>
      gen_15_cmp_pReg_22, a(21)=>gen_15_cmp_pReg_21, a(20)=>
      gen_15_cmp_pReg_20, a(19)=>gen_15_cmp_pReg_19, a(18)=>
      gen_15_cmp_pReg_18, a(17)=>gen_15_cmp_pReg_17, a(16)=>
      gen_15_cmp_pReg_16, a(15)=>gen_15_cmp_pReg_15, a(14)=>
      gen_15_cmp_pReg_14, a(13)=>gen_15_cmp_pReg_13, a(12)=>
      gen_15_cmp_pReg_12, a(11)=>gen_15_cmp_pReg_11, a(10)=>
      gen_15_cmp_pReg_10, a(9)=>gen_15_cmp_pReg_9, a(8)=>gen_15_cmp_pReg_8, 
      a(7)=>gen_15_cmp_pReg_7, a(6)=>gen_15_cmp_pReg_6, a(5)=>
      gen_15_cmp_pReg_5, a(4)=>gen_15_cmp_pReg_4, a(3)=>gen_15_cmp_pReg_3, 
      a(2)=>gen_15_cmp_pReg_2, a(1)=>gen_15_cmp_pReg_1, a(0)=>
      gen_15_cmp_pReg_0, b(32)=>working, b(31)=>working, b(30)=>working, 
      b(29)=>working, b(28)=>working, b(27)=>working, b(26)=>working, b(25)
      =>working, b(24)=>working, b(23)=>working, b(22)=>working, b(21)=>
      working, b(20)=>working, b(19)=>working, b(18)=>working, b(17)=>
      working, b(16)=>working, b(15)=>working, b(14)=>working, b(13)=>
      working, b(12)=>working, b(11)=>working, b(10)=>working, b(9)=>working, 
      b(8)=>filter_15_7, b(7)=>filter_15_6, b(6)=>filter_15_5, b(5)=>
      filter_15_4, b(4)=>filter_15_3, b(3)=>filter_15_2, b(2)=>filter_15_1, 
      b(1)=>filter_15_0, b(0)=>working, sel=>nx11179, f(32)=>DANGLING(47), 
      f(31)=>DANGLING(48), f(30)=>gen_15_cmp_pMux_30, f(29)=>
      gen_15_cmp_pMux_29, f(28)=>gen_15_cmp_pMux_28, f(27)=>
      gen_15_cmp_pMux_27, f(26)=>gen_15_cmp_pMux_26, f(25)=>
      gen_15_cmp_pMux_25, f(24)=>gen_15_cmp_pMux_24, f(23)=>
      gen_15_cmp_pMux_23, f(22)=>gen_15_cmp_pMux_22, f(21)=>
      gen_15_cmp_pMux_21, f(20)=>gen_15_cmp_pMux_20, f(19)=>
      gen_15_cmp_pMux_19, f(18)=>gen_15_cmp_pMux_18, f(17)=>
      gen_15_cmp_pMux_17, f(16)=>gen_15_cmp_pMux_16, f(15)=>
      gen_15_cmp_pMux_15, f(14)=>gen_15_cmp_pMux_14, f(13)=>
      gen_15_cmp_pMux_13, f(12)=>gen_15_cmp_pMux_12, f(11)=>
      gen_15_cmp_pMux_11, f(10)=>gen_15_cmp_pMux_10, f(9)=>gen_15_cmp_pMux_9, 
      f(8)=>gen_15_cmp_pMux_8, f(7)=>gen_15_cmp_pMux_7, f(6)=>
      gen_15_cmp_pMux_6, f(5)=>gen_15_cmp_pMux_5, f(4)=>gen_15_cmp_pMux_4, 
      f(3)=>gen_15_cmp_pMux_3, f(2)=>gen_15_cmp_pMux_2, f(1)=>
      gen_15_cmp_pMux_1, f(0)=>gen_15_cmp_pMux_0);
   gen_15_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>working, a(22)
      =>working, a(21)=>gen_15_cmp_pMux_30, a(20)=>gen_15_cmp_pMux_29, a(19)
      =>gen_15_cmp_pMux_28, a(18)=>gen_15_cmp_pMux_27, a(17)=>
      gen_15_cmp_pMux_26, a(16)=>gen_15_cmp_pMux_25, a(15)=>
      gen_15_cmp_pMux_24, a(14)=>gen_15_cmp_pMux_23, a(13)=>
      gen_15_cmp_pMux_22, a(12)=>gen_15_cmp_pMux_21, a(11)=>
      gen_15_cmp_pMux_20, a(10)=>gen_15_cmp_pMux_19, a(9)=>
      gen_15_cmp_pMux_18, a(8)=>gen_15_cmp_pMux_17, a(7)=>gen_15_cmp_pMux_16, 
      a(6)=>gen_15_cmp_pMux_15, a(5)=>gen_15_cmp_pMux_14, a(4)=>
      gen_15_cmp_pMux_13, a(3)=>gen_15_cmp_pMux_12, a(2)=>gen_15_cmp_pMux_11, 
      a(1)=>gen_15_cmp_pMux_10, a(0)=>gen_15_cmp_pMux_9, b(23)=>nx9811, 
      b(22)=>nx9811, b(21)=>nx9809, b(20)=>nx9817, b(19)=>nx9815, b(18)=>
      nx9813, b(17)=>nx9811, b(16)=>nx9809, b(15)=>gen_15_cmp_BSCmp_op2_15, 
      b(14)=>gen_15_cmp_BSCmp_op2_14, b(13)=>gen_15_cmp_BSCmp_op2_13, b(12)
      =>gen_15_cmp_BSCmp_op2_12, b(11)=>gen_15_cmp_BSCmp_op2_11, b(10)=>
      gen_15_cmp_BSCmp_op2_10, b(9)=>gen_15_cmp_BSCmp_op2_9, b(8)=>
      gen_15_cmp_BSCmp_op2_8, b(7)=>gen_15_cmp_BSCmp_op2_7, b(6)=>
      gen_15_cmp_BSCmp_op2_6, b(5)=>gen_15_cmp_BSCmp_op2_5, b(4)=>
      gen_15_cmp_BSCmp_op2_4, b(3)=>gen_15_cmp_BSCmp_op2_3, b(2)=>
      gen_15_cmp_BSCmp_op2_2, b(1)=>gen_15_cmp_BSCmp_op2_1, b(0)=>
      gen_15_cmp_BSCmp_op2_0, carryIn=>gen_15_cmp_BSCmp_carryIn, sum(23)=>
      gen_15_cmp_pBs_30, sum(22)=>gen_15_cmp_pBs_29, sum(21)=>
      gen_15_cmp_pBs_28, sum(20)=>gen_15_cmp_pBs_27, sum(19)=>
      gen_15_cmp_pBs_26, sum(18)=>gen_15_cmp_pBs_25, sum(17)=>
      gen_15_cmp_pBs_24, sum(16)=>gen_15_cmp_pBs_23, sum(15)=>outputs_15_15, 
      sum(14)=>outputs_15_14, sum(13)=>outputs_15_13, sum(12)=>outputs_15_12, 
      sum(11)=>outputs_15_11, sum(10)=>outputs_15_10, sum(9)=>outputs_15_9, 
      sum(8)=>outputs_15_8, sum(7)=>outputs_15_7, sum(6)=>outputs_15_6, 
      sum(5)=>outputs_15_5, sum(4)=>outputs_15_4, sum(3)=>outputs_15_3, 
      sum(2)=>outputs_15_2, sum(1)=>outputs_15_1, sum(0)=>outputs_15_0, 
      carryOut=>DANGLING(49));
   gen_14_cmp_pRegCmp : Reg_33 port map ( D(32)=>working, D(31)=>working, 
      D(30)=>gen_14_cmp_pBs_30, D(29)=>gen_14_cmp_pBs_29, D(28)=>
      gen_14_cmp_pBs_28, D(27)=>gen_14_cmp_pBs_27, D(26)=>gen_14_cmp_pBs_26, 
      D(25)=>gen_14_cmp_pBs_25, D(24)=>gen_14_cmp_pBs_24, D(23)=>
      gen_14_cmp_pBs_23, D(22)=>outputs_14_15, D(21)=>outputs_14_14, D(20)=>
      outputs_14_13, D(19)=>outputs_14_12, D(18)=>outputs_14_11, D(17)=>
      outputs_14_10, D(16)=>outputs_14_9, D(15)=>outputs_14_8, D(14)=>
      outputs_14_7, D(13)=>outputs_14_6, D(12)=>outputs_14_5, D(11)=>
      outputs_14_4, D(10)=>outputs_14_3, D(9)=>outputs_14_2, D(8)=>
      outputs_14_1, D(7)=>outputs_14_0, D(6)=>gen_14_cmp_pMux_8, D(5)=>
      gen_14_cmp_pMux_7, D(4)=>gen_14_cmp_pMux_6, D(3)=>gen_14_cmp_pMux_5, 
      D(2)=>gen_14_cmp_pMux_4, D(1)=>gen_14_cmp_pMux_3, D(0)=>nx9519, en=>
      nx11165, clk=>nx9393, rst=>rst, Q(32)=>DANGLING(50), Q(31)=>DANGLING(
      51), Q(30)=>gen_14_cmp_pReg_30, Q(29)=>gen_14_cmp_pReg_29, Q(28)=>
      gen_14_cmp_pReg_28, Q(27)=>gen_14_cmp_pReg_27, Q(26)=>
      gen_14_cmp_pReg_26, Q(25)=>gen_14_cmp_pReg_25, Q(24)=>
      gen_14_cmp_pReg_24, Q(23)=>gen_14_cmp_pReg_23, Q(22)=>
      gen_14_cmp_pReg_22, Q(21)=>gen_14_cmp_pReg_21, Q(20)=>
      gen_14_cmp_pReg_20, Q(19)=>gen_14_cmp_pReg_19, Q(18)=>
      gen_14_cmp_pReg_18, Q(17)=>gen_14_cmp_pReg_17, Q(16)=>
      gen_14_cmp_pReg_16, Q(15)=>gen_14_cmp_pReg_15, Q(14)=>
      gen_14_cmp_pReg_14, Q(13)=>gen_14_cmp_pReg_13, Q(12)=>
      gen_14_cmp_pReg_12, Q(11)=>gen_14_cmp_pReg_11, Q(10)=>
      gen_14_cmp_pReg_10, Q(9)=>gen_14_cmp_pReg_9, Q(8)=>gen_14_cmp_pReg_8, 
      Q(7)=>gen_14_cmp_pReg_7, Q(6)=>gen_14_cmp_pReg_6, Q(5)=>
      gen_14_cmp_pReg_5, Q(4)=>gen_14_cmp_pReg_4, Q(3)=>gen_14_cmp_pReg_3, 
      Q(2)=>gen_14_cmp_pReg_2, Q(1)=>gen_14_cmp_pReg_1, Q(0)=>
      gen_14_cmp_pReg_0);
   gen_14_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>working, a(31)=>
      working, a(30)=>gen_14_cmp_pReg_30, a(29)=>gen_14_cmp_pReg_29, a(28)=>
      gen_14_cmp_pReg_28, a(27)=>gen_14_cmp_pReg_27, a(26)=>
      gen_14_cmp_pReg_26, a(25)=>gen_14_cmp_pReg_25, a(24)=>
      gen_14_cmp_pReg_24, a(23)=>gen_14_cmp_pReg_23, a(22)=>
      gen_14_cmp_pReg_22, a(21)=>gen_14_cmp_pReg_21, a(20)=>
      gen_14_cmp_pReg_20, a(19)=>gen_14_cmp_pReg_19, a(18)=>
      gen_14_cmp_pReg_18, a(17)=>gen_14_cmp_pReg_17, a(16)=>
      gen_14_cmp_pReg_16, a(15)=>gen_14_cmp_pReg_15, a(14)=>
      gen_14_cmp_pReg_14, a(13)=>gen_14_cmp_pReg_13, a(12)=>
      gen_14_cmp_pReg_12, a(11)=>gen_14_cmp_pReg_11, a(10)=>
      gen_14_cmp_pReg_10, a(9)=>gen_14_cmp_pReg_9, a(8)=>gen_14_cmp_pReg_8, 
      a(7)=>gen_14_cmp_pReg_7, a(6)=>gen_14_cmp_pReg_6, a(5)=>
      gen_14_cmp_pReg_5, a(4)=>gen_14_cmp_pReg_4, a(3)=>gen_14_cmp_pReg_3, 
      a(2)=>gen_14_cmp_pReg_2, a(1)=>gen_14_cmp_pReg_1, a(0)=>
      gen_14_cmp_pReg_0, b(32)=>working, b(31)=>working, b(30)=>working, 
      b(29)=>working, b(28)=>working, b(27)=>working, b(26)=>working, b(25)
      =>working, b(24)=>working, b(23)=>working, b(22)=>working, b(21)=>
      working, b(20)=>working, b(19)=>working, b(18)=>working, b(17)=>
      working, b(16)=>working, b(15)=>working, b(14)=>working, b(13)=>
      working, b(12)=>working, b(11)=>working, b(10)=>working, b(9)=>working, 
      b(8)=>filter_14_7, b(7)=>filter_14_6, b(6)=>filter_14_5, b(5)=>
      filter_14_4, b(4)=>filter_14_3, b(3)=>filter_14_2, b(2)=>filter_14_1, 
      b(1)=>filter_14_0, b(0)=>working, sel=>nx11181, f(32)=>DANGLING(52), 
      f(31)=>DANGLING(53), f(30)=>gen_14_cmp_pMux_30, f(29)=>
      gen_14_cmp_pMux_29, f(28)=>gen_14_cmp_pMux_28, f(27)=>
      gen_14_cmp_pMux_27, f(26)=>gen_14_cmp_pMux_26, f(25)=>
      gen_14_cmp_pMux_25, f(24)=>gen_14_cmp_pMux_24, f(23)=>
      gen_14_cmp_pMux_23, f(22)=>gen_14_cmp_pMux_22, f(21)=>
      gen_14_cmp_pMux_21, f(20)=>gen_14_cmp_pMux_20, f(19)=>
      gen_14_cmp_pMux_19, f(18)=>gen_14_cmp_pMux_18, f(17)=>
      gen_14_cmp_pMux_17, f(16)=>gen_14_cmp_pMux_16, f(15)=>
      gen_14_cmp_pMux_15, f(14)=>gen_14_cmp_pMux_14, f(13)=>
      gen_14_cmp_pMux_13, f(12)=>gen_14_cmp_pMux_12, f(11)=>
      gen_14_cmp_pMux_11, f(10)=>gen_14_cmp_pMux_10, f(9)=>gen_14_cmp_pMux_9, 
      f(8)=>gen_14_cmp_pMux_8, f(7)=>gen_14_cmp_pMux_7, f(6)=>
      gen_14_cmp_pMux_6, f(5)=>gen_14_cmp_pMux_5, f(4)=>gen_14_cmp_pMux_4, 
      f(3)=>gen_14_cmp_pMux_3, f(2)=>gen_14_cmp_pMux_2, f(1)=>
      gen_14_cmp_pMux_1, f(0)=>gen_14_cmp_pMux_0);
   gen_14_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>working, a(22)
      =>working, a(21)=>gen_14_cmp_pMux_30, a(20)=>gen_14_cmp_pMux_29, a(19)
      =>gen_14_cmp_pMux_28, a(18)=>gen_14_cmp_pMux_27, a(17)=>
      gen_14_cmp_pMux_26, a(16)=>gen_14_cmp_pMux_25, a(15)=>
      gen_14_cmp_pMux_24, a(14)=>gen_14_cmp_pMux_23, a(13)=>
      gen_14_cmp_pMux_22, a(12)=>gen_14_cmp_pMux_21, a(11)=>
      gen_14_cmp_pMux_20, a(10)=>gen_14_cmp_pMux_19, a(9)=>
      gen_14_cmp_pMux_18, a(8)=>gen_14_cmp_pMux_17, a(7)=>gen_14_cmp_pMux_16, 
      a(6)=>gen_14_cmp_pMux_15, a(5)=>gen_14_cmp_pMux_14, a(4)=>
      gen_14_cmp_pMux_13, a(3)=>gen_14_cmp_pMux_12, a(2)=>gen_14_cmp_pMux_11, 
      a(1)=>gen_14_cmp_pMux_10, a(0)=>gen_14_cmp_pMux_9, b(23)=>nx9823, 
      b(22)=>nx9823, b(21)=>nx9821, b(20)=>nx9829, b(19)=>nx9827, b(18)=>
      nx9825, b(17)=>nx9823, b(16)=>nx9821, b(15)=>gen_14_cmp_BSCmp_op2_15, 
      b(14)=>gen_14_cmp_BSCmp_op2_14, b(13)=>gen_14_cmp_BSCmp_op2_13, b(12)
      =>gen_14_cmp_BSCmp_op2_12, b(11)=>gen_14_cmp_BSCmp_op2_11, b(10)=>
      gen_14_cmp_BSCmp_op2_10, b(9)=>gen_14_cmp_BSCmp_op2_9, b(8)=>
      gen_14_cmp_BSCmp_op2_8, b(7)=>gen_14_cmp_BSCmp_op2_7, b(6)=>
      gen_14_cmp_BSCmp_op2_6, b(5)=>gen_14_cmp_BSCmp_op2_5, b(4)=>
      gen_14_cmp_BSCmp_op2_4, b(3)=>gen_14_cmp_BSCmp_op2_3, b(2)=>
      gen_14_cmp_BSCmp_op2_2, b(1)=>gen_14_cmp_BSCmp_op2_1, b(0)=>
      gen_14_cmp_BSCmp_op2_0, carryIn=>gen_14_cmp_BSCmp_carryIn, sum(23)=>
      gen_14_cmp_pBs_30, sum(22)=>gen_14_cmp_pBs_29, sum(21)=>
      gen_14_cmp_pBs_28, sum(20)=>gen_14_cmp_pBs_27, sum(19)=>
      gen_14_cmp_pBs_26, sum(18)=>gen_14_cmp_pBs_25, sum(17)=>
      gen_14_cmp_pBs_24, sum(16)=>gen_14_cmp_pBs_23, sum(15)=>outputs_14_15, 
      sum(14)=>outputs_14_14, sum(13)=>outputs_14_13, sum(12)=>outputs_14_12, 
      sum(11)=>outputs_14_11, sum(10)=>outputs_14_10, sum(9)=>outputs_14_9, 
      sum(8)=>outputs_14_8, sum(7)=>outputs_14_7, sum(6)=>outputs_14_6, 
      sum(5)=>outputs_14_5, sum(4)=>outputs_14_4, sum(3)=>outputs_14_3, 
      sum(2)=>outputs_14_2, sum(1)=>outputs_14_1, sum(0)=>outputs_14_0, 
      carryOut=>DANGLING(54));
   gen_13_cmp_pRegCmp : Reg_33 port map ( D(32)=>working, D(31)=>working, 
      D(30)=>gen_13_cmp_pBs_30, D(29)=>gen_13_cmp_pBs_29, D(28)=>
      gen_13_cmp_pBs_28, D(27)=>gen_13_cmp_pBs_27, D(26)=>gen_13_cmp_pBs_26, 
      D(25)=>gen_13_cmp_pBs_25, D(24)=>gen_13_cmp_pBs_24, D(23)=>
      gen_13_cmp_pBs_23, D(22)=>outputs_13_15, D(21)=>outputs_13_14, D(20)=>
      outputs_13_13, D(19)=>outputs_13_12, D(18)=>outputs_13_11, D(17)=>
      outputs_13_10, D(16)=>outputs_13_9, D(15)=>outputs_13_8, D(14)=>
      outputs_13_7, D(13)=>outputs_13_6, D(12)=>outputs_13_5, D(11)=>
      outputs_13_4, D(10)=>outputs_13_3, D(9)=>outputs_13_2, D(8)=>
      outputs_13_1, D(7)=>outputs_13_0, D(6)=>gen_13_cmp_pMux_8, D(5)=>
      gen_13_cmp_pMux_7, D(4)=>gen_13_cmp_pMux_6, D(3)=>gen_13_cmp_pMux_5, 
      D(2)=>gen_13_cmp_pMux_4, D(1)=>gen_13_cmp_pMux_3, D(0)=>nx9531, en=>
      nx11165, clk=>nx9393, rst=>rst, Q(32)=>DANGLING(55), Q(31)=>DANGLING(
      56), Q(30)=>gen_13_cmp_pReg_30, Q(29)=>gen_13_cmp_pReg_29, Q(28)=>
      gen_13_cmp_pReg_28, Q(27)=>gen_13_cmp_pReg_27, Q(26)=>
      gen_13_cmp_pReg_26, Q(25)=>gen_13_cmp_pReg_25, Q(24)=>
      gen_13_cmp_pReg_24, Q(23)=>gen_13_cmp_pReg_23, Q(22)=>
      gen_13_cmp_pReg_22, Q(21)=>gen_13_cmp_pReg_21, Q(20)=>
      gen_13_cmp_pReg_20, Q(19)=>gen_13_cmp_pReg_19, Q(18)=>
      gen_13_cmp_pReg_18, Q(17)=>gen_13_cmp_pReg_17, Q(16)=>
      gen_13_cmp_pReg_16, Q(15)=>gen_13_cmp_pReg_15, Q(14)=>
      gen_13_cmp_pReg_14, Q(13)=>gen_13_cmp_pReg_13, Q(12)=>
      gen_13_cmp_pReg_12, Q(11)=>gen_13_cmp_pReg_11, Q(10)=>
      gen_13_cmp_pReg_10, Q(9)=>gen_13_cmp_pReg_9, Q(8)=>gen_13_cmp_pReg_8, 
      Q(7)=>gen_13_cmp_pReg_7, Q(6)=>gen_13_cmp_pReg_6, Q(5)=>
      gen_13_cmp_pReg_5, Q(4)=>gen_13_cmp_pReg_4, Q(3)=>gen_13_cmp_pReg_3, 
      Q(2)=>gen_13_cmp_pReg_2, Q(1)=>gen_13_cmp_pReg_1, Q(0)=>
      gen_13_cmp_pReg_0);
   gen_13_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>working, a(31)=>
      working, a(30)=>gen_13_cmp_pReg_30, a(29)=>gen_13_cmp_pReg_29, a(28)=>
      gen_13_cmp_pReg_28, a(27)=>gen_13_cmp_pReg_27, a(26)=>
      gen_13_cmp_pReg_26, a(25)=>gen_13_cmp_pReg_25, a(24)=>
      gen_13_cmp_pReg_24, a(23)=>gen_13_cmp_pReg_23, a(22)=>
      gen_13_cmp_pReg_22, a(21)=>gen_13_cmp_pReg_21, a(20)=>
      gen_13_cmp_pReg_20, a(19)=>gen_13_cmp_pReg_19, a(18)=>
      gen_13_cmp_pReg_18, a(17)=>gen_13_cmp_pReg_17, a(16)=>
      gen_13_cmp_pReg_16, a(15)=>gen_13_cmp_pReg_15, a(14)=>
      gen_13_cmp_pReg_14, a(13)=>gen_13_cmp_pReg_13, a(12)=>
      gen_13_cmp_pReg_12, a(11)=>gen_13_cmp_pReg_11, a(10)=>
      gen_13_cmp_pReg_10, a(9)=>gen_13_cmp_pReg_9, a(8)=>gen_13_cmp_pReg_8, 
      a(7)=>gen_13_cmp_pReg_7, a(6)=>gen_13_cmp_pReg_6, a(5)=>
      gen_13_cmp_pReg_5, a(4)=>gen_13_cmp_pReg_4, a(3)=>gen_13_cmp_pReg_3, 
      a(2)=>gen_13_cmp_pReg_2, a(1)=>gen_13_cmp_pReg_1, a(0)=>
      gen_13_cmp_pReg_0, b(32)=>working, b(31)=>working, b(30)=>working, 
      b(29)=>working, b(28)=>working, b(27)=>working, b(26)=>working, b(25)
      =>working, b(24)=>working, b(23)=>working, b(22)=>working, b(21)=>
      working, b(20)=>working, b(19)=>working, b(18)=>working, b(17)=>
      working, b(16)=>working, b(15)=>working, b(14)=>working, b(13)=>
      working, b(12)=>working, b(11)=>working, b(10)=>working, b(9)=>working, 
      b(8)=>filter_13_7, b(7)=>filter_13_6, b(6)=>filter_13_5, b(5)=>
      filter_13_4, b(4)=>filter_13_3, b(3)=>filter_13_2, b(2)=>filter_13_1, 
      b(1)=>filter_13_0, b(0)=>working, sel=>nx11181, f(32)=>DANGLING(57), 
      f(31)=>DANGLING(58), f(30)=>gen_13_cmp_pMux_30, f(29)=>
      gen_13_cmp_pMux_29, f(28)=>gen_13_cmp_pMux_28, f(27)=>
      gen_13_cmp_pMux_27, f(26)=>gen_13_cmp_pMux_26, f(25)=>
      gen_13_cmp_pMux_25, f(24)=>gen_13_cmp_pMux_24, f(23)=>
      gen_13_cmp_pMux_23, f(22)=>gen_13_cmp_pMux_22, f(21)=>
      gen_13_cmp_pMux_21, f(20)=>gen_13_cmp_pMux_20, f(19)=>
      gen_13_cmp_pMux_19, f(18)=>gen_13_cmp_pMux_18, f(17)=>
      gen_13_cmp_pMux_17, f(16)=>gen_13_cmp_pMux_16, f(15)=>
      gen_13_cmp_pMux_15, f(14)=>gen_13_cmp_pMux_14, f(13)=>
      gen_13_cmp_pMux_13, f(12)=>gen_13_cmp_pMux_12, f(11)=>
      gen_13_cmp_pMux_11, f(10)=>gen_13_cmp_pMux_10, f(9)=>gen_13_cmp_pMux_9, 
      f(8)=>gen_13_cmp_pMux_8, f(7)=>gen_13_cmp_pMux_7, f(6)=>
      gen_13_cmp_pMux_6, f(5)=>gen_13_cmp_pMux_5, f(4)=>gen_13_cmp_pMux_4, 
      f(3)=>gen_13_cmp_pMux_3, f(2)=>gen_13_cmp_pMux_2, f(1)=>
      gen_13_cmp_pMux_1, f(0)=>gen_13_cmp_pMux_0);
   gen_13_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>working, a(22)
      =>working, a(21)=>gen_13_cmp_pMux_30, a(20)=>gen_13_cmp_pMux_29, a(19)
      =>gen_13_cmp_pMux_28, a(18)=>gen_13_cmp_pMux_27, a(17)=>
      gen_13_cmp_pMux_26, a(16)=>gen_13_cmp_pMux_25, a(15)=>
      gen_13_cmp_pMux_24, a(14)=>gen_13_cmp_pMux_23, a(13)=>
      gen_13_cmp_pMux_22, a(12)=>gen_13_cmp_pMux_21, a(11)=>
      gen_13_cmp_pMux_20, a(10)=>gen_13_cmp_pMux_19, a(9)=>
      gen_13_cmp_pMux_18, a(8)=>gen_13_cmp_pMux_17, a(7)=>gen_13_cmp_pMux_16, 
      a(6)=>gen_13_cmp_pMux_15, a(5)=>gen_13_cmp_pMux_14, a(4)=>
      gen_13_cmp_pMux_13, a(3)=>gen_13_cmp_pMux_12, a(2)=>gen_13_cmp_pMux_11, 
      a(1)=>gen_13_cmp_pMux_10, a(0)=>gen_13_cmp_pMux_9, b(23)=>nx9835, 
      b(22)=>nx9835, b(21)=>nx9833, b(20)=>nx9841, b(19)=>nx9839, b(18)=>
      nx9837, b(17)=>nx9835, b(16)=>nx9833, b(15)=>gen_13_cmp_BSCmp_op2_15, 
      b(14)=>gen_13_cmp_BSCmp_op2_14, b(13)=>gen_13_cmp_BSCmp_op2_13, b(12)
      =>gen_13_cmp_BSCmp_op2_12, b(11)=>gen_13_cmp_BSCmp_op2_11, b(10)=>
      gen_13_cmp_BSCmp_op2_10, b(9)=>gen_13_cmp_BSCmp_op2_9, b(8)=>
      gen_13_cmp_BSCmp_op2_8, b(7)=>gen_13_cmp_BSCmp_op2_7, b(6)=>
      gen_13_cmp_BSCmp_op2_6, b(5)=>gen_13_cmp_BSCmp_op2_5, b(4)=>
      gen_13_cmp_BSCmp_op2_4, b(3)=>gen_13_cmp_BSCmp_op2_3, b(2)=>
      gen_13_cmp_BSCmp_op2_2, b(1)=>gen_13_cmp_BSCmp_op2_1, b(0)=>
      gen_13_cmp_BSCmp_op2_0, carryIn=>gen_13_cmp_BSCmp_carryIn, sum(23)=>
      gen_13_cmp_pBs_30, sum(22)=>gen_13_cmp_pBs_29, sum(21)=>
      gen_13_cmp_pBs_28, sum(20)=>gen_13_cmp_pBs_27, sum(19)=>
      gen_13_cmp_pBs_26, sum(18)=>gen_13_cmp_pBs_25, sum(17)=>
      gen_13_cmp_pBs_24, sum(16)=>gen_13_cmp_pBs_23, sum(15)=>outputs_13_15, 
      sum(14)=>outputs_13_14, sum(13)=>outputs_13_13, sum(12)=>outputs_13_12, 
      sum(11)=>outputs_13_11, sum(10)=>outputs_13_10, sum(9)=>outputs_13_9, 
      sum(8)=>outputs_13_8, sum(7)=>outputs_13_7, sum(6)=>outputs_13_6, 
      sum(5)=>outputs_13_5, sum(4)=>outputs_13_4, sum(3)=>outputs_13_3, 
      sum(2)=>outputs_13_2, sum(1)=>outputs_13_1, sum(0)=>outputs_13_0, 
      carryOut=>DANGLING(59));
   gen_12_cmp_pRegCmp : Reg_33 port map ( D(32)=>working, D(31)=>working, 
      D(30)=>gen_12_cmp_pBs_30, D(29)=>gen_12_cmp_pBs_29, D(28)=>
      gen_12_cmp_pBs_28, D(27)=>gen_12_cmp_pBs_27, D(26)=>gen_12_cmp_pBs_26, 
      D(25)=>gen_12_cmp_pBs_25, D(24)=>gen_12_cmp_pBs_24, D(23)=>
      gen_12_cmp_pBs_23, D(22)=>outputs_12_15, D(21)=>outputs_12_14, D(20)=>
      outputs_12_13, D(19)=>outputs_12_12, D(18)=>outputs_12_11, D(17)=>
      outputs_12_10, D(16)=>outputs_12_9, D(15)=>outputs_12_8, D(14)=>
      outputs_12_7, D(13)=>outputs_12_6, D(12)=>outputs_12_5, D(11)=>
      outputs_12_4, D(10)=>outputs_12_3, D(9)=>outputs_12_2, D(8)=>
      outputs_12_1, D(7)=>outputs_12_0, D(6)=>gen_12_cmp_pMux_8, D(5)=>
      gen_12_cmp_pMux_7, D(4)=>gen_12_cmp_pMux_6, D(3)=>gen_12_cmp_pMux_5, 
      D(2)=>gen_12_cmp_pMux_4, D(1)=>gen_12_cmp_pMux_3, D(0)=>nx9543, en=>
      nx11165, clk=>nx9393, rst=>rst, Q(32)=>DANGLING(60), Q(31)=>DANGLING(
      61), Q(30)=>gen_12_cmp_pReg_30, Q(29)=>gen_12_cmp_pReg_29, Q(28)=>
      gen_12_cmp_pReg_28, Q(27)=>gen_12_cmp_pReg_27, Q(26)=>
      gen_12_cmp_pReg_26, Q(25)=>gen_12_cmp_pReg_25, Q(24)=>
      gen_12_cmp_pReg_24, Q(23)=>gen_12_cmp_pReg_23, Q(22)=>
      gen_12_cmp_pReg_22, Q(21)=>gen_12_cmp_pReg_21, Q(20)=>
      gen_12_cmp_pReg_20, Q(19)=>gen_12_cmp_pReg_19, Q(18)=>
      gen_12_cmp_pReg_18, Q(17)=>gen_12_cmp_pReg_17, Q(16)=>
      gen_12_cmp_pReg_16, Q(15)=>gen_12_cmp_pReg_15, Q(14)=>
      gen_12_cmp_pReg_14, Q(13)=>gen_12_cmp_pReg_13, Q(12)=>
      gen_12_cmp_pReg_12, Q(11)=>gen_12_cmp_pReg_11, Q(10)=>
      gen_12_cmp_pReg_10, Q(9)=>gen_12_cmp_pReg_9, Q(8)=>gen_12_cmp_pReg_8, 
      Q(7)=>gen_12_cmp_pReg_7, Q(6)=>gen_12_cmp_pReg_6, Q(5)=>
      gen_12_cmp_pReg_5, Q(4)=>gen_12_cmp_pReg_4, Q(3)=>gen_12_cmp_pReg_3, 
      Q(2)=>gen_12_cmp_pReg_2, Q(1)=>gen_12_cmp_pReg_1, Q(0)=>
      gen_12_cmp_pReg_0);
   gen_12_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>working, a(31)=>
      working, a(30)=>gen_12_cmp_pReg_30, a(29)=>gen_12_cmp_pReg_29, a(28)=>
      gen_12_cmp_pReg_28, a(27)=>gen_12_cmp_pReg_27, a(26)=>
      gen_12_cmp_pReg_26, a(25)=>gen_12_cmp_pReg_25, a(24)=>
      gen_12_cmp_pReg_24, a(23)=>gen_12_cmp_pReg_23, a(22)=>
      gen_12_cmp_pReg_22, a(21)=>gen_12_cmp_pReg_21, a(20)=>
      gen_12_cmp_pReg_20, a(19)=>gen_12_cmp_pReg_19, a(18)=>
      gen_12_cmp_pReg_18, a(17)=>gen_12_cmp_pReg_17, a(16)=>
      gen_12_cmp_pReg_16, a(15)=>gen_12_cmp_pReg_15, a(14)=>
      gen_12_cmp_pReg_14, a(13)=>gen_12_cmp_pReg_13, a(12)=>
      gen_12_cmp_pReg_12, a(11)=>gen_12_cmp_pReg_11, a(10)=>
      gen_12_cmp_pReg_10, a(9)=>gen_12_cmp_pReg_9, a(8)=>gen_12_cmp_pReg_8, 
      a(7)=>gen_12_cmp_pReg_7, a(6)=>gen_12_cmp_pReg_6, a(5)=>
      gen_12_cmp_pReg_5, a(4)=>gen_12_cmp_pReg_4, a(3)=>gen_12_cmp_pReg_3, 
      a(2)=>gen_12_cmp_pReg_2, a(1)=>gen_12_cmp_pReg_1, a(0)=>
      gen_12_cmp_pReg_0, b(32)=>working, b(31)=>working, b(30)=>working, 
      b(29)=>working, b(28)=>working, b(27)=>working, b(26)=>working, b(25)
      =>working, b(24)=>working, b(23)=>working, b(22)=>working, b(21)=>
      working, b(20)=>working, b(19)=>working, b(18)=>working, b(17)=>
      working, b(16)=>working, b(15)=>working, b(14)=>working, b(13)=>
      working, b(12)=>working, b(11)=>working, b(10)=>working, b(9)=>working, 
      b(8)=>filter_12_7, b(7)=>filter_12_6, b(6)=>filter_12_5, b(5)=>
      filter_12_4, b(4)=>filter_12_3, b(3)=>filter_12_2, b(2)=>filter_12_1, 
      b(1)=>filter_12_0, b(0)=>working, sel=>nx11181, f(32)=>DANGLING(62), 
      f(31)=>DANGLING(63), f(30)=>gen_12_cmp_pMux_30, f(29)=>
      gen_12_cmp_pMux_29, f(28)=>gen_12_cmp_pMux_28, f(27)=>
      gen_12_cmp_pMux_27, f(26)=>gen_12_cmp_pMux_26, f(25)=>
      gen_12_cmp_pMux_25, f(24)=>gen_12_cmp_pMux_24, f(23)=>
      gen_12_cmp_pMux_23, f(22)=>gen_12_cmp_pMux_22, f(21)=>
      gen_12_cmp_pMux_21, f(20)=>gen_12_cmp_pMux_20, f(19)=>
      gen_12_cmp_pMux_19, f(18)=>gen_12_cmp_pMux_18, f(17)=>
      gen_12_cmp_pMux_17, f(16)=>gen_12_cmp_pMux_16, f(15)=>
      gen_12_cmp_pMux_15, f(14)=>gen_12_cmp_pMux_14, f(13)=>
      gen_12_cmp_pMux_13, f(12)=>gen_12_cmp_pMux_12, f(11)=>
      gen_12_cmp_pMux_11, f(10)=>gen_12_cmp_pMux_10, f(9)=>gen_12_cmp_pMux_9, 
      f(8)=>gen_12_cmp_pMux_8, f(7)=>gen_12_cmp_pMux_7, f(6)=>
      gen_12_cmp_pMux_6, f(5)=>gen_12_cmp_pMux_5, f(4)=>gen_12_cmp_pMux_4, 
      f(3)=>gen_12_cmp_pMux_3, f(2)=>gen_12_cmp_pMux_2, f(1)=>
      gen_12_cmp_pMux_1, f(0)=>gen_12_cmp_pMux_0);
   gen_12_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>working, a(22)
      =>working, a(21)=>gen_12_cmp_pMux_30, a(20)=>gen_12_cmp_pMux_29, a(19)
      =>gen_12_cmp_pMux_28, a(18)=>gen_12_cmp_pMux_27, a(17)=>
      gen_12_cmp_pMux_26, a(16)=>gen_12_cmp_pMux_25, a(15)=>
      gen_12_cmp_pMux_24, a(14)=>gen_12_cmp_pMux_23, a(13)=>
      gen_12_cmp_pMux_22, a(12)=>gen_12_cmp_pMux_21, a(11)=>
      gen_12_cmp_pMux_20, a(10)=>gen_12_cmp_pMux_19, a(9)=>
      gen_12_cmp_pMux_18, a(8)=>gen_12_cmp_pMux_17, a(7)=>gen_12_cmp_pMux_16, 
      a(6)=>gen_12_cmp_pMux_15, a(5)=>gen_12_cmp_pMux_14, a(4)=>
      gen_12_cmp_pMux_13, a(3)=>gen_12_cmp_pMux_12, a(2)=>gen_12_cmp_pMux_11, 
      a(1)=>gen_12_cmp_pMux_10, a(0)=>gen_12_cmp_pMux_9, b(23)=>nx9847, 
      b(22)=>nx9847, b(21)=>nx9845, b(20)=>nx9853, b(19)=>nx9851, b(18)=>
      nx9849, b(17)=>nx9847, b(16)=>nx9845, b(15)=>gen_12_cmp_BSCmp_op2_15, 
      b(14)=>gen_12_cmp_BSCmp_op2_14, b(13)=>gen_12_cmp_BSCmp_op2_13, b(12)
      =>gen_12_cmp_BSCmp_op2_12, b(11)=>gen_12_cmp_BSCmp_op2_11, b(10)=>
      gen_12_cmp_BSCmp_op2_10, b(9)=>gen_12_cmp_BSCmp_op2_9, b(8)=>
      gen_12_cmp_BSCmp_op2_8, b(7)=>gen_12_cmp_BSCmp_op2_7, b(6)=>
      gen_12_cmp_BSCmp_op2_6, b(5)=>gen_12_cmp_BSCmp_op2_5, b(4)=>
      gen_12_cmp_BSCmp_op2_4, b(3)=>gen_12_cmp_BSCmp_op2_3, b(2)=>
      gen_12_cmp_BSCmp_op2_2, b(1)=>gen_12_cmp_BSCmp_op2_1, b(0)=>
      gen_12_cmp_BSCmp_op2_0, carryIn=>gen_12_cmp_BSCmp_carryIn, sum(23)=>
      gen_12_cmp_pBs_30, sum(22)=>gen_12_cmp_pBs_29, sum(21)=>
      gen_12_cmp_pBs_28, sum(20)=>gen_12_cmp_pBs_27, sum(19)=>
      gen_12_cmp_pBs_26, sum(18)=>gen_12_cmp_pBs_25, sum(17)=>
      gen_12_cmp_pBs_24, sum(16)=>gen_12_cmp_pBs_23, sum(15)=>outputs_12_15, 
      sum(14)=>outputs_12_14, sum(13)=>outputs_12_13, sum(12)=>outputs_12_12, 
      sum(11)=>outputs_12_11, sum(10)=>outputs_12_10, sum(9)=>outputs_12_9, 
      sum(8)=>outputs_12_8, sum(7)=>outputs_12_7, sum(6)=>outputs_12_6, 
      sum(5)=>outputs_12_5, sum(4)=>outputs_12_4, sum(3)=>outputs_12_3, 
      sum(2)=>outputs_12_2, sum(1)=>outputs_12_1, sum(0)=>outputs_12_0, 
      carryOut=>DANGLING(64));
   gen_11_cmp_pRegCmp : Reg_33 port map ( D(32)=>working, D(31)=>working, 
      D(30)=>gen_11_cmp_pBs_30, D(29)=>gen_11_cmp_pBs_29, D(28)=>
      gen_11_cmp_pBs_28, D(27)=>gen_11_cmp_pBs_27, D(26)=>gen_11_cmp_pBs_26, 
      D(25)=>gen_11_cmp_pBs_25, D(24)=>gen_11_cmp_pBs_24, D(23)=>
      gen_11_cmp_pBs_23, D(22)=>outputs_11_15, D(21)=>outputs_11_14, D(20)=>
      outputs_11_13, D(19)=>outputs_11_12, D(18)=>outputs_11_11, D(17)=>
      outputs_11_10, D(16)=>outputs_11_9, D(15)=>outputs_11_8, D(14)=>
      outputs_11_7, D(13)=>outputs_11_6, D(12)=>outputs_11_5, D(11)=>
      outputs_11_4, D(10)=>outputs_11_3, D(9)=>outputs_11_2, D(8)=>
      outputs_11_1, D(7)=>outputs_11_0, D(6)=>gen_11_cmp_pMux_8, D(5)=>
      gen_11_cmp_pMux_7, D(4)=>gen_11_cmp_pMux_6, D(3)=>gen_11_cmp_pMux_5, 
      D(2)=>gen_11_cmp_pMux_4, D(1)=>gen_11_cmp_pMux_3, D(0)=>nx9555, en=>
      nx9377, clk=>nx9393, rst=>rst, Q(32)=>DANGLING(65), Q(31)=>DANGLING(66
      ), Q(30)=>gen_11_cmp_pReg_30, Q(29)=>gen_11_cmp_pReg_29, Q(28)=>
      gen_11_cmp_pReg_28, Q(27)=>gen_11_cmp_pReg_27, Q(26)=>
      gen_11_cmp_pReg_26, Q(25)=>gen_11_cmp_pReg_25, Q(24)=>
      gen_11_cmp_pReg_24, Q(23)=>gen_11_cmp_pReg_23, Q(22)=>
      gen_11_cmp_pReg_22, Q(21)=>gen_11_cmp_pReg_21, Q(20)=>
      gen_11_cmp_pReg_20, Q(19)=>gen_11_cmp_pReg_19, Q(18)=>
      gen_11_cmp_pReg_18, Q(17)=>gen_11_cmp_pReg_17, Q(16)=>
      gen_11_cmp_pReg_16, Q(15)=>gen_11_cmp_pReg_15, Q(14)=>
      gen_11_cmp_pReg_14, Q(13)=>gen_11_cmp_pReg_13, Q(12)=>
      gen_11_cmp_pReg_12, Q(11)=>gen_11_cmp_pReg_11, Q(10)=>
      gen_11_cmp_pReg_10, Q(9)=>gen_11_cmp_pReg_9, Q(8)=>gen_11_cmp_pReg_8, 
      Q(7)=>gen_11_cmp_pReg_7, Q(6)=>gen_11_cmp_pReg_6, Q(5)=>
      gen_11_cmp_pReg_5, Q(4)=>gen_11_cmp_pReg_4, Q(3)=>gen_11_cmp_pReg_3, 
      Q(2)=>gen_11_cmp_pReg_2, Q(1)=>gen_11_cmp_pReg_1, Q(0)=>
      gen_11_cmp_pReg_0);
   gen_11_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>working, a(31)=>
      working, a(30)=>gen_11_cmp_pReg_30, a(29)=>gen_11_cmp_pReg_29, a(28)=>
      gen_11_cmp_pReg_28, a(27)=>gen_11_cmp_pReg_27, a(26)=>
      gen_11_cmp_pReg_26, a(25)=>gen_11_cmp_pReg_25, a(24)=>
      gen_11_cmp_pReg_24, a(23)=>gen_11_cmp_pReg_23, a(22)=>
      gen_11_cmp_pReg_22, a(21)=>gen_11_cmp_pReg_21, a(20)=>
      gen_11_cmp_pReg_20, a(19)=>gen_11_cmp_pReg_19, a(18)=>
      gen_11_cmp_pReg_18, a(17)=>gen_11_cmp_pReg_17, a(16)=>
      gen_11_cmp_pReg_16, a(15)=>gen_11_cmp_pReg_15, a(14)=>
      gen_11_cmp_pReg_14, a(13)=>gen_11_cmp_pReg_13, a(12)=>
      gen_11_cmp_pReg_12, a(11)=>gen_11_cmp_pReg_11, a(10)=>
      gen_11_cmp_pReg_10, a(9)=>gen_11_cmp_pReg_9, a(8)=>gen_11_cmp_pReg_8, 
      a(7)=>gen_11_cmp_pReg_7, a(6)=>gen_11_cmp_pReg_6, a(5)=>
      gen_11_cmp_pReg_5, a(4)=>gen_11_cmp_pReg_4, a(3)=>gen_11_cmp_pReg_3, 
      a(2)=>gen_11_cmp_pReg_2, a(1)=>gen_11_cmp_pReg_1, a(0)=>
      gen_11_cmp_pReg_0, b(32)=>working, b(31)=>working, b(30)=>working, 
      b(29)=>working, b(28)=>working, b(27)=>working, b(26)=>working, b(25)
      =>working, b(24)=>working, b(23)=>working, b(22)=>working, b(21)=>
      working, b(20)=>working, b(19)=>working, b(18)=>working, b(17)=>
      working, b(16)=>working, b(15)=>working, b(14)=>working, b(13)=>
      working, b(12)=>working, b(11)=>working, b(10)=>working, b(9)=>working, 
      b(8)=>filter_11_7, b(7)=>filter_11_6, b(6)=>filter_11_5, b(5)=>
      filter_11_4, b(4)=>filter_11_3, b(3)=>filter_11_2, b(2)=>filter_11_1, 
      b(1)=>filter_11_0, b(0)=>working, sel=>nx11183, f(32)=>DANGLING(67), 
      f(31)=>DANGLING(68), f(30)=>gen_11_cmp_pMux_30, f(29)=>
      gen_11_cmp_pMux_29, f(28)=>gen_11_cmp_pMux_28, f(27)=>
      gen_11_cmp_pMux_27, f(26)=>gen_11_cmp_pMux_26, f(25)=>
      gen_11_cmp_pMux_25, f(24)=>gen_11_cmp_pMux_24, f(23)=>
      gen_11_cmp_pMux_23, f(22)=>gen_11_cmp_pMux_22, f(21)=>
      gen_11_cmp_pMux_21, f(20)=>gen_11_cmp_pMux_20, f(19)=>
      gen_11_cmp_pMux_19, f(18)=>gen_11_cmp_pMux_18, f(17)=>
      gen_11_cmp_pMux_17, f(16)=>gen_11_cmp_pMux_16, f(15)=>
      gen_11_cmp_pMux_15, f(14)=>gen_11_cmp_pMux_14, f(13)=>
      gen_11_cmp_pMux_13, f(12)=>gen_11_cmp_pMux_12, f(11)=>
      gen_11_cmp_pMux_11, f(10)=>gen_11_cmp_pMux_10, f(9)=>gen_11_cmp_pMux_9, 
      f(8)=>gen_11_cmp_pMux_8, f(7)=>gen_11_cmp_pMux_7, f(6)=>
      gen_11_cmp_pMux_6, f(5)=>gen_11_cmp_pMux_5, f(4)=>gen_11_cmp_pMux_4, 
      f(3)=>gen_11_cmp_pMux_3, f(2)=>gen_11_cmp_pMux_2, f(1)=>
      gen_11_cmp_pMux_1, f(0)=>gen_11_cmp_pMux_0);
   gen_11_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>working, a(22)
      =>working, a(21)=>gen_11_cmp_pMux_30, a(20)=>gen_11_cmp_pMux_29, a(19)
      =>gen_11_cmp_pMux_28, a(18)=>gen_11_cmp_pMux_27, a(17)=>
      gen_11_cmp_pMux_26, a(16)=>gen_11_cmp_pMux_25, a(15)=>
      gen_11_cmp_pMux_24, a(14)=>gen_11_cmp_pMux_23, a(13)=>
      gen_11_cmp_pMux_22, a(12)=>gen_11_cmp_pMux_21, a(11)=>
      gen_11_cmp_pMux_20, a(10)=>gen_11_cmp_pMux_19, a(9)=>
      gen_11_cmp_pMux_18, a(8)=>gen_11_cmp_pMux_17, a(7)=>gen_11_cmp_pMux_16, 
      a(6)=>gen_11_cmp_pMux_15, a(5)=>gen_11_cmp_pMux_14, a(4)=>
      gen_11_cmp_pMux_13, a(3)=>gen_11_cmp_pMux_12, a(2)=>gen_11_cmp_pMux_11, 
      a(1)=>gen_11_cmp_pMux_10, a(0)=>gen_11_cmp_pMux_9, b(23)=>nx9859, 
      b(22)=>nx9859, b(21)=>nx9857, b(20)=>nx9865, b(19)=>nx9863, b(18)=>
      nx9861, b(17)=>nx9859, b(16)=>nx9857, b(15)=>gen_11_cmp_BSCmp_op2_15, 
      b(14)=>gen_11_cmp_BSCmp_op2_14, b(13)=>gen_11_cmp_BSCmp_op2_13, b(12)
      =>gen_11_cmp_BSCmp_op2_12, b(11)=>gen_11_cmp_BSCmp_op2_11, b(10)=>
      gen_11_cmp_BSCmp_op2_10, b(9)=>gen_11_cmp_BSCmp_op2_9, b(8)=>
      gen_11_cmp_BSCmp_op2_8, b(7)=>gen_11_cmp_BSCmp_op2_7, b(6)=>
      gen_11_cmp_BSCmp_op2_6, b(5)=>gen_11_cmp_BSCmp_op2_5, b(4)=>
      gen_11_cmp_BSCmp_op2_4, b(3)=>gen_11_cmp_BSCmp_op2_3, b(2)=>
      gen_11_cmp_BSCmp_op2_2, b(1)=>gen_11_cmp_BSCmp_op2_1, b(0)=>
      gen_11_cmp_BSCmp_op2_0, carryIn=>gen_11_cmp_BSCmp_carryIn, sum(23)=>
      gen_11_cmp_pBs_30, sum(22)=>gen_11_cmp_pBs_29, sum(21)=>
      gen_11_cmp_pBs_28, sum(20)=>gen_11_cmp_pBs_27, sum(19)=>
      gen_11_cmp_pBs_26, sum(18)=>gen_11_cmp_pBs_25, sum(17)=>
      gen_11_cmp_pBs_24, sum(16)=>gen_11_cmp_pBs_23, sum(15)=>outputs_11_15, 
      sum(14)=>outputs_11_14, sum(13)=>outputs_11_13, sum(12)=>outputs_11_12, 
      sum(11)=>outputs_11_11, sum(10)=>outputs_11_10, sum(9)=>outputs_11_9, 
      sum(8)=>outputs_11_8, sum(7)=>outputs_11_7, sum(6)=>outputs_11_6, 
      sum(5)=>outputs_11_5, sum(4)=>outputs_11_4, sum(3)=>outputs_11_3, 
      sum(2)=>outputs_11_2, sum(1)=>outputs_11_1, sum(0)=>outputs_11_0, 
      carryOut=>DANGLING(69));
   gen_10_cmp_pRegCmp : Reg_33 port map ( D(32)=>working, D(31)=>working, 
      D(30)=>gen_10_cmp_pBs_30, D(29)=>gen_10_cmp_pBs_29, D(28)=>
      gen_10_cmp_pBs_28, D(27)=>gen_10_cmp_pBs_27, D(26)=>gen_10_cmp_pBs_26, 
      D(25)=>gen_10_cmp_pBs_25, D(24)=>gen_10_cmp_pBs_24, D(23)=>
      gen_10_cmp_pBs_23, D(22)=>outputs_10_15, D(21)=>outputs_10_14, D(20)=>
      outputs_10_13, D(19)=>outputs_10_12, D(18)=>outputs_10_11, D(17)=>
      outputs_10_10, D(16)=>outputs_10_9, D(15)=>outputs_10_8, D(14)=>
      outputs_10_7, D(13)=>outputs_10_6, D(12)=>outputs_10_5, D(11)=>
      outputs_10_4, D(10)=>outputs_10_3, D(9)=>outputs_10_2, D(8)=>
      outputs_10_1, D(7)=>outputs_10_0, D(6)=>gen_10_cmp_pMux_8, D(5)=>
      gen_10_cmp_pMux_7, D(4)=>gen_10_cmp_pMux_6, D(3)=>gen_10_cmp_pMux_5, 
      D(2)=>gen_10_cmp_pMux_4, D(1)=>gen_10_cmp_pMux_3, D(0)=>nx9567, en=>
      nx11167, clk=>nx9395, rst=>rst, Q(32)=>DANGLING(70), Q(31)=>DANGLING(
      71), Q(30)=>gen_10_cmp_pReg_30, Q(29)=>gen_10_cmp_pReg_29, Q(28)=>
      gen_10_cmp_pReg_28, Q(27)=>gen_10_cmp_pReg_27, Q(26)=>
      gen_10_cmp_pReg_26, Q(25)=>gen_10_cmp_pReg_25, Q(24)=>
      gen_10_cmp_pReg_24, Q(23)=>gen_10_cmp_pReg_23, Q(22)=>
      gen_10_cmp_pReg_22, Q(21)=>gen_10_cmp_pReg_21, Q(20)=>
      gen_10_cmp_pReg_20, Q(19)=>gen_10_cmp_pReg_19, Q(18)=>
      gen_10_cmp_pReg_18, Q(17)=>gen_10_cmp_pReg_17, Q(16)=>
      gen_10_cmp_pReg_16, Q(15)=>gen_10_cmp_pReg_15, Q(14)=>
      gen_10_cmp_pReg_14, Q(13)=>gen_10_cmp_pReg_13, Q(12)=>
      gen_10_cmp_pReg_12, Q(11)=>gen_10_cmp_pReg_11, Q(10)=>
      gen_10_cmp_pReg_10, Q(9)=>gen_10_cmp_pReg_9, Q(8)=>gen_10_cmp_pReg_8, 
      Q(7)=>gen_10_cmp_pReg_7, Q(6)=>gen_10_cmp_pReg_6, Q(5)=>
      gen_10_cmp_pReg_5, Q(4)=>gen_10_cmp_pReg_4, Q(3)=>gen_10_cmp_pReg_3, 
      Q(2)=>gen_10_cmp_pReg_2, Q(1)=>gen_10_cmp_pReg_1, Q(0)=>
      gen_10_cmp_pReg_0);
   gen_10_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>working, a(31)=>
      working, a(30)=>gen_10_cmp_pReg_30, a(29)=>gen_10_cmp_pReg_29, a(28)=>
      gen_10_cmp_pReg_28, a(27)=>gen_10_cmp_pReg_27, a(26)=>
      gen_10_cmp_pReg_26, a(25)=>gen_10_cmp_pReg_25, a(24)=>
      gen_10_cmp_pReg_24, a(23)=>gen_10_cmp_pReg_23, a(22)=>
      gen_10_cmp_pReg_22, a(21)=>gen_10_cmp_pReg_21, a(20)=>
      gen_10_cmp_pReg_20, a(19)=>gen_10_cmp_pReg_19, a(18)=>
      gen_10_cmp_pReg_18, a(17)=>gen_10_cmp_pReg_17, a(16)=>
      gen_10_cmp_pReg_16, a(15)=>gen_10_cmp_pReg_15, a(14)=>
      gen_10_cmp_pReg_14, a(13)=>gen_10_cmp_pReg_13, a(12)=>
      gen_10_cmp_pReg_12, a(11)=>gen_10_cmp_pReg_11, a(10)=>
      gen_10_cmp_pReg_10, a(9)=>gen_10_cmp_pReg_9, a(8)=>gen_10_cmp_pReg_8, 
      a(7)=>gen_10_cmp_pReg_7, a(6)=>gen_10_cmp_pReg_6, a(5)=>
      gen_10_cmp_pReg_5, a(4)=>gen_10_cmp_pReg_4, a(3)=>gen_10_cmp_pReg_3, 
      a(2)=>gen_10_cmp_pReg_2, a(1)=>gen_10_cmp_pReg_1, a(0)=>
      gen_10_cmp_pReg_0, b(32)=>working, b(31)=>working, b(30)=>working, 
      b(29)=>working, b(28)=>working, b(27)=>working, b(26)=>working, b(25)
      =>working, b(24)=>working, b(23)=>working, b(22)=>working, b(21)=>
      working, b(20)=>working, b(19)=>working, b(18)=>working, b(17)=>
      working, b(16)=>working, b(15)=>working, b(14)=>working, b(13)=>
      working, b(12)=>working, b(11)=>working, b(10)=>working, b(9)=>working, 
      b(8)=>filter_10_7, b(7)=>filter_10_6, b(6)=>filter_10_5, b(5)=>
      filter_10_4, b(4)=>filter_10_3, b(3)=>filter_10_2, b(2)=>filter_10_1, 
      b(1)=>filter_10_0, b(0)=>working, sel=>nx11185, f(32)=>DANGLING(72), 
      f(31)=>DANGLING(73), f(30)=>gen_10_cmp_pMux_30, f(29)=>
      gen_10_cmp_pMux_29, f(28)=>gen_10_cmp_pMux_28, f(27)=>
      gen_10_cmp_pMux_27, f(26)=>gen_10_cmp_pMux_26, f(25)=>
      gen_10_cmp_pMux_25, f(24)=>gen_10_cmp_pMux_24, f(23)=>
      gen_10_cmp_pMux_23, f(22)=>gen_10_cmp_pMux_22, f(21)=>
      gen_10_cmp_pMux_21, f(20)=>gen_10_cmp_pMux_20, f(19)=>
      gen_10_cmp_pMux_19, f(18)=>gen_10_cmp_pMux_18, f(17)=>
      gen_10_cmp_pMux_17, f(16)=>gen_10_cmp_pMux_16, f(15)=>
      gen_10_cmp_pMux_15, f(14)=>gen_10_cmp_pMux_14, f(13)=>
      gen_10_cmp_pMux_13, f(12)=>gen_10_cmp_pMux_12, f(11)=>
      gen_10_cmp_pMux_11, f(10)=>gen_10_cmp_pMux_10, f(9)=>gen_10_cmp_pMux_9, 
      f(8)=>gen_10_cmp_pMux_8, f(7)=>gen_10_cmp_pMux_7, f(6)=>
      gen_10_cmp_pMux_6, f(5)=>gen_10_cmp_pMux_5, f(4)=>gen_10_cmp_pMux_4, 
      f(3)=>gen_10_cmp_pMux_3, f(2)=>gen_10_cmp_pMux_2, f(1)=>
      gen_10_cmp_pMux_1, f(0)=>gen_10_cmp_pMux_0);
   gen_10_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>working, a(22)
      =>working, a(21)=>gen_10_cmp_pMux_30, a(20)=>gen_10_cmp_pMux_29, a(19)
      =>gen_10_cmp_pMux_28, a(18)=>gen_10_cmp_pMux_27, a(17)=>
      gen_10_cmp_pMux_26, a(16)=>gen_10_cmp_pMux_25, a(15)=>
      gen_10_cmp_pMux_24, a(14)=>gen_10_cmp_pMux_23, a(13)=>
      gen_10_cmp_pMux_22, a(12)=>gen_10_cmp_pMux_21, a(11)=>
      gen_10_cmp_pMux_20, a(10)=>gen_10_cmp_pMux_19, a(9)=>
      gen_10_cmp_pMux_18, a(8)=>gen_10_cmp_pMux_17, a(7)=>gen_10_cmp_pMux_16, 
      a(6)=>gen_10_cmp_pMux_15, a(5)=>gen_10_cmp_pMux_14, a(4)=>
      gen_10_cmp_pMux_13, a(3)=>gen_10_cmp_pMux_12, a(2)=>gen_10_cmp_pMux_11, 
      a(1)=>gen_10_cmp_pMux_10, a(0)=>gen_10_cmp_pMux_9, b(23)=>nx9871, 
      b(22)=>nx9871, b(21)=>nx9869, b(20)=>nx9877, b(19)=>nx9875, b(18)=>
      nx9873, b(17)=>nx9871, b(16)=>nx9869, b(15)=>gen_10_cmp_BSCmp_op2_15, 
      b(14)=>gen_10_cmp_BSCmp_op2_14, b(13)=>gen_10_cmp_BSCmp_op2_13, b(12)
      =>gen_10_cmp_BSCmp_op2_12, b(11)=>gen_10_cmp_BSCmp_op2_11, b(10)=>
      gen_10_cmp_BSCmp_op2_10, b(9)=>gen_10_cmp_BSCmp_op2_9, b(8)=>
      gen_10_cmp_BSCmp_op2_8, b(7)=>gen_10_cmp_BSCmp_op2_7, b(6)=>
      gen_10_cmp_BSCmp_op2_6, b(5)=>gen_10_cmp_BSCmp_op2_5, b(4)=>
      gen_10_cmp_BSCmp_op2_4, b(3)=>gen_10_cmp_BSCmp_op2_3, b(2)=>
      gen_10_cmp_BSCmp_op2_2, b(1)=>gen_10_cmp_BSCmp_op2_1, b(0)=>
      gen_10_cmp_BSCmp_op2_0, carryIn=>gen_10_cmp_BSCmp_carryIn, sum(23)=>
      gen_10_cmp_pBs_30, sum(22)=>gen_10_cmp_pBs_29, sum(21)=>
      gen_10_cmp_pBs_28, sum(20)=>gen_10_cmp_pBs_27, sum(19)=>
      gen_10_cmp_pBs_26, sum(18)=>gen_10_cmp_pBs_25, sum(17)=>
      gen_10_cmp_pBs_24, sum(16)=>gen_10_cmp_pBs_23, sum(15)=>outputs_10_15, 
      sum(14)=>outputs_10_14, sum(13)=>outputs_10_13, sum(12)=>outputs_10_12, 
      sum(11)=>outputs_10_11, sum(10)=>outputs_10_10, sum(9)=>outputs_10_9, 
      sum(8)=>outputs_10_8, sum(7)=>outputs_10_7, sum(6)=>outputs_10_6, 
      sum(5)=>outputs_10_5, sum(4)=>outputs_10_4, sum(3)=>outputs_10_3, 
      sum(2)=>outputs_10_2, sum(1)=>outputs_10_1, sum(0)=>outputs_10_0, 
      carryOut=>DANGLING(74));
   gen_9_cmp_pRegCmp : Reg_33 port map ( D(32)=>working, D(31)=>working, 
      D(30)=>gen_9_cmp_pBs_30, D(29)=>gen_9_cmp_pBs_29, D(28)=>
      gen_9_cmp_pBs_28, D(27)=>gen_9_cmp_pBs_27, D(26)=>gen_9_cmp_pBs_26, 
      D(25)=>gen_9_cmp_pBs_25, D(24)=>gen_9_cmp_pBs_24, D(23)=>
      gen_9_cmp_pBs_23, D(22)=>outputs_9_15, D(21)=>outputs_9_14, D(20)=>
      outputs_9_13, D(19)=>outputs_9_12, D(18)=>outputs_9_11, D(17)=>
      outputs_9_10, D(16)=>outputs_9_9, D(15)=>outputs_9_8, D(14)=>
      outputs_9_7, D(13)=>outputs_9_6, D(12)=>outputs_9_5, D(11)=>
      outputs_9_4, D(10)=>outputs_9_3, D(9)=>outputs_9_2, D(8)=>outputs_9_1, 
      D(7)=>outputs_9_0, D(6)=>gen_9_cmp_pMux_8, D(5)=>gen_9_cmp_pMux_7, 
      D(4)=>gen_9_cmp_pMux_6, D(3)=>gen_9_cmp_pMux_5, D(2)=>gen_9_cmp_pMux_4, 
      D(1)=>gen_9_cmp_pMux_3, D(0)=>nx9579, en=>nx11167, clk=>nx9395, rst=>
      rst, Q(32)=>DANGLING(75), Q(31)=>DANGLING(76), Q(30)=>
      gen_9_cmp_pReg_30, Q(29)=>gen_9_cmp_pReg_29, Q(28)=>gen_9_cmp_pReg_28, 
      Q(27)=>gen_9_cmp_pReg_27, Q(26)=>gen_9_cmp_pReg_26, Q(25)=>
      gen_9_cmp_pReg_25, Q(24)=>gen_9_cmp_pReg_24, Q(23)=>gen_9_cmp_pReg_23, 
      Q(22)=>gen_9_cmp_pReg_22, Q(21)=>gen_9_cmp_pReg_21, Q(20)=>
      gen_9_cmp_pReg_20, Q(19)=>gen_9_cmp_pReg_19, Q(18)=>gen_9_cmp_pReg_18, 
      Q(17)=>gen_9_cmp_pReg_17, Q(16)=>gen_9_cmp_pReg_16, Q(15)=>
      gen_9_cmp_pReg_15, Q(14)=>gen_9_cmp_pReg_14, Q(13)=>gen_9_cmp_pReg_13, 
      Q(12)=>gen_9_cmp_pReg_12, Q(11)=>gen_9_cmp_pReg_11, Q(10)=>
      gen_9_cmp_pReg_10, Q(9)=>gen_9_cmp_pReg_9, Q(8)=>gen_9_cmp_pReg_8, 
      Q(7)=>gen_9_cmp_pReg_7, Q(6)=>gen_9_cmp_pReg_6, Q(5)=>gen_9_cmp_pReg_5, 
      Q(4)=>gen_9_cmp_pReg_4, Q(3)=>gen_9_cmp_pReg_3, Q(2)=>gen_9_cmp_pReg_2, 
      Q(1)=>gen_9_cmp_pReg_1, Q(0)=>gen_9_cmp_pReg_0);
   gen_9_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>working, a(31)=>working, 
      a(30)=>gen_9_cmp_pReg_30, a(29)=>gen_9_cmp_pReg_29, a(28)=>
      gen_9_cmp_pReg_28, a(27)=>gen_9_cmp_pReg_27, a(26)=>gen_9_cmp_pReg_26, 
      a(25)=>gen_9_cmp_pReg_25, a(24)=>gen_9_cmp_pReg_24, a(23)=>
      gen_9_cmp_pReg_23, a(22)=>gen_9_cmp_pReg_22, a(21)=>gen_9_cmp_pReg_21, 
      a(20)=>gen_9_cmp_pReg_20, a(19)=>gen_9_cmp_pReg_19, a(18)=>
      gen_9_cmp_pReg_18, a(17)=>gen_9_cmp_pReg_17, a(16)=>gen_9_cmp_pReg_16, 
      a(15)=>gen_9_cmp_pReg_15, a(14)=>gen_9_cmp_pReg_14, a(13)=>
      gen_9_cmp_pReg_13, a(12)=>gen_9_cmp_pReg_12, a(11)=>gen_9_cmp_pReg_11, 
      a(10)=>gen_9_cmp_pReg_10, a(9)=>gen_9_cmp_pReg_9, a(8)=>
      gen_9_cmp_pReg_8, a(7)=>gen_9_cmp_pReg_7, a(6)=>gen_9_cmp_pReg_6, a(5)
      =>gen_9_cmp_pReg_5, a(4)=>gen_9_cmp_pReg_4, a(3)=>gen_9_cmp_pReg_3, 
      a(2)=>gen_9_cmp_pReg_2, a(1)=>gen_9_cmp_pReg_1, a(0)=>gen_9_cmp_pReg_0, 
      b(32)=>working, b(31)=>working, b(30)=>working, b(29)=>working, b(28)
      =>working, b(27)=>working, b(26)=>working, b(25)=>working, b(24)=>
      working, b(23)=>working, b(22)=>working, b(21)=>working, b(20)=>
      working, b(19)=>working, b(18)=>working, b(17)=>working, b(16)=>
      working, b(15)=>working, b(14)=>working, b(13)=>working, b(12)=>
      working, b(11)=>working, b(10)=>working, b(9)=>working, b(8)=>
      filter_9_7, b(7)=>filter_9_6, b(6)=>filter_9_5, b(5)=>filter_9_4, b(4)
      =>filter_9_3, b(3)=>filter_9_2, b(2)=>filter_9_1, b(1)=>filter_9_0, 
      b(0)=>working, sel=>nx11185, f(32)=>DANGLING(77), f(31)=>DANGLING(78), 
      f(30)=>gen_9_cmp_pMux_30, f(29)=>gen_9_cmp_pMux_29, f(28)=>
      gen_9_cmp_pMux_28, f(27)=>gen_9_cmp_pMux_27, f(26)=>gen_9_cmp_pMux_26, 
      f(25)=>gen_9_cmp_pMux_25, f(24)=>gen_9_cmp_pMux_24, f(23)=>
      gen_9_cmp_pMux_23, f(22)=>gen_9_cmp_pMux_22, f(21)=>gen_9_cmp_pMux_21, 
      f(20)=>gen_9_cmp_pMux_20, f(19)=>gen_9_cmp_pMux_19, f(18)=>
      gen_9_cmp_pMux_18, f(17)=>gen_9_cmp_pMux_17, f(16)=>gen_9_cmp_pMux_16, 
      f(15)=>gen_9_cmp_pMux_15, f(14)=>gen_9_cmp_pMux_14, f(13)=>
      gen_9_cmp_pMux_13, f(12)=>gen_9_cmp_pMux_12, f(11)=>gen_9_cmp_pMux_11, 
      f(10)=>gen_9_cmp_pMux_10, f(9)=>gen_9_cmp_pMux_9, f(8)=>
      gen_9_cmp_pMux_8, f(7)=>gen_9_cmp_pMux_7, f(6)=>gen_9_cmp_pMux_6, f(5)
      =>gen_9_cmp_pMux_5, f(4)=>gen_9_cmp_pMux_4, f(3)=>gen_9_cmp_pMux_3, 
      f(2)=>gen_9_cmp_pMux_2, f(1)=>gen_9_cmp_pMux_1, f(0)=>gen_9_cmp_pMux_0
   );
   gen_9_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>working, a(22)
      =>working, a(21)=>gen_9_cmp_pMux_30, a(20)=>gen_9_cmp_pMux_29, a(19)=>
      gen_9_cmp_pMux_28, a(18)=>gen_9_cmp_pMux_27, a(17)=>gen_9_cmp_pMux_26, 
      a(16)=>gen_9_cmp_pMux_25, a(15)=>gen_9_cmp_pMux_24, a(14)=>
      gen_9_cmp_pMux_23, a(13)=>gen_9_cmp_pMux_22, a(12)=>gen_9_cmp_pMux_21, 
      a(11)=>gen_9_cmp_pMux_20, a(10)=>gen_9_cmp_pMux_19, a(9)=>
      gen_9_cmp_pMux_18, a(8)=>gen_9_cmp_pMux_17, a(7)=>gen_9_cmp_pMux_16, 
      a(6)=>gen_9_cmp_pMux_15, a(5)=>gen_9_cmp_pMux_14, a(4)=>
      gen_9_cmp_pMux_13, a(3)=>gen_9_cmp_pMux_12, a(2)=>gen_9_cmp_pMux_11, 
      a(1)=>gen_9_cmp_pMux_10, a(0)=>gen_9_cmp_pMux_9, b(23)=>nx9883, b(22)
      =>nx9883, b(21)=>nx9881, b(20)=>nx9889, b(19)=>nx9887, b(18)=>nx9885, 
      b(17)=>nx9883, b(16)=>nx9881, b(15)=>gen_9_cmp_BSCmp_op2_15, b(14)=>
      gen_9_cmp_BSCmp_op2_14, b(13)=>gen_9_cmp_BSCmp_op2_13, b(12)=>
      gen_9_cmp_BSCmp_op2_12, b(11)=>gen_9_cmp_BSCmp_op2_11, b(10)=>
      gen_9_cmp_BSCmp_op2_10, b(9)=>gen_9_cmp_BSCmp_op2_9, b(8)=>
      gen_9_cmp_BSCmp_op2_8, b(7)=>gen_9_cmp_BSCmp_op2_7, b(6)=>
      gen_9_cmp_BSCmp_op2_6, b(5)=>gen_9_cmp_BSCmp_op2_5, b(4)=>
      gen_9_cmp_BSCmp_op2_4, b(3)=>gen_9_cmp_BSCmp_op2_3, b(2)=>
      gen_9_cmp_BSCmp_op2_2, b(1)=>gen_9_cmp_BSCmp_op2_1, b(0)=>
      gen_9_cmp_BSCmp_op2_0, carryIn=>gen_9_cmp_BSCmp_carryIn, sum(23)=>
      gen_9_cmp_pBs_30, sum(22)=>gen_9_cmp_pBs_29, sum(21)=>gen_9_cmp_pBs_28, 
      sum(20)=>gen_9_cmp_pBs_27, sum(19)=>gen_9_cmp_pBs_26, sum(18)=>
      gen_9_cmp_pBs_25, sum(17)=>gen_9_cmp_pBs_24, sum(16)=>gen_9_cmp_pBs_23, 
      sum(15)=>outputs_9_15, sum(14)=>outputs_9_14, sum(13)=>outputs_9_13, 
      sum(12)=>outputs_9_12, sum(11)=>outputs_9_11, sum(10)=>outputs_9_10, 
      sum(9)=>outputs_9_9, sum(8)=>outputs_9_8, sum(7)=>outputs_9_7, sum(6)
      =>outputs_9_6, sum(5)=>outputs_9_5, sum(4)=>outputs_9_4, sum(3)=>
      outputs_9_3, sum(2)=>outputs_9_2, sum(1)=>outputs_9_1, sum(0)=>
      outputs_9_0, carryOut=>DANGLING(79));
   gen_8_cmp_pRegCmp : Reg_33 port map ( D(32)=>working, D(31)=>working, 
      D(30)=>gen_8_cmp_pBs_30, D(29)=>gen_8_cmp_pBs_29, D(28)=>
      gen_8_cmp_pBs_28, D(27)=>gen_8_cmp_pBs_27, D(26)=>gen_8_cmp_pBs_26, 
      D(25)=>gen_8_cmp_pBs_25, D(24)=>gen_8_cmp_pBs_24, D(23)=>
      gen_8_cmp_pBs_23, D(22)=>outputs_8_15, D(21)=>outputs_8_14, D(20)=>
      outputs_8_13, D(19)=>outputs_8_12, D(18)=>outputs_8_11, D(17)=>
      outputs_8_10, D(16)=>outputs_8_9, D(15)=>outputs_8_8, D(14)=>
      outputs_8_7, D(13)=>outputs_8_6, D(12)=>outputs_8_5, D(11)=>
      outputs_8_4, D(10)=>outputs_8_3, D(9)=>outputs_8_2, D(8)=>outputs_8_1, 
      D(7)=>outputs_8_0, D(6)=>gen_8_cmp_pMux_8, D(5)=>gen_8_cmp_pMux_7, 
      D(4)=>gen_8_cmp_pMux_6, D(3)=>gen_8_cmp_pMux_5, D(2)=>gen_8_cmp_pMux_4, 
      D(1)=>gen_8_cmp_pMux_3, D(0)=>nx9591, en=>nx11167, clk=>nx9395, rst=>
      rst, Q(32)=>DANGLING(80), Q(31)=>DANGLING(81), Q(30)=>
      gen_8_cmp_pReg_30, Q(29)=>gen_8_cmp_pReg_29, Q(28)=>gen_8_cmp_pReg_28, 
      Q(27)=>gen_8_cmp_pReg_27, Q(26)=>gen_8_cmp_pReg_26, Q(25)=>
      gen_8_cmp_pReg_25, Q(24)=>gen_8_cmp_pReg_24, Q(23)=>gen_8_cmp_pReg_23, 
      Q(22)=>gen_8_cmp_pReg_22, Q(21)=>gen_8_cmp_pReg_21, Q(20)=>
      gen_8_cmp_pReg_20, Q(19)=>gen_8_cmp_pReg_19, Q(18)=>gen_8_cmp_pReg_18, 
      Q(17)=>gen_8_cmp_pReg_17, Q(16)=>gen_8_cmp_pReg_16, Q(15)=>
      gen_8_cmp_pReg_15, Q(14)=>gen_8_cmp_pReg_14, Q(13)=>gen_8_cmp_pReg_13, 
      Q(12)=>gen_8_cmp_pReg_12, Q(11)=>gen_8_cmp_pReg_11, Q(10)=>
      gen_8_cmp_pReg_10, Q(9)=>gen_8_cmp_pReg_9, Q(8)=>gen_8_cmp_pReg_8, 
      Q(7)=>gen_8_cmp_pReg_7, Q(6)=>gen_8_cmp_pReg_6, Q(5)=>gen_8_cmp_pReg_5, 
      Q(4)=>gen_8_cmp_pReg_4, Q(3)=>gen_8_cmp_pReg_3, Q(2)=>gen_8_cmp_pReg_2, 
      Q(1)=>gen_8_cmp_pReg_1, Q(0)=>gen_8_cmp_pReg_0);
   gen_8_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>working, a(31)=>working, 
      a(30)=>gen_8_cmp_pReg_30, a(29)=>gen_8_cmp_pReg_29, a(28)=>
      gen_8_cmp_pReg_28, a(27)=>gen_8_cmp_pReg_27, a(26)=>gen_8_cmp_pReg_26, 
      a(25)=>gen_8_cmp_pReg_25, a(24)=>gen_8_cmp_pReg_24, a(23)=>
      gen_8_cmp_pReg_23, a(22)=>gen_8_cmp_pReg_22, a(21)=>gen_8_cmp_pReg_21, 
      a(20)=>gen_8_cmp_pReg_20, a(19)=>gen_8_cmp_pReg_19, a(18)=>
      gen_8_cmp_pReg_18, a(17)=>gen_8_cmp_pReg_17, a(16)=>gen_8_cmp_pReg_16, 
      a(15)=>gen_8_cmp_pReg_15, a(14)=>gen_8_cmp_pReg_14, a(13)=>
      gen_8_cmp_pReg_13, a(12)=>gen_8_cmp_pReg_12, a(11)=>gen_8_cmp_pReg_11, 
      a(10)=>gen_8_cmp_pReg_10, a(9)=>gen_8_cmp_pReg_9, a(8)=>
      gen_8_cmp_pReg_8, a(7)=>gen_8_cmp_pReg_7, a(6)=>gen_8_cmp_pReg_6, a(5)
      =>gen_8_cmp_pReg_5, a(4)=>gen_8_cmp_pReg_4, a(3)=>gen_8_cmp_pReg_3, 
      a(2)=>gen_8_cmp_pReg_2, a(1)=>gen_8_cmp_pReg_1, a(0)=>gen_8_cmp_pReg_0, 
      b(32)=>working, b(31)=>working, b(30)=>working, b(29)=>working, b(28)
      =>working, b(27)=>working, b(26)=>working, b(25)=>working, b(24)=>
      working, b(23)=>working, b(22)=>working, b(21)=>working, b(20)=>
      working, b(19)=>working, b(18)=>working, b(17)=>working, b(16)=>
      working, b(15)=>working, b(14)=>working, b(13)=>working, b(12)=>
      working, b(11)=>working, b(10)=>working, b(9)=>working, b(8)=>
      filter_8_7, b(7)=>filter_8_6, b(6)=>filter_8_5, b(5)=>filter_8_4, b(4)
      =>filter_8_3, b(3)=>filter_8_2, b(2)=>filter_8_1, b(1)=>filter_8_0, 
      b(0)=>working, sel=>nx11185, f(32)=>DANGLING(82), f(31)=>DANGLING(83), 
      f(30)=>gen_8_cmp_pMux_30, f(29)=>gen_8_cmp_pMux_29, f(28)=>
      gen_8_cmp_pMux_28, f(27)=>gen_8_cmp_pMux_27, f(26)=>gen_8_cmp_pMux_26, 
      f(25)=>gen_8_cmp_pMux_25, f(24)=>gen_8_cmp_pMux_24, f(23)=>
      gen_8_cmp_pMux_23, f(22)=>gen_8_cmp_pMux_22, f(21)=>gen_8_cmp_pMux_21, 
      f(20)=>gen_8_cmp_pMux_20, f(19)=>gen_8_cmp_pMux_19, f(18)=>
      gen_8_cmp_pMux_18, f(17)=>gen_8_cmp_pMux_17, f(16)=>gen_8_cmp_pMux_16, 
      f(15)=>gen_8_cmp_pMux_15, f(14)=>gen_8_cmp_pMux_14, f(13)=>
      gen_8_cmp_pMux_13, f(12)=>gen_8_cmp_pMux_12, f(11)=>gen_8_cmp_pMux_11, 
      f(10)=>gen_8_cmp_pMux_10, f(9)=>gen_8_cmp_pMux_9, f(8)=>
      gen_8_cmp_pMux_8, f(7)=>gen_8_cmp_pMux_7, f(6)=>gen_8_cmp_pMux_6, f(5)
      =>gen_8_cmp_pMux_5, f(4)=>gen_8_cmp_pMux_4, f(3)=>gen_8_cmp_pMux_3, 
      f(2)=>gen_8_cmp_pMux_2, f(1)=>gen_8_cmp_pMux_1, f(0)=>gen_8_cmp_pMux_0
   );
   gen_8_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>working, a(22)
      =>working, a(21)=>gen_8_cmp_pMux_30, a(20)=>gen_8_cmp_pMux_29, a(19)=>
      gen_8_cmp_pMux_28, a(18)=>gen_8_cmp_pMux_27, a(17)=>gen_8_cmp_pMux_26, 
      a(16)=>gen_8_cmp_pMux_25, a(15)=>gen_8_cmp_pMux_24, a(14)=>
      gen_8_cmp_pMux_23, a(13)=>gen_8_cmp_pMux_22, a(12)=>gen_8_cmp_pMux_21, 
      a(11)=>gen_8_cmp_pMux_20, a(10)=>gen_8_cmp_pMux_19, a(9)=>
      gen_8_cmp_pMux_18, a(8)=>gen_8_cmp_pMux_17, a(7)=>gen_8_cmp_pMux_16, 
      a(6)=>gen_8_cmp_pMux_15, a(5)=>gen_8_cmp_pMux_14, a(4)=>
      gen_8_cmp_pMux_13, a(3)=>gen_8_cmp_pMux_12, a(2)=>gen_8_cmp_pMux_11, 
      a(1)=>gen_8_cmp_pMux_10, a(0)=>gen_8_cmp_pMux_9, b(23)=>nx9895, b(22)
      =>nx9895, b(21)=>nx9893, b(20)=>nx9901, b(19)=>nx9899, b(18)=>nx9897, 
      b(17)=>nx9895, b(16)=>nx9893, b(15)=>gen_8_cmp_BSCmp_op2_15, b(14)=>
      gen_8_cmp_BSCmp_op2_14, b(13)=>gen_8_cmp_BSCmp_op2_13, b(12)=>
      gen_8_cmp_BSCmp_op2_12, b(11)=>gen_8_cmp_BSCmp_op2_11, b(10)=>
      gen_8_cmp_BSCmp_op2_10, b(9)=>gen_8_cmp_BSCmp_op2_9, b(8)=>
      gen_8_cmp_BSCmp_op2_8, b(7)=>gen_8_cmp_BSCmp_op2_7, b(6)=>
      gen_8_cmp_BSCmp_op2_6, b(5)=>gen_8_cmp_BSCmp_op2_5, b(4)=>
      gen_8_cmp_BSCmp_op2_4, b(3)=>gen_8_cmp_BSCmp_op2_3, b(2)=>
      gen_8_cmp_BSCmp_op2_2, b(1)=>gen_8_cmp_BSCmp_op2_1, b(0)=>
      gen_8_cmp_BSCmp_op2_0, carryIn=>gen_8_cmp_BSCmp_carryIn, sum(23)=>
      gen_8_cmp_pBs_30, sum(22)=>gen_8_cmp_pBs_29, sum(21)=>gen_8_cmp_pBs_28, 
      sum(20)=>gen_8_cmp_pBs_27, sum(19)=>gen_8_cmp_pBs_26, sum(18)=>
      gen_8_cmp_pBs_25, sum(17)=>gen_8_cmp_pBs_24, sum(16)=>gen_8_cmp_pBs_23, 
      sum(15)=>outputs_8_15, sum(14)=>outputs_8_14, sum(13)=>outputs_8_13, 
      sum(12)=>outputs_8_12, sum(11)=>outputs_8_11, sum(10)=>outputs_8_10, 
      sum(9)=>outputs_8_9, sum(8)=>outputs_8_8, sum(7)=>outputs_8_7, sum(6)
      =>outputs_8_6, sum(5)=>outputs_8_5, sum(4)=>outputs_8_4, sum(3)=>
      outputs_8_3, sum(2)=>outputs_8_2, sum(1)=>outputs_8_1, sum(0)=>
      outputs_8_0, carryOut=>DANGLING(84));
   gen_7_cmp_pRegCmp : Reg_33 port map ( D(32)=>working, D(31)=>working, 
      D(30)=>gen_7_cmp_pBs_30, D(29)=>gen_7_cmp_pBs_29, D(28)=>
      gen_7_cmp_pBs_28, D(27)=>gen_7_cmp_pBs_27, D(26)=>gen_7_cmp_pBs_26, 
      D(25)=>gen_7_cmp_pBs_25, D(24)=>gen_7_cmp_pBs_24, D(23)=>
      gen_7_cmp_pBs_23, D(22)=>outputs_7_15, D(21)=>outputs_7_14, D(20)=>
      outputs_7_13, D(19)=>outputs_7_12, D(18)=>outputs_7_11, D(17)=>
      outputs_7_10, D(16)=>outputs_7_9, D(15)=>outputs_7_8, D(14)=>
      outputs_7_7, D(13)=>outputs_7_6, D(12)=>outputs_7_5, D(11)=>
      outputs_7_4, D(10)=>outputs_7_3, D(9)=>outputs_7_2, D(8)=>outputs_7_1, 
      D(7)=>outputs_7_0, D(6)=>gen_7_cmp_pMux_8, D(5)=>gen_7_cmp_pMux_7, 
      D(4)=>gen_7_cmp_pMux_6, D(3)=>gen_7_cmp_pMux_5, D(2)=>gen_7_cmp_pMux_4, 
      D(1)=>gen_7_cmp_pMux_3, D(0)=>nx9603, en=>nx11169, clk=>nx9395, rst=>
      rst, Q(32)=>DANGLING(85), Q(31)=>DANGLING(86), Q(30)=>
      gen_7_cmp_pReg_30, Q(29)=>gen_7_cmp_pReg_29, Q(28)=>gen_7_cmp_pReg_28, 
      Q(27)=>gen_7_cmp_pReg_27, Q(26)=>gen_7_cmp_pReg_26, Q(25)=>
      gen_7_cmp_pReg_25, Q(24)=>gen_7_cmp_pReg_24, Q(23)=>gen_7_cmp_pReg_23, 
      Q(22)=>gen_7_cmp_pReg_22, Q(21)=>gen_7_cmp_pReg_21, Q(20)=>
      gen_7_cmp_pReg_20, Q(19)=>gen_7_cmp_pReg_19, Q(18)=>gen_7_cmp_pReg_18, 
      Q(17)=>gen_7_cmp_pReg_17, Q(16)=>gen_7_cmp_pReg_16, Q(15)=>
      gen_7_cmp_pReg_15, Q(14)=>gen_7_cmp_pReg_14, Q(13)=>gen_7_cmp_pReg_13, 
      Q(12)=>gen_7_cmp_pReg_12, Q(11)=>gen_7_cmp_pReg_11, Q(10)=>
      gen_7_cmp_pReg_10, Q(9)=>gen_7_cmp_pReg_9, Q(8)=>gen_7_cmp_pReg_8, 
      Q(7)=>gen_7_cmp_pReg_7, Q(6)=>gen_7_cmp_pReg_6, Q(5)=>gen_7_cmp_pReg_5, 
      Q(4)=>gen_7_cmp_pReg_4, Q(3)=>gen_7_cmp_pReg_3, Q(2)=>gen_7_cmp_pReg_2, 
      Q(1)=>gen_7_cmp_pReg_1, Q(0)=>gen_7_cmp_pReg_0);
   gen_7_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>working, a(31)=>working, 
      a(30)=>gen_7_cmp_pReg_30, a(29)=>gen_7_cmp_pReg_29, a(28)=>
      gen_7_cmp_pReg_28, a(27)=>gen_7_cmp_pReg_27, a(26)=>gen_7_cmp_pReg_26, 
      a(25)=>gen_7_cmp_pReg_25, a(24)=>gen_7_cmp_pReg_24, a(23)=>
      gen_7_cmp_pReg_23, a(22)=>gen_7_cmp_pReg_22, a(21)=>gen_7_cmp_pReg_21, 
      a(20)=>gen_7_cmp_pReg_20, a(19)=>gen_7_cmp_pReg_19, a(18)=>
      gen_7_cmp_pReg_18, a(17)=>gen_7_cmp_pReg_17, a(16)=>gen_7_cmp_pReg_16, 
      a(15)=>gen_7_cmp_pReg_15, a(14)=>gen_7_cmp_pReg_14, a(13)=>
      gen_7_cmp_pReg_13, a(12)=>gen_7_cmp_pReg_12, a(11)=>gen_7_cmp_pReg_11, 
      a(10)=>gen_7_cmp_pReg_10, a(9)=>gen_7_cmp_pReg_9, a(8)=>
      gen_7_cmp_pReg_8, a(7)=>gen_7_cmp_pReg_7, a(6)=>gen_7_cmp_pReg_6, a(5)
      =>gen_7_cmp_pReg_5, a(4)=>gen_7_cmp_pReg_4, a(3)=>gen_7_cmp_pReg_3, 
      a(2)=>gen_7_cmp_pReg_2, a(1)=>gen_7_cmp_pReg_1, a(0)=>gen_7_cmp_pReg_0, 
      b(32)=>working, b(31)=>working, b(30)=>working, b(29)=>working, b(28)
      =>working, b(27)=>working, b(26)=>working, b(25)=>working, b(24)=>
      working, b(23)=>working, b(22)=>working, b(21)=>working, b(20)=>
      working, b(19)=>working, b(18)=>working, b(17)=>working, b(16)=>
      working, b(15)=>working, b(14)=>working, b(13)=>working, b(12)=>
      working, b(11)=>working, b(10)=>working, b(9)=>working, b(8)=>
      filter_7_7, b(7)=>filter_7_6, b(6)=>filter_7_5, b(5)=>filter_7_4, b(4)
      =>filter_7_3, b(3)=>filter_7_2, b(2)=>filter_7_1, b(1)=>filter_7_0, 
      b(0)=>working, sel=>nx11187, f(32)=>DANGLING(87), f(31)=>DANGLING(88), 
      f(30)=>gen_7_cmp_pMux_30, f(29)=>gen_7_cmp_pMux_29, f(28)=>
      gen_7_cmp_pMux_28, f(27)=>gen_7_cmp_pMux_27, f(26)=>gen_7_cmp_pMux_26, 
      f(25)=>gen_7_cmp_pMux_25, f(24)=>gen_7_cmp_pMux_24, f(23)=>
      gen_7_cmp_pMux_23, f(22)=>gen_7_cmp_pMux_22, f(21)=>gen_7_cmp_pMux_21, 
      f(20)=>gen_7_cmp_pMux_20, f(19)=>gen_7_cmp_pMux_19, f(18)=>
      gen_7_cmp_pMux_18, f(17)=>gen_7_cmp_pMux_17, f(16)=>gen_7_cmp_pMux_16, 
      f(15)=>gen_7_cmp_pMux_15, f(14)=>gen_7_cmp_pMux_14, f(13)=>
      gen_7_cmp_pMux_13, f(12)=>gen_7_cmp_pMux_12, f(11)=>gen_7_cmp_pMux_11, 
      f(10)=>gen_7_cmp_pMux_10, f(9)=>gen_7_cmp_pMux_9, f(8)=>
      gen_7_cmp_pMux_8, f(7)=>gen_7_cmp_pMux_7, f(6)=>gen_7_cmp_pMux_6, f(5)
      =>gen_7_cmp_pMux_5, f(4)=>gen_7_cmp_pMux_4, f(3)=>gen_7_cmp_pMux_3, 
      f(2)=>gen_7_cmp_pMux_2, f(1)=>gen_7_cmp_pMux_1, f(0)=>gen_7_cmp_pMux_0
   );
   gen_7_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>working, a(22)
      =>working, a(21)=>gen_7_cmp_pMux_30, a(20)=>gen_7_cmp_pMux_29, a(19)=>
      gen_7_cmp_pMux_28, a(18)=>gen_7_cmp_pMux_27, a(17)=>gen_7_cmp_pMux_26, 
      a(16)=>gen_7_cmp_pMux_25, a(15)=>gen_7_cmp_pMux_24, a(14)=>
      gen_7_cmp_pMux_23, a(13)=>gen_7_cmp_pMux_22, a(12)=>gen_7_cmp_pMux_21, 
      a(11)=>gen_7_cmp_pMux_20, a(10)=>gen_7_cmp_pMux_19, a(9)=>
      gen_7_cmp_pMux_18, a(8)=>gen_7_cmp_pMux_17, a(7)=>gen_7_cmp_pMux_16, 
      a(6)=>gen_7_cmp_pMux_15, a(5)=>gen_7_cmp_pMux_14, a(4)=>
      gen_7_cmp_pMux_13, a(3)=>gen_7_cmp_pMux_12, a(2)=>gen_7_cmp_pMux_11, 
      a(1)=>gen_7_cmp_pMux_10, a(0)=>gen_7_cmp_pMux_9, b(23)=>nx9907, b(22)
      =>nx9907, b(21)=>nx9905, b(20)=>nx9913, b(19)=>nx9911, b(18)=>nx9909, 
      b(17)=>nx9907, b(16)=>nx9905, b(15)=>gen_7_cmp_BSCmp_op2_15, b(14)=>
      gen_7_cmp_BSCmp_op2_14, b(13)=>gen_7_cmp_BSCmp_op2_13, b(12)=>
      gen_7_cmp_BSCmp_op2_12, b(11)=>gen_7_cmp_BSCmp_op2_11, b(10)=>
      gen_7_cmp_BSCmp_op2_10, b(9)=>gen_7_cmp_BSCmp_op2_9, b(8)=>
      gen_7_cmp_BSCmp_op2_8, b(7)=>gen_7_cmp_BSCmp_op2_7, b(6)=>
      gen_7_cmp_BSCmp_op2_6, b(5)=>gen_7_cmp_BSCmp_op2_5, b(4)=>
      gen_7_cmp_BSCmp_op2_4, b(3)=>gen_7_cmp_BSCmp_op2_3, b(2)=>
      gen_7_cmp_BSCmp_op2_2, b(1)=>gen_7_cmp_BSCmp_op2_1, b(0)=>
      gen_7_cmp_BSCmp_op2_0, carryIn=>gen_7_cmp_BSCmp_carryIn, sum(23)=>
      gen_7_cmp_pBs_30, sum(22)=>gen_7_cmp_pBs_29, sum(21)=>gen_7_cmp_pBs_28, 
      sum(20)=>gen_7_cmp_pBs_27, sum(19)=>gen_7_cmp_pBs_26, sum(18)=>
      gen_7_cmp_pBs_25, sum(17)=>gen_7_cmp_pBs_24, sum(16)=>gen_7_cmp_pBs_23, 
      sum(15)=>outputs_7_15, sum(14)=>outputs_7_14, sum(13)=>outputs_7_13, 
      sum(12)=>outputs_7_12, sum(11)=>outputs_7_11, sum(10)=>outputs_7_10, 
      sum(9)=>outputs_7_9, sum(8)=>outputs_7_8, sum(7)=>outputs_7_7, sum(6)
      =>outputs_7_6, sum(5)=>outputs_7_5, sum(4)=>outputs_7_4, sum(3)=>
      outputs_7_3, sum(2)=>outputs_7_2, sum(1)=>outputs_7_1, sum(0)=>
      outputs_7_0, carryOut=>DANGLING(89));
   gen_6_cmp_pRegCmp : Reg_33 port map ( D(32)=>working, D(31)=>working, 
      D(30)=>gen_6_cmp_pBs_30, D(29)=>gen_6_cmp_pBs_29, D(28)=>
      gen_6_cmp_pBs_28, D(27)=>gen_6_cmp_pBs_27, D(26)=>gen_6_cmp_pBs_26, 
      D(25)=>gen_6_cmp_pBs_25, D(24)=>gen_6_cmp_pBs_24, D(23)=>
      gen_6_cmp_pBs_23, D(22)=>outputs_6_15, D(21)=>outputs_6_14, D(20)=>
      outputs_6_13, D(19)=>outputs_6_12, D(18)=>outputs_6_11, D(17)=>
      outputs_6_10, D(16)=>outputs_6_9, D(15)=>outputs_6_8, D(14)=>
      outputs_6_7, D(13)=>outputs_6_6, D(12)=>outputs_6_5, D(11)=>
      outputs_6_4, D(10)=>outputs_6_3, D(9)=>outputs_6_2, D(8)=>outputs_6_1, 
      D(7)=>outputs_6_0, D(6)=>gen_6_cmp_pMux_8, D(5)=>gen_6_cmp_pMux_7, 
      D(4)=>gen_6_cmp_pMux_6, D(3)=>gen_6_cmp_pMux_5, D(2)=>gen_6_cmp_pMux_4, 
      D(1)=>gen_6_cmp_pMux_3, D(0)=>nx9615, en=>nx11169, clk=>nx9395, rst=>
      rst, Q(32)=>DANGLING(90), Q(31)=>DANGLING(91), Q(30)=>
      gen_6_cmp_pReg_30, Q(29)=>gen_6_cmp_pReg_29, Q(28)=>gen_6_cmp_pReg_28, 
      Q(27)=>gen_6_cmp_pReg_27, Q(26)=>gen_6_cmp_pReg_26, Q(25)=>
      gen_6_cmp_pReg_25, Q(24)=>gen_6_cmp_pReg_24, Q(23)=>gen_6_cmp_pReg_23, 
      Q(22)=>gen_6_cmp_pReg_22, Q(21)=>gen_6_cmp_pReg_21, Q(20)=>
      gen_6_cmp_pReg_20, Q(19)=>gen_6_cmp_pReg_19, Q(18)=>gen_6_cmp_pReg_18, 
      Q(17)=>gen_6_cmp_pReg_17, Q(16)=>gen_6_cmp_pReg_16, Q(15)=>
      gen_6_cmp_pReg_15, Q(14)=>gen_6_cmp_pReg_14, Q(13)=>gen_6_cmp_pReg_13, 
      Q(12)=>gen_6_cmp_pReg_12, Q(11)=>gen_6_cmp_pReg_11, Q(10)=>
      gen_6_cmp_pReg_10, Q(9)=>gen_6_cmp_pReg_9, Q(8)=>gen_6_cmp_pReg_8, 
      Q(7)=>gen_6_cmp_pReg_7, Q(6)=>gen_6_cmp_pReg_6, Q(5)=>gen_6_cmp_pReg_5, 
      Q(4)=>gen_6_cmp_pReg_4, Q(3)=>gen_6_cmp_pReg_3, Q(2)=>gen_6_cmp_pReg_2, 
      Q(1)=>gen_6_cmp_pReg_1, Q(0)=>gen_6_cmp_pReg_0);
   gen_6_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>working, a(31)=>working, 
      a(30)=>gen_6_cmp_pReg_30, a(29)=>gen_6_cmp_pReg_29, a(28)=>
      gen_6_cmp_pReg_28, a(27)=>gen_6_cmp_pReg_27, a(26)=>gen_6_cmp_pReg_26, 
      a(25)=>gen_6_cmp_pReg_25, a(24)=>gen_6_cmp_pReg_24, a(23)=>
      gen_6_cmp_pReg_23, a(22)=>gen_6_cmp_pReg_22, a(21)=>gen_6_cmp_pReg_21, 
      a(20)=>gen_6_cmp_pReg_20, a(19)=>gen_6_cmp_pReg_19, a(18)=>
      gen_6_cmp_pReg_18, a(17)=>gen_6_cmp_pReg_17, a(16)=>gen_6_cmp_pReg_16, 
      a(15)=>gen_6_cmp_pReg_15, a(14)=>gen_6_cmp_pReg_14, a(13)=>
      gen_6_cmp_pReg_13, a(12)=>gen_6_cmp_pReg_12, a(11)=>gen_6_cmp_pReg_11, 
      a(10)=>gen_6_cmp_pReg_10, a(9)=>gen_6_cmp_pReg_9, a(8)=>
      gen_6_cmp_pReg_8, a(7)=>gen_6_cmp_pReg_7, a(6)=>gen_6_cmp_pReg_6, a(5)
      =>gen_6_cmp_pReg_5, a(4)=>gen_6_cmp_pReg_4, a(3)=>gen_6_cmp_pReg_3, 
      a(2)=>gen_6_cmp_pReg_2, a(1)=>gen_6_cmp_pReg_1, a(0)=>gen_6_cmp_pReg_0, 
      b(32)=>working, b(31)=>working, b(30)=>working, b(29)=>working, b(28)
      =>working, b(27)=>working, b(26)=>working, b(25)=>working, b(24)=>
      working, b(23)=>working, b(22)=>working, b(21)=>working, b(20)=>
      working, b(19)=>working, b(18)=>working, b(17)=>working, b(16)=>
      working, b(15)=>working, b(14)=>working, b(13)=>working, b(12)=>
      working, b(11)=>working, b(10)=>working, b(9)=>working, b(8)=>
      filter_6_7, b(7)=>filter_6_6, b(6)=>filter_6_5, b(5)=>filter_6_4, b(4)
      =>filter_6_3, b(3)=>filter_6_2, b(2)=>filter_6_1, b(1)=>filter_6_0, 
      b(0)=>working, sel=>nx11187, f(32)=>DANGLING(92), f(31)=>DANGLING(93), 
      f(30)=>gen_6_cmp_pMux_30, f(29)=>gen_6_cmp_pMux_29, f(28)=>
      gen_6_cmp_pMux_28, f(27)=>gen_6_cmp_pMux_27, f(26)=>gen_6_cmp_pMux_26, 
      f(25)=>gen_6_cmp_pMux_25, f(24)=>gen_6_cmp_pMux_24, f(23)=>
      gen_6_cmp_pMux_23, f(22)=>gen_6_cmp_pMux_22, f(21)=>gen_6_cmp_pMux_21, 
      f(20)=>gen_6_cmp_pMux_20, f(19)=>gen_6_cmp_pMux_19, f(18)=>
      gen_6_cmp_pMux_18, f(17)=>gen_6_cmp_pMux_17, f(16)=>gen_6_cmp_pMux_16, 
      f(15)=>gen_6_cmp_pMux_15, f(14)=>gen_6_cmp_pMux_14, f(13)=>
      gen_6_cmp_pMux_13, f(12)=>gen_6_cmp_pMux_12, f(11)=>gen_6_cmp_pMux_11, 
      f(10)=>gen_6_cmp_pMux_10, f(9)=>gen_6_cmp_pMux_9, f(8)=>
      gen_6_cmp_pMux_8, f(7)=>gen_6_cmp_pMux_7, f(6)=>gen_6_cmp_pMux_6, f(5)
      =>gen_6_cmp_pMux_5, f(4)=>gen_6_cmp_pMux_4, f(3)=>gen_6_cmp_pMux_3, 
      f(2)=>gen_6_cmp_pMux_2, f(1)=>gen_6_cmp_pMux_1, f(0)=>gen_6_cmp_pMux_0
   );
   gen_6_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>working, a(22)
      =>working, a(21)=>gen_6_cmp_pMux_30, a(20)=>gen_6_cmp_pMux_29, a(19)=>
      gen_6_cmp_pMux_28, a(18)=>gen_6_cmp_pMux_27, a(17)=>gen_6_cmp_pMux_26, 
      a(16)=>gen_6_cmp_pMux_25, a(15)=>gen_6_cmp_pMux_24, a(14)=>
      gen_6_cmp_pMux_23, a(13)=>gen_6_cmp_pMux_22, a(12)=>gen_6_cmp_pMux_21, 
      a(11)=>gen_6_cmp_pMux_20, a(10)=>gen_6_cmp_pMux_19, a(9)=>
      gen_6_cmp_pMux_18, a(8)=>gen_6_cmp_pMux_17, a(7)=>gen_6_cmp_pMux_16, 
      a(6)=>gen_6_cmp_pMux_15, a(5)=>gen_6_cmp_pMux_14, a(4)=>
      gen_6_cmp_pMux_13, a(3)=>gen_6_cmp_pMux_12, a(2)=>gen_6_cmp_pMux_11, 
      a(1)=>gen_6_cmp_pMux_10, a(0)=>gen_6_cmp_pMux_9, b(23)=>nx9919, b(22)
      =>nx9919, b(21)=>nx9917, b(20)=>nx9925, b(19)=>nx9923, b(18)=>nx9921, 
      b(17)=>nx9919, b(16)=>nx9917, b(15)=>gen_6_cmp_BSCmp_op2_15, b(14)=>
      gen_6_cmp_BSCmp_op2_14, b(13)=>gen_6_cmp_BSCmp_op2_13, b(12)=>
      gen_6_cmp_BSCmp_op2_12, b(11)=>gen_6_cmp_BSCmp_op2_11, b(10)=>
      gen_6_cmp_BSCmp_op2_10, b(9)=>gen_6_cmp_BSCmp_op2_9, b(8)=>
      gen_6_cmp_BSCmp_op2_8, b(7)=>gen_6_cmp_BSCmp_op2_7, b(6)=>
      gen_6_cmp_BSCmp_op2_6, b(5)=>gen_6_cmp_BSCmp_op2_5, b(4)=>
      gen_6_cmp_BSCmp_op2_4, b(3)=>gen_6_cmp_BSCmp_op2_3, b(2)=>
      gen_6_cmp_BSCmp_op2_2, b(1)=>gen_6_cmp_BSCmp_op2_1, b(0)=>
      gen_6_cmp_BSCmp_op2_0, carryIn=>gen_6_cmp_BSCmp_carryIn, sum(23)=>
      gen_6_cmp_pBs_30, sum(22)=>gen_6_cmp_pBs_29, sum(21)=>gen_6_cmp_pBs_28, 
      sum(20)=>gen_6_cmp_pBs_27, sum(19)=>gen_6_cmp_pBs_26, sum(18)=>
      gen_6_cmp_pBs_25, sum(17)=>gen_6_cmp_pBs_24, sum(16)=>gen_6_cmp_pBs_23, 
      sum(15)=>outputs_6_15, sum(14)=>outputs_6_14, sum(13)=>outputs_6_13, 
      sum(12)=>outputs_6_12, sum(11)=>outputs_6_11, sum(10)=>outputs_6_10, 
      sum(9)=>outputs_6_9, sum(8)=>outputs_6_8, sum(7)=>outputs_6_7, sum(6)
      =>outputs_6_6, sum(5)=>outputs_6_5, sum(4)=>outputs_6_4, sum(3)=>
      outputs_6_3, sum(2)=>outputs_6_2, sum(1)=>outputs_6_1, sum(0)=>
      outputs_6_0, carryOut=>DANGLING(94));
   gen_5_cmp_pRegCmp : Reg_33 port map ( D(32)=>working, D(31)=>working, 
      D(30)=>gen_5_cmp_pBs_30, D(29)=>gen_5_cmp_pBs_29, D(28)=>
      gen_5_cmp_pBs_28, D(27)=>gen_5_cmp_pBs_27, D(26)=>gen_5_cmp_pBs_26, 
      D(25)=>gen_5_cmp_pBs_25, D(24)=>gen_5_cmp_pBs_24, D(23)=>
      gen_5_cmp_pBs_23, D(22)=>outputs_5_15, D(21)=>outputs_5_14, D(20)=>
      outputs_5_13, D(19)=>outputs_5_12, D(18)=>outputs_5_11, D(17)=>
      outputs_5_10, D(16)=>outputs_5_9, D(15)=>outputs_5_8, D(14)=>
      outputs_5_7, D(13)=>outputs_5_6, D(12)=>outputs_5_5, D(11)=>
      outputs_5_4, D(10)=>outputs_5_3, D(9)=>outputs_5_2, D(8)=>outputs_5_1, 
      D(7)=>outputs_5_0, D(6)=>gen_5_cmp_pMux_8, D(5)=>gen_5_cmp_pMux_7, 
      D(4)=>gen_5_cmp_pMux_6, D(3)=>gen_5_cmp_pMux_5, D(2)=>gen_5_cmp_pMux_4, 
      D(1)=>gen_5_cmp_pMux_3, D(0)=>nx9627, en=>nx11169, clk=>nx9395, rst=>
      rst, Q(32)=>DANGLING(95), Q(31)=>DANGLING(96), Q(30)=>
      gen_5_cmp_pReg_30, Q(29)=>gen_5_cmp_pReg_29, Q(28)=>gen_5_cmp_pReg_28, 
      Q(27)=>gen_5_cmp_pReg_27, Q(26)=>gen_5_cmp_pReg_26, Q(25)=>
      gen_5_cmp_pReg_25, Q(24)=>gen_5_cmp_pReg_24, Q(23)=>gen_5_cmp_pReg_23, 
      Q(22)=>gen_5_cmp_pReg_22, Q(21)=>gen_5_cmp_pReg_21, Q(20)=>
      gen_5_cmp_pReg_20, Q(19)=>gen_5_cmp_pReg_19, Q(18)=>gen_5_cmp_pReg_18, 
      Q(17)=>gen_5_cmp_pReg_17, Q(16)=>gen_5_cmp_pReg_16, Q(15)=>
      gen_5_cmp_pReg_15, Q(14)=>gen_5_cmp_pReg_14, Q(13)=>gen_5_cmp_pReg_13, 
      Q(12)=>gen_5_cmp_pReg_12, Q(11)=>gen_5_cmp_pReg_11, Q(10)=>
      gen_5_cmp_pReg_10, Q(9)=>gen_5_cmp_pReg_9, Q(8)=>gen_5_cmp_pReg_8, 
      Q(7)=>gen_5_cmp_pReg_7, Q(6)=>gen_5_cmp_pReg_6, Q(5)=>gen_5_cmp_pReg_5, 
      Q(4)=>gen_5_cmp_pReg_4, Q(3)=>gen_5_cmp_pReg_3, Q(2)=>gen_5_cmp_pReg_2, 
      Q(1)=>gen_5_cmp_pReg_1, Q(0)=>gen_5_cmp_pReg_0);
   gen_5_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>working, a(31)=>working, 
      a(30)=>gen_5_cmp_pReg_30, a(29)=>gen_5_cmp_pReg_29, a(28)=>
      gen_5_cmp_pReg_28, a(27)=>gen_5_cmp_pReg_27, a(26)=>gen_5_cmp_pReg_26, 
      a(25)=>gen_5_cmp_pReg_25, a(24)=>gen_5_cmp_pReg_24, a(23)=>
      gen_5_cmp_pReg_23, a(22)=>gen_5_cmp_pReg_22, a(21)=>gen_5_cmp_pReg_21, 
      a(20)=>gen_5_cmp_pReg_20, a(19)=>gen_5_cmp_pReg_19, a(18)=>
      gen_5_cmp_pReg_18, a(17)=>gen_5_cmp_pReg_17, a(16)=>gen_5_cmp_pReg_16, 
      a(15)=>gen_5_cmp_pReg_15, a(14)=>gen_5_cmp_pReg_14, a(13)=>
      gen_5_cmp_pReg_13, a(12)=>gen_5_cmp_pReg_12, a(11)=>gen_5_cmp_pReg_11, 
      a(10)=>gen_5_cmp_pReg_10, a(9)=>gen_5_cmp_pReg_9, a(8)=>
      gen_5_cmp_pReg_8, a(7)=>gen_5_cmp_pReg_7, a(6)=>gen_5_cmp_pReg_6, a(5)
      =>gen_5_cmp_pReg_5, a(4)=>gen_5_cmp_pReg_4, a(3)=>gen_5_cmp_pReg_3, 
      a(2)=>gen_5_cmp_pReg_2, a(1)=>gen_5_cmp_pReg_1, a(0)=>gen_5_cmp_pReg_0, 
      b(32)=>working, b(31)=>working, b(30)=>working, b(29)=>working, b(28)
      =>working, b(27)=>working, b(26)=>working, b(25)=>working, b(24)=>
      working, b(23)=>working, b(22)=>working, b(21)=>working, b(20)=>
      working, b(19)=>working, b(18)=>working, b(17)=>working, b(16)=>
      working, b(15)=>working, b(14)=>working, b(13)=>working, b(12)=>
      working, b(11)=>working, b(10)=>working, b(9)=>working, b(8)=>
      filter_5_7, b(7)=>filter_5_6, b(6)=>filter_5_5, b(5)=>filter_5_4, b(4)
      =>filter_5_3, b(3)=>filter_5_2, b(2)=>filter_5_1, b(1)=>filter_5_0, 
      b(0)=>working, sel=>nx11187, f(32)=>DANGLING(97), f(31)=>DANGLING(98), 
      f(30)=>gen_5_cmp_pMux_30, f(29)=>gen_5_cmp_pMux_29, f(28)=>
      gen_5_cmp_pMux_28, f(27)=>gen_5_cmp_pMux_27, f(26)=>gen_5_cmp_pMux_26, 
      f(25)=>gen_5_cmp_pMux_25, f(24)=>gen_5_cmp_pMux_24, f(23)=>
      gen_5_cmp_pMux_23, f(22)=>gen_5_cmp_pMux_22, f(21)=>gen_5_cmp_pMux_21, 
      f(20)=>gen_5_cmp_pMux_20, f(19)=>gen_5_cmp_pMux_19, f(18)=>
      gen_5_cmp_pMux_18, f(17)=>gen_5_cmp_pMux_17, f(16)=>gen_5_cmp_pMux_16, 
      f(15)=>gen_5_cmp_pMux_15, f(14)=>gen_5_cmp_pMux_14, f(13)=>
      gen_5_cmp_pMux_13, f(12)=>gen_5_cmp_pMux_12, f(11)=>gen_5_cmp_pMux_11, 
      f(10)=>gen_5_cmp_pMux_10, f(9)=>gen_5_cmp_pMux_9, f(8)=>
      gen_5_cmp_pMux_8, f(7)=>gen_5_cmp_pMux_7, f(6)=>gen_5_cmp_pMux_6, f(5)
      =>gen_5_cmp_pMux_5, f(4)=>gen_5_cmp_pMux_4, f(3)=>gen_5_cmp_pMux_3, 
      f(2)=>gen_5_cmp_pMux_2, f(1)=>gen_5_cmp_pMux_1, f(0)=>gen_5_cmp_pMux_0
   );
   gen_5_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>working, a(22)
      =>working, a(21)=>gen_5_cmp_pMux_30, a(20)=>gen_5_cmp_pMux_29, a(19)=>
      gen_5_cmp_pMux_28, a(18)=>gen_5_cmp_pMux_27, a(17)=>gen_5_cmp_pMux_26, 
      a(16)=>gen_5_cmp_pMux_25, a(15)=>gen_5_cmp_pMux_24, a(14)=>
      gen_5_cmp_pMux_23, a(13)=>gen_5_cmp_pMux_22, a(12)=>gen_5_cmp_pMux_21, 
      a(11)=>gen_5_cmp_pMux_20, a(10)=>gen_5_cmp_pMux_19, a(9)=>
      gen_5_cmp_pMux_18, a(8)=>gen_5_cmp_pMux_17, a(7)=>gen_5_cmp_pMux_16, 
      a(6)=>gen_5_cmp_pMux_15, a(5)=>gen_5_cmp_pMux_14, a(4)=>
      gen_5_cmp_pMux_13, a(3)=>gen_5_cmp_pMux_12, a(2)=>gen_5_cmp_pMux_11, 
      a(1)=>gen_5_cmp_pMux_10, a(0)=>gen_5_cmp_pMux_9, b(23)=>nx9931, b(22)
      =>nx9931, b(21)=>nx9929, b(20)=>nx9937, b(19)=>nx9935, b(18)=>nx9933, 
      b(17)=>nx9931, b(16)=>nx9929, b(15)=>gen_5_cmp_BSCmp_op2_15, b(14)=>
      gen_5_cmp_BSCmp_op2_14, b(13)=>gen_5_cmp_BSCmp_op2_13, b(12)=>
      gen_5_cmp_BSCmp_op2_12, b(11)=>gen_5_cmp_BSCmp_op2_11, b(10)=>
      gen_5_cmp_BSCmp_op2_10, b(9)=>gen_5_cmp_BSCmp_op2_9, b(8)=>
      gen_5_cmp_BSCmp_op2_8, b(7)=>gen_5_cmp_BSCmp_op2_7, b(6)=>
      gen_5_cmp_BSCmp_op2_6, b(5)=>gen_5_cmp_BSCmp_op2_5, b(4)=>
      gen_5_cmp_BSCmp_op2_4, b(3)=>gen_5_cmp_BSCmp_op2_3, b(2)=>
      gen_5_cmp_BSCmp_op2_2, b(1)=>gen_5_cmp_BSCmp_op2_1, b(0)=>
      gen_5_cmp_BSCmp_op2_0, carryIn=>gen_5_cmp_BSCmp_carryIn, sum(23)=>
      gen_5_cmp_pBs_30, sum(22)=>gen_5_cmp_pBs_29, sum(21)=>gen_5_cmp_pBs_28, 
      sum(20)=>gen_5_cmp_pBs_27, sum(19)=>gen_5_cmp_pBs_26, sum(18)=>
      gen_5_cmp_pBs_25, sum(17)=>gen_5_cmp_pBs_24, sum(16)=>gen_5_cmp_pBs_23, 
      sum(15)=>outputs_5_15, sum(14)=>outputs_5_14, sum(13)=>outputs_5_13, 
      sum(12)=>outputs_5_12, sum(11)=>outputs_5_11, sum(10)=>outputs_5_10, 
      sum(9)=>outputs_5_9, sum(8)=>outputs_5_8, sum(7)=>outputs_5_7, sum(6)
      =>outputs_5_6, sum(5)=>outputs_5_5, sum(4)=>outputs_5_4, sum(3)=>
      outputs_5_3, sum(2)=>outputs_5_2, sum(1)=>outputs_5_1, sum(0)=>
      outputs_5_0, carryOut=>DANGLING(99));
   gen_4_cmp_pRegCmp : Reg_33 port map ( D(32)=>working, D(31)=>working, 
      D(30)=>gen_4_cmp_pBs_30, D(29)=>gen_4_cmp_pBs_29, D(28)=>
      gen_4_cmp_pBs_28, D(27)=>gen_4_cmp_pBs_27, D(26)=>gen_4_cmp_pBs_26, 
      D(25)=>gen_4_cmp_pBs_25, D(24)=>gen_4_cmp_pBs_24, D(23)=>
      gen_4_cmp_pBs_23, D(22)=>outputs_4_15, D(21)=>outputs_4_14, D(20)=>
      outputs_4_13, D(19)=>outputs_4_12, D(18)=>outputs_4_11, D(17)=>
      outputs_4_10, D(16)=>outputs_4_9, D(15)=>outputs_4_8, D(14)=>
      outputs_4_7, D(13)=>outputs_4_6, D(12)=>outputs_4_5, D(11)=>
      outputs_4_4, D(10)=>outputs_4_3, D(9)=>outputs_4_2, D(8)=>outputs_4_1, 
      D(7)=>outputs_4_0, D(6)=>gen_4_cmp_pMux_8, D(5)=>gen_4_cmp_pMux_7, 
      D(4)=>gen_4_cmp_pMux_6, D(3)=>gen_4_cmp_pMux_5, D(2)=>gen_4_cmp_pMux_4, 
      D(1)=>gen_4_cmp_pMux_3, D(0)=>nx9639, en=>nx9379, clk=>nx9395, rst=>
      rst, Q(32)=>DANGLING(100), Q(31)=>DANGLING(101), Q(30)=>
      gen_4_cmp_pReg_30, Q(29)=>gen_4_cmp_pReg_29, Q(28)=>gen_4_cmp_pReg_28, 
      Q(27)=>gen_4_cmp_pReg_27, Q(26)=>gen_4_cmp_pReg_26, Q(25)=>
      gen_4_cmp_pReg_25, Q(24)=>gen_4_cmp_pReg_24, Q(23)=>gen_4_cmp_pReg_23, 
      Q(22)=>gen_4_cmp_pReg_22, Q(21)=>gen_4_cmp_pReg_21, Q(20)=>
      gen_4_cmp_pReg_20, Q(19)=>gen_4_cmp_pReg_19, Q(18)=>gen_4_cmp_pReg_18, 
      Q(17)=>gen_4_cmp_pReg_17, Q(16)=>gen_4_cmp_pReg_16, Q(15)=>
      gen_4_cmp_pReg_15, Q(14)=>gen_4_cmp_pReg_14, Q(13)=>gen_4_cmp_pReg_13, 
      Q(12)=>gen_4_cmp_pReg_12, Q(11)=>gen_4_cmp_pReg_11, Q(10)=>
      gen_4_cmp_pReg_10, Q(9)=>gen_4_cmp_pReg_9, Q(8)=>gen_4_cmp_pReg_8, 
      Q(7)=>gen_4_cmp_pReg_7, Q(6)=>gen_4_cmp_pReg_6, Q(5)=>gen_4_cmp_pReg_5, 
      Q(4)=>gen_4_cmp_pReg_4, Q(3)=>gen_4_cmp_pReg_3, Q(2)=>gen_4_cmp_pReg_2, 
      Q(1)=>gen_4_cmp_pReg_1, Q(0)=>gen_4_cmp_pReg_0);
   gen_4_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>working, a(31)=>working, 
      a(30)=>gen_4_cmp_pReg_30, a(29)=>gen_4_cmp_pReg_29, a(28)=>
      gen_4_cmp_pReg_28, a(27)=>gen_4_cmp_pReg_27, a(26)=>gen_4_cmp_pReg_26, 
      a(25)=>gen_4_cmp_pReg_25, a(24)=>gen_4_cmp_pReg_24, a(23)=>
      gen_4_cmp_pReg_23, a(22)=>gen_4_cmp_pReg_22, a(21)=>gen_4_cmp_pReg_21, 
      a(20)=>gen_4_cmp_pReg_20, a(19)=>gen_4_cmp_pReg_19, a(18)=>
      gen_4_cmp_pReg_18, a(17)=>gen_4_cmp_pReg_17, a(16)=>gen_4_cmp_pReg_16, 
      a(15)=>gen_4_cmp_pReg_15, a(14)=>gen_4_cmp_pReg_14, a(13)=>
      gen_4_cmp_pReg_13, a(12)=>gen_4_cmp_pReg_12, a(11)=>gen_4_cmp_pReg_11, 
      a(10)=>gen_4_cmp_pReg_10, a(9)=>gen_4_cmp_pReg_9, a(8)=>
      gen_4_cmp_pReg_8, a(7)=>gen_4_cmp_pReg_7, a(6)=>gen_4_cmp_pReg_6, a(5)
      =>gen_4_cmp_pReg_5, a(4)=>gen_4_cmp_pReg_4, a(3)=>gen_4_cmp_pReg_3, 
      a(2)=>gen_4_cmp_pReg_2, a(1)=>gen_4_cmp_pReg_1, a(0)=>gen_4_cmp_pReg_0, 
      b(32)=>working, b(31)=>working, b(30)=>working, b(29)=>working, b(28)
      =>working, b(27)=>working, b(26)=>working, b(25)=>working, b(24)=>
      working, b(23)=>working, b(22)=>working, b(21)=>working, b(20)=>
      working, b(19)=>working, b(18)=>working, b(17)=>working, b(16)=>
      working, b(15)=>working, b(14)=>working, b(13)=>working, b(12)=>
      working, b(11)=>working, b(10)=>working, b(9)=>working, b(8)=>
      filter_4_7, b(7)=>filter_4_6, b(6)=>filter_4_5, b(5)=>filter_4_4, b(4)
      =>filter_4_3, b(3)=>filter_4_2, b(2)=>filter_4_1, b(1)=>filter_4_0, 
      b(0)=>working, sel=>nx11189, f(32)=>DANGLING(102), f(31)=>DANGLING(103
      ), f(30)=>gen_4_cmp_pMux_30, f(29)=>gen_4_cmp_pMux_29, f(28)=>
      gen_4_cmp_pMux_28, f(27)=>gen_4_cmp_pMux_27, f(26)=>gen_4_cmp_pMux_26, 
      f(25)=>gen_4_cmp_pMux_25, f(24)=>gen_4_cmp_pMux_24, f(23)=>
      gen_4_cmp_pMux_23, f(22)=>gen_4_cmp_pMux_22, f(21)=>gen_4_cmp_pMux_21, 
      f(20)=>gen_4_cmp_pMux_20, f(19)=>gen_4_cmp_pMux_19, f(18)=>
      gen_4_cmp_pMux_18, f(17)=>gen_4_cmp_pMux_17, f(16)=>gen_4_cmp_pMux_16, 
      f(15)=>gen_4_cmp_pMux_15, f(14)=>gen_4_cmp_pMux_14, f(13)=>
      gen_4_cmp_pMux_13, f(12)=>gen_4_cmp_pMux_12, f(11)=>gen_4_cmp_pMux_11, 
      f(10)=>gen_4_cmp_pMux_10, f(9)=>gen_4_cmp_pMux_9, f(8)=>
      gen_4_cmp_pMux_8, f(7)=>gen_4_cmp_pMux_7, f(6)=>gen_4_cmp_pMux_6, f(5)
      =>gen_4_cmp_pMux_5, f(4)=>gen_4_cmp_pMux_4, f(3)=>gen_4_cmp_pMux_3, 
      f(2)=>gen_4_cmp_pMux_2, f(1)=>gen_4_cmp_pMux_1, f(0)=>gen_4_cmp_pMux_0
   );
   gen_4_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>working, a(22)
      =>working, a(21)=>gen_4_cmp_pMux_30, a(20)=>gen_4_cmp_pMux_29, a(19)=>
      gen_4_cmp_pMux_28, a(18)=>gen_4_cmp_pMux_27, a(17)=>gen_4_cmp_pMux_26, 
      a(16)=>gen_4_cmp_pMux_25, a(15)=>gen_4_cmp_pMux_24, a(14)=>
      gen_4_cmp_pMux_23, a(13)=>gen_4_cmp_pMux_22, a(12)=>gen_4_cmp_pMux_21, 
      a(11)=>gen_4_cmp_pMux_20, a(10)=>gen_4_cmp_pMux_19, a(9)=>
      gen_4_cmp_pMux_18, a(8)=>gen_4_cmp_pMux_17, a(7)=>gen_4_cmp_pMux_16, 
      a(6)=>gen_4_cmp_pMux_15, a(5)=>gen_4_cmp_pMux_14, a(4)=>
      gen_4_cmp_pMux_13, a(3)=>gen_4_cmp_pMux_12, a(2)=>gen_4_cmp_pMux_11, 
      a(1)=>gen_4_cmp_pMux_10, a(0)=>gen_4_cmp_pMux_9, b(23)=>nx9943, b(22)
      =>nx9943, b(21)=>nx9941, b(20)=>nx9949, b(19)=>nx9947, b(18)=>nx9945, 
      b(17)=>nx9943, b(16)=>nx9941, b(15)=>gen_4_cmp_BSCmp_op2_15, b(14)=>
      gen_4_cmp_BSCmp_op2_14, b(13)=>gen_4_cmp_BSCmp_op2_13, b(12)=>
      gen_4_cmp_BSCmp_op2_12, b(11)=>gen_4_cmp_BSCmp_op2_11, b(10)=>
      gen_4_cmp_BSCmp_op2_10, b(9)=>gen_4_cmp_BSCmp_op2_9, b(8)=>
      gen_4_cmp_BSCmp_op2_8, b(7)=>gen_4_cmp_BSCmp_op2_7, b(6)=>
      gen_4_cmp_BSCmp_op2_6, b(5)=>gen_4_cmp_BSCmp_op2_5, b(4)=>
      gen_4_cmp_BSCmp_op2_4, b(3)=>gen_4_cmp_BSCmp_op2_3, b(2)=>
      gen_4_cmp_BSCmp_op2_2, b(1)=>gen_4_cmp_BSCmp_op2_1, b(0)=>
      gen_4_cmp_BSCmp_op2_0, carryIn=>gen_4_cmp_BSCmp_carryIn, sum(23)=>
      gen_4_cmp_pBs_30, sum(22)=>gen_4_cmp_pBs_29, sum(21)=>gen_4_cmp_pBs_28, 
      sum(20)=>gen_4_cmp_pBs_27, sum(19)=>gen_4_cmp_pBs_26, sum(18)=>
      gen_4_cmp_pBs_25, sum(17)=>gen_4_cmp_pBs_24, sum(16)=>gen_4_cmp_pBs_23, 
      sum(15)=>outputs_4_15, sum(14)=>outputs_4_14, sum(13)=>outputs_4_13, 
      sum(12)=>outputs_4_12, sum(11)=>outputs_4_11, sum(10)=>outputs_4_10, 
      sum(9)=>outputs_4_9, sum(8)=>outputs_4_8, sum(7)=>outputs_4_7, sum(6)
      =>outputs_4_6, sum(5)=>outputs_4_5, sum(4)=>outputs_4_4, sum(3)=>
      outputs_4_3, sum(2)=>outputs_4_2, sum(1)=>outputs_4_1, sum(0)=>
      outputs_4_0, carryOut=>DANGLING(104));
   gen_3_cmp_pRegCmp : Reg_33 port map ( D(32)=>working, D(31)=>working, 
      D(30)=>gen_3_cmp_pBs_30, D(29)=>gen_3_cmp_pBs_29, D(28)=>
      gen_3_cmp_pBs_28, D(27)=>gen_3_cmp_pBs_27, D(26)=>gen_3_cmp_pBs_26, 
      D(25)=>gen_3_cmp_pBs_25, D(24)=>gen_3_cmp_pBs_24, D(23)=>
      gen_3_cmp_pBs_23, D(22)=>outputs_3_15, D(21)=>outputs_3_14, D(20)=>
      outputs_3_13, D(19)=>outputs_3_12, D(18)=>outputs_3_11, D(17)=>
      outputs_3_10, D(16)=>outputs_3_9, D(15)=>outputs_3_8, D(14)=>
      outputs_3_7, D(13)=>outputs_3_6, D(12)=>outputs_3_5, D(11)=>
      outputs_3_4, D(10)=>outputs_3_3, D(9)=>outputs_3_2, D(8)=>outputs_3_1, 
      D(7)=>outputs_3_0, D(6)=>gen_3_cmp_pMux_8, D(5)=>gen_3_cmp_pMux_7, 
      D(4)=>gen_3_cmp_pMux_6, D(3)=>gen_3_cmp_pMux_5, D(2)=>gen_3_cmp_pMux_4, 
      D(1)=>gen_3_cmp_pMux_3, D(0)=>nx9651, en=>nx11171, clk=>nx9397, rst=>
      rst, Q(32)=>DANGLING(105), Q(31)=>DANGLING(106), Q(30)=>
      gen_3_cmp_pReg_30, Q(29)=>gen_3_cmp_pReg_29, Q(28)=>gen_3_cmp_pReg_28, 
      Q(27)=>gen_3_cmp_pReg_27, Q(26)=>gen_3_cmp_pReg_26, Q(25)=>
      gen_3_cmp_pReg_25, Q(24)=>gen_3_cmp_pReg_24, Q(23)=>gen_3_cmp_pReg_23, 
      Q(22)=>gen_3_cmp_pReg_22, Q(21)=>gen_3_cmp_pReg_21, Q(20)=>
      gen_3_cmp_pReg_20, Q(19)=>gen_3_cmp_pReg_19, Q(18)=>gen_3_cmp_pReg_18, 
      Q(17)=>gen_3_cmp_pReg_17, Q(16)=>gen_3_cmp_pReg_16, Q(15)=>
      gen_3_cmp_pReg_15, Q(14)=>gen_3_cmp_pReg_14, Q(13)=>gen_3_cmp_pReg_13, 
      Q(12)=>gen_3_cmp_pReg_12, Q(11)=>gen_3_cmp_pReg_11, Q(10)=>
      gen_3_cmp_pReg_10, Q(9)=>gen_3_cmp_pReg_9, Q(8)=>gen_3_cmp_pReg_8, 
      Q(7)=>gen_3_cmp_pReg_7, Q(6)=>gen_3_cmp_pReg_6, Q(5)=>gen_3_cmp_pReg_5, 
      Q(4)=>gen_3_cmp_pReg_4, Q(3)=>gen_3_cmp_pReg_3, Q(2)=>gen_3_cmp_pReg_2, 
      Q(1)=>gen_3_cmp_pReg_1, Q(0)=>gen_3_cmp_pReg_0);
   gen_3_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>working, a(31)=>working, 
      a(30)=>gen_3_cmp_pReg_30, a(29)=>gen_3_cmp_pReg_29, a(28)=>
      gen_3_cmp_pReg_28, a(27)=>gen_3_cmp_pReg_27, a(26)=>gen_3_cmp_pReg_26, 
      a(25)=>gen_3_cmp_pReg_25, a(24)=>gen_3_cmp_pReg_24, a(23)=>
      gen_3_cmp_pReg_23, a(22)=>gen_3_cmp_pReg_22, a(21)=>gen_3_cmp_pReg_21, 
      a(20)=>gen_3_cmp_pReg_20, a(19)=>gen_3_cmp_pReg_19, a(18)=>
      gen_3_cmp_pReg_18, a(17)=>gen_3_cmp_pReg_17, a(16)=>gen_3_cmp_pReg_16, 
      a(15)=>gen_3_cmp_pReg_15, a(14)=>gen_3_cmp_pReg_14, a(13)=>
      gen_3_cmp_pReg_13, a(12)=>gen_3_cmp_pReg_12, a(11)=>gen_3_cmp_pReg_11, 
      a(10)=>gen_3_cmp_pReg_10, a(9)=>gen_3_cmp_pReg_9, a(8)=>
      gen_3_cmp_pReg_8, a(7)=>gen_3_cmp_pReg_7, a(6)=>gen_3_cmp_pReg_6, a(5)
      =>gen_3_cmp_pReg_5, a(4)=>gen_3_cmp_pReg_4, a(3)=>gen_3_cmp_pReg_3, 
      a(2)=>gen_3_cmp_pReg_2, a(1)=>gen_3_cmp_pReg_1, a(0)=>gen_3_cmp_pReg_0, 
      b(32)=>working, b(31)=>working, b(30)=>working, b(29)=>working, b(28)
      =>working, b(27)=>working, b(26)=>working, b(25)=>working, b(24)=>
      working, b(23)=>working, b(22)=>working, b(21)=>working, b(20)=>
      working, b(19)=>working, b(18)=>working, b(17)=>working, b(16)=>
      working, b(15)=>working, b(14)=>working, b(13)=>working, b(12)=>
      working, b(11)=>working, b(10)=>working, b(9)=>working, b(8)=>
      filter_3_7, b(7)=>filter_3_6, b(6)=>filter_3_5, b(5)=>filter_3_4, b(4)
      =>filter_3_3, b(3)=>filter_3_2, b(2)=>filter_3_1, b(1)=>filter_3_0, 
      b(0)=>working, sel=>nx11191, f(32)=>DANGLING(107), f(31)=>DANGLING(108
      ), f(30)=>gen_3_cmp_pMux_30, f(29)=>gen_3_cmp_pMux_29, f(28)=>
      gen_3_cmp_pMux_28, f(27)=>gen_3_cmp_pMux_27, f(26)=>gen_3_cmp_pMux_26, 
      f(25)=>gen_3_cmp_pMux_25, f(24)=>gen_3_cmp_pMux_24, f(23)=>
      gen_3_cmp_pMux_23, f(22)=>gen_3_cmp_pMux_22, f(21)=>gen_3_cmp_pMux_21, 
      f(20)=>gen_3_cmp_pMux_20, f(19)=>gen_3_cmp_pMux_19, f(18)=>
      gen_3_cmp_pMux_18, f(17)=>gen_3_cmp_pMux_17, f(16)=>gen_3_cmp_pMux_16, 
      f(15)=>gen_3_cmp_pMux_15, f(14)=>gen_3_cmp_pMux_14, f(13)=>
      gen_3_cmp_pMux_13, f(12)=>gen_3_cmp_pMux_12, f(11)=>gen_3_cmp_pMux_11, 
      f(10)=>gen_3_cmp_pMux_10, f(9)=>gen_3_cmp_pMux_9, f(8)=>
      gen_3_cmp_pMux_8, f(7)=>gen_3_cmp_pMux_7, f(6)=>gen_3_cmp_pMux_6, f(5)
      =>gen_3_cmp_pMux_5, f(4)=>gen_3_cmp_pMux_4, f(3)=>gen_3_cmp_pMux_3, 
      f(2)=>gen_3_cmp_pMux_2, f(1)=>gen_3_cmp_pMux_1, f(0)=>gen_3_cmp_pMux_0
   );
   gen_3_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>working, a(22)
      =>working, a(21)=>gen_3_cmp_pMux_30, a(20)=>gen_3_cmp_pMux_29, a(19)=>
      gen_3_cmp_pMux_28, a(18)=>gen_3_cmp_pMux_27, a(17)=>gen_3_cmp_pMux_26, 
      a(16)=>gen_3_cmp_pMux_25, a(15)=>gen_3_cmp_pMux_24, a(14)=>
      gen_3_cmp_pMux_23, a(13)=>gen_3_cmp_pMux_22, a(12)=>gen_3_cmp_pMux_21, 
      a(11)=>gen_3_cmp_pMux_20, a(10)=>gen_3_cmp_pMux_19, a(9)=>
      gen_3_cmp_pMux_18, a(8)=>gen_3_cmp_pMux_17, a(7)=>gen_3_cmp_pMux_16, 
      a(6)=>gen_3_cmp_pMux_15, a(5)=>gen_3_cmp_pMux_14, a(4)=>
      gen_3_cmp_pMux_13, a(3)=>gen_3_cmp_pMux_12, a(2)=>gen_3_cmp_pMux_11, 
      a(1)=>gen_3_cmp_pMux_10, a(0)=>gen_3_cmp_pMux_9, b(23)=>nx9955, b(22)
      =>nx9955, b(21)=>nx9953, b(20)=>nx9961, b(19)=>nx9959, b(18)=>nx9957, 
      b(17)=>nx9955, b(16)=>nx9953, b(15)=>gen_3_cmp_BSCmp_op2_15, b(14)=>
      gen_3_cmp_BSCmp_op2_14, b(13)=>gen_3_cmp_BSCmp_op2_13, b(12)=>
      gen_3_cmp_BSCmp_op2_12, b(11)=>gen_3_cmp_BSCmp_op2_11, b(10)=>
      gen_3_cmp_BSCmp_op2_10, b(9)=>gen_3_cmp_BSCmp_op2_9, b(8)=>
      gen_3_cmp_BSCmp_op2_8, b(7)=>gen_3_cmp_BSCmp_op2_7, b(6)=>
      gen_3_cmp_BSCmp_op2_6, b(5)=>gen_3_cmp_BSCmp_op2_5, b(4)=>
      gen_3_cmp_BSCmp_op2_4, b(3)=>gen_3_cmp_BSCmp_op2_3, b(2)=>
      gen_3_cmp_BSCmp_op2_2, b(1)=>gen_3_cmp_BSCmp_op2_1, b(0)=>
      gen_3_cmp_BSCmp_op2_0, carryIn=>gen_3_cmp_BSCmp_carryIn, sum(23)=>
      gen_3_cmp_pBs_30, sum(22)=>gen_3_cmp_pBs_29, sum(21)=>gen_3_cmp_pBs_28, 
      sum(20)=>gen_3_cmp_pBs_27, sum(19)=>gen_3_cmp_pBs_26, sum(18)=>
      gen_3_cmp_pBs_25, sum(17)=>gen_3_cmp_pBs_24, sum(16)=>gen_3_cmp_pBs_23, 
      sum(15)=>outputs_3_15, sum(14)=>outputs_3_14, sum(13)=>outputs_3_13, 
      sum(12)=>outputs_3_12, sum(11)=>outputs_3_11, sum(10)=>outputs_3_10, 
      sum(9)=>outputs_3_9, sum(8)=>outputs_3_8, sum(7)=>outputs_3_7, sum(6)
      =>outputs_3_6, sum(5)=>outputs_3_5, sum(4)=>outputs_3_4, sum(3)=>
      outputs_3_3, sum(2)=>outputs_3_2, sum(1)=>outputs_3_1, sum(0)=>
      outputs_3_0, carryOut=>DANGLING(109));
   gen_2_cmp_pRegCmp : Reg_33 port map ( D(32)=>working, D(31)=>working, 
      D(30)=>gen_2_cmp_pBs_30, D(29)=>gen_2_cmp_pBs_29, D(28)=>
      gen_2_cmp_pBs_28, D(27)=>gen_2_cmp_pBs_27, D(26)=>gen_2_cmp_pBs_26, 
      D(25)=>gen_2_cmp_pBs_25, D(24)=>gen_2_cmp_pBs_24, D(23)=>
      gen_2_cmp_pBs_23, D(22)=>outputs_2_15, D(21)=>outputs_2_14, D(20)=>
      outputs_2_13, D(19)=>outputs_2_12, D(18)=>outputs_2_11, D(17)=>
      outputs_2_10, D(16)=>outputs_2_9, D(15)=>outputs_2_8, D(14)=>
      outputs_2_7, D(13)=>outputs_2_6, D(12)=>outputs_2_5, D(11)=>
      outputs_2_4, D(10)=>outputs_2_3, D(9)=>outputs_2_2, D(8)=>outputs_2_1, 
      D(7)=>outputs_2_0, D(6)=>gen_2_cmp_pMux_8, D(5)=>gen_2_cmp_pMux_7, 
      D(4)=>gen_2_cmp_pMux_6, D(3)=>gen_2_cmp_pMux_5, D(2)=>gen_2_cmp_pMux_4, 
      D(1)=>gen_2_cmp_pMux_3, D(0)=>nx9663, en=>nx11171, clk=>nx9397, rst=>
      rst, Q(32)=>DANGLING(110), Q(31)=>DANGLING(111), Q(30)=>
      gen_2_cmp_pReg_30, Q(29)=>gen_2_cmp_pReg_29, Q(28)=>gen_2_cmp_pReg_28, 
      Q(27)=>gen_2_cmp_pReg_27, Q(26)=>gen_2_cmp_pReg_26, Q(25)=>
      gen_2_cmp_pReg_25, Q(24)=>gen_2_cmp_pReg_24, Q(23)=>gen_2_cmp_pReg_23, 
      Q(22)=>gen_2_cmp_pReg_22, Q(21)=>gen_2_cmp_pReg_21, Q(20)=>
      gen_2_cmp_pReg_20, Q(19)=>gen_2_cmp_pReg_19, Q(18)=>gen_2_cmp_pReg_18, 
      Q(17)=>gen_2_cmp_pReg_17, Q(16)=>gen_2_cmp_pReg_16, Q(15)=>
      gen_2_cmp_pReg_15, Q(14)=>gen_2_cmp_pReg_14, Q(13)=>gen_2_cmp_pReg_13, 
      Q(12)=>gen_2_cmp_pReg_12, Q(11)=>gen_2_cmp_pReg_11, Q(10)=>
      gen_2_cmp_pReg_10, Q(9)=>gen_2_cmp_pReg_9, Q(8)=>gen_2_cmp_pReg_8, 
      Q(7)=>gen_2_cmp_pReg_7, Q(6)=>gen_2_cmp_pReg_6, Q(5)=>gen_2_cmp_pReg_5, 
      Q(4)=>gen_2_cmp_pReg_4, Q(3)=>gen_2_cmp_pReg_3, Q(2)=>gen_2_cmp_pReg_2, 
      Q(1)=>gen_2_cmp_pReg_1, Q(0)=>gen_2_cmp_pReg_0);
   gen_2_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>working, a(31)=>working, 
      a(30)=>gen_2_cmp_pReg_30, a(29)=>gen_2_cmp_pReg_29, a(28)=>
      gen_2_cmp_pReg_28, a(27)=>gen_2_cmp_pReg_27, a(26)=>gen_2_cmp_pReg_26, 
      a(25)=>gen_2_cmp_pReg_25, a(24)=>gen_2_cmp_pReg_24, a(23)=>
      gen_2_cmp_pReg_23, a(22)=>gen_2_cmp_pReg_22, a(21)=>gen_2_cmp_pReg_21, 
      a(20)=>gen_2_cmp_pReg_20, a(19)=>gen_2_cmp_pReg_19, a(18)=>
      gen_2_cmp_pReg_18, a(17)=>gen_2_cmp_pReg_17, a(16)=>gen_2_cmp_pReg_16, 
      a(15)=>gen_2_cmp_pReg_15, a(14)=>gen_2_cmp_pReg_14, a(13)=>
      gen_2_cmp_pReg_13, a(12)=>gen_2_cmp_pReg_12, a(11)=>gen_2_cmp_pReg_11, 
      a(10)=>gen_2_cmp_pReg_10, a(9)=>gen_2_cmp_pReg_9, a(8)=>
      gen_2_cmp_pReg_8, a(7)=>gen_2_cmp_pReg_7, a(6)=>gen_2_cmp_pReg_6, a(5)
      =>gen_2_cmp_pReg_5, a(4)=>gen_2_cmp_pReg_4, a(3)=>gen_2_cmp_pReg_3, 
      a(2)=>gen_2_cmp_pReg_2, a(1)=>gen_2_cmp_pReg_1, a(0)=>gen_2_cmp_pReg_0, 
      b(32)=>working, b(31)=>working, b(30)=>working, b(29)=>working, b(28)
      =>working, b(27)=>working, b(26)=>working, b(25)=>working, b(24)=>
      working, b(23)=>working, b(22)=>working, b(21)=>working, b(20)=>
      working, b(19)=>working, b(18)=>working, b(17)=>working, b(16)=>
      working, b(15)=>working, b(14)=>working, b(13)=>working, b(12)=>
      working, b(11)=>working, b(10)=>working, b(9)=>working, b(8)=>
      filter_2_7, b(7)=>filter_2_6, b(6)=>filter_2_5, b(5)=>filter_2_4, b(4)
      =>filter_2_3, b(3)=>filter_2_2, b(2)=>filter_2_1, b(1)=>filter_2_0, 
      b(0)=>working, sel=>nx11191, f(32)=>DANGLING(112), f(31)=>DANGLING(113
      ), f(30)=>gen_2_cmp_pMux_30, f(29)=>gen_2_cmp_pMux_29, f(28)=>
      gen_2_cmp_pMux_28, f(27)=>gen_2_cmp_pMux_27, f(26)=>gen_2_cmp_pMux_26, 
      f(25)=>gen_2_cmp_pMux_25, f(24)=>gen_2_cmp_pMux_24, f(23)=>
      gen_2_cmp_pMux_23, f(22)=>gen_2_cmp_pMux_22, f(21)=>gen_2_cmp_pMux_21, 
      f(20)=>gen_2_cmp_pMux_20, f(19)=>gen_2_cmp_pMux_19, f(18)=>
      gen_2_cmp_pMux_18, f(17)=>gen_2_cmp_pMux_17, f(16)=>gen_2_cmp_pMux_16, 
      f(15)=>gen_2_cmp_pMux_15, f(14)=>gen_2_cmp_pMux_14, f(13)=>
      gen_2_cmp_pMux_13, f(12)=>gen_2_cmp_pMux_12, f(11)=>gen_2_cmp_pMux_11, 
      f(10)=>gen_2_cmp_pMux_10, f(9)=>gen_2_cmp_pMux_9, f(8)=>
      gen_2_cmp_pMux_8, f(7)=>gen_2_cmp_pMux_7, f(6)=>gen_2_cmp_pMux_6, f(5)
      =>gen_2_cmp_pMux_5, f(4)=>gen_2_cmp_pMux_4, f(3)=>gen_2_cmp_pMux_3, 
      f(2)=>gen_2_cmp_pMux_2, f(1)=>gen_2_cmp_pMux_1, f(0)=>gen_2_cmp_pMux_0
   );
   gen_2_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>working, a(22)
      =>working, a(21)=>gen_2_cmp_pMux_30, a(20)=>gen_2_cmp_pMux_29, a(19)=>
      gen_2_cmp_pMux_28, a(18)=>gen_2_cmp_pMux_27, a(17)=>gen_2_cmp_pMux_26, 
      a(16)=>gen_2_cmp_pMux_25, a(15)=>gen_2_cmp_pMux_24, a(14)=>
      gen_2_cmp_pMux_23, a(13)=>gen_2_cmp_pMux_22, a(12)=>gen_2_cmp_pMux_21, 
      a(11)=>gen_2_cmp_pMux_20, a(10)=>gen_2_cmp_pMux_19, a(9)=>
      gen_2_cmp_pMux_18, a(8)=>gen_2_cmp_pMux_17, a(7)=>gen_2_cmp_pMux_16, 
      a(6)=>gen_2_cmp_pMux_15, a(5)=>gen_2_cmp_pMux_14, a(4)=>
      gen_2_cmp_pMux_13, a(3)=>gen_2_cmp_pMux_12, a(2)=>gen_2_cmp_pMux_11, 
      a(1)=>gen_2_cmp_pMux_10, a(0)=>gen_2_cmp_pMux_9, b(23)=>nx9967, b(22)
      =>nx9967, b(21)=>nx9965, b(20)=>nx9973, b(19)=>nx9971, b(18)=>nx9969, 
      b(17)=>nx9967, b(16)=>nx9965, b(15)=>gen_2_cmp_BSCmp_op2_15, b(14)=>
      gen_2_cmp_BSCmp_op2_14, b(13)=>gen_2_cmp_BSCmp_op2_13, b(12)=>
      gen_2_cmp_BSCmp_op2_12, b(11)=>gen_2_cmp_BSCmp_op2_11, b(10)=>
      gen_2_cmp_BSCmp_op2_10, b(9)=>gen_2_cmp_BSCmp_op2_9, b(8)=>
      gen_2_cmp_BSCmp_op2_8, b(7)=>gen_2_cmp_BSCmp_op2_7, b(6)=>
      gen_2_cmp_BSCmp_op2_6, b(5)=>gen_2_cmp_BSCmp_op2_5, b(4)=>
      gen_2_cmp_BSCmp_op2_4, b(3)=>gen_2_cmp_BSCmp_op2_3, b(2)=>
      gen_2_cmp_BSCmp_op2_2, b(1)=>gen_2_cmp_BSCmp_op2_1, b(0)=>
      gen_2_cmp_BSCmp_op2_0, carryIn=>gen_2_cmp_BSCmp_carryIn, sum(23)=>
      gen_2_cmp_pBs_30, sum(22)=>gen_2_cmp_pBs_29, sum(21)=>gen_2_cmp_pBs_28, 
      sum(20)=>gen_2_cmp_pBs_27, sum(19)=>gen_2_cmp_pBs_26, sum(18)=>
      gen_2_cmp_pBs_25, sum(17)=>gen_2_cmp_pBs_24, sum(16)=>gen_2_cmp_pBs_23, 
      sum(15)=>outputs_2_15, sum(14)=>outputs_2_14, sum(13)=>outputs_2_13, 
      sum(12)=>outputs_2_12, sum(11)=>outputs_2_11, sum(10)=>outputs_2_10, 
      sum(9)=>outputs_2_9, sum(8)=>outputs_2_8, sum(7)=>outputs_2_7, sum(6)
      =>outputs_2_6, sum(5)=>outputs_2_5, sum(4)=>outputs_2_4, sum(3)=>
      outputs_2_3, sum(2)=>outputs_2_2, sum(1)=>outputs_2_1, sum(0)=>
      outputs_2_0, carryOut=>DANGLING(114));
   gen_1_cmp_pRegCmp : Reg_33 port map ( D(32)=>working, D(31)=>working, 
      D(30)=>gen_1_cmp_pBs_30, D(29)=>gen_1_cmp_pBs_29, D(28)=>
      gen_1_cmp_pBs_28, D(27)=>gen_1_cmp_pBs_27, D(26)=>gen_1_cmp_pBs_26, 
      D(25)=>gen_1_cmp_pBs_25, D(24)=>gen_1_cmp_pBs_24, D(23)=>
      gen_1_cmp_pBs_23, D(22)=>outputs_1_15, D(21)=>outputs_1_14, D(20)=>
      outputs_1_13, D(19)=>outputs_1_12, D(18)=>outputs_1_11, D(17)=>
      outputs_1_10, D(16)=>outputs_1_9, D(15)=>outputs_1_8, D(14)=>
      outputs_1_7, D(13)=>outputs_1_6, D(12)=>outputs_1_5, D(11)=>
      outputs_1_4, D(10)=>outputs_1_3, D(9)=>outputs_1_2, D(8)=>outputs_1_1, 
      D(7)=>outputs_1_0, D(6)=>gen_1_cmp_pMux_8, D(5)=>gen_1_cmp_pMux_7, 
      D(4)=>gen_1_cmp_pMux_6, D(3)=>gen_1_cmp_pMux_5, D(2)=>gen_1_cmp_pMux_4, 
      D(1)=>gen_1_cmp_pMux_3, D(0)=>nx9675, en=>nx11171, clk=>nx9397, rst=>
      rst, Q(32)=>DANGLING(115), Q(31)=>DANGLING(116), Q(30)=>
      gen_1_cmp_pReg_30, Q(29)=>gen_1_cmp_pReg_29, Q(28)=>gen_1_cmp_pReg_28, 
      Q(27)=>gen_1_cmp_pReg_27, Q(26)=>gen_1_cmp_pReg_26, Q(25)=>
      gen_1_cmp_pReg_25, Q(24)=>gen_1_cmp_pReg_24, Q(23)=>gen_1_cmp_pReg_23, 
      Q(22)=>gen_1_cmp_pReg_22, Q(21)=>gen_1_cmp_pReg_21, Q(20)=>
      gen_1_cmp_pReg_20, Q(19)=>gen_1_cmp_pReg_19, Q(18)=>gen_1_cmp_pReg_18, 
      Q(17)=>gen_1_cmp_pReg_17, Q(16)=>gen_1_cmp_pReg_16, Q(15)=>
      gen_1_cmp_pReg_15, Q(14)=>gen_1_cmp_pReg_14, Q(13)=>gen_1_cmp_pReg_13, 
      Q(12)=>gen_1_cmp_pReg_12, Q(11)=>gen_1_cmp_pReg_11, Q(10)=>
      gen_1_cmp_pReg_10, Q(9)=>gen_1_cmp_pReg_9, Q(8)=>gen_1_cmp_pReg_8, 
      Q(7)=>gen_1_cmp_pReg_7, Q(6)=>gen_1_cmp_pReg_6, Q(5)=>gen_1_cmp_pReg_5, 
      Q(4)=>gen_1_cmp_pReg_4, Q(3)=>gen_1_cmp_pReg_3, Q(2)=>gen_1_cmp_pReg_2, 
      Q(1)=>gen_1_cmp_pReg_1, Q(0)=>gen_1_cmp_pReg_0);
   gen_1_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>working, a(31)=>working, 
      a(30)=>gen_1_cmp_pReg_30, a(29)=>gen_1_cmp_pReg_29, a(28)=>
      gen_1_cmp_pReg_28, a(27)=>gen_1_cmp_pReg_27, a(26)=>gen_1_cmp_pReg_26, 
      a(25)=>gen_1_cmp_pReg_25, a(24)=>gen_1_cmp_pReg_24, a(23)=>
      gen_1_cmp_pReg_23, a(22)=>gen_1_cmp_pReg_22, a(21)=>gen_1_cmp_pReg_21, 
      a(20)=>gen_1_cmp_pReg_20, a(19)=>gen_1_cmp_pReg_19, a(18)=>
      gen_1_cmp_pReg_18, a(17)=>gen_1_cmp_pReg_17, a(16)=>gen_1_cmp_pReg_16, 
      a(15)=>gen_1_cmp_pReg_15, a(14)=>gen_1_cmp_pReg_14, a(13)=>
      gen_1_cmp_pReg_13, a(12)=>gen_1_cmp_pReg_12, a(11)=>gen_1_cmp_pReg_11, 
      a(10)=>gen_1_cmp_pReg_10, a(9)=>gen_1_cmp_pReg_9, a(8)=>
      gen_1_cmp_pReg_8, a(7)=>gen_1_cmp_pReg_7, a(6)=>gen_1_cmp_pReg_6, a(5)
      =>gen_1_cmp_pReg_5, a(4)=>gen_1_cmp_pReg_4, a(3)=>gen_1_cmp_pReg_3, 
      a(2)=>gen_1_cmp_pReg_2, a(1)=>gen_1_cmp_pReg_1, a(0)=>gen_1_cmp_pReg_0, 
      b(32)=>working, b(31)=>working, b(30)=>working, b(29)=>working, b(28)
      =>working, b(27)=>working, b(26)=>working, b(25)=>working, b(24)=>
      working, b(23)=>working, b(22)=>working, b(21)=>working, b(20)=>
      working, b(19)=>working, b(18)=>working, b(17)=>working, b(16)=>
      working, b(15)=>working, b(14)=>working, b(13)=>working, b(12)=>
      working, b(11)=>working, b(10)=>working, b(9)=>working, b(8)=>
      filter_1_7, b(7)=>filter_1_6, b(6)=>filter_1_5, b(5)=>filter_1_4, b(4)
      =>filter_1_3, b(3)=>filter_1_2, b(2)=>filter_1_1, b(1)=>filter_1_0, 
      b(0)=>working, sel=>nx9389, f(32)=>DANGLING(117), f(31)=>DANGLING(118), 
      f(30)=>gen_1_cmp_pMux_30, f(29)=>gen_1_cmp_pMux_29, f(28)=>
      gen_1_cmp_pMux_28, f(27)=>gen_1_cmp_pMux_27, f(26)=>gen_1_cmp_pMux_26, 
      f(25)=>gen_1_cmp_pMux_25, f(24)=>gen_1_cmp_pMux_24, f(23)=>
      gen_1_cmp_pMux_23, f(22)=>gen_1_cmp_pMux_22, f(21)=>gen_1_cmp_pMux_21, 
      f(20)=>gen_1_cmp_pMux_20, f(19)=>gen_1_cmp_pMux_19, f(18)=>
      gen_1_cmp_pMux_18, f(17)=>gen_1_cmp_pMux_17, f(16)=>gen_1_cmp_pMux_16, 
      f(15)=>gen_1_cmp_pMux_15, f(14)=>gen_1_cmp_pMux_14, f(13)=>
      gen_1_cmp_pMux_13, f(12)=>gen_1_cmp_pMux_12, f(11)=>gen_1_cmp_pMux_11, 
      f(10)=>gen_1_cmp_pMux_10, f(9)=>gen_1_cmp_pMux_9, f(8)=>
      gen_1_cmp_pMux_8, f(7)=>gen_1_cmp_pMux_7, f(6)=>gen_1_cmp_pMux_6, f(5)
      =>gen_1_cmp_pMux_5, f(4)=>gen_1_cmp_pMux_4, f(3)=>gen_1_cmp_pMux_3, 
      f(2)=>gen_1_cmp_pMux_2, f(1)=>gen_1_cmp_pMux_1, f(0)=>gen_1_cmp_pMux_0
   );
   gen_1_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>working, a(22)
      =>working, a(21)=>gen_1_cmp_pMux_30, a(20)=>gen_1_cmp_pMux_29, a(19)=>
      gen_1_cmp_pMux_28, a(18)=>gen_1_cmp_pMux_27, a(17)=>gen_1_cmp_pMux_26, 
      a(16)=>gen_1_cmp_pMux_25, a(15)=>gen_1_cmp_pMux_24, a(14)=>
      gen_1_cmp_pMux_23, a(13)=>gen_1_cmp_pMux_22, a(12)=>gen_1_cmp_pMux_21, 
      a(11)=>gen_1_cmp_pMux_20, a(10)=>gen_1_cmp_pMux_19, a(9)=>
      gen_1_cmp_pMux_18, a(8)=>gen_1_cmp_pMux_17, a(7)=>gen_1_cmp_pMux_16, 
      a(6)=>gen_1_cmp_pMux_15, a(5)=>gen_1_cmp_pMux_14, a(4)=>
      gen_1_cmp_pMux_13, a(3)=>gen_1_cmp_pMux_12, a(2)=>gen_1_cmp_pMux_11, 
      a(1)=>gen_1_cmp_pMux_10, a(0)=>gen_1_cmp_pMux_9, b(23)=>nx9979, b(22)
      =>nx9979, b(21)=>nx9977, b(20)=>nx9985, b(19)=>nx9983, b(18)=>nx9981, 
      b(17)=>nx9979, b(16)=>nx9977, b(15)=>gen_1_cmp_BSCmp_op2_15, b(14)=>
      gen_1_cmp_BSCmp_op2_14, b(13)=>gen_1_cmp_BSCmp_op2_13, b(12)=>
      gen_1_cmp_BSCmp_op2_12, b(11)=>gen_1_cmp_BSCmp_op2_11, b(10)=>
      gen_1_cmp_BSCmp_op2_10, b(9)=>gen_1_cmp_BSCmp_op2_9, b(8)=>
      gen_1_cmp_BSCmp_op2_8, b(7)=>gen_1_cmp_BSCmp_op2_7, b(6)=>
      gen_1_cmp_BSCmp_op2_6, b(5)=>gen_1_cmp_BSCmp_op2_5, b(4)=>
      gen_1_cmp_BSCmp_op2_4, b(3)=>gen_1_cmp_BSCmp_op2_3, b(2)=>
      gen_1_cmp_BSCmp_op2_2, b(1)=>gen_1_cmp_BSCmp_op2_1, b(0)=>
      gen_1_cmp_BSCmp_op2_0, carryIn=>gen_1_cmp_BSCmp_carryIn, sum(23)=>
      gen_1_cmp_pBs_30, sum(22)=>gen_1_cmp_pBs_29, sum(21)=>gen_1_cmp_pBs_28, 
      sum(20)=>gen_1_cmp_pBs_27, sum(19)=>gen_1_cmp_pBs_26, sum(18)=>
      gen_1_cmp_pBs_25, sum(17)=>gen_1_cmp_pBs_24, sum(16)=>gen_1_cmp_pBs_23, 
      sum(15)=>outputs_1_15, sum(14)=>outputs_1_14, sum(13)=>outputs_1_13, 
      sum(12)=>outputs_1_12, sum(11)=>outputs_1_11, sum(10)=>outputs_1_10, 
      sum(9)=>outputs_1_9, sum(8)=>outputs_1_8, sum(7)=>outputs_1_7, sum(6)
      =>outputs_1_6, sum(5)=>outputs_1_5, sum(4)=>outputs_1_4, sum(3)=>
      outputs_1_3, sum(2)=>outputs_1_2, sum(1)=>outputs_1_1, sum(0)=>
      outputs_1_0, carryOut=>DANGLING(119));
   gen_0_cmp_pRegCmp : Reg_33 port map ( D(32)=>working, D(31)=>working, 
      D(30)=>gen_0_cmp_pBs_30, D(29)=>gen_0_cmp_pBs_29, D(28)=>
      gen_0_cmp_pBs_28, D(27)=>gen_0_cmp_pBs_27, D(26)=>gen_0_cmp_pBs_26, 
      D(25)=>gen_0_cmp_pBs_25, D(24)=>gen_0_cmp_pBs_24, D(23)=>
      gen_0_cmp_pBs_23, D(22)=>outputs_0_15, D(21)=>outputs_0_14, D(20)=>
      outputs_0_13, D(19)=>outputs_0_12, D(18)=>outputs_0_11, D(17)=>
      outputs_0_10, D(16)=>outputs_0_9, D(15)=>outputs_0_8, D(14)=>
      outputs_0_7, D(13)=>outputs_0_6, D(12)=>outputs_0_5, D(11)=>
      outputs_0_4, D(10)=>outputs_0_3, D(9)=>outputs_0_2, D(8)=>outputs_0_1, 
      D(7)=>outputs_0_0, D(6)=>gen_0_cmp_pMux_8, D(5)=>gen_0_cmp_pMux_7, 
      D(4)=>gen_0_cmp_pMux_6, D(3)=>gen_0_cmp_pMux_5, D(2)=>gen_0_cmp_pMux_4, 
      D(1)=>gen_0_cmp_pMux_3, D(0)=>nx9687, en=>nx9381, clk=>nx9397, rst=>
      rst, Q(32)=>DANGLING(120), Q(31)=>DANGLING(121), Q(30)=>
      gen_0_cmp_pReg_30, Q(29)=>gen_0_cmp_pReg_29, Q(28)=>gen_0_cmp_pReg_28, 
      Q(27)=>gen_0_cmp_pReg_27, Q(26)=>gen_0_cmp_pReg_26, Q(25)=>
      gen_0_cmp_pReg_25, Q(24)=>gen_0_cmp_pReg_24, Q(23)=>gen_0_cmp_pReg_23, 
      Q(22)=>gen_0_cmp_pReg_22, Q(21)=>gen_0_cmp_pReg_21, Q(20)=>
      gen_0_cmp_pReg_20, Q(19)=>gen_0_cmp_pReg_19, Q(18)=>gen_0_cmp_pReg_18, 
      Q(17)=>gen_0_cmp_pReg_17, Q(16)=>gen_0_cmp_pReg_16, Q(15)=>
      gen_0_cmp_pReg_15, Q(14)=>gen_0_cmp_pReg_14, Q(13)=>gen_0_cmp_pReg_13, 
      Q(12)=>gen_0_cmp_pReg_12, Q(11)=>gen_0_cmp_pReg_11, Q(10)=>
      gen_0_cmp_pReg_10, Q(9)=>gen_0_cmp_pReg_9, Q(8)=>gen_0_cmp_pReg_8, 
      Q(7)=>gen_0_cmp_pReg_7, Q(6)=>gen_0_cmp_pReg_6, Q(5)=>gen_0_cmp_pReg_5, 
      Q(4)=>gen_0_cmp_pReg_4, Q(3)=>gen_0_cmp_pReg_3, Q(2)=>gen_0_cmp_pReg_2, 
      Q(1)=>gen_0_cmp_pReg_1, Q(0)=>gen_0_cmp_pReg_0);
   gen_0_cmp_MuxCmp : BinaryMux_33 port map ( a(32)=>working, a(31)=>working, 
      a(30)=>gen_0_cmp_pReg_30, a(29)=>gen_0_cmp_pReg_29, a(28)=>
      gen_0_cmp_pReg_28, a(27)=>gen_0_cmp_pReg_27, a(26)=>gen_0_cmp_pReg_26, 
      a(25)=>gen_0_cmp_pReg_25, a(24)=>gen_0_cmp_pReg_24, a(23)=>
      gen_0_cmp_pReg_23, a(22)=>gen_0_cmp_pReg_22, a(21)=>gen_0_cmp_pReg_21, 
      a(20)=>gen_0_cmp_pReg_20, a(19)=>gen_0_cmp_pReg_19, a(18)=>
      gen_0_cmp_pReg_18, a(17)=>gen_0_cmp_pReg_17, a(16)=>gen_0_cmp_pReg_16, 
      a(15)=>gen_0_cmp_pReg_15, a(14)=>gen_0_cmp_pReg_14, a(13)=>
      gen_0_cmp_pReg_13, a(12)=>gen_0_cmp_pReg_12, a(11)=>gen_0_cmp_pReg_11, 
      a(10)=>gen_0_cmp_pReg_10, a(9)=>gen_0_cmp_pReg_9, a(8)=>
      gen_0_cmp_pReg_8, a(7)=>gen_0_cmp_pReg_7, a(6)=>gen_0_cmp_pReg_6, a(5)
      =>gen_0_cmp_pReg_5, a(4)=>gen_0_cmp_pReg_4, a(3)=>gen_0_cmp_pReg_3, 
      a(2)=>gen_0_cmp_pReg_2, a(1)=>gen_0_cmp_pReg_1, a(0)=>gen_0_cmp_pReg_0, 
      b(32)=>working, b(31)=>working, b(30)=>working, b(29)=>working, b(28)
      =>working, b(27)=>working, b(26)=>working, b(25)=>working, b(24)=>
      working, b(23)=>working, b(22)=>working, b(21)=>working, b(20)=>
      working, b(19)=>working, b(18)=>working, b(17)=>working, b(16)=>
      working, b(15)=>working, b(14)=>working, b(13)=>working, b(12)=>
      working, b(11)=>working, b(10)=>working, b(9)=>working, b(8)=>
      filter_0_7, b(7)=>filter_0_6, b(6)=>filter_0_5, b(5)=>filter_0_4, b(4)
      =>filter_0_3, b(3)=>filter_0_2, b(2)=>filter_0_1, b(1)=>filter_0_0, 
      b(0)=>working, sel=>nx9389, f(32)=>DANGLING(122), f(31)=>DANGLING(123), 
      f(30)=>gen_0_cmp_pMux_30, f(29)=>gen_0_cmp_pMux_29, f(28)=>
      gen_0_cmp_pMux_28, f(27)=>gen_0_cmp_pMux_27, f(26)=>gen_0_cmp_pMux_26, 
      f(25)=>gen_0_cmp_pMux_25, f(24)=>gen_0_cmp_pMux_24, f(23)=>
      gen_0_cmp_pMux_23, f(22)=>gen_0_cmp_pMux_22, f(21)=>gen_0_cmp_pMux_21, 
      f(20)=>gen_0_cmp_pMux_20, f(19)=>gen_0_cmp_pMux_19, f(18)=>
      gen_0_cmp_pMux_18, f(17)=>gen_0_cmp_pMux_17, f(16)=>gen_0_cmp_pMux_16, 
      f(15)=>gen_0_cmp_pMux_15, f(14)=>gen_0_cmp_pMux_14, f(13)=>
      gen_0_cmp_pMux_13, f(12)=>gen_0_cmp_pMux_12, f(11)=>gen_0_cmp_pMux_11, 
      f(10)=>gen_0_cmp_pMux_10, f(9)=>gen_0_cmp_pMux_9, f(8)=>
      gen_0_cmp_pMux_8, f(7)=>gen_0_cmp_pMux_7, f(6)=>gen_0_cmp_pMux_6, f(5)
      =>gen_0_cmp_pMux_5, f(4)=>gen_0_cmp_pMux_4, f(3)=>gen_0_cmp_pMux_3, 
      f(2)=>gen_0_cmp_pMux_2, f(1)=>gen_0_cmp_pMux_1, f(0)=>gen_0_cmp_pMux_0
   );
   gen_0_cmp_BSCmp_AdderCmp : NBitAdder_24 port map ( a(23)=>working, a(22)
      =>working, a(21)=>gen_0_cmp_pMux_30, a(20)=>gen_0_cmp_pMux_29, a(19)=>
      gen_0_cmp_pMux_28, a(18)=>gen_0_cmp_pMux_27, a(17)=>gen_0_cmp_pMux_26, 
      a(16)=>gen_0_cmp_pMux_25, a(15)=>gen_0_cmp_pMux_24, a(14)=>
      gen_0_cmp_pMux_23, a(13)=>gen_0_cmp_pMux_22, a(12)=>gen_0_cmp_pMux_21, 
      a(11)=>gen_0_cmp_pMux_20, a(10)=>gen_0_cmp_pMux_19, a(9)=>
      gen_0_cmp_pMux_18, a(8)=>gen_0_cmp_pMux_17, a(7)=>gen_0_cmp_pMux_16, 
      a(6)=>gen_0_cmp_pMux_15, a(5)=>gen_0_cmp_pMux_14, a(4)=>
      gen_0_cmp_pMux_13, a(3)=>gen_0_cmp_pMux_12, a(2)=>gen_0_cmp_pMux_11, 
      a(1)=>gen_0_cmp_pMux_10, a(0)=>gen_0_cmp_pMux_9, b(23)=>nx9991, b(22)
      =>nx9991, b(21)=>nx9989, b(20)=>nx9997, b(19)=>nx9995, b(18)=>nx9993, 
      b(17)=>nx9991, b(16)=>nx9989, b(15)=>gen_0_cmp_BSCmp_op2_15, b(14)=>
      gen_0_cmp_BSCmp_op2_14, b(13)=>gen_0_cmp_BSCmp_op2_13, b(12)=>
      gen_0_cmp_BSCmp_op2_12, b(11)=>gen_0_cmp_BSCmp_op2_11, b(10)=>
      gen_0_cmp_BSCmp_op2_10, b(9)=>gen_0_cmp_BSCmp_op2_9, b(8)=>
      gen_0_cmp_BSCmp_op2_8, b(7)=>gen_0_cmp_BSCmp_op2_7, b(6)=>
      gen_0_cmp_BSCmp_op2_6, b(5)=>gen_0_cmp_BSCmp_op2_5, b(4)=>
      gen_0_cmp_BSCmp_op2_4, b(3)=>gen_0_cmp_BSCmp_op2_3, b(2)=>
      gen_0_cmp_BSCmp_op2_2, b(1)=>gen_0_cmp_BSCmp_op2_1, b(0)=>
      gen_0_cmp_BSCmp_op2_0, carryIn=>gen_0_cmp_BSCmp_carryIn, sum(23)=>
      gen_0_cmp_pBs_30, sum(22)=>gen_0_cmp_pBs_29, sum(21)=>gen_0_cmp_pBs_28, 
      sum(20)=>gen_0_cmp_pBs_27, sum(19)=>gen_0_cmp_pBs_26, sum(18)=>
      gen_0_cmp_pBs_25, sum(17)=>gen_0_cmp_pBs_24, sum(16)=>gen_0_cmp_pBs_23, 
      sum(15)=>outputs_0_15, sum(14)=>outputs_0_14, sum(13)=>outputs_0_13, 
      sum(12)=>outputs_0_12, sum(11)=>outputs_0_11, sum(10)=>outputs_0_10, 
      sum(9)=>outputs_0_9, sum(8)=>outputs_0_8, sum(7)=>outputs_0_7, sum(6)
      =>outputs_0_6, sum(5)=>outputs_0_5, sum(4)=>outputs_0_4, sum(3)=>
      outputs_0_3, sum(2)=>outputs_0_2, sum(1)=>outputs_0_1, sum(0)=>
      outputs_0_0, carryOut=>DANGLING(124));
   ix9651 : fake_vcc port map ( Y=>nx9650);
   ix2325 : fake_gnd port map ( Y=>working);
   ix67 : nand02 port map ( Y=>gen_0_cmp_BSCmp_op2_1, A0=>nx2853, A1=>nx2873
   );
   ix2854 : nor02_2x port map ( Y=>nx2853, A0=>nx62, A1=>nx58);
   ix63 : nor03_2x port map ( Y=>nx62, A0=>gen_0_cmp_mReg_0, A1=>nx9693, A2
      =>nx10151);
   gen_0_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_0_cmp_mReg_0, QB=>
      nx2859, D=>window_0_0, CLK=>start, R=>rst);
   ix2864 : inv01 port map ( Y=>nx2862, A=>gen_0_cmp_pMux_0);
   ix59 : nor03_2x port map ( Y=>nx58, A0=>nx2859, A1=>nx10157, A2=>nx10167
   );
   ix2872 : inv02 port map ( Y=>nx2871, A=>gen_0_cmp_pMux_2);
   ix2874 : nor02_2x port map ( Y=>nx2873, A0=>nx48, A1=>nx46);
   ix49 : nor03_2x port map ( Y=>nx48, A0=>nx2877, A1=>nx9687, A2=>nx10175);
   gen_0_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_0_cmp_mReg_1, QB=>
      nx2877, D=>window_0_1, CLK=>start, R=>rst);
   ix47 : nor03_2x port map ( Y=>nx46, A0=>gen_0_cmp_mReg_1, A1=>nx9999, A2
      =>nx10183);
   ix7 : nor03_2x port map ( Y=>nx6, A0=>nx9693, A1=>nx2871, A2=>
      gen_0_cmp_pMux_0);
   ix89 : nand02 port map ( Y=>gen_0_cmp_BSCmp_op2_2, A0=>nx2887, A1=>nx2893
   );
   ix2888 : nor02_2x port map ( Y=>nx2887, A0=>nx84, A1=>nx80);
   ix85 : nor03_2x port map ( Y=>nx84, A0=>gen_0_cmp_mReg_1, A1=>nx9693, A2
      =>nx10151);
   ix81 : nor03_2x port map ( Y=>nx80, A0=>nx2877, A1=>nx10157, A2=>nx10167
   );
   ix2894 : nor02_2x port map ( Y=>nx2893, A0=>nx76, A1=>nx74);
   ix77 : nor03_2x port map ( Y=>nx76, A0=>nx2897, A1=>nx9687, A2=>nx10175);
   gen_0_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_0_cmp_mReg_2, QB=>
      nx2897, D=>window_0_2, CLK=>start, R=>rst);
   ix75 : nor03_2x port map ( Y=>nx74, A0=>gen_0_cmp_mReg_2, A1=>nx9999, A2
      =>nx10183);
   ix111 : nand02 port map ( Y=>gen_0_cmp_BSCmp_op2_3, A0=>nx2903, A1=>
      nx2907);
   ix2904 : nor02_2x port map ( Y=>nx2903, A0=>nx106, A1=>nx102);
   ix107 : nor03_2x port map ( Y=>nx106, A0=>gen_0_cmp_mReg_2, A1=>nx9693, 
      A2=>nx10151);
   ix103 : nor03_2x port map ( Y=>nx102, A0=>nx2897, A1=>nx10157, A2=>
      nx10167);
   ix2908 : nor02_2x port map ( Y=>nx2907, A0=>nx98, A1=>nx96);
   ix99 : nor03_2x port map ( Y=>nx98, A0=>nx2911, A1=>nx9687, A2=>nx10175);
   gen_0_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_0_cmp_mReg_3, QB=>
      nx2911, D=>window_0_3, CLK=>start, R=>rst);
   ix97 : nor03_2x port map ( Y=>nx96, A0=>gen_0_cmp_mReg_3, A1=>nx9999, A2
      =>nx10183);
   ix133 : nand02 port map ( Y=>gen_0_cmp_BSCmp_op2_4, A0=>nx2917, A1=>
      nx2923);
   ix2918 : nor02_2x port map ( Y=>nx2917, A0=>nx128, A1=>nx124);
   ix129 : nor03_2x port map ( Y=>nx128, A0=>gen_0_cmp_mReg_3, A1=>nx9693, 
      A2=>nx10151);
   ix125 : nor03_2x port map ( Y=>nx124, A0=>nx2911, A1=>nx10157, A2=>
      nx10167);
   ix2924 : nor02_2x port map ( Y=>nx2923, A0=>nx120, A1=>nx118);
   ix121 : nor03_2x port map ( Y=>nx120, A0=>nx2926, A1=>nx9687, A2=>nx10175
   );
   gen_0_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_0_cmp_mReg_4, QB=>
      nx2926, D=>window_0_4, CLK=>start, R=>rst);
   ix119 : nor03_2x port map ( Y=>nx118, A0=>gen_0_cmp_mReg_4, A1=>nx9999, 
      A2=>nx10183);
   ix155 : nand02 port map ( Y=>gen_0_cmp_BSCmp_op2_5, A0=>nx2931, A1=>
      nx2937);
   ix2932 : nor02_2x port map ( Y=>nx2931, A0=>nx150, A1=>nx146);
   ix151 : nor03_2x port map ( Y=>nx150, A0=>gen_0_cmp_mReg_4, A1=>nx9693, 
      A2=>nx10151);
   ix147 : nor03_2x port map ( Y=>nx146, A0=>nx2926, A1=>nx10157, A2=>
      nx10167);
   ix2938 : nor02_2x port map ( Y=>nx2937, A0=>nx142, A1=>nx140);
   ix143 : nor03_2x port map ( Y=>nx142, A0=>nx2941, A1=>nx9689, A2=>nx10175
   );
   gen_0_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_0_cmp_mReg_5, QB=>
      nx2941, D=>window_0_5, CLK=>start, R=>rst);
   ix141 : nor03_2x port map ( Y=>nx140, A0=>gen_0_cmp_mReg_5, A1=>nx9999, 
      A2=>nx10183);
   ix177 : nand02 port map ( Y=>gen_0_cmp_BSCmp_op2_6, A0=>nx2947, A1=>
      nx2951);
   ix2948 : nor02_2x port map ( Y=>nx2947, A0=>nx172, A1=>nx168);
   ix173 : nor03_2x port map ( Y=>nx172, A0=>gen_0_cmp_mReg_5, A1=>nx9695, 
      A2=>nx10151);
   ix169 : nor03_2x port map ( Y=>nx168, A0=>nx2941, A1=>nx10157, A2=>
      nx10167);
   ix2952 : nor02_2x port map ( Y=>nx2951, A0=>nx164, A1=>nx162);
   ix165 : nor03_2x port map ( Y=>nx164, A0=>nx2955, A1=>nx9689, A2=>nx10175
   );
   gen_0_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_0_cmp_mReg_6, QB=>
      nx2955, D=>window_0_6, CLK=>start, R=>rst);
   ix163 : nor03_2x port map ( Y=>nx162, A0=>gen_0_cmp_mReg_6, A1=>nx9999, 
      A2=>nx10183);
   ix199 : nand02 port map ( Y=>gen_0_cmp_BSCmp_op2_7, A0=>nx2961, A1=>
      nx2967);
   ix2962 : nor02_2x port map ( Y=>nx2961, A0=>nx194, A1=>nx190);
   ix195 : nor03_2x port map ( Y=>nx194, A0=>gen_0_cmp_mReg_6, A1=>nx9695, 
      A2=>nx10153);
   ix191 : nor03_2x port map ( Y=>nx190, A0=>nx2955, A1=>nx10159, A2=>
      nx10169);
   ix2968 : nor02_2x port map ( Y=>nx2967, A0=>nx186, A1=>nx184);
   ix187 : nor03_2x port map ( Y=>nx186, A0=>nx2970, A1=>nx9689, A2=>nx10177
   );
   gen_0_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_0_cmp_mReg_7, QB=>
      nx2970, D=>window_0_7, CLK=>start, R=>rst);
   ix185 : nor03_2x port map ( Y=>nx184, A0=>gen_0_cmp_mReg_7, A1=>nx9999, 
      A2=>nx10185);
   ix221 : nand02 port map ( Y=>gen_0_cmp_BSCmp_op2_8, A0=>nx2975, A1=>
      nx2981);
   ix2976 : nor02_2x port map ( Y=>nx2975, A0=>nx216, A1=>nx212);
   ix217 : nor03_2x port map ( Y=>nx216, A0=>gen_0_cmp_mReg_7, A1=>nx9695, 
      A2=>nx10153);
   ix213 : nor03_2x port map ( Y=>nx212, A0=>nx2970, A1=>nx10159, A2=>
      nx10169);
   ix2982 : nor02_2x port map ( Y=>nx2981, A0=>nx208, A1=>nx206);
   ix209 : nor03_2x port map ( Y=>nx208, A0=>nx2985, A1=>nx9689, A2=>nx10177
   );
   gen_0_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_0_cmp_mReg_8, QB=>
      nx2985, D=>window_0_8, CLK=>start, R=>rst);
   ix207 : nor03_2x port map ( Y=>nx206, A0=>gen_0_cmp_mReg_8, A1=>nx10001, 
      A2=>nx10185);
   ix243 : nand02 port map ( Y=>gen_0_cmp_BSCmp_op2_9, A0=>nx2991, A1=>
      nx2995);
   ix2992 : nor02_2x port map ( Y=>nx2991, A0=>nx238, A1=>nx234);
   ix239 : nor03_2x port map ( Y=>nx238, A0=>gen_0_cmp_mReg_8, A1=>nx9695, 
      A2=>nx10153);
   ix235 : nor03_2x port map ( Y=>nx234, A0=>nx2985, A1=>nx10159, A2=>
      nx10169);
   ix2996 : nor02_2x port map ( Y=>nx2995, A0=>nx230, A1=>nx228);
   ix231 : nor03_2x port map ( Y=>nx230, A0=>nx2999, A1=>nx9689, A2=>nx10177
   );
   gen_0_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_0_cmp_mReg_9, QB=>
      nx2999, D=>window_0_9, CLK=>start, R=>rst);
   ix229 : nor03_2x port map ( Y=>nx228, A0=>gen_0_cmp_mReg_9, A1=>nx10001, 
      A2=>nx10185);
   ix265 : nand02 port map ( Y=>gen_0_cmp_BSCmp_op2_10, A0=>nx3005, A1=>
      nx3011);
   ix3006 : nor02_2x port map ( Y=>nx3005, A0=>nx260, A1=>nx256);
   ix261 : nor03_2x port map ( Y=>nx260, A0=>gen_0_cmp_mReg_9, A1=>nx9695, 
      A2=>nx10153);
   ix257 : nor03_2x port map ( Y=>nx256, A0=>nx2999, A1=>nx10159, A2=>
      nx10169);
   ix3012 : nor02_2x port map ( Y=>nx3011, A0=>nx252, A1=>nx250);
   ix253 : nor03_2x port map ( Y=>nx252, A0=>nx3014, A1=>nx9689, A2=>nx10177
   );
   gen_0_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_0_cmp_mReg_10, QB=>
      nx3014, D=>window_0_10, CLK=>start, R=>rst);
   ix251 : nor03_2x port map ( Y=>nx250, A0=>gen_0_cmp_mReg_10, A1=>nx10001, 
      A2=>nx10185);
   ix287 : nand02 port map ( Y=>gen_0_cmp_BSCmp_op2_11, A0=>nx3019, A1=>
      nx3025);
   ix3020 : nor02_2x port map ( Y=>nx3019, A0=>nx282, A1=>nx278);
   ix283 : nor03_2x port map ( Y=>nx282, A0=>gen_0_cmp_mReg_10, A1=>nx9695, 
      A2=>nx10153);
   ix279 : nor03_2x port map ( Y=>nx278, A0=>nx3014, A1=>nx10159, A2=>
      nx10169);
   ix3026 : nor02_2x port map ( Y=>nx3025, A0=>nx274, A1=>nx272);
   ix275 : nor03_2x port map ( Y=>nx274, A0=>nx3029, A1=>nx9689, A2=>nx10177
   );
   gen_0_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_0_cmp_mReg_11, QB=>
      nx3029, D=>window_0_11, CLK=>start, R=>rst);
   ix273 : nor03_2x port map ( Y=>nx272, A0=>gen_0_cmp_mReg_11, A1=>nx10001, 
      A2=>nx10185);
   ix309 : nand02 port map ( Y=>gen_0_cmp_BSCmp_op2_12, A0=>nx3035, A1=>
      nx3039);
   ix3036 : nor02_2x port map ( Y=>nx3035, A0=>nx304, A1=>nx300);
   ix305 : nor03_2x port map ( Y=>nx304, A0=>gen_0_cmp_mReg_11, A1=>nx9695, 
      A2=>nx10153);
   ix301 : nor03_2x port map ( Y=>nx300, A0=>nx3029, A1=>nx10159, A2=>
      nx10169);
   ix3040 : nor02_2x port map ( Y=>nx3039, A0=>nx296, A1=>nx294);
   ix297 : nor03_2x port map ( Y=>nx296, A0=>nx3043, A1=>nx9691, A2=>nx10177
   );
   gen_0_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_0_cmp_mReg_12, QB=>
      nx3043, D=>window_0_12, CLK=>start, R=>rst);
   ix295 : nor03_2x port map ( Y=>nx294, A0=>gen_0_cmp_mReg_12, A1=>nx10001, 
      A2=>nx10185);
   ix331 : nand02 port map ( Y=>gen_0_cmp_BSCmp_op2_13, A0=>nx3049, A1=>
      nx3055);
   ix3050 : nor02_2x port map ( Y=>nx3049, A0=>nx326, A1=>nx322);
   ix327 : nor03_2x port map ( Y=>nx326, A0=>gen_0_cmp_mReg_12, A1=>nx9697, 
      A2=>nx10155);
   ix323 : nor03_2x port map ( Y=>nx322, A0=>nx3043, A1=>nx10159, A2=>
      nx10171);
   ix3056 : nor02_2x port map ( Y=>nx3055, A0=>nx318, A1=>nx316);
   ix319 : nor03_2x port map ( Y=>nx318, A0=>nx3058, A1=>nx9691, A2=>nx10179
   );
   gen_0_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_0_cmp_mReg_13, QB=>
      nx3058, D=>window_0_13, CLK=>start, R=>rst);
   ix317 : nor03_2x port map ( Y=>nx316, A0=>gen_0_cmp_mReg_13, A1=>nx10001, 
      A2=>nx10187);
   ix353 : nand02 port map ( Y=>gen_0_cmp_BSCmp_op2_14, A0=>nx3063, A1=>
      nx3069);
   ix3064 : nor02_2x port map ( Y=>nx3063, A0=>nx348, A1=>nx344);
   ix349 : nor03_2x port map ( Y=>nx348, A0=>gen_0_cmp_mReg_13, A1=>nx9697, 
      A2=>nx10155);
   ix345 : nor03_2x port map ( Y=>nx344, A0=>nx3058, A1=>nx10161, A2=>
      nx10171);
   ix3070 : nor02_2x port map ( Y=>nx3069, A0=>nx340, A1=>nx338);
   ix341 : nor03_2x port map ( Y=>nx340, A0=>nx3073, A1=>nx9691, A2=>nx10179
   );
   gen_0_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_0_cmp_mReg_14, QB=>
      nx3073, D=>window_0_14, CLK=>start, R=>rst);
   ix339 : nor03_2x port map ( Y=>nx338, A0=>gen_0_cmp_mReg_14, A1=>nx10001, 
      A2=>nx10187);
   ix375 : nand02 port map ( Y=>gen_0_cmp_BSCmp_op2_15, A0=>nx3079, A1=>
      nx3083);
   ix3080 : nor02_2x port map ( Y=>nx3079, A0=>nx370, A1=>nx366);
   ix371 : nor03_2x port map ( Y=>nx370, A0=>gen_0_cmp_mReg_14, A1=>nx9697, 
      A2=>nx10155);
   ix367 : nor03_2x port map ( Y=>nx366, A0=>nx3073, A1=>nx10161, A2=>
      nx10171);
   ix3084 : nor02_2x port map ( Y=>nx3083, A0=>nx362, A1=>nx360);
   ix363 : nor03_2x port map ( Y=>nx362, A0=>nx3087, A1=>nx9691, A2=>nx10179
   );
   gen_0_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_0_cmp_mReg_15, QB=>
      nx3087, D=>window_0_15, CLK=>start, R=>rst);
   ix361 : nor03_2x port map ( Y=>nx360, A0=>gen_0_cmp_mReg_15, A1=>nx10003, 
      A2=>nx10187);
   ix385 : nand02 port map ( Y=>gen_0_cmp_BSCmp_op2_16, A0=>nx3093, A1=>
      nx3083);
   ix3094 : nor02_2x port map ( Y=>nx3093, A0=>nx380, A1=>nx376);
   ix381 : nor03_2x port map ( Y=>nx380, A0=>gen_0_cmp_mReg_15, A1=>nx9697, 
      A2=>nx10155);
   ix377 : nor03_2x port map ( Y=>nx376, A0=>nx3087, A1=>nx10161, A2=>
      nx10171);
   ix453 : nand02 port map ( Y=>gen_1_cmp_BSCmp_op2_1, A0=>nx3099, A1=>
      nx3117);
   ix3100 : nor02_2x port map ( Y=>nx3099, A0=>nx448, A1=>nx444);
   ix449 : nor03_2x port map ( Y=>nx448, A0=>gen_1_cmp_mReg_0, A1=>nx9681, 
      A2=>nx10191);
   gen_1_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_1_cmp_mReg_0, QB=>
      nx3103, D=>window_1_0, CLK=>start, R=>rst);
   ix3108 : inv01 port map ( Y=>nx3107, A=>gen_1_cmp_pMux_0);
   ix445 : nor03_2x port map ( Y=>nx444, A0=>nx3103, A1=>nx10197, A2=>
      nx10207);
   ix3116 : inv02 port map ( Y=>nx3115, A=>gen_1_cmp_pMux_2);
   ix3118 : nor02_2x port map ( Y=>nx3117, A0=>nx434, A1=>nx432);
   ix435 : nor03_2x port map ( Y=>nx434, A0=>nx3121, A1=>nx9675, A2=>nx10215
   );
   gen_1_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_1_cmp_mReg_1, QB=>
      nx3121, D=>window_1_1, CLK=>start, R=>rst);
   ix433 : nor03_2x port map ( Y=>nx432, A0=>gen_1_cmp_mReg_1, A1=>nx10005, 
      A2=>nx10223);
   ix393 : nor03_2x port map ( Y=>nx392, A0=>nx9681, A1=>nx3115, A2=>
      gen_1_cmp_pMux_0);
   ix475 : nand02 port map ( Y=>gen_1_cmp_BSCmp_op2_2, A0=>nx3132, A1=>
      nx3139);
   ix3134 : nor02_2x port map ( Y=>nx3132, A0=>nx470, A1=>nx466);
   ix471 : nor03_2x port map ( Y=>nx470, A0=>gen_1_cmp_mReg_1, A1=>nx9681, 
      A2=>nx10191);
   ix467 : nor03_2x port map ( Y=>nx466, A0=>nx3121, A1=>nx10197, A2=>
      nx10207);
   ix3140 : nor02_2x port map ( Y=>nx3139, A0=>nx462, A1=>nx460);
   ix463 : nor03_2x port map ( Y=>nx462, A0=>nx3143, A1=>nx9675, A2=>nx10215
   );
   gen_1_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_1_cmp_mReg_2, QB=>
      nx3143, D=>window_1_2, CLK=>start, R=>rst);
   ix461 : nor03_2x port map ( Y=>nx460, A0=>gen_1_cmp_mReg_2, A1=>nx10005, 
      A2=>nx10223);
   ix497 : nand02 port map ( Y=>gen_1_cmp_BSCmp_op2_3, A0=>nx3149, A1=>
      nx3155);
   ix3150 : nor02_2x port map ( Y=>nx3149, A0=>nx492, A1=>nx488);
   ix493 : nor03_2x port map ( Y=>nx492, A0=>gen_1_cmp_mReg_2, A1=>nx9681, 
      A2=>nx10191);
   ix489 : nor03_2x port map ( Y=>nx488, A0=>nx3143, A1=>nx10197, A2=>
      nx10207);
   ix3156 : nor02_2x port map ( Y=>nx3155, A0=>nx484, A1=>nx482);
   ix485 : nor03_2x port map ( Y=>nx484, A0=>nx3158, A1=>nx9675, A2=>nx10215
   );
   gen_1_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_1_cmp_mReg_3, QB=>
      nx3158, D=>window_1_3, CLK=>start, R=>rst);
   ix483 : nor03_2x port map ( Y=>nx482, A0=>gen_1_cmp_mReg_3, A1=>nx10005, 
      A2=>nx10223);
   ix519 : nand02 port map ( Y=>gen_1_cmp_BSCmp_op2_4, A0=>nx3163, A1=>
      nx3169);
   ix3164 : nor02_2x port map ( Y=>nx3163, A0=>nx514, A1=>nx510);
   ix515 : nor03_2x port map ( Y=>nx514, A0=>gen_1_cmp_mReg_3, A1=>nx9681, 
      A2=>nx10191);
   ix511 : nor03_2x port map ( Y=>nx510, A0=>nx3158, A1=>nx10197, A2=>
      nx10207);
   ix3170 : nor02_2x port map ( Y=>nx3169, A0=>nx506, A1=>nx504);
   ix507 : nor03_2x port map ( Y=>nx506, A0=>nx3173, A1=>nx9675, A2=>nx10215
   );
   gen_1_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_1_cmp_mReg_4, QB=>
      nx3173, D=>window_1_4, CLK=>start, R=>rst);
   ix505 : nor03_2x port map ( Y=>nx504, A0=>gen_1_cmp_mReg_4, A1=>nx10005, 
      A2=>nx10223);
   ix541 : nand02 port map ( Y=>gen_1_cmp_BSCmp_op2_5, A0=>nx3179, A1=>
      nx3183);
   ix3180 : nor02_2x port map ( Y=>nx3179, A0=>nx536, A1=>nx532);
   ix537 : nor03_2x port map ( Y=>nx536, A0=>gen_1_cmp_mReg_4, A1=>nx9681, 
      A2=>nx10191);
   ix533 : nor03_2x port map ( Y=>nx532, A0=>nx3173, A1=>nx10197, A2=>
      nx10207);
   ix3184 : nor02_2x port map ( Y=>nx3183, A0=>nx528, A1=>nx526);
   ix529 : nor03_2x port map ( Y=>nx528, A0=>nx3187, A1=>nx9677, A2=>nx10215
   );
   gen_1_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_1_cmp_mReg_5, QB=>
      nx3187, D=>window_1_5, CLK=>start, R=>rst);
   ix527 : nor03_2x port map ( Y=>nx526, A0=>gen_1_cmp_mReg_5, A1=>nx10005, 
      A2=>nx10223);
   ix563 : nand02 port map ( Y=>gen_1_cmp_BSCmp_op2_6, A0=>nx3193, A1=>
      nx3199);
   ix3194 : nor02_2x port map ( Y=>nx3193, A0=>nx558, A1=>nx554);
   ix559 : nor03_2x port map ( Y=>nx558, A0=>gen_1_cmp_mReg_5, A1=>nx9683, 
      A2=>nx10191);
   ix555 : nor03_2x port map ( Y=>nx554, A0=>nx3187, A1=>nx10197, A2=>
      nx10207);
   ix3200 : nor02_2x port map ( Y=>nx3199, A0=>nx550, A1=>nx548);
   ix551 : nor03_2x port map ( Y=>nx550, A0=>nx3202, A1=>nx9677, A2=>nx10215
   );
   gen_1_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_1_cmp_mReg_6, QB=>
      nx3202, D=>window_1_6, CLK=>start, R=>rst);
   ix549 : nor03_2x port map ( Y=>nx548, A0=>gen_1_cmp_mReg_6, A1=>nx10005, 
      A2=>nx10223);
   ix585 : nand02 port map ( Y=>gen_1_cmp_BSCmp_op2_7, A0=>nx3207, A1=>
      nx3213);
   ix3208 : nor02_2x port map ( Y=>nx3207, A0=>nx580, A1=>nx576);
   ix581 : nor03_2x port map ( Y=>nx580, A0=>gen_1_cmp_mReg_6, A1=>nx9683, 
      A2=>nx10193);
   ix577 : nor03_2x port map ( Y=>nx576, A0=>nx3202, A1=>nx10199, A2=>
      nx10209);
   ix3214 : nor02_2x port map ( Y=>nx3213, A0=>nx572, A1=>nx570);
   ix573 : nor03_2x port map ( Y=>nx572, A0=>nx3217, A1=>nx9677, A2=>nx10217
   );
   gen_1_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_1_cmp_mReg_7, QB=>
      nx3217, D=>window_1_7, CLK=>start, R=>rst);
   ix571 : nor03_2x port map ( Y=>nx570, A0=>gen_1_cmp_mReg_7, A1=>nx10005, 
      A2=>nx10225);
   ix607 : nand02 port map ( Y=>gen_1_cmp_BSCmp_op2_8, A0=>nx3223, A1=>
      nx3227);
   ix3224 : nor02_2x port map ( Y=>nx3223, A0=>nx602, A1=>nx598);
   ix603 : nor03_2x port map ( Y=>nx602, A0=>gen_1_cmp_mReg_7, A1=>nx9683, 
      A2=>nx10193);
   ix599 : nor03_2x port map ( Y=>nx598, A0=>nx3217, A1=>nx10199, A2=>
      nx10209);
   ix3228 : nor02_2x port map ( Y=>nx3227, A0=>nx594, A1=>nx592);
   ix595 : nor03_2x port map ( Y=>nx594, A0=>nx3231, A1=>nx9677, A2=>nx10217
   );
   gen_1_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_1_cmp_mReg_8, QB=>
      nx3231, D=>window_1_8, CLK=>start, R=>rst);
   ix593 : nor03_2x port map ( Y=>nx592, A0=>gen_1_cmp_mReg_8, A1=>nx10007, 
      A2=>nx10225);
   ix629 : nand02 port map ( Y=>gen_1_cmp_BSCmp_op2_9, A0=>nx3237, A1=>
      nx3243);
   ix3238 : nor02_2x port map ( Y=>nx3237, A0=>nx624, A1=>nx620);
   ix625 : nor03_2x port map ( Y=>nx624, A0=>gen_1_cmp_mReg_8, A1=>nx9683, 
      A2=>nx10193);
   ix621 : nor03_2x port map ( Y=>nx620, A0=>nx3231, A1=>nx10199, A2=>
      nx10209);
   ix3244 : nor02_2x port map ( Y=>nx3243, A0=>nx616, A1=>nx614);
   ix617 : nor03_2x port map ( Y=>nx616, A0=>nx3246, A1=>nx9677, A2=>nx10217
   );
   gen_1_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_1_cmp_mReg_9, QB=>
      nx3246, D=>window_1_9, CLK=>start, R=>rst);
   ix615 : nor03_2x port map ( Y=>nx614, A0=>gen_1_cmp_mReg_9, A1=>nx10007, 
      A2=>nx10225);
   ix651 : nand02 port map ( Y=>gen_1_cmp_BSCmp_op2_10, A0=>nx3251, A1=>
      nx3257);
   ix3252 : nor02_2x port map ( Y=>nx3251, A0=>nx646, A1=>nx642);
   ix647 : nor03_2x port map ( Y=>nx646, A0=>gen_1_cmp_mReg_9, A1=>nx9683, 
      A2=>nx10193);
   ix643 : nor03_2x port map ( Y=>nx642, A0=>nx3246, A1=>nx10199, A2=>
      nx10209);
   ix3258 : nor02_2x port map ( Y=>nx3257, A0=>nx638, A1=>nx636);
   ix639 : nor03_2x port map ( Y=>nx638, A0=>nx3261, A1=>nx9677, A2=>nx10217
   );
   gen_1_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_1_cmp_mReg_10, QB=>
      nx3261, D=>window_1_10, CLK=>start, R=>rst);
   ix637 : nor03_2x port map ( Y=>nx636, A0=>gen_1_cmp_mReg_10, A1=>nx10007, 
      A2=>nx10225);
   ix673 : nand02 port map ( Y=>gen_1_cmp_BSCmp_op2_11, A0=>nx3267, A1=>
      nx3271);
   ix3268 : nor02_2x port map ( Y=>nx3267, A0=>nx668, A1=>nx664);
   ix669 : nor03_2x port map ( Y=>nx668, A0=>gen_1_cmp_mReg_10, A1=>nx9683, 
      A2=>nx10193);
   ix665 : nor03_2x port map ( Y=>nx664, A0=>nx3261, A1=>nx10199, A2=>
      nx10209);
   ix3272 : nor02_2x port map ( Y=>nx3271, A0=>nx660, A1=>nx658);
   ix661 : nor03_2x port map ( Y=>nx660, A0=>nx3275, A1=>nx9677, A2=>nx10217
   );
   gen_1_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_1_cmp_mReg_11, QB=>
      nx3275, D=>window_1_11, CLK=>start, R=>rst);
   ix659 : nor03_2x port map ( Y=>nx658, A0=>gen_1_cmp_mReg_11, A1=>nx10007, 
      A2=>nx10225);
   ix695 : nand02 port map ( Y=>gen_1_cmp_BSCmp_op2_12, A0=>nx3281, A1=>
      nx3287);
   ix3282 : nor02_2x port map ( Y=>nx3281, A0=>nx690, A1=>nx686);
   ix691 : nor03_2x port map ( Y=>nx690, A0=>gen_1_cmp_mReg_11, A1=>nx9683, 
      A2=>nx10193);
   ix687 : nor03_2x port map ( Y=>nx686, A0=>nx3275, A1=>nx10199, A2=>
      nx10209);
   ix3288 : nor02_2x port map ( Y=>nx3287, A0=>nx682, A1=>nx680);
   ix683 : nor03_2x port map ( Y=>nx682, A0=>nx3290, A1=>nx9679, A2=>nx10217
   );
   gen_1_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_1_cmp_mReg_12, QB=>
      nx3290, D=>window_1_12, CLK=>start, R=>rst);
   ix681 : nor03_2x port map ( Y=>nx680, A0=>gen_1_cmp_mReg_12, A1=>nx10007, 
      A2=>nx10225);
   ix717 : nand02 port map ( Y=>gen_1_cmp_BSCmp_op2_13, A0=>nx3295, A1=>
      nx3301);
   ix3296 : nor02_2x port map ( Y=>nx3295, A0=>nx712, A1=>nx708);
   ix713 : nor03_2x port map ( Y=>nx712, A0=>gen_1_cmp_mReg_12, A1=>nx9685, 
      A2=>nx10195);
   ix709 : nor03_2x port map ( Y=>nx708, A0=>nx3290, A1=>nx10199, A2=>
      nx10211);
   ix3302 : nor02_2x port map ( Y=>nx3301, A0=>nx704, A1=>nx702);
   ix705 : nor03_2x port map ( Y=>nx704, A0=>nx3305, A1=>nx9679, A2=>nx10219
   );
   gen_1_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_1_cmp_mReg_13, QB=>
      nx3305, D=>window_1_13, CLK=>start, R=>rst);
   ix703 : nor03_2x port map ( Y=>nx702, A0=>gen_1_cmp_mReg_13, A1=>nx10007, 
      A2=>nx10227);
   ix739 : nand02 port map ( Y=>gen_1_cmp_BSCmp_op2_14, A0=>nx3311, A1=>
      nx3315);
   ix3312 : nor02_2x port map ( Y=>nx3311, A0=>nx734, A1=>nx730);
   ix735 : nor03_2x port map ( Y=>nx734, A0=>gen_1_cmp_mReg_13, A1=>nx9685, 
      A2=>nx10195);
   ix731 : nor03_2x port map ( Y=>nx730, A0=>nx3305, A1=>nx10201, A2=>
      nx10211);
   ix3316 : nor02_2x port map ( Y=>nx3315, A0=>nx726, A1=>nx724);
   ix727 : nor03_2x port map ( Y=>nx726, A0=>nx3319, A1=>nx9679, A2=>nx10219
   );
   gen_1_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_1_cmp_mReg_14, QB=>
      nx3319, D=>window_1_14, CLK=>start, R=>rst);
   ix725 : nor03_2x port map ( Y=>nx724, A0=>gen_1_cmp_mReg_14, A1=>nx10007, 
      A2=>nx10227);
   ix761 : nand02 port map ( Y=>gen_1_cmp_BSCmp_op2_15, A0=>nx3325, A1=>
      nx3331);
   ix3326 : nor02_2x port map ( Y=>nx3325, A0=>nx756, A1=>nx752);
   ix757 : nor03_2x port map ( Y=>nx756, A0=>gen_1_cmp_mReg_14, A1=>nx9685, 
      A2=>nx10195);
   ix753 : nor03_2x port map ( Y=>nx752, A0=>nx3319, A1=>nx10201, A2=>
      nx10211);
   ix3332 : nor02_2x port map ( Y=>nx3331, A0=>nx748, A1=>nx746);
   ix749 : nor03_2x port map ( Y=>nx748, A0=>nx3334, A1=>nx9679, A2=>nx10219
   );
   gen_1_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_1_cmp_mReg_15, QB=>
      nx3334, D=>window_1_15, CLK=>start, R=>rst);
   ix747 : nor03_2x port map ( Y=>nx746, A0=>gen_1_cmp_mReg_15, A1=>nx10009, 
      A2=>nx10227);
   ix771 : nand02 port map ( Y=>gen_1_cmp_BSCmp_op2_16, A0=>nx3339, A1=>
      nx3331);
   ix3340 : nor02_2x port map ( Y=>nx3339, A0=>nx766, A1=>nx762);
   ix767 : nor03_2x port map ( Y=>nx766, A0=>gen_1_cmp_mReg_15, A1=>nx9685, 
      A2=>nx10195);
   ix763 : nor03_2x port map ( Y=>nx762, A0=>nx3334, A1=>nx10201, A2=>
      nx10211);
   ix839 : nand02 port map ( Y=>gen_2_cmp_BSCmp_op2_1, A0=>nx3347, A1=>
      nx3365);
   ix3348 : nor02_2x port map ( Y=>nx3347, A0=>nx834, A1=>nx830);
   ix835 : nor03_2x port map ( Y=>nx834, A0=>gen_2_cmp_mReg_0, A1=>nx9669, 
      A2=>nx10231);
   gen_2_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_2_cmp_mReg_0, QB=>
      nx3353, D=>window_2_0, CLK=>start, R=>rst);
   ix3357 : inv01 port map ( Y=>nx3356, A=>gen_2_cmp_pMux_0);
   ix831 : nor03_2x port map ( Y=>nx830, A0=>nx3353, A1=>nx10237, A2=>
      nx10247);
   ix3364 : inv02 port map ( Y=>nx3363, A=>gen_2_cmp_pMux_2);
   ix3366 : nor02_2x port map ( Y=>nx3365, A0=>nx820, A1=>nx818);
   ix821 : nor03_2x port map ( Y=>nx820, A0=>nx3369, A1=>nx9663, A2=>nx10255
   );
   gen_2_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_2_cmp_mReg_1, QB=>
      nx3369, D=>window_2_1, CLK=>start, R=>rst);
   ix819 : nor03_2x port map ( Y=>nx818, A0=>gen_2_cmp_mReg_1, A1=>nx10011, 
      A2=>nx10263);
   ix779 : nor03_2x port map ( Y=>nx778, A0=>nx9669, A1=>nx3363, A2=>
      gen_2_cmp_pMux_0);
   ix861 : nand02 port map ( Y=>gen_2_cmp_BSCmp_op2_2, A0=>nx3380, A1=>
      nx3387);
   ix3382 : nor02_2x port map ( Y=>nx3380, A0=>nx856, A1=>nx852);
   ix857 : nor03_2x port map ( Y=>nx856, A0=>gen_2_cmp_mReg_1, A1=>nx9669, 
      A2=>nx10231);
   ix853 : nor03_2x port map ( Y=>nx852, A0=>nx3369, A1=>nx10237, A2=>
      nx10247);
   ix3388 : nor02_2x port map ( Y=>nx3387, A0=>nx848, A1=>nx846);
   ix849 : nor03_2x port map ( Y=>nx848, A0=>nx3391, A1=>nx9663, A2=>nx10255
   );
   gen_2_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_2_cmp_mReg_2, QB=>
      nx3391, D=>window_2_2, CLK=>start, R=>rst);
   ix847 : nor03_2x port map ( Y=>nx846, A0=>gen_2_cmp_mReg_2, A1=>nx10011, 
      A2=>nx10263);
   ix883 : nand02 port map ( Y=>gen_2_cmp_BSCmp_op2_3, A0=>nx3397, A1=>
      nx3401);
   ix3398 : nor02_2x port map ( Y=>nx3397, A0=>nx878, A1=>nx874);
   ix879 : nor03_2x port map ( Y=>nx878, A0=>gen_2_cmp_mReg_2, A1=>nx9669, 
      A2=>nx10231);
   ix875 : nor03_2x port map ( Y=>nx874, A0=>nx3391, A1=>nx10237, A2=>
      nx10247);
   ix3402 : nor02_2x port map ( Y=>nx3401, A0=>nx870, A1=>nx868);
   ix871 : nor03_2x port map ( Y=>nx870, A0=>nx3405, A1=>nx9663, A2=>nx10255
   );
   gen_2_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_2_cmp_mReg_3, QB=>
      nx3405, D=>window_2_3, CLK=>start, R=>rst);
   ix869 : nor03_2x port map ( Y=>nx868, A0=>gen_2_cmp_mReg_3, A1=>nx10011, 
      A2=>nx10263);
   ix905 : nand02 port map ( Y=>gen_2_cmp_BSCmp_op2_4, A0=>nx3411, A1=>
      nx3415);
   ix3412 : nor02_2x port map ( Y=>nx3411, A0=>nx900, A1=>nx896);
   ix901 : nor03_2x port map ( Y=>nx900, A0=>gen_2_cmp_mReg_3, A1=>nx9669, 
      A2=>nx10231);
   ix897 : nor03_2x port map ( Y=>nx896, A0=>nx3405, A1=>nx10237, A2=>
      nx10247);
   ix3416 : nor02_2x port map ( Y=>nx3415, A0=>nx892, A1=>nx890);
   ix893 : nor03_2x port map ( Y=>nx892, A0=>nx3419, A1=>nx9663, A2=>nx10255
   );
   gen_2_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_2_cmp_mReg_4, QB=>
      nx3419, D=>window_2_4, CLK=>start, R=>rst);
   ix891 : nor03_2x port map ( Y=>nx890, A0=>gen_2_cmp_mReg_4, A1=>nx10011, 
      A2=>nx10263);
   ix927 : nand02 port map ( Y=>gen_2_cmp_BSCmp_op2_5, A0=>nx3423, A1=>
      nx3429);
   ix3424 : nor02_2x port map ( Y=>nx3423, A0=>nx922, A1=>nx918);
   ix923 : nor03_2x port map ( Y=>nx922, A0=>gen_2_cmp_mReg_4, A1=>nx9669, 
      A2=>nx10231);
   ix919 : nor03_2x port map ( Y=>nx918, A0=>nx3419, A1=>nx10237, A2=>
      nx10247);
   ix3430 : nor02_2x port map ( Y=>nx3429, A0=>nx914, A1=>nx912);
   ix915 : nor03_2x port map ( Y=>nx914, A0=>nx3433, A1=>nx9665, A2=>nx10255
   );
   gen_2_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_2_cmp_mReg_5, QB=>
      nx3433, D=>window_2_5, CLK=>start, R=>rst);
   ix913 : nor03_2x port map ( Y=>nx912, A0=>gen_2_cmp_mReg_5, A1=>nx10011, 
      A2=>nx10263);
   ix949 : nand02 port map ( Y=>gen_2_cmp_BSCmp_op2_6, A0=>nx3437, A1=>
      nx3443);
   ix3438 : nor02_2x port map ( Y=>nx3437, A0=>nx944, A1=>nx940);
   ix945 : nor03_2x port map ( Y=>nx944, A0=>gen_2_cmp_mReg_5, A1=>nx9671, 
      A2=>nx10231);
   ix941 : nor03_2x port map ( Y=>nx940, A0=>nx3433, A1=>nx10237, A2=>
      nx10247);
   ix3444 : nor02_2x port map ( Y=>nx3443, A0=>nx936, A1=>nx934);
   ix937 : nor03_2x port map ( Y=>nx936, A0=>nx3446, A1=>nx9665, A2=>nx10255
   );
   gen_2_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_2_cmp_mReg_6, QB=>
      nx3446, D=>window_2_6, CLK=>start, R=>rst);
   ix935 : nor03_2x port map ( Y=>nx934, A0=>gen_2_cmp_mReg_6, A1=>nx10011, 
      A2=>nx10263);
   ix971 : nand02 port map ( Y=>gen_2_cmp_BSCmp_op2_7, A0=>nx3453, A1=>
      nx3459);
   ix3454 : nor02_2x port map ( Y=>nx3453, A0=>nx966, A1=>nx962);
   ix967 : nor03_2x port map ( Y=>nx966, A0=>gen_2_cmp_mReg_6, A1=>nx9671, 
      A2=>nx10233);
   ix963 : nor03_2x port map ( Y=>nx962, A0=>nx3446, A1=>nx10239, A2=>
      nx10249);
   ix3460 : nor02_2x port map ( Y=>nx3459, A0=>nx958, A1=>nx956);
   ix959 : nor03_2x port map ( Y=>nx958, A0=>nx3463, A1=>nx9665, A2=>nx10257
   );
   gen_2_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_2_cmp_mReg_7, QB=>
      nx3463, D=>window_2_7, CLK=>start, R=>rst);
   ix957 : nor03_2x port map ( Y=>nx956, A0=>gen_2_cmp_mReg_7, A1=>nx10011, 
      A2=>nx10265);
   ix993 : nand02 port map ( Y=>gen_2_cmp_BSCmp_op2_8, A0=>nx3469, A1=>
      nx3475);
   ix3470 : nor02_2x port map ( Y=>nx3469, A0=>nx988, A1=>nx984);
   ix989 : nor03_2x port map ( Y=>nx988, A0=>gen_2_cmp_mReg_7, A1=>nx9671, 
      A2=>nx10233);
   ix985 : nor03_2x port map ( Y=>nx984, A0=>nx3463, A1=>nx10239, A2=>
      nx10249);
   ix3476 : nor02_2x port map ( Y=>nx3475, A0=>nx980, A1=>nx978);
   ix981 : nor03_2x port map ( Y=>nx980, A0=>nx3479, A1=>nx9665, A2=>nx10257
   );
   gen_2_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_2_cmp_mReg_8, QB=>
      nx3479, D=>window_2_8, CLK=>start, R=>rst);
   ix979 : nor03_2x port map ( Y=>nx978, A0=>gen_2_cmp_mReg_8, A1=>nx10013, 
      A2=>nx10265);
   ix1015 : nand02 port map ( Y=>gen_2_cmp_BSCmp_op2_9, A0=>nx3484, A1=>
      nx3488);
   ix3485 : nor02_2x port map ( Y=>nx3484, A0=>nx1010, A1=>nx1006);
   ix1011 : nor03_2x port map ( Y=>nx1010, A0=>gen_2_cmp_mReg_8, A1=>nx9671, 
      A2=>nx10233);
   ix1007 : nor03_2x port map ( Y=>nx1006, A0=>nx3479, A1=>nx10239, A2=>
      nx10249);
   ix3489 : nor02_2x port map ( Y=>nx3488, A0=>nx1002, A1=>nx1000);
   ix1003 : nor03_2x port map ( Y=>nx1002, A0=>nx3491, A1=>nx9665, A2=>
      nx10257);
   gen_2_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_2_cmp_mReg_9, QB=>
      nx3491, D=>window_2_9, CLK=>start, R=>rst);
   ix1001 : nor03_2x port map ( Y=>nx1000, A0=>gen_2_cmp_mReg_9, A1=>nx10013, 
      A2=>nx10265);
   ix1037 : nand02 port map ( Y=>gen_2_cmp_BSCmp_op2_10, A0=>nx3497, A1=>
      nx3503);
   ix3498 : nor02_2x port map ( Y=>nx3497, A0=>nx1032, A1=>nx1028);
   ix1033 : nor03_2x port map ( Y=>nx1032, A0=>gen_2_cmp_mReg_9, A1=>nx9671, 
      A2=>nx10233);
   ix1029 : nor03_2x port map ( Y=>nx1028, A0=>nx3491, A1=>nx10239, A2=>
      nx10249);
   ix3504 : nor02_2x port map ( Y=>nx3503, A0=>nx1024, A1=>nx1022);
   ix1025 : nor03_2x port map ( Y=>nx1024, A0=>nx3507, A1=>nx9665, A2=>
      nx10257);
   gen_2_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_2_cmp_mReg_10, QB=>
      nx3507, D=>window_2_10, CLK=>start, R=>rst);
   ix1023 : nor03_2x port map ( Y=>nx1022, A0=>gen_2_cmp_mReg_10, A1=>
      nx10013, A2=>nx10265);
   ix1059 : nand02 port map ( Y=>gen_2_cmp_BSCmp_op2_11, A0=>nx3513, A1=>
      nx3517);
   ix3514 : nor02_2x port map ( Y=>nx3513, A0=>nx1054, A1=>nx1050);
   ix1055 : nor03_2x port map ( Y=>nx1054, A0=>gen_2_cmp_mReg_10, A1=>nx9671, 
      A2=>nx10233);
   ix1051 : nor03_2x port map ( Y=>nx1050, A0=>nx3507, A1=>nx10239, A2=>
      nx10249);
   ix3518 : nor02_2x port map ( Y=>nx3517, A0=>nx1046, A1=>nx1044);
   ix1047 : nor03_2x port map ( Y=>nx1046, A0=>nx3521, A1=>nx9665, A2=>
      nx10257);
   gen_2_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_2_cmp_mReg_11, QB=>
      nx3521, D=>window_2_11, CLK=>start, R=>rst);
   ix1045 : nor03_2x port map ( Y=>nx1044, A0=>gen_2_cmp_mReg_11, A1=>
      nx10013, A2=>nx10265);
   ix1081 : nand02 port map ( Y=>gen_2_cmp_BSCmp_op2_12, A0=>nx3527, A1=>
      nx3533);
   ix3528 : nor02_2x port map ( Y=>nx3527, A0=>nx1076, A1=>nx1072);
   ix1077 : nor03_2x port map ( Y=>nx1076, A0=>gen_2_cmp_mReg_11, A1=>nx9671, 
      A2=>nx10233);
   ix1073 : nor03_2x port map ( Y=>nx1072, A0=>nx3521, A1=>nx10239, A2=>
      nx10249);
   ix3534 : nor02_2x port map ( Y=>nx3533, A0=>nx1068, A1=>nx1066);
   ix1069 : nor03_2x port map ( Y=>nx1068, A0=>nx3537, A1=>nx9667, A2=>
      nx10257);
   gen_2_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_2_cmp_mReg_12, QB=>
      nx3537, D=>window_2_12, CLK=>start, R=>rst);
   ix1067 : nor03_2x port map ( Y=>nx1066, A0=>gen_2_cmp_mReg_12, A1=>
      nx10013, A2=>nx10265);
   ix1103 : nand02 port map ( Y=>gen_2_cmp_BSCmp_op2_13, A0=>nx3543, A1=>
      nx3547);
   ix3544 : nor02_2x port map ( Y=>nx3543, A0=>nx1098, A1=>nx1094);
   ix1099 : nor03_2x port map ( Y=>nx1098, A0=>gen_2_cmp_mReg_12, A1=>nx9673, 
      A2=>nx10235);
   ix1095 : nor03_2x port map ( Y=>nx1094, A0=>nx3537, A1=>nx10239, A2=>
      nx10251);
   ix3548 : nor02_2x port map ( Y=>nx3547, A0=>nx1090, A1=>nx1088);
   ix1091 : nor03_2x port map ( Y=>nx1090, A0=>nx3551, A1=>nx9667, A2=>
      nx10259);
   gen_2_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_2_cmp_mReg_13, QB=>
      nx3551, D=>window_2_13, CLK=>start, R=>rst);
   ix1089 : nor03_2x port map ( Y=>nx1088, A0=>gen_2_cmp_mReg_13, A1=>
      nx10013, A2=>nx10267);
   ix1125 : nand02 port map ( Y=>gen_2_cmp_BSCmp_op2_14, A0=>nx3557, A1=>
      nx3563);
   ix3558 : nor02_2x port map ( Y=>nx3557, A0=>nx1120, A1=>nx1116);
   ix1121 : nor03_2x port map ( Y=>nx1120, A0=>gen_2_cmp_mReg_13, A1=>nx9673, 
      A2=>nx10235);
   ix1117 : nor03_2x port map ( Y=>nx1116, A0=>nx3551, A1=>nx10241, A2=>
      nx10251);
   ix3564 : nor02_2x port map ( Y=>nx3563, A0=>nx1112, A1=>nx1110);
   ix1113 : nor03_2x port map ( Y=>nx1112, A0=>nx3566, A1=>nx9667, A2=>
      nx10259);
   gen_2_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_2_cmp_mReg_14, QB=>
      nx3566, D=>window_2_14, CLK=>start, R=>rst);
   ix1111 : nor03_2x port map ( Y=>nx1110, A0=>gen_2_cmp_mReg_14, A1=>
      nx10013, A2=>nx10267);
   ix1147 : nand02 port map ( Y=>gen_2_cmp_BSCmp_op2_15, A0=>nx3571, A1=>
      nx3577);
   ix3572 : nor02_2x port map ( Y=>nx3571, A0=>nx1142, A1=>nx1138);
   ix1143 : nor03_2x port map ( Y=>nx1142, A0=>gen_2_cmp_mReg_14, A1=>nx9673, 
      A2=>nx10235);
   ix1139 : nor03_2x port map ( Y=>nx1138, A0=>nx3566, A1=>nx10241, A2=>
      nx10251);
   ix3578 : nor02_2x port map ( Y=>nx3577, A0=>nx1134, A1=>nx1132);
   ix1135 : nor03_2x port map ( Y=>nx1134, A0=>nx3581, A1=>nx9667, A2=>
      nx10259);
   gen_2_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_2_cmp_mReg_15, QB=>
      nx3581, D=>window_2_15, CLK=>start, R=>rst);
   ix1133 : nor03_2x port map ( Y=>nx1132, A0=>gen_2_cmp_mReg_15, A1=>
      nx10015, A2=>nx10267);
   ix1157 : nand02 port map ( Y=>gen_2_cmp_BSCmp_op2_16, A0=>nx3587, A1=>
      nx3577);
   ix3588 : nor02_2x port map ( Y=>nx3587, A0=>nx1152, A1=>nx1148);
   ix1153 : nor03_2x port map ( Y=>nx1152, A0=>gen_2_cmp_mReg_15, A1=>nx9673, 
      A2=>nx10235);
   ix1149 : nor03_2x port map ( Y=>nx1148, A0=>nx3581, A1=>nx10241, A2=>
      nx10251);
   ix1225 : nand02 port map ( Y=>gen_3_cmp_BSCmp_op2_1, A0=>nx3593, A1=>
      nx3613);
   ix3594 : nor02_2x port map ( Y=>nx3593, A0=>nx1220, A1=>nx1216);
   ix1221 : nor03_2x port map ( Y=>nx1220, A0=>gen_3_cmp_mReg_0, A1=>nx9657, 
      A2=>nx10271);
   gen_3_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_3_cmp_mReg_0, QB=>
      nx3599, D=>window_3_0, CLK=>start, R=>rst);
   ix3604 : inv01 port map ( Y=>nx3603, A=>gen_3_cmp_pMux_0);
   ix1217 : nor03_2x port map ( Y=>nx1216, A0=>nx3599, A1=>nx10277, A2=>
      nx10287);
   ix3612 : inv02 port map ( Y=>nx3611, A=>gen_3_cmp_pMux_2);
   ix3614 : nor02_2x port map ( Y=>nx3613, A0=>nx1206, A1=>nx1204);
   ix1207 : nor03_2x port map ( Y=>nx1206, A0=>nx3617, A1=>nx9651, A2=>
      nx10295);
   gen_3_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_3_cmp_mReg_1, QB=>
      nx3617, D=>window_3_1, CLK=>start, R=>rst);
   ix1205 : nor03_2x port map ( Y=>nx1204, A0=>gen_3_cmp_mReg_1, A1=>nx10017, 
      A2=>nx10303);
   ix1165 : nor03_2x port map ( Y=>nx1164, A0=>nx9657, A1=>nx3611, A2=>
      gen_3_cmp_pMux_0);
   ix1247 : nand02 port map ( Y=>gen_3_cmp_BSCmp_op2_2, A0=>nx3629, A1=>
      nx3633);
   ix3630 : nor02_2x port map ( Y=>nx3629, A0=>nx1242, A1=>nx1238);
   ix1243 : nor03_2x port map ( Y=>nx1242, A0=>gen_3_cmp_mReg_1, A1=>nx9657, 
      A2=>nx10271);
   ix1239 : nor03_2x port map ( Y=>nx1238, A0=>nx3617, A1=>nx10277, A2=>
      nx10287);
   ix3634 : nor02_2x port map ( Y=>nx3633, A0=>nx1234, A1=>nx1232);
   ix1235 : nor03_2x port map ( Y=>nx1234, A0=>nx3637, A1=>nx9651, A2=>
      nx10295);
   gen_3_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_3_cmp_mReg_2, QB=>
      nx3637, D=>window_3_2, CLK=>start, R=>rst);
   ix1233 : nor03_2x port map ( Y=>nx1232, A0=>gen_3_cmp_mReg_2, A1=>nx10017, 
      A2=>nx10303);
   ix1269 : nand02 port map ( Y=>gen_3_cmp_BSCmp_op2_3, A0=>nx3643, A1=>
      nx3647);
   ix3644 : nor02_2x port map ( Y=>nx3643, A0=>nx1264, A1=>nx1260);
   ix1265 : nor03_2x port map ( Y=>nx1264, A0=>gen_3_cmp_mReg_2, A1=>nx9657, 
      A2=>nx10271);
   ix1261 : nor03_2x port map ( Y=>nx1260, A0=>nx3637, A1=>nx10277, A2=>
      nx10287);
   ix3648 : nor02_2x port map ( Y=>nx3647, A0=>nx1256, A1=>nx1254);
   ix1257 : nor03_2x port map ( Y=>nx1256, A0=>nx3651, A1=>nx9651, A2=>
      nx10295);
   gen_3_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_3_cmp_mReg_3, QB=>
      nx3651, D=>window_3_3, CLK=>start, R=>rst);
   ix1255 : nor03_2x port map ( Y=>nx1254, A0=>gen_3_cmp_mReg_3, A1=>nx10017, 
      A2=>nx10303);
   ix1291 : nand02 port map ( Y=>gen_3_cmp_BSCmp_op2_4, A0=>nx3655, A1=>
      nx3661);
   ix3656 : nor02_2x port map ( Y=>nx3655, A0=>nx1286, A1=>nx1282);
   ix1287 : nor03_2x port map ( Y=>nx1286, A0=>gen_3_cmp_mReg_3, A1=>nx9657, 
      A2=>nx10271);
   ix1283 : nor03_2x port map ( Y=>nx1282, A0=>nx3651, A1=>nx10277, A2=>
      nx10287);
   ix3662 : nor02_2x port map ( Y=>nx3661, A0=>nx1278, A1=>nx1276);
   ix1279 : nor03_2x port map ( Y=>nx1278, A0=>nx3665, A1=>nx9651, A2=>
      nx10295);
   gen_3_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_3_cmp_mReg_4, QB=>
      nx3665, D=>window_3_4, CLK=>start, R=>rst);
   ix1277 : nor03_2x port map ( Y=>nx1276, A0=>gen_3_cmp_mReg_4, A1=>nx10017, 
      A2=>nx10303);
   ix1313 : nand02 port map ( Y=>gen_3_cmp_BSCmp_op2_5, A0=>nx3669, A1=>
      nx3675);
   ix3670 : nor02_2x port map ( Y=>nx3669, A0=>nx1308, A1=>nx1304);
   ix1309 : nor03_2x port map ( Y=>nx1308, A0=>gen_3_cmp_mReg_4, A1=>nx9657, 
      A2=>nx10271);
   ix1305 : nor03_2x port map ( Y=>nx1304, A0=>nx3665, A1=>nx10277, A2=>
      nx10287);
   ix3676 : nor02_2x port map ( Y=>nx3675, A0=>nx1300, A1=>nx1298);
   ix1301 : nor03_2x port map ( Y=>nx1300, A0=>nx3678, A1=>nx9653, A2=>
      nx10295);
   gen_3_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_3_cmp_mReg_5, QB=>
      nx3678, D=>window_3_5, CLK=>start, R=>rst);
   ix1299 : nor03_2x port map ( Y=>nx1298, A0=>gen_3_cmp_mReg_5, A1=>nx10017, 
      A2=>nx10303);
   ix1335 : nand02 port map ( Y=>gen_3_cmp_BSCmp_op2_6, A0=>nx3685, A1=>
      nx3691);
   ix3686 : nor02_2x port map ( Y=>nx3685, A0=>nx1330, A1=>nx1326);
   ix1331 : nor03_2x port map ( Y=>nx1330, A0=>gen_3_cmp_mReg_5, A1=>nx9659, 
      A2=>nx10271);
   ix1327 : nor03_2x port map ( Y=>nx1326, A0=>nx3678, A1=>nx10277, A2=>
      nx10287);
   ix3692 : nor02_2x port map ( Y=>nx3691, A0=>nx1322, A1=>nx1320);
   ix1323 : nor03_2x port map ( Y=>nx1322, A0=>nx3695, A1=>nx9653, A2=>
      nx10295);
   gen_3_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_3_cmp_mReg_6, QB=>
      nx3695, D=>window_3_6, CLK=>start, R=>rst);
   ix1321 : nor03_2x port map ( Y=>nx1320, A0=>gen_3_cmp_mReg_6, A1=>nx10017, 
      A2=>nx10303);
   ix1357 : nand02 port map ( Y=>gen_3_cmp_BSCmp_op2_7, A0=>nx3699, A1=>
      nx3705);
   ix3700 : nor02_2x port map ( Y=>nx3699, A0=>nx1352, A1=>nx1348);
   ix1353 : nor03_2x port map ( Y=>nx1352, A0=>gen_3_cmp_mReg_6, A1=>nx9659, 
      A2=>nx10273);
   ix1349 : nor03_2x port map ( Y=>nx1348, A0=>nx3695, A1=>nx10279, A2=>
      nx10289);
   ix3706 : nor02_2x port map ( Y=>nx3705, A0=>nx1344, A1=>nx1342);
   ix1345 : nor03_2x port map ( Y=>nx1344, A0=>nx3709, A1=>nx9653, A2=>
      nx10297);
   gen_3_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_3_cmp_mReg_7, QB=>
      nx3709, D=>window_3_7, CLK=>start, R=>rst);
   ix1343 : nor03_2x port map ( Y=>nx1342, A0=>gen_3_cmp_mReg_7, A1=>nx10017, 
      A2=>nx10305);
   ix1379 : nand02 port map ( Y=>gen_3_cmp_BSCmp_op2_8, A0=>nx3713, A1=>
      nx3719);
   ix3714 : nor02_2x port map ( Y=>nx3713, A0=>nx1374, A1=>nx1370);
   ix1375 : nor03_2x port map ( Y=>nx1374, A0=>gen_3_cmp_mReg_7, A1=>nx9659, 
      A2=>nx10273);
   ix1371 : nor03_2x port map ( Y=>nx1370, A0=>nx3709, A1=>nx10279, A2=>
      nx10289);
   ix3720 : nor02_2x port map ( Y=>nx3719, A0=>nx1366, A1=>nx1364);
   ix1367 : nor03_2x port map ( Y=>nx1366, A0=>nx3722, A1=>nx9653, A2=>
      nx10297);
   gen_3_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_3_cmp_mReg_8, QB=>
      nx3722, D=>window_3_8, CLK=>start, R=>rst);
   ix1365 : nor03_2x port map ( Y=>nx1364, A0=>gen_3_cmp_mReg_8, A1=>nx10019, 
      A2=>nx10305);
   ix1401 : nand02 port map ( Y=>gen_3_cmp_BSCmp_op2_9, A0=>nx3729, A1=>
      nx3735);
   ix3730 : nor02_2x port map ( Y=>nx3729, A0=>nx1396, A1=>nx1392);
   ix1397 : nor03_2x port map ( Y=>nx1396, A0=>gen_3_cmp_mReg_8, A1=>nx9659, 
      A2=>nx10273);
   ix1393 : nor03_2x port map ( Y=>nx1392, A0=>nx3722, A1=>nx10279, A2=>
      nx10289);
   ix3736 : nor02_2x port map ( Y=>nx3735, A0=>nx1388, A1=>nx1386);
   ix1389 : nor03_2x port map ( Y=>nx1388, A0=>nx3739, A1=>nx9653, A2=>
      nx10297);
   gen_3_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_3_cmp_mReg_9, QB=>
      nx3739, D=>window_3_9, CLK=>start, R=>rst);
   ix1387 : nor03_2x port map ( Y=>nx1386, A0=>gen_3_cmp_mReg_9, A1=>nx10019, 
      A2=>nx10305);
   ix1423 : nand02 port map ( Y=>gen_3_cmp_BSCmp_op2_10, A0=>nx3743, A1=>
      nx3749);
   ix3744 : nor02_2x port map ( Y=>nx3743, A0=>nx1418, A1=>nx1414);
   ix1419 : nor03_2x port map ( Y=>nx1418, A0=>gen_3_cmp_mReg_9, A1=>nx9659, 
      A2=>nx10273);
   ix1415 : nor03_2x port map ( Y=>nx1414, A0=>nx3739, A1=>nx10279, A2=>
      nx10289);
   ix3750 : nor02_2x port map ( Y=>nx3749, A0=>nx1410, A1=>nx1408);
   ix1411 : nor03_2x port map ( Y=>nx1410, A0=>nx3753, A1=>nx9653, A2=>
      nx10297);
   gen_3_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_3_cmp_mReg_10, QB=>
      nx3753, D=>window_3_10, CLK=>start, R=>rst);
   ix1409 : nor03_2x port map ( Y=>nx1408, A0=>gen_3_cmp_mReg_10, A1=>
      nx10019, A2=>nx10305);
   ix1445 : nand02 port map ( Y=>gen_3_cmp_BSCmp_op2_11, A0=>nx3757, A1=>
      nx3763);
   ix3758 : nor02_2x port map ( Y=>nx3757, A0=>nx1440, A1=>nx1436);
   ix1441 : nor03_2x port map ( Y=>nx1440, A0=>gen_3_cmp_mReg_10, A1=>nx9659, 
      A2=>nx10273);
   ix1437 : nor03_2x port map ( Y=>nx1436, A0=>nx3753, A1=>nx10279, A2=>
      nx10289);
   ix3764 : nor02_2x port map ( Y=>nx3763, A0=>nx1432, A1=>nx1430);
   ix1433 : nor03_2x port map ( Y=>nx1432, A0=>nx3766, A1=>nx9653, A2=>
      nx10297);
   gen_3_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_3_cmp_mReg_11, QB=>
      nx3766, D=>window_3_11, CLK=>start, R=>rst);
   ix1431 : nor03_2x port map ( Y=>nx1430, A0=>gen_3_cmp_mReg_11, A1=>
      nx10019, A2=>nx10305);
   ix1467 : nand02 port map ( Y=>gen_3_cmp_BSCmp_op2_12, A0=>nx3773, A1=>
      nx3779);
   ix3774 : nor02_2x port map ( Y=>nx3773, A0=>nx1462, A1=>nx1458);
   ix1463 : nor03_2x port map ( Y=>nx1462, A0=>gen_3_cmp_mReg_11, A1=>nx9659, 
      A2=>nx10273);
   ix1459 : nor03_2x port map ( Y=>nx1458, A0=>nx3766, A1=>nx10279, A2=>
      nx10289);
   ix3780 : nor02_2x port map ( Y=>nx3779, A0=>nx1454, A1=>nx1452);
   ix1455 : nor03_2x port map ( Y=>nx1454, A0=>nx3783, A1=>nx9655, A2=>
      nx10297);
   gen_3_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_3_cmp_mReg_12, QB=>
      nx3783, D=>window_3_12, CLK=>start, R=>rst);
   ix1453 : nor03_2x port map ( Y=>nx1452, A0=>gen_3_cmp_mReg_12, A1=>
      nx10019, A2=>nx10305);
   ix1489 : nand02 port map ( Y=>gen_3_cmp_BSCmp_op2_13, A0=>nx3787, A1=>
      nx3793);
   ix3788 : nor02_2x port map ( Y=>nx3787, A0=>nx1484, A1=>nx1480);
   ix1485 : nor03_2x port map ( Y=>nx1484, A0=>gen_3_cmp_mReg_12, A1=>nx9661, 
      A2=>nx10275);
   ix1481 : nor03_2x port map ( Y=>nx1480, A0=>nx3783, A1=>nx10279, A2=>
      nx10291);
   ix3794 : nor02_2x port map ( Y=>nx3793, A0=>nx1476, A1=>nx1474);
   ix1477 : nor03_2x port map ( Y=>nx1476, A0=>nx3797, A1=>nx9655, A2=>
      nx10299);
   gen_3_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_3_cmp_mReg_13, QB=>
      nx3797, D=>window_3_13, CLK=>start, R=>rst);
   ix1475 : nor03_2x port map ( Y=>nx1474, A0=>gen_3_cmp_mReg_13, A1=>
      nx10019, A2=>nx10307);
   ix1511 : nand02 port map ( Y=>gen_3_cmp_BSCmp_op2_14, A0=>nx3801, A1=>
      nx3807);
   ix3802 : nor02_2x port map ( Y=>nx3801, A0=>nx1506, A1=>nx1502);
   ix1507 : nor03_2x port map ( Y=>nx1506, A0=>gen_3_cmp_mReg_13, A1=>nx9661, 
      A2=>nx10275);
   ix1503 : nor03_2x port map ( Y=>nx1502, A0=>nx3797, A1=>nx10281, A2=>
      nx10291);
   ix3808 : nor02_2x port map ( Y=>nx3807, A0=>nx1498, A1=>nx1496);
   ix1499 : nor03_2x port map ( Y=>nx1498, A0=>nx3810, A1=>nx9655, A2=>
      nx10299);
   gen_3_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_3_cmp_mReg_14, QB=>
      nx3810, D=>window_3_14, CLK=>start, R=>rst);
   ix1497 : nor03_2x port map ( Y=>nx1496, A0=>gen_3_cmp_mReg_14, A1=>
      nx10019, A2=>nx10307);
   ix1533 : nand02 port map ( Y=>gen_3_cmp_BSCmp_op2_15, A0=>nx3817, A1=>
      nx3823);
   ix3818 : nor02_2x port map ( Y=>nx3817, A0=>nx1528, A1=>nx1524);
   ix1529 : nor03_2x port map ( Y=>nx1528, A0=>gen_3_cmp_mReg_14, A1=>nx9661, 
      A2=>nx10275);
   ix1525 : nor03_2x port map ( Y=>nx1524, A0=>nx3810, A1=>nx10281, A2=>
      nx10291);
   ix3824 : nor02_2x port map ( Y=>nx3823, A0=>nx1520, A1=>nx1518);
   ix1521 : nor03_2x port map ( Y=>nx1520, A0=>nx3827, A1=>nx9655, A2=>
      nx10299);
   gen_3_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_3_cmp_mReg_15, QB=>
      nx3827, D=>window_3_15, CLK=>start, R=>rst);
   ix1519 : nor03_2x port map ( Y=>nx1518, A0=>gen_3_cmp_mReg_15, A1=>
      nx10021, A2=>nx10307);
   ix1543 : nand02 port map ( Y=>gen_3_cmp_BSCmp_op2_16, A0=>nx3831, A1=>
      nx3823);
   ix3832 : nor02_2x port map ( Y=>nx3831, A0=>nx1538, A1=>nx1534);
   ix1539 : nor03_2x port map ( Y=>nx1538, A0=>gen_3_cmp_mReg_15, A1=>nx9661, 
      A2=>nx10275);
   ix1535 : nor03_2x port map ( Y=>nx1534, A0=>nx3827, A1=>nx10281, A2=>
      nx10291);
   ix1611 : nand02 port map ( Y=>gen_4_cmp_BSCmp_op2_1, A0=>nx3839, A1=>
      nx3859);
   ix3840 : nor02_2x port map ( Y=>nx3839, A0=>nx1606, A1=>nx1602);
   ix1607 : nor03_2x port map ( Y=>nx1606, A0=>gen_4_cmp_mReg_0, A1=>nx9645, 
      A2=>nx10311);
   gen_4_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_4_cmp_mReg_0, QB=>
      nx3845, D=>window_4_0, CLK=>start, R=>rst);
   ix3850 : inv01 port map ( Y=>nx3849, A=>gen_4_cmp_pMux_0);
   ix1603 : nor03_2x port map ( Y=>nx1602, A0=>nx3845, A1=>nx10317, A2=>
      nx10327);
   ix3858 : inv02 port map ( Y=>nx3857, A=>gen_4_cmp_pMux_2);
   ix3860 : nor02_2x port map ( Y=>nx3859, A0=>nx1592, A1=>nx1590);
   ix1593 : nor03_2x port map ( Y=>nx1592, A0=>nx3863, A1=>nx9639, A2=>
      nx10335);
   gen_4_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_4_cmp_mReg_1, QB=>
      nx3863, D=>window_4_1, CLK=>start, R=>rst);
   ix1591 : nor03_2x port map ( Y=>nx1590, A0=>gen_4_cmp_mReg_1, A1=>nx10023, 
      A2=>nx10343);
   ix1551 : nor03_2x port map ( Y=>nx1550, A0=>nx9645, A1=>nx3857, A2=>
      gen_4_cmp_pMux_0);
   ix1633 : nand02 port map ( Y=>gen_4_cmp_BSCmp_op2_2, A0=>nx3873, A1=>
      nx3877);
   ix3874 : nor02_2x port map ( Y=>nx3873, A0=>nx1628, A1=>nx1624);
   ix1629 : nor03_2x port map ( Y=>nx1628, A0=>gen_4_cmp_mReg_1, A1=>nx9645, 
      A2=>nx10311);
   ix1625 : nor03_2x port map ( Y=>nx1624, A0=>nx3863, A1=>nx10317, A2=>
      nx10327);
   ix3878 : nor02_2x port map ( Y=>nx3877, A0=>nx1620, A1=>nx1618);
   ix1621 : nor03_2x port map ( Y=>nx1620, A0=>nx3881, A1=>nx9639, A2=>
      nx10335);
   gen_4_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_4_cmp_mReg_2, QB=>
      nx3881, D=>window_4_2, CLK=>start, R=>rst);
   ix1619 : nor03_2x port map ( Y=>nx1618, A0=>gen_4_cmp_mReg_2, A1=>nx10023, 
      A2=>nx10343);
   ix1655 : nand02 port map ( Y=>gen_4_cmp_BSCmp_op2_3, A0=>nx3887, A1=>
      nx3893);
   ix3888 : nor02_2x port map ( Y=>nx3887, A0=>nx1650, A1=>nx1646);
   ix1651 : nor03_2x port map ( Y=>nx1650, A0=>gen_4_cmp_mReg_2, A1=>nx9645, 
      A2=>nx10311);
   ix1647 : nor03_2x port map ( Y=>nx1646, A0=>nx3881, A1=>nx10317, A2=>
      nx10327);
   ix3894 : nor02_2x port map ( Y=>nx3893, A0=>nx1642, A1=>nx1640);
   ix1643 : nor03_2x port map ( Y=>nx1642, A0=>nx3897, A1=>nx9639, A2=>
      nx10335);
   gen_4_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_4_cmp_mReg_3, QB=>
      nx3897, D=>window_4_3, CLK=>start, R=>rst);
   ix1641 : nor03_2x port map ( Y=>nx1640, A0=>gen_4_cmp_mReg_3, A1=>nx10023, 
      A2=>nx10343);
   ix1677 : nand02 port map ( Y=>gen_4_cmp_BSCmp_op2_4, A0=>nx3902, A1=>
      nx3907);
   ix3903 : nor02_2x port map ( Y=>nx3902, A0=>nx1672, A1=>nx1668);
   ix1673 : nor03_2x port map ( Y=>nx1672, A0=>gen_4_cmp_mReg_3, A1=>nx9645, 
      A2=>nx10311);
   ix1669 : nor03_2x port map ( Y=>nx1668, A0=>nx3897, A1=>nx10317, A2=>
      nx10327);
   ix3908 : nor02_2x port map ( Y=>nx3907, A0=>nx1664, A1=>nx1662);
   ix1665 : nor03_2x port map ( Y=>nx1664, A0=>nx3911, A1=>nx9639, A2=>
      nx10335);
   gen_4_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_4_cmp_mReg_4, QB=>
      nx3911, D=>window_4_4, CLK=>start, R=>rst);
   ix1663 : nor03_2x port map ( Y=>nx1662, A0=>gen_4_cmp_mReg_4, A1=>nx10023, 
      A2=>nx10343);
   ix1699 : nand02 port map ( Y=>gen_4_cmp_BSCmp_op2_5, A0=>nx3915, A1=>
      nx3921);
   ix3916 : nor02_2x port map ( Y=>nx3915, A0=>nx1694, A1=>nx1690);
   ix1695 : nor03_2x port map ( Y=>nx1694, A0=>gen_4_cmp_mReg_4, A1=>nx9645, 
      A2=>nx10311);
   ix1691 : nor03_2x port map ( Y=>nx1690, A0=>nx3911, A1=>nx10317, A2=>
      nx10327);
   ix3922 : nor02_2x port map ( Y=>nx3921, A0=>nx1686, A1=>nx1684);
   ix1687 : nor03_2x port map ( Y=>nx1686, A0=>nx3925, A1=>nx9641, A2=>
      nx10335);
   gen_4_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_4_cmp_mReg_5, QB=>
      nx3925, D=>window_4_5, CLK=>start, R=>rst);
   ix1685 : nor03_2x port map ( Y=>nx1684, A0=>gen_4_cmp_mReg_5, A1=>nx10023, 
      A2=>nx10343);
   ix1721 : nand02 port map ( Y=>gen_4_cmp_BSCmp_op2_6, A0=>nx3930, A1=>
      nx3935);
   ix3931 : nor02_2x port map ( Y=>nx3930, A0=>nx1716, A1=>nx1712);
   ix1717 : nor03_2x port map ( Y=>nx1716, A0=>gen_4_cmp_mReg_5, A1=>nx9647, 
      A2=>nx10311);
   ix1713 : nor03_2x port map ( Y=>nx1712, A0=>nx3925, A1=>nx10317, A2=>
      nx10327);
   ix3936 : nor02_2x port map ( Y=>nx3935, A0=>nx1708, A1=>nx1706);
   ix1709 : nor03_2x port map ( Y=>nx1708, A0=>nx3939, A1=>nx9641, A2=>
      nx10335);
   gen_4_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_4_cmp_mReg_6, QB=>
      nx3939, D=>window_4_6, CLK=>start, R=>rst);
   ix1707 : nor03_2x port map ( Y=>nx1706, A0=>gen_4_cmp_mReg_6, A1=>nx10023, 
      A2=>nx10343);
   ix1743 : nand02 port map ( Y=>gen_4_cmp_BSCmp_op2_7, A0=>nx3945, A1=>
      nx3951);
   ix3946 : nor02_2x port map ( Y=>nx3945, A0=>nx1738, A1=>nx1734);
   ix1739 : nor03_2x port map ( Y=>nx1738, A0=>gen_4_cmp_mReg_6, A1=>nx9647, 
      A2=>nx10313);
   ix1735 : nor03_2x port map ( Y=>nx1734, A0=>nx3939, A1=>nx10319, A2=>
      nx10329);
   ix3952 : nor02_2x port map ( Y=>nx3951, A0=>nx1730, A1=>nx1728);
   ix1731 : nor03_2x port map ( Y=>nx1730, A0=>nx3954, A1=>nx9641, A2=>
      nx10337);
   gen_4_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_4_cmp_mReg_7, QB=>
      nx3954, D=>window_4_7, CLK=>start, R=>rst);
   ix1729 : nor03_2x port map ( Y=>nx1728, A0=>gen_4_cmp_mReg_7, A1=>nx10023, 
      A2=>nx10345);
   ix1765 : nand02 port map ( Y=>gen_4_cmp_BSCmp_op2_8, A0=>nx3961, A1=>
      nx3967);
   ix3962 : nor02_2x port map ( Y=>nx3961, A0=>nx1760, A1=>nx1756);
   ix1761 : nor03_2x port map ( Y=>nx1760, A0=>gen_4_cmp_mReg_7, A1=>nx9647, 
      A2=>nx10313);
   ix1757 : nor03_2x port map ( Y=>nx1756, A0=>nx3954, A1=>nx10319, A2=>
      nx10329);
   ix3968 : nor02_2x port map ( Y=>nx3967, A0=>nx1752, A1=>nx1750);
   ix1753 : nor03_2x port map ( Y=>nx1752, A0=>nx3971, A1=>nx9641, A2=>
      nx10337);
   gen_4_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_4_cmp_mReg_8, QB=>
      nx3971, D=>window_4_8, CLK=>start, R=>rst);
   ix1751 : nor03_2x port map ( Y=>nx1750, A0=>gen_4_cmp_mReg_8, A1=>nx10025, 
      A2=>nx10345);
   ix1787 : nand02 port map ( Y=>gen_4_cmp_BSCmp_op2_9, A0=>nx3975, A1=>
      nx3981);
   ix3976 : nor02_2x port map ( Y=>nx3975, A0=>nx1782, A1=>nx1778);
   ix1783 : nor03_2x port map ( Y=>nx1782, A0=>gen_4_cmp_mReg_8, A1=>nx9647, 
      A2=>nx10313);
   ix1779 : nor03_2x port map ( Y=>nx1778, A0=>nx3971, A1=>nx10319, A2=>
      nx10329);
   ix3982 : nor02_2x port map ( Y=>nx3981, A0=>nx1774, A1=>nx1772);
   ix1775 : nor03_2x port map ( Y=>nx1774, A0=>nx3985, A1=>nx9641, A2=>
      nx10337);
   gen_4_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_4_cmp_mReg_9, QB=>
      nx3985, D=>window_4_9, CLK=>start, R=>rst);
   ix1773 : nor03_2x port map ( Y=>nx1772, A0=>gen_4_cmp_mReg_9, A1=>nx10025, 
      A2=>nx10345);
   ix1809 : nand02 port map ( Y=>gen_4_cmp_BSCmp_op2_10, A0=>nx3989, A1=>
      nx3995);
   ix3990 : nor02_2x port map ( Y=>nx3989, A0=>nx1804, A1=>nx1800);
   ix1805 : nor03_2x port map ( Y=>nx1804, A0=>gen_4_cmp_mReg_9, A1=>nx9647, 
      A2=>nx10313);
   ix1801 : nor03_2x port map ( Y=>nx1800, A0=>nx3985, A1=>nx10319, A2=>
      nx10329);
   ix3996 : nor02_2x port map ( Y=>nx3995, A0=>nx1796, A1=>nx1794);
   ix1797 : nor03_2x port map ( Y=>nx1796, A0=>nx3998, A1=>nx9641, A2=>
      nx10337);
   gen_4_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_4_cmp_mReg_10, QB=>
      nx3998, D=>window_4_10, CLK=>start, R=>rst);
   ix1795 : nor03_2x port map ( Y=>nx1794, A0=>gen_4_cmp_mReg_10, A1=>
      nx10025, A2=>nx10345);
   ix1831 : nand02 port map ( Y=>gen_4_cmp_BSCmp_op2_11, A0=>nx4005, A1=>
      nx4011);
   ix4006 : nor02_2x port map ( Y=>nx4005, A0=>nx1826, A1=>nx1822);
   ix1827 : nor03_2x port map ( Y=>nx1826, A0=>gen_4_cmp_mReg_10, A1=>nx9647, 
      A2=>nx10313);
   ix1823 : nor03_2x port map ( Y=>nx1822, A0=>nx3998, A1=>nx10319, A2=>
      nx10329);
   ix4012 : nor02_2x port map ( Y=>nx4011, A0=>nx1818, A1=>nx1816);
   ix1819 : nor03_2x port map ( Y=>nx1818, A0=>nx4015, A1=>nx9641, A2=>
      nx10337);
   gen_4_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_4_cmp_mReg_11, QB=>
      nx4015, D=>window_4_11, CLK=>start, R=>rst);
   ix1817 : nor03_2x port map ( Y=>nx1816, A0=>gen_4_cmp_mReg_11, A1=>
      nx10025, A2=>nx10345);
   ix1853 : nand02 port map ( Y=>gen_4_cmp_BSCmp_op2_12, A0=>nx4019, A1=>
      nx4025);
   ix4020 : nor02_2x port map ( Y=>nx4019, A0=>nx1848, A1=>nx1844);
   ix1849 : nor03_2x port map ( Y=>nx1848, A0=>gen_4_cmp_mReg_11, A1=>nx9647, 
      A2=>nx10313);
   ix1845 : nor03_2x port map ( Y=>nx1844, A0=>nx4015, A1=>nx10319, A2=>
      nx10329);
   ix4026 : nor02_2x port map ( Y=>nx4025, A0=>nx1840, A1=>nx1838);
   ix1841 : nor03_2x port map ( Y=>nx1840, A0=>nx4029, A1=>nx9643, A2=>
      nx10337);
   gen_4_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_4_cmp_mReg_12, QB=>
      nx4029, D=>window_4_12, CLK=>start, R=>rst);
   ix1839 : nor03_2x port map ( Y=>nx1838, A0=>gen_4_cmp_mReg_12, A1=>
      nx10025, A2=>nx10345);
   ix1875 : nand02 port map ( Y=>gen_4_cmp_BSCmp_op2_13, A0=>nx4033, A1=>
      nx4039);
   ix4034 : nor02_2x port map ( Y=>nx4033, A0=>nx1870, A1=>nx1866);
   ix1871 : nor03_2x port map ( Y=>nx1870, A0=>gen_4_cmp_mReg_12, A1=>nx9649, 
      A2=>nx10315);
   ix1867 : nor03_2x port map ( Y=>nx1866, A0=>nx4029, A1=>nx10319, A2=>
      nx10331);
   ix4040 : nor02_2x port map ( Y=>nx4039, A0=>nx1862, A1=>nx1860);
   ix1863 : nor03_2x port map ( Y=>nx1862, A0=>nx4042, A1=>nx9643, A2=>
      nx10339);
   gen_4_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_4_cmp_mReg_13, QB=>
      nx4042, D=>window_4_13, CLK=>start, R=>rst);
   ix1861 : nor03_2x port map ( Y=>nx1860, A0=>gen_4_cmp_mReg_13, A1=>
      nx10025, A2=>nx10347);
   ix1897 : nand02 port map ( Y=>gen_4_cmp_BSCmp_op2_14, A0=>nx4049, A1=>
      nx4055);
   ix4050 : nor02_2x port map ( Y=>nx4049, A0=>nx1892, A1=>nx1888);
   ix1893 : nor03_2x port map ( Y=>nx1892, A0=>gen_4_cmp_mReg_13, A1=>nx9649, 
      A2=>nx10315);
   ix1889 : nor03_2x port map ( Y=>nx1888, A0=>nx4042, A1=>nx10321, A2=>
      nx10331);
   ix4056 : nor02_2x port map ( Y=>nx4055, A0=>nx1884, A1=>nx1882);
   ix1885 : nor03_2x port map ( Y=>nx1884, A0=>nx4059, A1=>nx9643, A2=>
      nx10339);
   gen_4_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_4_cmp_mReg_14, QB=>
      nx4059, D=>window_4_14, CLK=>start, R=>rst);
   ix1883 : nor03_2x port map ( Y=>nx1882, A0=>gen_4_cmp_mReg_14, A1=>
      nx10025, A2=>nx10347);
   ix1919 : nand02 port map ( Y=>gen_4_cmp_BSCmp_op2_15, A0=>nx4063, A1=>
      nx4069);
   ix4064 : nor02_2x port map ( Y=>nx4063, A0=>nx1914, A1=>nx1910);
   ix1915 : nor03_2x port map ( Y=>nx1914, A0=>gen_4_cmp_mReg_14, A1=>nx9649, 
      A2=>nx10315);
   ix1911 : nor03_2x port map ( Y=>nx1910, A0=>nx4059, A1=>nx10321, A2=>
      nx10331);
   ix4070 : nor02_2x port map ( Y=>nx4069, A0=>nx1906, A1=>nx1904);
   ix1907 : nor03_2x port map ( Y=>nx1906, A0=>nx4073, A1=>nx9643, A2=>
      nx10339);
   gen_4_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_4_cmp_mReg_15, QB=>
      nx4073, D=>window_4_15, CLK=>start, R=>rst);
   ix1905 : nor03_2x port map ( Y=>nx1904, A0=>gen_4_cmp_mReg_15, A1=>
      nx10027, A2=>nx10347);
   ix1929 : nand02 port map ( Y=>gen_4_cmp_BSCmp_op2_16, A0=>nx4077, A1=>
      nx4069);
   ix4078 : nor02_2x port map ( Y=>nx4077, A0=>nx1924, A1=>nx1920);
   ix1925 : nor03_2x port map ( Y=>nx1924, A0=>gen_4_cmp_mReg_15, A1=>nx9649, 
      A2=>nx10315);
   ix1921 : nor03_2x port map ( Y=>nx1920, A0=>nx4073, A1=>nx10321, A2=>
      nx10331);
   ix1997 : nand02 port map ( Y=>gen_5_cmp_BSCmp_op2_1, A0=>nx4084, A1=>
      nx4103);
   ix4085 : nor02_2x port map ( Y=>nx4084, A0=>nx1992, A1=>nx1988);
   ix1993 : nor03_2x port map ( Y=>nx1992, A0=>gen_5_cmp_mReg_0, A1=>nx9633, 
      A2=>nx10351);
   gen_5_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_5_cmp_mReg_0, QB=>
      nx4089, D=>window_5_0, CLK=>start, R=>rst);
   ix4094 : inv01 port map ( Y=>nx4093, A=>gen_5_cmp_pMux_0);
   ix1989 : nor03_2x port map ( Y=>nx1988, A0=>nx4089, A1=>nx10357, A2=>
      nx10367);
   ix4102 : inv02 port map ( Y=>nx4101, A=>gen_5_cmp_pMux_2);
   ix4104 : nor02_2x port map ( Y=>nx4103, A0=>nx1978, A1=>nx1976);
   ix1979 : nor03_2x port map ( Y=>nx1978, A0=>nx4106, A1=>nx9627, A2=>
      nx10375);
   gen_5_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_5_cmp_mReg_1, QB=>
      nx4106, D=>window_5_1, CLK=>start, R=>rst);
   ix1977 : nor03_2x port map ( Y=>nx1976, A0=>gen_5_cmp_mReg_1, A1=>nx10029, 
      A2=>nx10383);
   ix1937 : nor03_2x port map ( Y=>nx1936, A0=>nx9633, A1=>nx4101, A2=>
      gen_5_cmp_pMux_0);
   ix2019 : nand02 port map ( Y=>gen_5_cmp_BSCmp_op2_2, A0=>nx4119, A1=>
      nx4125);
   ix4120 : nor02_2x port map ( Y=>nx4119, A0=>nx2014, A1=>nx2010);
   ix2015 : nor03_2x port map ( Y=>nx2014, A0=>gen_5_cmp_mReg_1, A1=>nx9633, 
      A2=>nx10351);
   ix2011 : nor03_2x port map ( Y=>nx2010, A0=>nx4106, A1=>nx10357, A2=>
      nx10367);
   ix4126 : nor02_2x port map ( Y=>nx4125, A0=>nx2006, A1=>nx2004);
   ix2007 : nor03_2x port map ( Y=>nx2006, A0=>nx4128, A1=>nx9627, A2=>
      nx10375);
   gen_5_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_5_cmp_mReg_2, QB=>
      nx4128, D=>window_5_2, CLK=>start, R=>rst);
   ix2005 : nor03_2x port map ( Y=>nx2004, A0=>gen_5_cmp_mReg_2, A1=>nx10029, 
      A2=>nx10383);
   ix2041 : nand02 port map ( Y=>gen_5_cmp_BSCmp_op2_3, A0=>nx4133, A1=>
      nx4139);
   ix4134 : nor02_2x port map ( Y=>nx4133, A0=>nx2036, A1=>nx2032);
   ix2037 : nor03_2x port map ( Y=>nx2036, A0=>gen_5_cmp_mReg_2, A1=>nx9633, 
      A2=>nx10351);
   ix2033 : nor03_2x port map ( Y=>nx2032, A0=>nx4128, A1=>nx10357, A2=>
      nx10367);
   ix4140 : nor02_2x port map ( Y=>nx4139, A0=>nx2028, A1=>nx2026);
   ix2029 : nor03_2x port map ( Y=>nx2028, A0=>nx4143, A1=>nx9627, A2=>
      nx10375);
   gen_5_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_5_cmp_mReg_3, QB=>
      nx4143, D=>window_5_3, CLK=>start, R=>rst);
   ix2027 : nor03_2x port map ( Y=>nx2026, A0=>gen_5_cmp_mReg_3, A1=>nx10029, 
      A2=>nx10383);
   ix2063 : nand02 port map ( Y=>gen_5_cmp_BSCmp_op2_4, A0=>nx4149, A1=>
      nx4153);
   ix4150 : nor02_2x port map ( Y=>nx4149, A0=>nx2058, A1=>nx2054);
   ix2059 : nor03_2x port map ( Y=>nx2058, A0=>gen_5_cmp_mReg_3, A1=>nx9633, 
      A2=>nx10351);
   ix2055 : nor03_2x port map ( Y=>nx2054, A0=>nx4143, A1=>nx10357, A2=>
      nx10367);
   ix4154 : nor02_2x port map ( Y=>nx4153, A0=>nx2050, A1=>nx2048);
   ix2051 : nor03_2x port map ( Y=>nx2050, A0=>nx4157, A1=>nx9627, A2=>
      nx10375);
   gen_5_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_5_cmp_mReg_4, QB=>
      nx4157, D=>window_5_4, CLK=>start, R=>rst);
   ix2049 : nor03_2x port map ( Y=>nx2048, A0=>gen_5_cmp_mReg_4, A1=>nx10029, 
      A2=>nx10383);
   ix2085 : nand02 port map ( Y=>gen_5_cmp_BSCmp_op2_5, A0=>nx4163, A1=>
      nx4169);
   ix4164 : nor02_2x port map ( Y=>nx4163, A0=>nx2080, A1=>nx2076);
   ix2081 : nor03_2x port map ( Y=>nx2080, A0=>gen_5_cmp_mReg_4, A1=>nx9633, 
      A2=>nx10351);
   ix2077 : nor03_2x port map ( Y=>nx2076, A0=>nx4157, A1=>nx10357, A2=>
      nx10367);
   ix4170 : nor02_2x port map ( Y=>nx4169, A0=>nx2072, A1=>nx2070);
   ix2073 : nor03_2x port map ( Y=>nx2072, A0=>nx4172, A1=>nx9629, A2=>
      nx10375);
   gen_5_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_5_cmp_mReg_5, QB=>
      nx4172, D=>window_5_5, CLK=>start, R=>rst);
   ix2071 : nor03_2x port map ( Y=>nx2070, A0=>gen_5_cmp_mReg_5, A1=>nx10029, 
      A2=>nx10383);
   ix2107 : nand02 port map ( Y=>gen_5_cmp_BSCmp_op2_6, A0=>nx4177, A1=>
      nx4183);
   ix4178 : nor02_2x port map ( Y=>nx4177, A0=>nx2102, A1=>nx2098);
   ix2103 : nor03_2x port map ( Y=>nx2102, A0=>gen_5_cmp_mReg_5, A1=>nx9635, 
      A2=>nx10351);
   ix2099 : nor03_2x port map ( Y=>nx2098, A0=>nx4172, A1=>nx10357, A2=>
      nx10367);
   ix4184 : nor02_2x port map ( Y=>nx4183, A0=>nx2094, A1=>nx2092);
   ix2095 : nor03_2x port map ( Y=>nx2094, A0=>nx4187, A1=>nx9629, A2=>
      nx10375);
   gen_5_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_5_cmp_mReg_6, QB=>
      nx4187, D=>window_5_6, CLK=>start, R=>rst);
   ix2093 : nor03_2x port map ( Y=>nx2092, A0=>gen_5_cmp_mReg_6, A1=>nx10029, 
      A2=>nx10383);
   ix2129 : nand02 port map ( Y=>gen_5_cmp_BSCmp_op2_7, A0=>nx4193, A1=>
      nx4197);
   ix4194 : nor02_2x port map ( Y=>nx4193, A0=>nx2124, A1=>nx2120);
   ix2125 : nor03_2x port map ( Y=>nx2124, A0=>gen_5_cmp_mReg_6, A1=>nx9635, 
      A2=>nx10353);
   ix2121 : nor03_2x port map ( Y=>nx2120, A0=>nx4187, A1=>nx10359, A2=>
      nx10369);
   ix4198 : nor02_2x port map ( Y=>nx4197, A0=>nx2116, A1=>nx2114);
   ix2117 : nor03_2x port map ( Y=>nx2116, A0=>nx4201, A1=>nx9629, A2=>
      nx10377);
   gen_5_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_5_cmp_mReg_7, QB=>
      nx4201, D=>window_5_7, CLK=>start, R=>rst);
   ix2115 : nor03_2x port map ( Y=>nx2114, A0=>gen_5_cmp_mReg_7, A1=>nx10029, 
      A2=>nx10385);
   ix2151 : nand02 port map ( Y=>gen_5_cmp_BSCmp_op2_8, A0=>nx4207, A1=>
      nx4213);
   ix4208 : nor02_2x port map ( Y=>nx4207, A0=>nx2146, A1=>nx2142);
   ix2147 : nor03_2x port map ( Y=>nx2146, A0=>gen_5_cmp_mReg_7, A1=>nx9635, 
      A2=>nx10353);
   ix2143 : nor03_2x port map ( Y=>nx2142, A0=>nx4201, A1=>nx10359, A2=>
      nx10369);
   ix4214 : nor02_2x port map ( Y=>nx4213, A0=>nx2138, A1=>nx2136);
   ix2139 : nor03_2x port map ( Y=>nx2138, A0=>nx4216, A1=>nx9629, A2=>
      nx10377);
   gen_5_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_5_cmp_mReg_8, QB=>
      nx4216, D=>window_5_8, CLK=>start, R=>rst);
   ix2137 : nor03_2x port map ( Y=>nx2136, A0=>gen_5_cmp_mReg_8, A1=>nx10031, 
      A2=>nx10385);
   ix2173 : nand02 port map ( Y=>gen_5_cmp_BSCmp_op2_9, A0=>nx4221, A1=>
      nx4227);
   ix4222 : nor02_2x port map ( Y=>nx4221, A0=>nx2168, A1=>nx2164);
   ix2169 : nor03_2x port map ( Y=>nx2168, A0=>gen_5_cmp_mReg_8, A1=>nx9635, 
      A2=>nx10353);
   ix2165 : nor03_2x port map ( Y=>nx2164, A0=>nx4216, A1=>nx10359, A2=>
      nx10369);
   ix4228 : nor02_2x port map ( Y=>nx4227, A0=>nx2160, A1=>nx2158);
   ix2161 : nor03_2x port map ( Y=>nx2160, A0=>nx4231, A1=>nx9629, A2=>
      nx10377);
   gen_5_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_5_cmp_mReg_9, QB=>
      nx4231, D=>window_5_9, CLK=>start, R=>rst);
   ix2159 : nor03_2x port map ( Y=>nx2158, A0=>gen_5_cmp_mReg_9, A1=>nx10031, 
      A2=>nx10385);
   ix2195 : nand02 port map ( Y=>gen_5_cmp_BSCmp_op2_10, A0=>nx4237, A1=>
      nx4241);
   ix4238 : nor02_2x port map ( Y=>nx4237, A0=>nx2190, A1=>nx2186);
   ix2191 : nor03_2x port map ( Y=>nx2190, A0=>gen_5_cmp_mReg_9, A1=>nx9635, 
      A2=>nx10353);
   ix2187 : nor03_2x port map ( Y=>nx2186, A0=>nx4231, A1=>nx10359, A2=>
      nx10369);
   ix4242 : nor02_2x port map ( Y=>nx4241, A0=>nx2182, A1=>nx2180);
   ix2183 : nor03_2x port map ( Y=>nx2182, A0=>nx4245, A1=>nx9629, A2=>
      nx10377);
   gen_5_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_5_cmp_mReg_10, QB=>
      nx4245, D=>window_5_10, CLK=>start, R=>rst);
   ix2181 : nor03_2x port map ( Y=>nx2180, A0=>gen_5_cmp_mReg_10, A1=>
      nx10031, A2=>nx10385);
   ix2217 : nand02 port map ( Y=>gen_5_cmp_BSCmp_op2_11, A0=>nx4251, A1=>
      nx4256);
   ix4252 : nor02_2x port map ( Y=>nx4251, A0=>nx2212, A1=>nx2208);
   ix2213 : nor03_2x port map ( Y=>nx2212, A0=>gen_5_cmp_mReg_10, A1=>nx9635, 
      A2=>nx10353);
   ix2209 : nor03_2x port map ( Y=>nx2208, A0=>nx4245, A1=>nx10359, A2=>
      nx10369);
   ix4257 : nor02_2x port map ( Y=>nx4256, A0=>nx2204, A1=>nx2202);
   ix2205 : nor03_2x port map ( Y=>nx2204, A0=>nx4259, A1=>nx9629, A2=>
      nx10377);
   gen_5_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_5_cmp_mReg_11, QB=>
      nx4259, D=>window_5_11, CLK=>start, R=>rst);
   ix2203 : nor03_2x port map ( Y=>nx2202, A0=>gen_5_cmp_mReg_11, A1=>
      nx10031, A2=>nx10385);
   ix2239 : nand02 port map ( Y=>gen_5_cmp_BSCmp_op2_12, A0=>nx4263, A1=>
      nx4269);
   ix4264 : nor02_2x port map ( Y=>nx4263, A0=>nx2234, A1=>nx2230);
   ix2235 : nor03_2x port map ( Y=>nx2234, A0=>gen_5_cmp_mReg_11, A1=>nx9635, 
      A2=>nx10353);
   ix2231 : nor03_2x port map ( Y=>nx2230, A0=>nx4259, A1=>nx10359, A2=>
      nx10369);
   ix4270 : nor02_2x port map ( Y=>nx4269, A0=>nx2226, A1=>nx2224);
   ix2227 : nor03_2x port map ( Y=>nx2226, A0=>nx4273, A1=>nx9631, A2=>
      nx10377);
   gen_5_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_5_cmp_mReg_12, QB=>
      nx4273, D=>window_5_12, CLK=>start, R=>rst);
   ix2225 : nor03_2x port map ( Y=>nx2224, A0=>gen_5_cmp_mReg_12, A1=>
      nx10031, A2=>nx10385);
   ix2261 : nand02 port map ( Y=>gen_5_cmp_BSCmp_op2_13, A0=>nx4279, A1=>
      nx4285);
   ix4280 : nor02_2x port map ( Y=>nx4279, A0=>nx2256, A1=>nx2252);
   ix2257 : nor03_2x port map ( Y=>nx2256, A0=>gen_5_cmp_mReg_12, A1=>nx9637, 
      A2=>nx10355);
   ix2253 : nor03_2x port map ( Y=>nx2252, A0=>nx4273, A1=>nx10359, A2=>
      nx10371);
   ix4286 : nor02_2x port map ( Y=>nx4285, A0=>nx2248, A1=>nx2246);
   ix2249 : nor03_2x port map ( Y=>nx2248, A0=>nx4288, A1=>nx9631, A2=>
      nx10379);
   gen_5_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_5_cmp_mReg_13, QB=>
      nx4288, D=>window_5_13, CLK=>start, R=>rst);
   ix2247 : nor03_2x port map ( Y=>nx2246, A0=>gen_5_cmp_mReg_13, A1=>
      nx10031, A2=>nx10387);
   ix2283 : nand02 port map ( Y=>gen_5_cmp_BSCmp_op2_14, A0=>nx4293, A1=>
      nx4299);
   ix4294 : nor02_2x port map ( Y=>nx4293, A0=>nx2278, A1=>nx2274);
   ix2279 : nor03_2x port map ( Y=>nx2278, A0=>gen_5_cmp_mReg_13, A1=>nx9637, 
      A2=>nx10355);
   ix2275 : nor03_2x port map ( Y=>nx2274, A0=>nx4288, A1=>nx10361, A2=>
      nx10371);
   ix4300 : nor02_2x port map ( Y=>nx4299, A0=>nx2270, A1=>nx2268);
   ix2271 : nor03_2x port map ( Y=>nx2270, A0=>nx4303, A1=>nx9631, A2=>
      nx10379);
   gen_5_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_5_cmp_mReg_14, QB=>
      nx4303, D=>window_5_14, CLK=>start, R=>rst);
   ix2269 : nor03_2x port map ( Y=>nx2268, A0=>gen_5_cmp_mReg_14, A1=>
      nx10031, A2=>nx10387);
   ix2305 : nand02 port map ( Y=>gen_5_cmp_BSCmp_op2_15, A0=>nx4309, A1=>
      nx4315);
   ix4310 : nor02_2x port map ( Y=>nx4309, A0=>nx2300, A1=>nx2296);
   ix2301 : nor03_2x port map ( Y=>nx2300, A0=>gen_5_cmp_mReg_14, A1=>nx9637, 
      A2=>nx10355);
   ix2297 : nor03_2x port map ( Y=>nx2296, A0=>nx4303, A1=>nx10361, A2=>
      nx10371);
   ix4316 : nor02_2x port map ( Y=>nx4315, A0=>nx2292, A1=>nx2290);
   ix2293 : nor03_2x port map ( Y=>nx2292, A0=>nx4318, A1=>nx9631, A2=>
      nx10379);
   gen_5_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_5_cmp_mReg_15, QB=>
      nx4318, D=>window_5_15, CLK=>start, R=>rst);
   ix2291 : nor03_2x port map ( Y=>nx2290, A0=>gen_5_cmp_mReg_15, A1=>
      nx10033, A2=>nx10387);
   ix2315 : nand02 port map ( Y=>gen_5_cmp_BSCmp_op2_16, A0=>nx4325, A1=>
      nx4315);
   ix4326 : nor02_2x port map ( Y=>nx4325, A0=>nx2310, A1=>nx2306);
   ix2311 : nor03_2x port map ( Y=>nx2310, A0=>gen_5_cmp_mReg_15, A1=>nx9637, 
      A2=>nx10355);
   ix2307 : nor03_2x port map ( Y=>nx2306, A0=>nx4318, A1=>nx10361, A2=>
      nx10371);
   ix2383 : nand02 port map ( Y=>gen_6_cmp_BSCmp_op2_1, A0=>nx4331, A1=>
      nx4351);
   ix4332 : nor02_2x port map ( Y=>nx4331, A0=>nx2378, A1=>nx2374);
   ix2379 : nor03_2x port map ( Y=>nx2378, A0=>gen_6_cmp_mReg_0, A1=>nx9621, 
      A2=>nx10391);
   gen_6_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_6_cmp_mReg_0, QB=>
      nx4337, D=>window_6_0, CLK=>start, R=>rst);
   ix4342 : inv01 port map ( Y=>nx4340, A=>gen_6_cmp_pMux_0);
   ix2375 : nor03_2x port map ( Y=>nx2374, A0=>nx4337, A1=>nx10397, A2=>
      nx10407);
   ix4350 : inv02 port map ( Y=>nx4349, A=>gen_6_cmp_pMux_2);
   ix4352 : nor02_2x port map ( Y=>nx4351, A0=>nx2364, A1=>nx2362);
   ix2365 : nor03_2x port map ( Y=>nx2364, A0=>nx4355, A1=>nx9615, A2=>
      nx10415);
   gen_6_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_6_cmp_mReg_1, QB=>
      nx4355, D=>window_6_1, CLK=>start, R=>rst);
   ix2363 : nor03_2x port map ( Y=>nx2362, A0=>gen_6_cmp_mReg_1, A1=>nx10035, 
      A2=>nx10423);
   ix2326 : nor03_2x port map ( Y=>nx2322, A0=>nx9621, A1=>nx4349, A2=>
      gen_6_cmp_pMux_0);
   ix2405 : nand02 port map ( Y=>gen_6_cmp_BSCmp_op2_2, A0=>nx4365, A1=>
      nx4371);
   ix4366 : nor02_2x port map ( Y=>nx4365, A0=>nx2400, A1=>nx2396);
   ix2401 : nor03_2x port map ( Y=>nx2400, A0=>gen_6_cmp_mReg_1, A1=>nx9621, 
      A2=>nx10391);
   ix2397 : nor03_2x port map ( Y=>nx2396, A0=>nx4355, A1=>nx10397, A2=>
      nx10407);
   ix4372 : nor02_2x port map ( Y=>nx4371, A0=>nx2392, A1=>nx2390);
   ix2393 : nor03_2x port map ( Y=>nx2392, A0=>nx4375, A1=>nx9615, A2=>
      nx10415);
   gen_6_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_6_cmp_mReg_2, QB=>
      nx4375, D=>window_6_2, CLK=>start, R=>rst);
   ix2391 : nor03_2x port map ( Y=>nx2390, A0=>gen_6_cmp_mReg_2, A1=>nx10035, 
      A2=>nx10423);
   ix2427 : nand02 port map ( Y=>gen_6_cmp_BSCmp_op2_3, A0=>nx4381, A1=>
      nx4385);
   ix4382 : nor02_2x port map ( Y=>nx4381, A0=>nx2422, A1=>nx2418);
   ix2423 : nor03_2x port map ( Y=>nx2422, A0=>gen_6_cmp_mReg_2, A1=>nx9621, 
      A2=>nx10391);
   ix2419 : nor03_2x port map ( Y=>nx2418, A0=>nx4375, A1=>nx10397, A2=>
      nx10407);
   ix4386 : nor02_2x port map ( Y=>nx4385, A0=>nx2414, A1=>nx2412);
   ix2415 : nor03_2x port map ( Y=>nx2414, A0=>nx4389, A1=>nx9615, A2=>
      nx10415);
   gen_6_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_6_cmp_mReg_3, QB=>
      nx4389, D=>window_6_3, CLK=>start, R=>rst);
   ix2413 : nor03_2x port map ( Y=>nx2412, A0=>gen_6_cmp_mReg_3, A1=>nx10035, 
      A2=>nx10423);
   ix2449 : nand02 port map ( Y=>gen_6_cmp_BSCmp_op2_4, A0=>nx4395, A1=>
      nx4401);
   ix4396 : nor02_2x port map ( Y=>nx4395, A0=>nx2444, A1=>nx2440);
   ix2445 : nor03_2x port map ( Y=>nx2444, A0=>gen_6_cmp_mReg_3, A1=>nx9621, 
      A2=>nx10391);
   ix2441 : nor03_2x port map ( Y=>nx2440, A0=>nx4389, A1=>nx10397, A2=>
      nx10407);
   ix4402 : nor02_2x port map ( Y=>nx4401, A0=>nx2436, A1=>nx2434);
   ix2437 : nor03_2x port map ( Y=>nx2436, A0=>nx4404, A1=>nx9615, A2=>
      nx10415);
   gen_6_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_6_cmp_mReg_4, QB=>
      nx4404, D=>window_6_4, CLK=>start, R=>rst);
   ix2435 : nor03_2x port map ( Y=>nx2434, A0=>gen_6_cmp_mReg_4, A1=>nx10035, 
      A2=>nx10423);
   ix2471 : nand02 port map ( Y=>gen_6_cmp_BSCmp_op2_5, A0=>nx4409, A1=>
      nx4415);
   ix4410 : nor02_2x port map ( Y=>nx4409, A0=>nx2466, A1=>nx2462);
   ix2467 : nor03_2x port map ( Y=>nx2466, A0=>gen_6_cmp_mReg_4, A1=>nx9621, 
      A2=>nx10391);
   ix2463 : nor03_2x port map ( Y=>nx2462, A0=>nx4404, A1=>nx10397, A2=>
      nx10407);
   ix4416 : nor02_2x port map ( Y=>nx4415, A0=>nx2458, A1=>nx2456);
   ix2459 : nor03_2x port map ( Y=>nx2458, A0=>nx4419, A1=>nx9617, A2=>
      nx10415);
   gen_6_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_6_cmp_mReg_5, QB=>
      nx4419, D=>window_6_5, CLK=>start, R=>rst);
   ix2457 : nor03_2x port map ( Y=>nx2456, A0=>gen_6_cmp_mReg_5, A1=>nx10035, 
      A2=>nx10423);
   ix2493 : nand02 port map ( Y=>gen_6_cmp_BSCmp_op2_6, A0=>nx4425, A1=>
      nx4429);
   ix4426 : nor02_2x port map ( Y=>nx4425, A0=>nx2488, A1=>nx2484);
   ix2489 : nor03_2x port map ( Y=>nx2488, A0=>gen_6_cmp_mReg_5, A1=>nx9623, 
      A2=>nx10391);
   ix2485 : nor03_2x port map ( Y=>nx2484, A0=>nx4419, A1=>nx10397, A2=>
      nx10407);
   ix4430 : nor02_2x port map ( Y=>nx4429, A0=>nx2480, A1=>nx2478);
   ix2481 : nor03_2x port map ( Y=>nx2480, A0=>nx4433, A1=>nx9617, A2=>
      nx10415);
   gen_6_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_6_cmp_mReg_6, QB=>
      nx4433, D=>window_6_6, CLK=>start, R=>rst);
   ix2479 : nor03_2x port map ( Y=>nx2478, A0=>gen_6_cmp_mReg_6, A1=>nx10035, 
      A2=>nx10423);
   ix2515 : nand02 port map ( Y=>gen_6_cmp_BSCmp_op2_7, A0=>nx4439, A1=>
      nx4445);
   ix4440 : nor02_2x port map ( Y=>nx4439, A0=>nx2510, A1=>nx2506);
   ix2511 : nor03_2x port map ( Y=>nx2510, A0=>gen_6_cmp_mReg_6, A1=>nx9623, 
      A2=>nx10393);
   ix2507 : nor03_2x port map ( Y=>nx2506, A0=>nx4433, A1=>nx10399, A2=>
      nx10409);
   ix4446 : nor02_2x port map ( Y=>nx4445, A0=>nx2502, A1=>nx2500);
   ix2503 : nor03_2x port map ( Y=>nx2502, A0=>nx4448, A1=>nx9617, A2=>
      nx10417);
   gen_6_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_6_cmp_mReg_7, QB=>
      nx4448, D=>window_6_7, CLK=>start, R=>rst);
   ix2501 : nor03_2x port map ( Y=>nx2500, A0=>gen_6_cmp_mReg_7, A1=>nx10035, 
      A2=>nx10425);
   ix2537 : nand02 port map ( Y=>gen_6_cmp_BSCmp_op2_8, A0=>nx4453, A1=>
      nx4459);
   ix4454 : nor02_2x port map ( Y=>nx4453, A0=>nx2532, A1=>nx2528);
   ix2533 : nor03_2x port map ( Y=>nx2532, A0=>gen_6_cmp_mReg_7, A1=>nx9623, 
      A2=>nx10393);
   ix2529 : nor03_2x port map ( Y=>nx2528, A0=>nx4448, A1=>nx10399, A2=>
      nx10409);
   ix4460 : nor02_2x port map ( Y=>nx4459, A0=>nx2524, A1=>nx2522);
   ix2525 : nor03_2x port map ( Y=>nx2524, A0=>nx4463, A1=>nx9617, A2=>
      nx10417);
   gen_6_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_6_cmp_mReg_8, QB=>
      nx4463, D=>window_6_8, CLK=>start, R=>rst);
   ix2523 : nor03_2x port map ( Y=>nx2522, A0=>gen_6_cmp_mReg_8, A1=>nx10037, 
      A2=>nx10425);
   ix2559 : nand02 port map ( Y=>gen_6_cmp_BSCmp_op2_9, A0=>nx4469, A1=>
      nx4473);
   ix4470 : nor02_2x port map ( Y=>nx4469, A0=>nx2554, A1=>nx2550);
   ix2555 : nor03_2x port map ( Y=>nx2554, A0=>gen_6_cmp_mReg_8, A1=>nx9623, 
      A2=>nx10393);
   ix2551 : nor03_2x port map ( Y=>nx2550, A0=>nx4463, A1=>nx10399, A2=>
      nx10409);
   ix4474 : nor02_2x port map ( Y=>nx4473, A0=>nx2546, A1=>nx2544);
   ix2547 : nor03_2x port map ( Y=>nx2546, A0=>nx4477, A1=>nx9617, A2=>
      nx10417);
   gen_6_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_6_cmp_mReg_9, QB=>
      nx4477, D=>window_6_9, CLK=>start, R=>rst);
   ix2545 : nor03_2x port map ( Y=>nx2544, A0=>gen_6_cmp_mReg_9, A1=>nx10037, 
      A2=>nx10425);
   ix2581 : nand02 port map ( Y=>gen_6_cmp_BSCmp_op2_10, A0=>nx4483, A1=>
      nx4489);
   ix4484 : nor02_2x port map ( Y=>nx4483, A0=>nx2576, A1=>nx2572);
   ix2577 : nor03_2x port map ( Y=>nx2576, A0=>gen_6_cmp_mReg_9, A1=>nx9623, 
      A2=>nx10393);
   ix2573 : nor03_2x port map ( Y=>nx2572, A0=>nx4477, A1=>nx10399, A2=>
      nx10409);
   ix4490 : nor02_2x port map ( Y=>nx4489, A0=>nx2568, A1=>nx2566);
   ix2569 : nor03_2x port map ( Y=>nx2568, A0=>nx4492, A1=>nx9617, A2=>
      nx10417);
   gen_6_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_6_cmp_mReg_10, QB=>
      nx4492, D=>window_6_10, CLK=>start, R=>rst);
   ix2567 : nor03_2x port map ( Y=>nx2566, A0=>gen_6_cmp_mReg_10, A1=>
      nx10037, A2=>nx10425);
   ix2603 : nand02 port map ( Y=>gen_6_cmp_BSCmp_op2_11, A0=>nx4497, A1=>
      nx4503);
   ix4498 : nor02_2x port map ( Y=>nx4497, A0=>nx2598, A1=>nx2594);
   ix2599 : nor03_2x port map ( Y=>nx2598, A0=>gen_6_cmp_mReg_10, A1=>nx9623, 
      A2=>nx10393);
   ix2595 : nor03_2x port map ( Y=>nx2594, A0=>nx4492, A1=>nx10399, A2=>
      nx10409);
   ix4504 : nor02_2x port map ( Y=>nx4503, A0=>nx2590, A1=>nx2588);
   ix2591 : nor03_2x port map ( Y=>nx2590, A0=>nx4507, A1=>nx9617, A2=>
      nx10417);
   gen_6_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_6_cmp_mReg_11, QB=>
      nx4507, D=>window_6_11, CLK=>start, R=>rst);
   ix2589 : nor03_2x port map ( Y=>nx2588, A0=>gen_6_cmp_mReg_11, A1=>
      nx10037, A2=>nx10425);
   ix2625 : nand02 port map ( Y=>gen_6_cmp_BSCmp_op2_12, A0=>nx4513, A1=>
      nx4517);
   ix4514 : nor02_2x port map ( Y=>nx4513, A0=>nx2620, A1=>nx2616);
   ix2621 : nor03_2x port map ( Y=>nx2620, A0=>gen_6_cmp_mReg_11, A1=>nx9623, 
      A2=>nx10393);
   ix2617 : nor03_2x port map ( Y=>nx2616, A0=>nx4507, A1=>nx10399, A2=>
      nx10409);
   ix4518 : nor02_2x port map ( Y=>nx4517, A0=>nx2612, A1=>nx2610);
   ix2613 : nor03_2x port map ( Y=>nx2612, A0=>nx4521, A1=>nx9619, A2=>
      nx10417);
   gen_6_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_6_cmp_mReg_12, QB=>
      nx4521, D=>window_6_12, CLK=>start, R=>rst);
   ix2611 : nor03_2x port map ( Y=>nx2610, A0=>gen_6_cmp_mReg_12, A1=>
      nx10037, A2=>nx10425);
   ix2647 : nand02 port map ( Y=>gen_6_cmp_BSCmp_op2_13, A0=>nx4527, A1=>
      nx4533);
   ix4528 : nor02_2x port map ( Y=>nx4527, A0=>nx2642, A1=>nx2638);
   ix2643 : nor03_2x port map ( Y=>nx2642, A0=>gen_6_cmp_mReg_12, A1=>nx9625, 
      A2=>nx10395);
   ix2639 : nor03_2x port map ( Y=>nx2638, A0=>nx4521, A1=>nx10399, A2=>
      nx10411);
   ix4534 : nor02_2x port map ( Y=>nx4533, A0=>nx2634, A1=>nx2632);
   ix2635 : nor03_2x port map ( Y=>nx2634, A0=>nx4536, A1=>nx9619, A2=>
      nx10419);
   gen_6_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_6_cmp_mReg_13, QB=>
      nx4536, D=>window_6_13, CLK=>start, R=>rst);
   ix2633 : nor03_2x port map ( Y=>nx2632, A0=>gen_6_cmp_mReg_13, A1=>
      nx10037, A2=>nx10427);
   ix2669 : nand02 port map ( Y=>gen_6_cmp_BSCmp_op2_14, A0=>nx4541, A1=>
      nx4547);
   ix4542 : nor02_2x port map ( Y=>nx4541, A0=>nx2664, A1=>nx2660);
   ix2665 : nor03_2x port map ( Y=>nx2664, A0=>gen_6_cmp_mReg_13, A1=>nx9625, 
      A2=>nx10395);
   ix2661 : nor03_2x port map ( Y=>nx2660, A0=>nx4536, A1=>nx10401, A2=>
      nx10411);
   ix4548 : nor02_2x port map ( Y=>nx4547, A0=>nx2656, A1=>nx2654);
   ix2657 : nor03_2x port map ( Y=>nx2656, A0=>nx4551, A1=>nx9619, A2=>
      nx10419);
   gen_6_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_6_cmp_mReg_14, QB=>
      nx4551, D=>window_6_14, CLK=>start, R=>rst);
   ix2655 : nor03_2x port map ( Y=>nx2654, A0=>gen_6_cmp_mReg_14, A1=>
      nx10037, A2=>nx10427);
   ix2691 : nand02 port map ( Y=>gen_6_cmp_BSCmp_op2_15, A0=>nx4557, A1=>
      nx4561);
   ix4558 : nor02_2x port map ( Y=>nx4557, A0=>nx2686, A1=>nx2682);
   ix2687 : nor03_2x port map ( Y=>nx2686, A0=>gen_6_cmp_mReg_14, A1=>nx9625, 
      A2=>nx10395);
   ix2683 : nor03_2x port map ( Y=>nx2682, A0=>nx4551, A1=>nx10401, A2=>
      nx10411);
   ix4562 : nor02_2x port map ( Y=>nx4561, A0=>nx2678, A1=>nx2676);
   ix2679 : nor03_2x port map ( Y=>nx2678, A0=>nx4565, A1=>nx9619, A2=>
      nx10419);
   gen_6_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_6_cmp_mReg_15, QB=>
      nx4565, D=>window_6_15, CLK=>start, R=>rst);
   ix2677 : nor03_2x port map ( Y=>nx2676, A0=>gen_6_cmp_mReg_15, A1=>
      nx10039, A2=>nx10427);
   ix2701 : nand02 port map ( Y=>gen_6_cmp_BSCmp_op2_16, A0=>nx4571, A1=>
      nx4561);
   ix4572 : nor02_2x port map ( Y=>nx4571, A0=>nx2696, A1=>nx2692);
   ix2697 : nor03_2x port map ( Y=>nx2696, A0=>gen_6_cmp_mReg_15, A1=>nx9625, 
      A2=>nx10395);
   ix2693 : nor03_2x port map ( Y=>nx2692, A0=>nx4565, A1=>nx10401, A2=>
      nx10411);
   ix2769 : nand02 port map ( Y=>gen_7_cmp_BSCmp_op2_1, A0=>nx4579, A1=>
      nx4597);
   ix4580 : nor02_2x port map ( Y=>nx4579, A0=>nx2764, A1=>nx2760);
   ix2765 : nor03_2x port map ( Y=>nx2764, A0=>gen_7_cmp_mReg_0, A1=>nx9609, 
      A2=>nx10431);
   gen_7_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_7_cmp_mReg_0, QB=>
      nx4583, D=>window_7_0, CLK=>start, R=>rst);
   ix4588 : inv01 port map ( Y=>nx4587, A=>gen_7_cmp_pMux_0);
   ix2761 : nor03_2x port map ( Y=>nx2760, A0=>nx4583, A1=>nx10437, A2=>
      nx10447);
   ix4596 : inv02 port map ( Y=>nx4595, A=>gen_7_cmp_pMux_2);
   ix4598 : nor02_2x port map ( Y=>nx4597, A0=>nx2750, A1=>nx2748);
   ix2751 : nor03_2x port map ( Y=>nx2750, A0=>nx4601, A1=>nx9603, A2=>
      nx10455);
   gen_7_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_7_cmp_mReg_1, QB=>
      nx4601, D=>window_7_1, CLK=>start, R=>rst);
   ix2749 : nor03_2x port map ( Y=>nx2748, A0=>gen_7_cmp_mReg_1, A1=>nx10041, 
      A2=>nx10463);
   ix2709 : nor03_2x port map ( Y=>nx2708, A0=>nx9609, A1=>nx4595, A2=>
      gen_7_cmp_pMux_0);
   ix2791 : nand02 port map ( Y=>gen_7_cmp_BSCmp_op2_2, A0=>nx4613, A1=>
      nx4617);
   ix4614 : nor02_2x port map ( Y=>nx4613, A0=>nx2786, A1=>nx2782);
   ix2787 : nor03_2x port map ( Y=>nx2786, A0=>gen_7_cmp_mReg_1, A1=>nx9609, 
      A2=>nx10431);
   ix2783 : nor03_2x port map ( Y=>nx2782, A0=>nx4601, A1=>nx10437, A2=>
      nx10447);
   ix4618 : nor02_2x port map ( Y=>nx4617, A0=>nx2778, A1=>nx2776);
   ix2779 : nor03_2x port map ( Y=>nx2778, A0=>nx4621, A1=>nx9603, A2=>
      nx10455);
   gen_7_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_7_cmp_mReg_2, QB=>
      nx4621, D=>window_7_2, CLK=>start, R=>rst);
   ix2777 : nor03_2x port map ( Y=>nx2776, A0=>gen_7_cmp_mReg_2, A1=>nx10041, 
      A2=>nx10463);
   ix2813 : nand02 port map ( Y=>gen_7_cmp_BSCmp_op2_3, A0=>nx4627, A1=>
      nx4633);
   ix4628 : nor02_2x port map ( Y=>nx4627, A0=>nx2808, A1=>nx2804);
   ix2809 : nor03_2x port map ( Y=>nx2808, A0=>gen_7_cmp_mReg_2, A1=>nx9609, 
      A2=>nx10431);
   ix2805 : nor03_2x port map ( Y=>nx2804, A0=>nx4621, A1=>nx10437, A2=>
      nx10447);
   ix4634 : nor02_2x port map ( Y=>nx4633, A0=>nx2800, A1=>nx2798);
   ix2801 : nor03_2x port map ( Y=>nx2800, A0=>nx4637, A1=>nx9603, A2=>
      nx10455);
   gen_7_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_7_cmp_mReg_3, QB=>
      nx4637, D=>window_7_3, CLK=>start, R=>rst);
   ix2799 : nor03_2x port map ( Y=>nx2798, A0=>gen_7_cmp_mReg_3, A1=>nx10041, 
      A2=>nx10463);
   ix2835 : nand02 port map ( Y=>gen_7_cmp_BSCmp_op2_4, A0=>nx4642, A1=>
      nx4646);
   ix4643 : nor02_2x port map ( Y=>nx4642, A0=>nx2830, A1=>nx2826);
   ix2831 : nor03_2x port map ( Y=>nx2830, A0=>gen_7_cmp_mReg_3, A1=>nx9609, 
      A2=>nx10431);
   ix2827 : nor03_2x port map ( Y=>nx2826, A0=>nx4637, A1=>nx10437, A2=>
      nx10447);
   ix4647 : nor02_2x port map ( Y=>nx4646, A0=>nx2822, A1=>nx2820);
   ix2823 : nor03_2x port map ( Y=>nx2822, A0=>nx4649, A1=>nx9603, A2=>
      nx10455);
   gen_7_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_7_cmp_mReg_4, QB=>
      nx4649, D=>window_7_4, CLK=>start, R=>rst);
   ix2821 : nor03_2x port map ( Y=>nx2820, A0=>gen_7_cmp_mReg_4, A1=>nx10041, 
      A2=>nx10463);
   ix2857 : nand02 port map ( Y=>gen_7_cmp_BSCmp_op2_5, A0=>nx4655, A1=>
      nx4661);
   ix4656 : nor02_2x port map ( Y=>nx4655, A0=>nx2852, A1=>nx2848);
   ix2853 : nor03_2x port map ( Y=>nx2852, A0=>gen_7_cmp_mReg_4, A1=>nx9609, 
      A2=>nx10431);
   ix2849 : nor03_2x port map ( Y=>nx2848, A0=>nx4649, A1=>nx10437, A2=>
      nx10447);
   ix4662 : nor02_2x port map ( Y=>nx4661, A0=>nx2844, A1=>nx2842);
   ix2845 : nor03_2x port map ( Y=>nx2844, A0=>nx4665, A1=>nx9605, A2=>
      nx10455);
   gen_7_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_7_cmp_mReg_5, QB=>
      nx4665, D=>window_7_5, CLK=>start, R=>rst);
   ix2843 : nor03_2x port map ( Y=>nx2842, A0=>gen_7_cmp_mReg_5, A1=>nx10041, 
      A2=>nx10463);
   ix2879 : nand02 port map ( Y=>gen_7_cmp_BSCmp_op2_6, A0=>nx4671, A1=>
      nx4675);
   ix4672 : nor02_2x port map ( Y=>nx4671, A0=>nx2874, A1=>nx2870);
   ix2875 : nor03_2x port map ( Y=>nx2874, A0=>gen_7_cmp_mReg_5, A1=>nx9611, 
      A2=>nx10431);
   ix2871 : nor03_2x port map ( Y=>nx2870, A0=>nx4665, A1=>nx10437, A2=>
      nx10447);
   ix4676 : nor02_2x port map ( Y=>nx4675, A0=>nx2866, A1=>nx2864);
   ix2867 : nor03_2x port map ( Y=>nx2866, A0=>nx4679, A1=>nx9605, A2=>
      nx10455);
   gen_7_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_7_cmp_mReg_6, QB=>
      nx4679, D=>window_7_6, CLK=>start, R=>rst);
   ix2865 : nor03_2x port map ( Y=>nx2864, A0=>gen_7_cmp_mReg_6, A1=>nx10041, 
      A2=>nx10463);
   ix2901 : nand02 port map ( Y=>gen_7_cmp_BSCmp_op2_7, A0=>nx4685, A1=>
      nx4691);
   ix4686 : nor02_2x port map ( Y=>nx4685, A0=>nx2896, A1=>nx2892);
   ix2897 : nor03_2x port map ( Y=>nx2896, A0=>gen_7_cmp_mReg_6, A1=>nx9611, 
      A2=>nx10433);
   ix2893 : nor03_2x port map ( Y=>nx2892, A0=>nx4679, A1=>nx10439, A2=>
      nx10449);
   ix4692 : nor02_2x port map ( Y=>nx4691, A0=>nx2888, A1=>nx2886);
   ix2889 : nor03_2x port map ( Y=>nx2888, A0=>nx4695, A1=>nx9605, A2=>
      nx10457);
   gen_7_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_7_cmp_mReg_7, QB=>
      nx4695, D=>window_7_7, CLK=>start, R=>rst);
   ix2887 : nor03_2x port map ( Y=>nx2886, A0=>gen_7_cmp_mReg_7, A1=>nx10041, 
      A2=>nx10465);
   ix2923 : nand02 port map ( Y=>gen_7_cmp_BSCmp_op2_8, A0=>nx4701, A1=>
      nx4705);
   ix4702 : nor02_2x port map ( Y=>nx4701, A0=>nx2918, A1=>nx2914);
   ix2919 : nor03_2x port map ( Y=>nx2918, A0=>gen_7_cmp_mReg_7, A1=>nx9611, 
      A2=>nx10433);
   ix2915 : nor03_2x port map ( Y=>nx2914, A0=>nx4695, A1=>nx10439, A2=>
      nx10449);
   ix4706 : nor02_2x port map ( Y=>nx4705, A0=>nx2910, A1=>nx2908);
   ix2911 : nor03_2x port map ( Y=>nx2910, A0=>nx4709, A1=>nx9605, A2=>
      nx10457);
   gen_7_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_7_cmp_mReg_8, QB=>
      nx4709, D=>window_7_8, CLK=>start, R=>rst);
   ix2909 : nor03_2x port map ( Y=>nx2908, A0=>gen_7_cmp_mReg_8, A1=>nx10043, 
      A2=>nx10465);
   ix2945 : nand02 port map ( Y=>gen_7_cmp_BSCmp_op2_9, A0=>nx4715, A1=>
      nx4721);
   ix4716 : nor02_2x port map ( Y=>nx4715, A0=>nx2940, A1=>nx2936);
   ix2941 : nor03_2x port map ( Y=>nx2940, A0=>gen_7_cmp_mReg_8, A1=>nx9611, 
      A2=>nx10433);
   ix2937 : nor03_2x port map ( Y=>nx2936, A0=>nx4709, A1=>nx10439, A2=>
      nx10449);
   ix4722 : nor02_2x port map ( Y=>nx4721, A0=>nx2932, A1=>nx2930);
   ix2933 : nor03_2x port map ( Y=>nx2932, A0=>nx4724, A1=>nx9605, A2=>
      nx10457);
   gen_7_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_7_cmp_mReg_9, QB=>
      nx4724, D=>window_7_9, CLK=>start, R=>rst);
   ix2931 : nor03_2x port map ( Y=>nx2930, A0=>gen_7_cmp_mReg_9, A1=>nx10043, 
      A2=>nx10465);
   ix2967 : nand02 port map ( Y=>gen_7_cmp_BSCmp_op2_10, A0=>nx4729, A1=>
      nx4735);
   ix4730 : nor02_2x port map ( Y=>nx4729, A0=>nx2962, A1=>nx2958);
   ix2963 : nor03_2x port map ( Y=>nx2962, A0=>gen_7_cmp_mReg_9, A1=>nx9611, 
      A2=>nx10433);
   ix2959 : nor03_2x port map ( Y=>nx2958, A0=>nx4724, A1=>nx10439, A2=>
      nx10449);
   ix4736 : nor02_2x port map ( Y=>nx4735, A0=>nx2954, A1=>nx2952);
   ix2955 : nor03_2x port map ( Y=>nx2954, A0=>nx4739, A1=>nx9605, A2=>
      nx10457);
   gen_7_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_7_cmp_mReg_10, QB=>
      nx4739, D=>window_7_10, CLK=>start, R=>rst);
   ix2953 : nor03_2x port map ( Y=>nx2952, A0=>gen_7_cmp_mReg_10, A1=>
      nx10043, A2=>nx10465);
   ix2989 : nand02 port map ( Y=>gen_7_cmp_BSCmp_op2_11, A0=>nx4745, A1=>
      nx4749);
   ix4746 : nor02_2x port map ( Y=>nx4745, A0=>nx2984, A1=>nx2980);
   ix2985 : nor03_2x port map ( Y=>nx2984, A0=>gen_7_cmp_mReg_10, A1=>nx9611, 
      A2=>nx10433);
   ix2981 : nor03_2x port map ( Y=>nx2980, A0=>nx4739, A1=>nx10439, A2=>
      nx10449);
   ix4750 : nor02_2x port map ( Y=>nx4749, A0=>nx2976, A1=>nx2974);
   ix2977 : nor03_2x port map ( Y=>nx2976, A0=>nx4753, A1=>nx9605, A2=>
      nx10457);
   gen_7_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_7_cmp_mReg_11, QB=>
      nx4753, D=>window_7_11, CLK=>start, R=>rst);
   ix2975 : nor03_2x port map ( Y=>nx2974, A0=>gen_7_cmp_mReg_11, A1=>
      nx10043, A2=>nx10465);
   ix3011 : nand02 port map ( Y=>gen_7_cmp_BSCmp_op2_12, A0=>nx4759, A1=>
      nx4765);
   ix4760 : nor02_2x port map ( Y=>nx4759, A0=>nx3006, A1=>nx3002);
   ix3007 : nor03_2x port map ( Y=>nx3006, A0=>gen_7_cmp_mReg_11, A1=>nx9611, 
      A2=>nx10433);
   ix3003 : nor03_2x port map ( Y=>nx3002, A0=>nx4753, A1=>nx10439, A2=>
      nx10449);
   ix4766 : nor02_2x port map ( Y=>nx4765, A0=>nx2998, A1=>nx2996);
   ix2999 : nor03_2x port map ( Y=>nx2998, A0=>nx4768, A1=>nx9607, A2=>
      nx10457);
   gen_7_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_7_cmp_mReg_12, QB=>
      nx4768, D=>window_7_12, CLK=>start, R=>rst);
   ix2997 : nor03_2x port map ( Y=>nx2996, A0=>gen_7_cmp_mReg_12, A1=>
      nx10043, A2=>nx10465);
   ix3033 : nand02 port map ( Y=>gen_7_cmp_BSCmp_op2_13, A0=>nx4773, A1=>
      nx4779);
   ix4774 : nor02_2x port map ( Y=>nx4773, A0=>nx3028, A1=>nx3024);
   ix3029 : nor03_2x port map ( Y=>nx3028, A0=>gen_7_cmp_mReg_12, A1=>nx9613, 
      A2=>nx10435);
   ix3025 : nor03_2x port map ( Y=>nx3024, A0=>nx4768, A1=>nx10439, A2=>
      nx10451);
   ix4780 : nor02_2x port map ( Y=>nx4779, A0=>nx3020, A1=>nx3018);
   ix3021 : nor03_2x port map ( Y=>nx3020, A0=>nx4783, A1=>nx9607, A2=>
      nx10459);
   gen_7_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_7_cmp_mReg_13, QB=>
      nx4783, D=>window_7_13, CLK=>start, R=>rst);
   ix3019 : nor03_2x port map ( Y=>nx3018, A0=>gen_7_cmp_mReg_13, A1=>
      nx10043, A2=>nx10467);
   ix3055 : nand02 port map ( Y=>gen_7_cmp_BSCmp_op2_14, A0=>nx4789, A1=>
      nx4793);
   ix4790 : nor02_2x port map ( Y=>nx4789, A0=>nx3050, A1=>nx3046);
   ix3051 : nor03_2x port map ( Y=>nx3050, A0=>gen_7_cmp_mReg_13, A1=>nx9613, 
      A2=>nx10435);
   ix3047 : nor03_2x port map ( Y=>nx3046, A0=>nx4783, A1=>nx10441, A2=>
      nx10451);
   ix4794 : nor02_2x port map ( Y=>nx4793, A0=>nx3042, A1=>nx3040);
   ix3043 : nor03_2x port map ( Y=>nx3042, A0=>nx4797, A1=>nx9607, A2=>
      nx10459);
   gen_7_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_7_cmp_mReg_14, QB=>
      nx4797, D=>window_7_14, CLK=>start, R=>rst);
   ix3041 : nor03_2x port map ( Y=>nx3040, A0=>gen_7_cmp_mReg_14, A1=>
      nx10043, A2=>nx10467);
   ix3077 : nand02 port map ( Y=>gen_7_cmp_BSCmp_op2_15, A0=>nx4803, A1=>
      nx4809);
   ix4804 : nor02_2x port map ( Y=>nx4803, A0=>nx3072, A1=>nx3068);
   ix3073 : nor03_2x port map ( Y=>nx3072, A0=>gen_7_cmp_mReg_14, A1=>nx9613, 
      A2=>nx10435);
   ix3069 : nor03_2x port map ( Y=>nx3068, A0=>nx4797, A1=>nx10441, A2=>
      nx10451);
   ix4810 : nor02_2x port map ( Y=>nx4809, A0=>nx3064, A1=>nx3062);
   ix3065 : nor03_2x port map ( Y=>nx3064, A0=>nx4812, A1=>nx9607, A2=>
      nx10459);
   gen_7_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_7_cmp_mReg_15, QB=>
      nx4812, D=>window_7_15, CLK=>start, R=>rst);
   ix3063 : nor03_2x port map ( Y=>nx3062, A0=>gen_7_cmp_mReg_15, A1=>
      nx10045, A2=>nx10467);
   ix3087 : nand02 port map ( Y=>gen_7_cmp_BSCmp_op2_16, A0=>nx4817, A1=>
      nx4809);
   ix4818 : nor02_2x port map ( Y=>nx4817, A0=>nx3082, A1=>nx3078);
   ix3083 : nor03_2x port map ( Y=>nx3082, A0=>gen_7_cmp_mReg_15, A1=>nx9613, 
      A2=>nx10435);
   ix3079 : nor03_2x port map ( Y=>nx3078, A0=>nx4812, A1=>nx10441, A2=>
      nx10451);
   ix3155 : nand02 port map ( Y=>gen_8_cmp_BSCmp_op2_1, A0=>nx4825, A1=>
      nx4843);
   ix4826 : nor02_2x port map ( Y=>nx4825, A0=>nx3150, A1=>nx3146);
   ix3151 : nor03_2x port map ( Y=>nx3150, A0=>gen_8_cmp_mReg_0, A1=>nx9597, 
      A2=>nx10471);
   gen_8_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_8_cmp_mReg_0, QB=>
      nx4831, D=>window_8_0, CLK=>start, R=>rst);
   ix4835 : inv01 port map ( Y=>nx4834, A=>gen_8_cmp_pMux_0);
   ix3147 : nor03_2x port map ( Y=>nx3146, A0=>nx4831, A1=>nx10477, A2=>
      nx10487);
   ix4842 : inv02 port map ( Y=>nx4841, A=>gen_8_cmp_pMux_2);
   ix4844 : nor02_2x port map ( Y=>nx4843, A0=>nx3136, A1=>nx3134);
   ix3137 : nor03_2x port map ( Y=>nx3136, A0=>nx4847, A1=>nx9591, A2=>
      nx10495);
   gen_8_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_8_cmp_mReg_1, QB=>
      nx4847, D=>window_8_1, CLK=>start, R=>rst);
   ix3135 : nor03_2x port map ( Y=>nx3134, A0=>gen_8_cmp_mReg_1, A1=>nx10047, 
      A2=>nx10503);
   ix3095 : nor03_2x port map ( Y=>nx3094, A0=>nx9597, A1=>nx4841, A2=>
      gen_8_cmp_pMux_0);
   ix3177 : nand02 port map ( Y=>gen_8_cmp_BSCmp_op2_2, A0=>nx4858, A1=>
      nx4865);
   ix4860 : nor02_2x port map ( Y=>nx4858, A0=>nx3172, A1=>nx3168);
   ix3173 : nor03_2x port map ( Y=>nx3172, A0=>gen_8_cmp_mReg_1, A1=>nx9597, 
      A2=>nx10471);
   ix3169 : nor03_2x port map ( Y=>nx3168, A0=>nx4847, A1=>nx10477, A2=>
      nx10487);
   ix4866 : nor02_2x port map ( Y=>nx4865, A0=>nx3164, A1=>nx3162);
   ix3165 : nor03_2x port map ( Y=>nx3164, A0=>nx4869, A1=>nx9591, A2=>
      nx10495);
   gen_8_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_8_cmp_mReg_2, QB=>
      nx4869, D=>window_8_2, CLK=>start, R=>rst);
   ix3163 : nor03_2x port map ( Y=>nx3162, A0=>gen_8_cmp_mReg_2, A1=>nx10047, 
      A2=>nx10503);
   ix3199 : nand02 port map ( Y=>gen_8_cmp_BSCmp_op2_3, A0=>nx4875, A1=>
      nx4879);
   ix4876 : nor02_2x port map ( Y=>nx4875, A0=>nx3194, A1=>nx3190);
   ix3195 : nor03_2x port map ( Y=>nx3194, A0=>gen_8_cmp_mReg_2, A1=>nx9597, 
      A2=>nx10471);
   ix3191 : nor03_2x port map ( Y=>nx3190, A0=>nx4869, A1=>nx10477, A2=>
      nx10487);
   ix4880 : nor02_2x port map ( Y=>nx4879, A0=>nx3186, A1=>nx3184);
   ix3187 : nor03_2x port map ( Y=>nx3186, A0=>nx4883, A1=>nx9591, A2=>
      nx10495);
   gen_8_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_8_cmp_mReg_3, QB=>
      nx4883, D=>window_8_3, CLK=>start, R=>rst);
   ix3185 : nor03_2x port map ( Y=>nx3184, A0=>gen_8_cmp_mReg_3, A1=>nx10047, 
      A2=>nx10503);
   ix3221 : nand02 port map ( Y=>gen_8_cmp_BSCmp_op2_4, A0=>nx4889, A1=>
      nx4893);
   ix4890 : nor02_2x port map ( Y=>nx4889, A0=>nx3216, A1=>nx3212);
   ix3217 : nor03_2x port map ( Y=>nx3216, A0=>gen_8_cmp_mReg_3, A1=>nx9597, 
      A2=>nx10471);
   ix3213 : nor03_2x port map ( Y=>nx3212, A0=>nx4883, A1=>nx10477, A2=>
      nx10487);
   ix4894 : nor02_2x port map ( Y=>nx4893, A0=>nx3208, A1=>nx3206);
   ix3209 : nor03_2x port map ( Y=>nx3208, A0=>nx4897, A1=>nx9591, A2=>
      nx10495);
   gen_8_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_8_cmp_mReg_4, QB=>
      nx4897, D=>window_8_4, CLK=>start, R=>rst);
   ix3207 : nor03_2x port map ( Y=>nx3206, A0=>gen_8_cmp_mReg_4, A1=>nx10047, 
      A2=>nx10503);
   ix3243 : nand02 port map ( Y=>gen_8_cmp_BSCmp_op2_5, A0=>nx4901, A1=>
      nx4907);
   ix4902 : nor02_2x port map ( Y=>nx4901, A0=>nx3238, A1=>nx3234);
   ix3239 : nor03_2x port map ( Y=>nx3238, A0=>gen_8_cmp_mReg_4, A1=>nx9597, 
      A2=>nx10471);
   ix3235 : nor03_2x port map ( Y=>nx3234, A0=>nx4897, A1=>nx10477, A2=>
      nx10487);
   ix4908 : nor02_2x port map ( Y=>nx4907, A0=>nx3230, A1=>nx3228);
   ix3231 : nor03_2x port map ( Y=>nx3230, A0=>nx4911, A1=>nx9593, A2=>
      nx10495);
   gen_8_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_8_cmp_mReg_5, QB=>
      nx4911, D=>window_8_5, CLK=>start, R=>rst);
   ix3229 : nor03_2x port map ( Y=>nx3228, A0=>gen_8_cmp_mReg_5, A1=>nx10047, 
      A2=>nx10503);
   ix3265 : nand02 port map ( Y=>gen_8_cmp_BSCmp_op2_6, A0=>nx4915, A1=>
      nx4921);
   ix4916 : nor02_2x port map ( Y=>nx4915, A0=>nx3260, A1=>nx3256);
   ix3261 : nor03_2x port map ( Y=>nx3260, A0=>gen_8_cmp_mReg_5, A1=>nx9599, 
      A2=>nx10471);
   ix3257 : nor03_2x port map ( Y=>nx3256, A0=>nx4911, A1=>nx10477, A2=>
      nx10487);
   ix4922 : nor02_2x port map ( Y=>nx4921, A0=>nx3252, A1=>nx3250);
   ix3253 : nor03_2x port map ( Y=>nx3252, A0=>nx4924, A1=>nx9593, A2=>
      nx10495);
   gen_8_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_8_cmp_mReg_6, QB=>
      nx4924, D=>window_8_6, CLK=>start, R=>rst);
   ix3251 : nor03_2x port map ( Y=>nx3250, A0=>gen_8_cmp_mReg_6, A1=>nx10047, 
      A2=>nx10503);
   ix3287 : nand02 port map ( Y=>gen_8_cmp_BSCmp_op2_7, A0=>nx4931, A1=>
      nx4937);
   ix4932 : nor02_2x port map ( Y=>nx4931, A0=>nx3282, A1=>nx3278);
   ix3283 : nor03_2x port map ( Y=>nx3282, A0=>gen_8_cmp_mReg_6, A1=>nx9599, 
      A2=>nx10473);
   ix3279 : nor03_2x port map ( Y=>nx3278, A0=>nx4924, A1=>nx10479, A2=>
      nx10489);
   ix4938 : nor02_2x port map ( Y=>nx4937, A0=>nx3274, A1=>nx3272);
   ix3275 : nor03_2x port map ( Y=>nx3274, A0=>nx4941, A1=>nx9593, A2=>
      nx10497);
   gen_8_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_8_cmp_mReg_7, QB=>
      nx4941, D=>window_8_7, CLK=>start, R=>rst);
   ix3273 : nor03_2x port map ( Y=>nx3272, A0=>gen_8_cmp_mReg_7, A1=>nx10047, 
      A2=>nx10505);
   ix3309 : nand02 port map ( Y=>gen_8_cmp_BSCmp_op2_8, A0=>nx4945, A1=>
      nx4951);
   ix4946 : nor02_2x port map ( Y=>nx4945, A0=>nx3304, A1=>nx3300);
   ix3305 : nor03_2x port map ( Y=>nx3304, A0=>gen_8_cmp_mReg_7, A1=>nx9599, 
      A2=>nx10473);
   ix3301 : nor03_2x port map ( Y=>nx3300, A0=>nx4941, A1=>nx10479, A2=>
      nx10489);
   ix4952 : nor02_2x port map ( Y=>nx4951, A0=>nx3296, A1=>nx3294);
   ix3297 : nor03_2x port map ( Y=>nx3296, A0=>nx4955, A1=>nx9593, A2=>
      nx10497);
   gen_8_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_8_cmp_mReg_8, QB=>
      nx4955, D=>window_8_8, CLK=>start, R=>rst);
   ix3295 : nor03_2x port map ( Y=>nx3294, A0=>gen_8_cmp_mReg_8, A1=>nx10049, 
      A2=>nx10505);
   ix3331 : nand02 port map ( Y=>gen_8_cmp_BSCmp_op2_9, A0=>nx4959, A1=>
      nx4965);
   ix4960 : nor02_2x port map ( Y=>nx4959, A0=>nx3326, A1=>nx3322);
   ix3327 : nor03_2x port map ( Y=>nx3326, A0=>gen_8_cmp_mReg_8, A1=>nx9599, 
      A2=>nx10473);
   ix3323 : nor03_2x port map ( Y=>nx3322, A0=>nx4955, A1=>nx10479, A2=>
      nx10489);
   ix4966 : nor02_2x port map ( Y=>nx4965, A0=>nx3318, A1=>nx3316);
   ix3319 : nor03_2x port map ( Y=>nx3318, A0=>nx4968, A1=>nx9593, A2=>
      nx10497);
   gen_8_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_8_cmp_mReg_9, QB=>
      nx4968, D=>window_8_9, CLK=>start, R=>rst);
   ix3317 : nor03_2x port map ( Y=>nx3316, A0=>gen_8_cmp_mReg_9, A1=>nx10049, 
      A2=>nx10505);
   ix3353 : nand02 port map ( Y=>gen_8_cmp_BSCmp_op2_10, A0=>nx4975, A1=>
      nx4981);
   ix4976 : nor02_2x port map ( Y=>nx4975, A0=>nx3348, A1=>nx3344);
   ix3349 : nor03_2x port map ( Y=>nx3348, A0=>gen_8_cmp_mReg_9, A1=>nx9599, 
      A2=>nx10473);
   ix3345 : nor03_2x port map ( Y=>nx3344, A0=>nx4968, A1=>nx10479, A2=>
      nx10489);
   ix4982 : nor02_2x port map ( Y=>nx4981, A0=>nx3340, A1=>nx3338);
   ix3341 : nor03_2x port map ( Y=>nx3340, A0=>nx4985, A1=>nx9593, A2=>
      nx10497);
   gen_8_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_8_cmp_mReg_10, QB=>
      nx4985, D=>window_8_10, CLK=>start, R=>rst);
   ix3339 : nor03_2x port map ( Y=>nx3338, A0=>gen_8_cmp_mReg_10, A1=>
      nx10049, A2=>nx10505);
   ix3375 : nand02 port map ( Y=>gen_8_cmp_BSCmp_op2_11, A0=>nx4989, A1=>
      nx4995);
   ix4990 : nor02_2x port map ( Y=>nx4989, A0=>nx3370, A1=>nx3366);
   ix3371 : nor03_2x port map ( Y=>nx3370, A0=>gen_8_cmp_mReg_10, A1=>nx9599, 
      A2=>nx10473);
   ix3367 : nor03_2x port map ( Y=>nx3366, A0=>nx4985, A1=>nx10479, A2=>
      nx10489);
   ix4996 : nor02_2x port map ( Y=>nx4995, A0=>nx3362, A1=>nx3360);
   ix3363 : nor03_2x port map ( Y=>nx3362, A0=>nx4999, A1=>nx9593, A2=>
      nx10497);
   gen_8_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_8_cmp_mReg_11, QB=>
      nx4999, D=>window_8_11, CLK=>start, R=>rst);
   ix3361 : nor03_2x port map ( Y=>nx3360, A0=>gen_8_cmp_mReg_11, A1=>
      nx10049, A2=>nx10505);
   ix3397 : nand02 port map ( Y=>gen_8_cmp_BSCmp_op2_12, A0=>nx5003, A1=>
      nx5009);
   ix5004 : nor02_2x port map ( Y=>nx5003, A0=>nx3392, A1=>nx3388);
   ix3393 : nor03_2x port map ( Y=>nx3392, A0=>gen_8_cmp_mReg_11, A1=>nx9599, 
      A2=>nx10473);
   ix3389 : nor03_2x port map ( Y=>nx3388, A0=>nx4999, A1=>nx10479, A2=>
      nx10489);
   ix5010 : nor02_2x port map ( Y=>nx5009, A0=>nx3384, A1=>nx3382);
   ix3385 : nor03_2x port map ( Y=>nx3384, A0=>nx5013, A1=>nx9595, A2=>
      nx10497);
   gen_8_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_8_cmp_mReg_12, QB=>
      nx5013, D=>window_8_12, CLK=>start, R=>rst);
   ix3383 : nor03_2x port map ( Y=>nx3382, A0=>gen_8_cmp_mReg_12, A1=>
      nx10049, A2=>nx10505);
   ix3419 : nand02 port map ( Y=>gen_8_cmp_BSCmp_op2_13, A0=>nx5019, A1=>
      nx5025);
   ix5020 : nor02_2x port map ( Y=>nx5019, A0=>nx3414, A1=>nx3410);
   ix3415 : nor03_2x port map ( Y=>nx3414, A0=>gen_8_cmp_mReg_12, A1=>nx9601, 
      A2=>nx10475);
   ix3411 : nor03_2x port map ( Y=>nx3410, A0=>nx5013, A1=>nx10479, A2=>
      nx10491);
   ix5026 : nor02_2x port map ( Y=>nx5025, A0=>nx3406, A1=>nx3404);
   ix3407 : nor03_2x port map ( Y=>nx3406, A0=>nx5028, A1=>nx9595, A2=>
      nx10499);
   gen_8_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_8_cmp_mReg_13, QB=>
      nx5028, D=>window_8_13, CLK=>start, R=>rst);
   ix3405 : nor03_2x port map ( Y=>nx3404, A0=>gen_8_cmp_mReg_13, A1=>
      nx10049, A2=>nx10507);
   ix3441 : nand02 port map ( Y=>gen_8_cmp_BSCmp_op2_14, A0=>nx5032, A1=>
      nx5037);
   ix5033 : nor02_2x port map ( Y=>nx5032, A0=>nx3436, A1=>nx3432);
   ix3437 : nor03_2x port map ( Y=>nx3436, A0=>gen_8_cmp_mReg_13, A1=>nx9601, 
      A2=>nx10475);
   ix3433 : nor03_2x port map ( Y=>nx3432, A0=>nx5028, A1=>nx10481, A2=>
      nx10491);
   ix5038 : nor02_2x port map ( Y=>nx5037, A0=>nx3428, A1=>nx3426);
   ix3429 : nor03_2x port map ( Y=>nx3428, A0=>nx5041, A1=>nx9595, A2=>
      nx10499);
   gen_8_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_8_cmp_mReg_14, QB=>
      nx5041, D=>window_8_14, CLK=>start, R=>rst);
   ix3427 : nor03_2x port map ( Y=>nx3426, A0=>gen_8_cmp_mReg_14, A1=>
      nx10049, A2=>nx10507);
   ix3463 : nand02 port map ( Y=>gen_8_cmp_BSCmp_op2_15, A0=>nx5047, A1=>
      nx5053);
   ix5048 : nor02_2x port map ( Y=>nx5047, A0=>nx3458, A1=>nx3454);
   ix3459 : nor03_2x port map ( Y=>nx3458, A0=>gen_8_cmp_mReg_14, A1=>nx9601, 
      A2=>nx10475);
   ix3455 : nor03_2x port map ( Y=>nx3454, A0=>nx5041, A1=>nx10481, A2=>
      nx10491);
   ix5054 : nor02_2x port map ( Y=>nx5053, A0=>nx3450, A1=>nx3448);
   ix3451 : nor03_2x port map ( Y=>nx3450, A0=>nx5057, A1=>nx9595, A2=>
      nx10499);
   gen_8_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_8_cmp_mReg_15, QB=>
      nx5057, D=>window_8_15, CLK=>start, R=>rst);
   ix3449 : nor03_2x port map ( Y=>nx3448, A0=>gen_8_cmp_mReg_15, A1=>
      nx10051, A2=>nx10507);
   ix3473 : nand02 port map ( Y=>gen_8_cmp_BSCmp_op2_16, A0=>nx5061, A1=>
      nx5053);
   ix5062 : nor02_2x port map ( Y=>nx5061, A0=>nx3468, A1=>nx3464);
   ix3469 : nor03_2x port map ( Y=>nx3468, A0=>gen_8_cmp_mReg_15, A1=>nx9601, 
      A2=>nx10475);
   ix3465 : nor03_2x port map ( Y=>nx3464, A0=>nx5057, A1=>nx10481, A2=>
      nx10491);
   ix3541 : nand02 port map ( Y=>gen_9_cmp_BSCmp_op2_1, A0=>nx5069, A1=>
      nx5087);
   ix5070 : nor02_2x port map ( Y=>nx5069, A0=>nx3536, A1=>nx3532);
   ix3537 : nor03_2x port map ( Y=>nx3536, A0=>gen_9_cmp_mReg_0, A1=>nx9585, 
      A2=>nx10511);
   gen_9_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_9_cmp_mReg_0, QB=>
      nx5073, D=>window_9_0, CLK=>start, R=>rst);
   ix5078 : inv01 port map ( Y=>nx5077, A=>gen_9_cmp_pMux_0);
   ix3533 : nor03_2x port map ( Y=>nx3532, A0=>nx5073, A1=>nx10517, A2=>
      nx10527);
   ix5086 : inv02 port map ( Y=>nx5085, A=>gen_9_cmp_pMux_2);
   ix5088 : nor02_2x port map ( Y=>nx5087, A0=>nx3522, A1=>nx3520);
   ix3523 : nor03_2x port map ( Y=>nx3522, A0=>nx5090, A1=>nx9579, A2=>
      nx10535);
   gen_9_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_9_cmp_mReg_1, QB=>
      nx5090, D=>window_9_1, CLK=>start, R=>rst);
   ix3521 : nor03_2x port map ( Y=>nx3520, A0=>gen_9_cmp_mReg_1, A1=>nx10053, 
      A2=>nx10543);
   ix3481 : nor03_2x port map ( Y=>nx3480, A0=>nx9585, A1=>nx5085, A2=>
      gen_9_cmp_pMux_0);
   ix3563 : nand02 port map ( Y=>gen_9_cmp_BSCmp_op2_2, A0=>nx5103, A1=>
      nx5109);
   ix5104 : nor02_2x port map ( Y=>nx5103, A0=>nx3558, A1=>nx3554);
   ix3559 : nor03_2x port map ( Y=>nx3558, A0=>gen_9_cmp_mReg_1, A1=>nx9585, 
      A2=>nx10511);
   ix3555 : nor03_2x port map ( Y=>nx3554, A0=>nx5090, A1=>nx10517, A2=>
      nx10527);
   ix5110 : nor02_2x port map ( Y=>nx5109, A0=>nx3550, A1=>nx3548);
   ix3551 : nor03_2x port map ( Y=>nx3550, A0=>nx5112, A1=>nx9579, A2=>
      nx10535);
   gen_9_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_9_cmp_mReg_2, QB=>
      nx5112, D=>window_9_2, CLK=>start, R=>rst);
   ix3549 : nor03_2x port map ( Y=>nx3548, A0=>gen_9_cmp_mReg_2, A1=>nx10053, 
      A2=>nx10543);
   ix3585 : nand02 port map ( Y=>gen_9_cmp_BSCmp_op2_3, A0=>nx5119, A1=>
      nx5125);
   ix5120 : nor02_2x port map ( Y=>nx5119, A0=>nx3580, A1=>nx3576);
   ix3581 : nor03_2x port map ( Y=>nx3580, A0=>gen_9_cmp_mReg_2, A1=>nx9585, 
      A2=>nx10511);
   ix3577 : nor03_2x port map ( Y=>nx3576, A0=>nx5112, A1=>nx10517, A2=>
      nx10527);
   ix5126 : nor02_2x port map ( Y=>nx5125, A0=>nx3572, A1=>nx3570);
   ix3573 : nor03_2x port map ( Y=>nx3572, A0=>nx5129, A1=>nx9579, A2=>
      nx10535);
   gen_9_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_9_cmp_mReg_3, QB=>
      nx5129, D=>window_9_3, CLK=>start, R=>rst);
   ix3571 : nor03_2x port map ( Y=>nx3570, A0=>gen_9_cmp_mReg_3, A1=>nx10053, 
      A2=>nx10543);
   ix3607 : nand02 port map ( Y=>gen_9_cmp_BSCmp_op2_4, A0=>nx5133, A1=>
      nx5139);
   ix5134 : nor02_2x port map ( Y=>nx5133, A0=>nx3602, A1=>nx3598);
   ix3603 : nor03_2x port map ( Y=>nx3602, A0=>gen_9_cmp_mReg_3, A1=>nx9585, 
      A2=>nx10511);
   ix3599 : nor03_2x port map ( Y=>nx3598, A0=>nx5129, A1=>nx10517, A2=>
      nx10527);
   ix5140 : nor02_2x port map ( Y=>nx5139, A0=>nx3594, A1=>nx3592);
   ix3595 : nor03_2x port map ( Y=>nx3594, A0=>nx5143, A1=>nx9579, A2=>
      nx10535);
   gen_9_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_9_cmp_mReg_4, QB=>
      nx5143, D=>window_9_4, CLK=>start, R=>rst);
   ix3593 : nor03_2x port map ( Y=>nx3592, A0=>gen_9_cmp_mReg_4, A1=>nx10053, 
      A2=>nx10543);
   ix3629 : nand02 port map ( Y=>gen_9_cmp_BSCmp_op2_5, A0=>nx5147, A1=>
      nx5153);
   ix5148 : nor02_2x port map ( Y=>nx5147, A0=>nx3624, A1=>nx3620);
   ix3625 : nor03_2x port map ( Y=>nx3624, A0=>gen_9_cmp_mReg_4, A1=>nx9585, 
      A2=>nx10511);
   ix3621 : nor03_2x port map ( Y=>nx3620, A0=>nx5143, A1=>nx10517, A2=>
      nx10527);
   ix5154 : nor02_2x port map ( Y=>nx5153, A0=>nx3616, A1=>nx3614);
   ix3617 : nor03_2x port map ( Y=>nx3616, A0=>nx5156, A1=>nx9581, A2=>
      nx10535);
   gen_9_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_9_cmp_mReg_5, QB=>
      nx5156, D=>window_9_5, CLK=>start, R=>rst);
   ix3615 : nor03_2x port map ( Y=>nx3614, A0=>gen_9_cmp_mReg_5, A1=>nx10053, 
      A2=>nx10543);
   ix3651 : nand02 port map ( Y=>gen_9_cmp_BSCmp_op2_6, A0=>nx5163, A1=>
      nx5169);
   ix5164 : nor02_2x port map ( Y=>nx5163, A0=>nx3646, A1=>nx3642);
   ix3647 : nor03_2x port map ( Y=>nx3646, A0=>gen_9_cmp_mReg_5, A1=>nx9587, 
      A2=>nx10511);
   ix3643 : nor03_2x port map ( Y=>nx3642, A0=>nx5156, A1=>nx10517, A2=>
      nx10527);
   ix5170 : nor02_2x port map ( Y=>nx5169, A0=>nx3638, A1=>nx3636);
   ix3639 : nor03_2x port map ( Y=>nx3638, A0=>nx5173, A1=>nx9581, A2=>
      nx10535);
   gen_9_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_9_cmp_mReg_6, QB=>
      nx5173, D=>window_9_6, CLK=>start, R=>rst);
   ix3637 : nor03_2x port map ( Y=>nx3636, A0=>gen_9_cmp_mReg_6, A1=>nx10053, 
      A2=>nx10543);
   ix3673 : nand02 port map ( Y=>gen_9_cmp_BSCmp_op2_7, A0=>nx5177, A1=>
      nx5183);
   ix5178 : nor02_2x port map ( Y=>nx5177, A0=>nx3668, A1=>nx3664);
   ix3669 : nor03_2x port map ( Y=>nx3668, A0=>gen_9_cmp_mReg_6, A1=>nx9587, 
      A2=>nx10513);
   ix3665 : nor03_2x port map ( Y=>nx3664, A0=>nx5173, A1=>nx10519, A2=>
      nx10529);
   ix5184 : nor02_2x port map ( Y=>nx5183, A0=>nx3660, A1=>nx3658);
   ix3661 : nor03_2x port map ( Y=>nx3660, A0=>nx5187, A1=>nx9581, A2=>
      nx10537);
   gen_9_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_9_cmp_mReg_7, QB=>
      nx5187, D=>window_9_7, CLK=>start, R=>rst);
   ix3659 : nor03_2x port map ( Y=>nx3658, A0=>gen_9_cmp_mReg_7, A1=>nx10053, 
      A2=>nx10545);
   ix3695 : nand02 port map ( Y=>gen_9_cmp_BSCmp_op2_8, A0=>nx5191, A1=>
      nx5197);
   ix5192 : nor02_2x port map ( Y=>nx5191, A0=>nx3690, A1=>nx3686);
   ix3691 : nor03_2x port map ( Y=>nx3690, A0=>gen_9_cmp_mReg_7, A1=>nx9587, 
      A2=>nx10513);
   ix3687 : nor03_2x port map ( Y=>nx3686, A0=>nx5187, A1=>nx10519, A2=>
      nx10529);
   ix5198 : nor02_2x port map ( Y=>nx5197, A0=>nx3682, A1=>nx3680);
   ix3683 : nor03_2x port map ( Y=>nx3682, A0=>nx5200, A1=>nx9581, A2=>
      nx10537);
   gen_9_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_9_cmp_mReg_8, QB=>
      nx5200, D=>window_9_8, CLK=>start, R=>rst);
   ix3681 : nor03_2x port map ( Y=>nx3680, A0=>gen_9_cmp_mReg_8, A1=>nx10055, 
      A2=>nx10545);
   ix3717 : nand02 port map ( Y=>gen_9_cmp_BSCmp_op2_9, A0=>nx5207, A1=>
      nx5213);
   ix5208 : nor02_2x port map ( Y=>nx5207, A0=>nx3712, A1=>nx3708);
   ix3713 : nor03_2x port map ( Y=>nx3712, A0=>gen_9_cmp_mReg_8, A1=>nx9587, 
      A2=>nx10513);
   ix3709 : nor03_2x port map ( Y=>nx3708, A0=>nx5200, A1=>nx10519, A2=>
      nx10529);
   ix5214 : nor02_2x port map ( Y=>nx5213, A0=>nx3704, A1=>nx3702);
   ix3705 : nor03_2x port map ( Y=>nx3704, A0=>nx5217, A1=>nx9581, A2=>
      nx10537);
   gen_9_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_9_cmp_mReg_9, QB=>
      nx5217, D=>window_9_9, CLK=>start, R=>rst);
   ix3703 : nor03_2x port map ( Y=>nx3702, A0=>gen_9_cmp_mReg_9, A1=>nx10055, 
      A2=>nx10545);
   ix3739 : nand02 port map ( Y=>gen_9_cmp_BSCmp_op2_10, A0=>nx5221, A1=>
      nx5227);
   ix5222 : nor02_2x port map ( Y=>nx5221, A0=>nx3734, A1=>nx3730);
   ix3735 : nor03_2x port map ( Y=>nx3734, A0=>gen_9_cmp_mReg_9, A1=>nx9587, 
      A2=>nx10513);
   ix3731 : nor03_2x port map ( Y=>nx3730, A0=>nx5217, A1=>nx10519, A2=>
      nx10529);
   ix5228 : nor02_2x port map ( Y=>nx5227, A0=>nx3726, A1=>nx3724);
   ix3727 : nor03_2x port map ( Y=>nx3726, A0=>nx5231, A1=>nx9581, A2=>
      nx10537);
   gen_9_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_9_cmp_mReg_10, QB=>
      nx5231, D=>window_9_10, CLK=>start, R=>rst);
   ix3725 : nor03_2x port map ( Y=>nx3724, A0=>gen_9_cmp_mReg_10, A1=>
      nx10055, A2=>nx10545);
   ix3761 : nand02 port map ( Y=>gen_9_cmp_BSCmp_op2_11, A0=>nx5235, A1=>
      nx5241);
   ix5236 : nor02_2x port map ( Y=>nx5235, A0=>nx3756, A1=>nx3752);
   ix3757 : nor03_2x port map ( Y=>nx3756, A0=>gen_9_cmp_mReg_10, A1=>nx9587, 
      A2=>nx10513);
   ix3753 : nor03_2x port map ( Y=>nx3752, A0=>nx5231, A1=>nx10519, A2=>
      nx10529);
   ix5242 : nor02_2x port map ( Y=>nx5241, A0=>nx3748, A1=>nx3746);
   ix3749 : nor03_2x port map ( Y=>nx3748, A0=>nx5244, A1=>nx9581, A2=>
      nx10537);
   gen_9_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_9_cmp_mReg_11, QB=>
      nx5244, D=>window_9_11, CLK=>start, R=>rst);
   ix3747 : nor03_2x port map ( Y=>nx3746, A0=>gen_9_cmp_mReg_11, A1=>
      nx10055, A2=>nx10545);
   ix3783 : nand02 port map ( Y=>gen_9_cmp_BSCmp_op2_12, A0=>nx5251, A1=>
      nx5257);
   ix5252 : nor02_2x port map ( Y=>nx5251, A0=>nx3778, A1=>nx3774);
   ix3779 : nor03_2x port map ( Y=>nx3778, A0=>gen_9_cmp_mReg_11, A1=>nx9587, 
      A2=>nx10513);
   ix3775 : nor03_2x port map ( Y=>nx3774, A0=>nx5244, A1=>nx10519, A2=>
      nx10529);
   ix5258 : nor02_2x port map ( Y=>nx5257, A0=>nx3770, A1=>nx3768);
   ix3771 : nor03_2x port map ( Y=>nx3770, A0=>nx5261, A1=>nx9583, A2=>
      nx10537);
   gen_9_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_9_cmp_mReg_12, QB=>
      nx5261, D=>window_9_12, CLK=>start, R=>rst);
   ix3769 : nor03_2x port map ( Y=>nx3768, A0=>gen_9_cmp_mReg_12, A1=>
      nx10055, A2=>nx10545);
   ix3805 : nand02 port map ( Y=>gen_9_cmp_BSCmp_op2_13, A0=>nx5265, A1=>
      nx5271);
   ix5266 : nor02_2x port map ( Y=>nx5265, A0=>nx3800, A1=>nx3796);
   ix3801 : nor03_2x port map ( Y=>nx3800, A0=>gen_9_cmp_mReg_12, A1=>nx9589, 
      A2=>nx10515);
   ix3797 : nor03_2x port map ( Y=>nx3796, A0=>nx5261, A1=>nx10519, A2=>
      nx10531);
   ix5272 : nor02_2x port map ( Y=>nx5271, A0=>nx3792, A1=>nx3790);
   ix3793 : nor03_2x port map ( Y=>nx3792, A0=>nx5275, A1=>nx9583, A2=>
      nx10539);
   gen_9_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_9_cmp_mReg_13, QB=>
      nx5275, D=>window_9_13, CLK=>start, R=>rst);
   ix3791 : nor03_2x port map ( Y=>nx3790, A0=>gen_9_cmp_mReg_13, A1=>
      nx10055, A2=>nx10547);
   ix3827 : nand02 port map ( Y=>gen_9_cmp_BSCmp_op2_14, A0=>nx5279, A1=>
      nx5285);
   ix5280 : nor02_2x port map ( Y=>nx5279, A0=>nx3822, A1=>nx3818);
   ix3823 : nor03_2x port map ( Y=>nx3822, A0=>gen_9_cmp_mReg_13, A1=>nx9589, 
      A2=>nx10515);
   ix3819 : nor03_2x port map ( Y=>nx3818, A0=>nx5275, A1=>nx10521, A2=>
      nx10531);
   ix5286 : nor02_2x port map ( Y=>nx5285, A0=>nx3814, A1=>nx3812);
   ix3815 : nor03_2x port map ( Y=>nx3814, A0=>nx5288, A1=>nx9583, A2=>
      nx10539);
   gen_9_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_9_cmp_mReg_14, QB=>
      nx5288, D=>window_9_14, CLK=>start, R=>rst);
   ix3813 : nor03_2x port map ( Y=>nx3812, A0=>gen_9_cmp_mReg_14, A1=>
      nx10055, A2=>nx10547);
   ix3849 : nand02 port map ( Y=>gen_9_cmp_BSCmp_op2_15, A0=>nx5295, A1=>
      nx5301);
   ix5296 : nor02_2x port map ( Y=>nx5295, A0=>nx3844, A1=>nx3840);
   ix3845 : nor03_2x port map ( Y=>nx3844, A0=>gen_9_cmp_mReg_14, A1=>nx9589, 
      A2=>nx10515);
   ix3841 : nor03_2x port map ( Y=>nx3840, A0=>nx5288, A1=>nx10521, A2=>
      nx10531);
   ix5302 : nor02_2x port map ( Y=>nx5301, A0=>nx3836, A1=>nx3834);
   ix3837 : nor03_2x port map ( Y=>nx3836, A0=>nx5305, A1=>nx9583, A2=>
      nx10539);
   gen_9_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_9_cmp_mReg_15, QB=>
      nx5305, D=>window_9_15, CLK=>start, R=>rst);
   ix3835 : nor03_2x port map ( Y=>nx3834, A0=>gen_9_cmp_mReg_15, A1=>
      nx10057, A2=>nx10547);
   ix3859 : nand02 port map ( Y=>gen_9_cmp_BSCmp_op2_16, A0=>nx5309, A1=>
      nx5301);
   ix5310 : nor02_2x port map ( Y=>nx5309, A0=>nx3854, A1=>nx3850);
   ix3855 : nor03_2x port map ( Y=>nx3854, A0=>gen_9_cmp_mReg_15, A1=>nx9589, 
      A2=>nx10515);
   ix3851 : nor03_2x port map ( Y=>nx3850, A0=>nx5305, A1=>nx10521, A2=>
      nx10531);
   ix3927 : nand02 port map ( Y=>gen_10_cmp_BSCmp_op2_1, A0=>nx5317, A1=>
      nx5337);
   ix5318 : nor02_2x port map ( Y=>nx5317, A0=>nx3922, A1=>nx3918);
   ix3923 : nor03_2x port map ( Y=>nx3922, A0=>gen_10_cmp_mReg_0, A1=>nx9573, 
      A2=>nx10551);
   gen_10_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_10_cmp_mReg_0, QB=>
      nx5323, D=>window_10_0, CLK=>start, R=>rst);
   ix5328 : inv01 port map ( Y=>nx5327, A=>gen_10_cmp_pMux_0);
   ix3919 : nor03_2x port map ( Y=>nx3918, A0=>nx5323, A1=>nx10557, A2=>
      nx10567);
   ix5336 : inv02 port map ( Y=>nx5335, A=>gen_10_cmp_pMux_2);
   ix5338 : nor02_2x port map ( Y=>nx5337, A0=>nx3908, A1=>nx3906);
   ix3909 : nor03_2x port map ( Y=>nx3908, A0=>nx5341, A1=>nx9567, A2=>
      nx10575);
   gen_10_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_10_cmp_mReg_1, QB=>
      nx5341, D=>window_10_1, CLK=>start, R=>rst);
   ix3907 : nor03_2x port map ( Y=>nx3906, A0=>gen_10_cmp_mReg_1, A1=>
      nx10059, A2=>nx10583);
   ix3867 : nor03_2x port map ( Y=>nx3866, A0=>nx9573, A1=>nx5335, A2=>
      gen_10_cmp_pMux_0);
   ix3949 : nand02 port map ( Y=>gen_10_cmp_BSCmp_op2_2, A0=>nx5352, A1=>
      nx5357);
   ix5353 : nor02_2x port map ( Y=>nx5352, A0=>nx3944, A1=>nx3940);
   ix3945 : nor03_2x port map ( Y=>nx3944, A0=>gen_10_cmp_mReg_1, A1=>nx9573, 
      A2=>nx10551);
   ix3941 : nor03_2x port map ( Y=>nx3940, A0=>nx5341, A1=>nx10557, A2=>
      nx10567);
   ix5358 : nor02_2x port map ( Y=>nx5357, A0=>nx3936, A1=>nx3934);
   ix3937 : nor03_2x port map ( Y=>nx3936, A0=>nx5361, A1=>nx9567, A2=>
      nx10575);
   gen_10_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_10_cmp_mReg_2, QB=>
      nx5361, D=>window_10_2, CLK=>start, R=>rst);
   ix3935 : nor03_2x port map ( Y=>nx3934, A0=>gen_10_cmp_mReg_2, A1=>
      nx10059, A2=>nx10583);
   ix3971 : nand02 port map ( Y=>gen_10_cmp_BSCmp_op2_3, A0=>nx5367, A1=>
      nx5373);
   ix5368 : nor02_2x port map ( Y=>nx5367, A0=>nx3966, A1=>nx3962);
   ix3967 : nor03_2x port map ( Y=>nx3966, A0=>gen_10_cmp_mReg_2, A1=>nx9573, 
      A2=>nx10551);
   ix3963 : nor03_2x port map ( Y=>nx3962, A0=>nx5361, A1=>nx10557, A2=>
      nx10567);
   ix5374 : nor02_2x port map ( Y=>nx5373, A0=>nx3958, A1=>nx3956);
   ix3959 : nor03_2x port map ( Y=>nx3958, A0=>nx5376, A1=>nx9567, A2=>
      nx10575);
   gen_10_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_10_cmp_mReg_3, QB=>
      nx5376, D=>window_10_3, CLK=>start, R=>rst);
   ix3957 : nor03_2x port map ( Y=>nx3956, A0=>gen_10_cmp_mReg_3, A1=>
      nx10059, A2=>nx10583);
   ix3993 : nand02 port map ( Y=>gen_10_cmp_BSCmp_op2_4, A0=>nx5383, A1=>
      nx5389);
   ix5384 : nor02_2x port map ( Y=>nx5383, A0=>nx3988, A1=>nx3984);
   ix3989 : nor03_2x port map ( Y=>nx3988, A0=>gen_10_cmp_mReg_3, A1=>nx9573, 
      A2=>nx10551);
   ix3985 : nor03_2x port map ( Y=>nx3984, A0=>nx5376, A1=>nx10557, A2=>
      nx10567);
   ix5390 : nor02_2x port map ( Y=>nx5389, A0=>nx3980, A1=>nx3978);
   ix3981 : nor03_2x port map ( Y=>nx3980, A0=>nx5393, A1=>nx9567, A2=>
      nx10575);
   gen_10_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_10_cmp_mReg_4, QB=>
      nx5393, D=>window_10_4, CLK=>start, R=>rst);
   ix3979 : nor03_2x port map ( Y=>nx3978, A0=>gen_10_cmp_mReg_4, A1=>
      nx10059, A2=>nx10583);
   ix4015 : nand02 port map ( Y=>gen_10_cmp_BSCmp_op2_5, A0=>nx5399, A1=>
      nx5405);
   ix5400 : nor02_2x port map ( Y=>nx5399, A0=>nx4010, A1=>nx4006);
   ix4011 : nor03_2x port map ( Y=>nx4010, A0=>gen_10_cmp_mReg_4, A1=>nx9573, 
      A2=>nx10551);
   ix4007 : nor03_2x port map ( Y=>nx4006, A0=>nx5393, A1=>nx10557, A2=>
      nx10567);
   ix5406 : nor02_2x port map ( Y=>nx5405, A0=>nx4002, A1=>nx4000);
   ix4003 : nor03_2x port map ( Y=>nx4002, A0=>nx5409, A1=>nx9569, A2=>
      nx10575);
   gen_10_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_10_cmp_mReg_5, QB=>
      nx5409, D=>window_10_5, CLK=>start, R=>rst);
   ix4001 : nor03_2x port map ( Y=>nx4000, A0=>gen_10_cmp_mReg_5, A1=>
      nx10059, A2=>nx10583);
   ix4037 : nand02 port map ( Y=>gen_10_cmp_BSCmp_op2_6, A0=>nx5414, A1=>
      nx5418);
   ix5415 : nor02_2x port map ( Y=>nx5414, A0=>nx4032, A1=>nx4028);
   ix4033 : nor03_2x port map ( Y=>nx4032, A0=>gen_10_cmp_mReg_5, A1=>nx9575, 
      A2=>nx10551);
   ix4029 : nor03_2x port map ( Y=>nx4028, A0=>nx5409, A1=>nx10557, A2=>
      nx10567);
   ix5419 : nor02_2x port map ( Y=>nx5418, A0=>nx4024, A1=>nx4022);
   ix4025 : nor03_2x port map ( Y=>nx4024, A0=>nx5421, A1=>nx9569, A2=>
      nx10575);
   gen_10_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_10_cmp_mReg_6, QB=>
      nx5421, D=>window_10_6, CLK=>start, R=>rst);
   ix4023 : nor03_2x port map ( Y=>nx4022, A0=>gen_10_cmp_mReg_6, A1=>
      nx10059, A2=>nx10583);
   ix4059 : nand02 port map ( Y=>gen_10_cmp_BSCmp_op2_7, A0=>nx5427, A1=>
      nx5433);
   ix5428 : nor02_2x port map ( Y=>nx5427, A0=>nx4054, A1=>nx4050);
   ix4055 : nor03_2x port map ( Y=>nx4054, A0=>gen_10_cmp_mReg_6, A1=>nx9575, 
      A2=>nx10553);
   ix4051 : nor03_2x port map ( Y=>nx4050, A0=>nx5421, A1=>nx10559, A2=>
      nx10569);
   ix5434 : nor02_2x port map ( Y=>nx5433, A0=>nx4046, A1=>nx4044);
   ix4047 : nor03_2x port map ( Y=>nx4046, A0=>nx5437, A1=>nx9569, A2=>
      nx10577);
   gen_10_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_10_cmp_mReg_7, QB=>
      nx5437, D=>window_10_7, CLK=>start, R=>rst);
   ix4045 : nor03_2x port map ( Y=>nx4044, A0=>gen_10_cmp_mReg_7, A1=>
      nx10059, A2=>nx10585);
   ix4081 : nand02 port map ( Y=>gen_10_cmp_BSCmp_op2_8, A0=>nx5443, A1=>
      nx5447);
   ix5444 : nor02_2x port map ( Y=>nx5443, A0=>nx4076, A1=>nx4072);
   ix4077 : nor03_2x port map ( Y=>nx4076, A0=>gen_10_cmp_mReg_7, A1=>nx9575, 
      A2=>nx10553);
   ix4073 : nor03_2x port map ( Y=>nx4072, A0=>nx5437, A1=>nx10559, A2=>
      nx10569);
   ix5448 : nor02_2x port map ( Y=>nx5447, A0=>nx4068, A1=>nx4066);
   ix4069 : nor03_2x port map ( Y=>nx4068, A0=>nx5451, A1=>nx9569, A2=>
      nx10577);
   gen_10_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_10_cmp_mReg_8, QB=>
      nx5451, D=>window_10_8, CLK=>start, R=>rst);
   ix4067 : nor03_2x port map ( Y=>nx4066, A0=>gen_10_cmp_mReg_8, A1=>
      nx10061, A2=>nx10585);
   ix4103 : nand02 port map ( Y=>gen_10_cmp_BSCmp_op2_9, A0=>nx5457, A1=>
      nx5463);
   ix5458 : nor02_2x port map ( Y=>nx5457, A0=>nx4098, A1=>nx4094);
   ix4099 : nor03_2x port map ( Y=>nx4098, A0=>gen_10_cmp_mReg_8, A1=>nx9575, 
      A2=>nx10553);
   ix4095 : nor03_2x port map ( Y=>nx4094, A0=>nx5451, A1=>nx10559, A2=>
      nx10569);
   ix5464 : nor02_2x port map ( Y=>nx5463, A0=>nx4090, A1=>nx4088);
   ix4091 : nor03_2x port map ( Y=>nx4090, A0=>nx5467, A1=>nx9569, A2=>
      nx10577);
   gen_10_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_10_cmp_mReg_9, QB=>
      nx5467, D=>window_10_9, CLK=>start, R=>rst);
   ix4089 : nor03_2x port map ( Y=>nx4088, A0=>gen_10_cmp_mReg_9, A1=>
      nx10061, A2=>nx10585);
   ix4125 : nand02 port map ( Y=>gen_10_cmp_BSCmp_op2_10, A0=>nx5473, A1=>
      nx5477);
   ix5474 : nor02_2x port map ( Y=>nx5473, A0=>nx4120, A1=>nx4116);
   ix4121 : nor03_2x port map ( Y=>nx4120, A0=>gen_10_cmp_mReg_9, A1=>nx9575, 
      A2=>nx10553);
   ix4117 : nor03_2x port map ( Y=>nx4116, A0=>nx5467, A1=>nx10559, A2=>
      nx10569);
   ix5478 : nor02_2x port map ( Y=>nx5477, A0=>nx4112, A1=>nx4110);
   ix4113 : nor03_2x port map ( Y=>nx4112, A0=>nx5481, A1=>nx9569, A2=>
      nx10577);
   gen_10_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_10_cmp_mReg_10, QB=>
      nx5481, D=>window_10_10, CLK=>start, R=>rst);
   ix4111 : nor03_2x port map ( Y=>nx4110, A0=>gen_10_cmp_mReg_10, A1=>
      nx10061, A2=>nx10585);
   ix4147 : nand02 port map ( Y=>gen_10_cmp_BSCmp_op2_11, A0=>nx5487, A1=>
      nx5493);
   ix5488 : nor02_2x port map ( Y=>nx5487, A0=>nx4142, A1=>nx4138);
   ix4143 : nor03_2x port map ( Y=>nx4142, A0=>gen_10_cmp_mReg_10, A1=>
      nx9575, A2=>nx10553);
   ix4139 : nor03_2x port map ( Y=>nx4138, A0=>nx5481, A1=>nx10559, A2=>
      nx10569);
   ix5494 : nor02_2x port map ( Y=>nx5493, A0=>nx4134, A1=>nx4132);
   ix4135 : nor03_2x port map ( Y=>nx4134, A0=>nx5496, A1=>nx9569, A2=>
      nx10577);
   gen_10_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_10_cmp_mReg_11, QB=>
      nx5496, D=>window_10_11, CLK=>start, R=>rst);
   ix4133 : nor03_2x port map ( Y=>nx4132, A0=>gen_10_cmp_mReg_11, A1=>
      nx10061, A2=>nx10585);
   ix4169 : nand02 port map ( Y=>gen_10_cmp_BSCmp_op2_12, A0=>nx5501, A1=>
      nx5507);
   ix5502 : nor02_2x port map ( Y=>nx5501, A0=>nx4164, A1=>nx4160);
   ix4165 : nor03_2x port map ( Y=>nx4164, A0=>gen_10_cmp_mReg_11, A1=>
      nx9575, A2=>nx10553);
   ix4161 : nor03_2x port map ( Y=>nx4160, A0=>nx5496, A1=>nx10559, A2=>
      nx10569);
   ix5508 : nor02_2x port map ( Y=>nx5507, A0=>nx4156, A1=>nx4154);
   ix4157 : nor03_2x port map ( Y=>nx4156, A0=>nx5511, A1=>nx9571, A2=>
      nx10577);
   gen_10_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_10_cmp_mReg_12, QB=>
      nx5511, D=>window_10_12, CLK=>start, R=>rst);
   ix4155 : nor03_2x port map ( Y=>nx4154, A0=>gen_10_cmp_mReg_12, A1=>
      nx10061, A2=>nx10585);
   ix4191 : nand02 port map ( Y=>gen_10_cmp_BSCmp_op2_13, A0=>nx5517, A1=>
      nx5521);
   ix5518 : nor02_2x port map ( Y=>nx5517, A0=>nx4186, A1=>nx4182);
   ix4187 : nor03_2x port map ( Y=>nx4186, A0=>gen_10_cmp_mReg_12, A1=>
      nx9577, A2=>nx10555);
   ix4183 : nor03_2x port map ( Y=>nx4182, A0=>nx5511, A1=>nx10559, A2=>
      nx10571);
   ix5522 : nor02_2x port map ( Y=>nx5521, A0=>nx4178, A1=>nx4176);
   ix4179 : nor03_2x port map ( Y=>nx4178, A0=>nx5525, A1=>nx9571, A2=>
      nx10579);
   gen_10_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_10_cmp_mReg_13, QB=>
      nx5525, D=>window_10_13, CLK=>start, R=>rst);
   ix4177 : nor03_2x port map ( Y=>nx4176, A0=>gen_10_cmp_mReg_13, A1=>
      nx10061, A2=>nx10587);
   ix4213 : nand02 port map ( Y=>gen_10_cmp_BSCmp_op2_14, A0=>nx5531, A1=>
      nx5537);
   ix5532 : nor02_2x port map ( Y=>nx5531, A0=>nx4208, A1=>nx4204);
   ix4209 : nor03_2x port map ( Y=>nx4208, A0=>gen_10_cmp_mReg_13, A1=>
      nx9577, A2=>nx10555);
   ix4205 : nor03_2x port map ( Y=>nx4204, A0=>nx5525, A1=>nx10561, A2=>
      nx10571);
   ix5538 : nor02_2x port map ( Y=>nx5537, A0=>nx4200, A1=>nx4198);
   ix4201 : nor03_2x port map ( Y=>nx4200, A0=>nx5540, A1=>nx9571, A2=>
      nx10579);
   gen_10_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_10_cmp_mReg_14, QB=>
      nx5540, D=>window_10_14, CLK=>start, R=>rst);
   ix4199 : nor03_2x port map ( Y=>nx4198, A0=>gen_10_cmp_mReg_14, A1=>
      nx10061, A2=>nx10587);
   ix4235 : nand02 port map ( Y=>gen_10_cmp_BSCmp_op2_15, A0=>nx5545, A1=>
      nx5551);
   ix5546 : nor02_2x port map ( Y=>nx5545, A0=>nx4230, A1=>nx4226);
   ix4231 : nor03_2x port map ( Y=>nx4230, A0=>gen_10_cmp_mReg_14, A1=>
      nx9577, A2=>nx10555);
   ix4227 : nor03_2x port map ( Y=>nx4226, A0=>nx5540, A1=>nx10561, A2=>
      nx10571);
   ix5552 : nor02_2x port map ( Y=>nx5551, A0=>nx4222, A1=>nx4220);
   ix4223 : nor03_2x port map ( Y=>nx4222, A0=>nx5555, A1=>nx9571, A2=>
      nx10579);
   gen_10_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_10_cmp_mReg_15, QB=>
      nx5555, D=>window_10_15, CLK=>start, R=>rst);
   ix4221 : nor03_2x port map ( Y=>nx4220, A0=>gen_10_cmp_mReg_15, A1=>
      nx10063, A2=>nx10587);
   ix4245 : nand02 port map ( Y=>gen_10_cmp_BSCmp_op2_16, A0=>nx5561, A1=>
      nx5551);
   ix5562 : nor02_2x port map ( Y=>nx5561, A0=>nx4240, A1=>nx4236);
   ix4241 : nor03_2x port map ( Y=>nx4240, A0=>gen_10_cmp_mReg_15, A1=>
      nx9577, A2=>nx10555);
   ix4237 : nor03_2x port map ( Y=>nx4236, A0=>nx5555, A1=>nx10561, A2=>
      nx10571);
   ix4313 : nand02 port map ( Y=>gen_11_cmp_BSCmp_op2_1, A0=>nx5567, A1=>
      nx5587);
   ix5568 : nor02_2x port map ( Y=>nx5567, A0=>nx4308, A1=>nx4304);
   ix4309 : nor03_2x port map ( Y=>nx4308, A0=>gen_11_cmp_mReg_0, A1=>nx9561, 
      A2=>nx10591);
   gen_11_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_11_cmp_mReg_0, QB=>
      nx5573, D=>window_11_0, CLK=>start, R=>rst);
   ix5578 : inv01 port map ( Y=>nx5577, A=>gen_11_cmp_pMux_0);
   ix4305 : nor03_2x port map ( Y=>nx4304, A0=>nx5573, A1=>nx10597, A2=>
      nx10607);
   ix5586 : inv02 port map ( Y=>nx5585, A=>gen_11_cmp_pMux_2);
   ix5588 : nor02_2x port map ( Y=>nx5587, A0=>nx4294, A1=>nx4292);
   ix4295 : nor03_2x port map ( Y=>nx4294, A0=>nx5591, A1=>nx9555, A2=>
      nx10615);
   gen_11_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_11_cmp_mReg_1, QB=>
      nx5591, D=>window_11_1, CLK=>start, R=>rst);
   ix4293 : nor03_2x port map ( Y=>nx4292, A0=>gen_11_cmp_mReg_1, A1=>
      nx10065, A2=>nx10623);
   ix4253 : nor03_2x port map ( Y=>nx4252, A0=>nx9561, A1=>nx5585, A2=>
      gen_11_cmp_pMux_0);
   ix4335 : nand02 port map ( Y=>gen_11_cmp_BSCmp_op2_2, A0=>nx5603, A1=>
      nx5607);
   ix5604 : nor02_2x port map ( Y=>nx5603, A0=>nx4330, A1=>nx4326);
   ix4331 : nor03_2x port map ( Y=>nx4330, A0=>gen_11_cmp_mReg_1, A1=>nx9561, 
      A2=>nx10591);
   ix4327 : nor03_2x port map ( Y=>nx4326, A0=>nx5591, A1=>nx10597, A2=>
      nx10607);
   ix5608 : nor02_2x port map ( Y=>nx5607, A0=>nx4322, A1=>nx4320);
   ix4323 : nor03_2x port map ( Y=>nx4322, A0=>nx5611, A1=>nx9555, A2=>
      nx10615);
   gen_11_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_11_cmp_mReg_2, QB=>
      nx5611, D=>window_11_2, CLK=>start, R=>rst);
   ix4321 : nor03_2x port map ( Y=>nx4320, A0=>gen_11_cmp_mReg_2, A1=>
      nx10065, A2=>nx10623);
   ix4357 : nand02 port map ( Y=>gen_11_cmp_BSCmp_op2_3, A0=>nx5617, A1=>
      nx5621);
   ix5618 : nor02_2x port map ( Y=>nx5617, A0=>nx4352, A1=>nx4348);
   ix4353 : nor03_2x port map ( Y=>nx4352, A0=>gen_11_cmp_mReg_2, A1=>nx9561, 
      A2=>nx10591);
   ix4349 : nor03_2x port map ( Y=>nx4348, A0=>nx5611, A1=>nx10597, A2=>
      nx10607);
   ix5622 : nor02_2x port map ( Y=>nx5621, A0=>nx4344, A1=>nx4342);
   ix4345 : nor03_2x port map ( Y=>nx4344, A0=>nx5625, A1=>nx9555, A2=>
      nx10615);
   gen_11_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_11_cmp_mReg_3, QB=>
      nx5625, D=>window_11_3, CLK=>start, R=>rst);
   ix4343 : nor03_2x port map ( Y=>nx4342, A0=>gen_11_cmp_mReg_3, A1=>
      nx10065, A2=>nx10623);
   ix4379 : nand02 port map ( Y=>gen_11_cmp_BSCmp_op2_4, A0=>nx5629, A1=>
      nx5635);
   ix5630 : nor02_2x port map ( Y=>nx5629, A0=>nx4374, A1=>nx4370);
   ix4375 : nor03_2x port map ( Y=>nx4374, A0=>gen_11_cmp_mReg_3, A1=>nx9561, 
      A2=>nx10591);
   ix4371 : nor03_2x port map ( Y=>nx4370, A0=>nx5625, A1=>nx10597, A2=>
      nx10607);
   ix5636 : nor02_2x port map ( Y=>nx5635, A0=>nx4366, A1=>nx4364);
   ix4367 : nor03_2x port map ( Y=>nx4366, A0=>nx5639, A1=>nx9555, A2=>
      nx10615);
   gen_11_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_11_cmp_mReg_4, QB=>
      nx5639, D=>window_11_4, CLK=>start, R=>rst);
   ix4365 : nor03_2x port map ( Y=>nx4364, A0=>gen_11_cmp_mReg_4, A1=>
      nx10065, A2=>nx10623);
   ix4401 : nand02 port map ( Y=>gen_11_cmp_BSCmp_op2_5, A0=>nx5643, A1=>
      nx5649);
   ix5644 : nor02_2x port map ( Y=>nx5643, A0=>nx4396, A1=>nx4392);
   ix4397 : nor03_2x port map ( Y=>nx4396, A0=>gen_11_cmp_mReg_4, A1=>nx9561, 
      A2=>nx10591);
   ix4393 : nor03_2x port map ( Y=>nx4392, A0=>nx5639, A1=>nx10597, A2=>
      nx10607);
   ix5650 : nor02_2x port map ( Y=>nx5649, A0=>nx4388, A1=>nx4386);
   ix4389 : nor03_2x port map ( Y=>nx4388, A0=>nx5652, A1=>nx9557, A2=>
      nx10615);
   gen_11_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_11_cmp_mReg_5, QB=>
      nx5652, D=>window_11_5, CLK=>start, R=>rst);
   ix4387 : nor03_2x port map ( Y=>nx4386, A0=>gen_11_cmp_mReg_5, A1=>
      nx10065, A2=>nx10623);
   ix4423 : nand02 port map ( Y=>gen_11_cmp_BSCmp_op2_6, A0=>nx5659, A1=>
      nx5665);
   ix5660 : nor02_2x port map ( Y=>nx5659, A0=>nx4418, A1=>nx4414);
   ix4419 : nor03_2x port map ( Y=>nx4418, A0=>gen_11_cmp_mReg_5, A1=>nx9563, 
      A2=>nx10591);
   ix4415 : nor03_2x port map ( Y=>nx4414, A0=>nx5652, A1=>nx10597, A2=>
      nx10607);
   ix5666 : nor02_2x port map ( Y=>nx5665, A0=>nx4410, A1=>nx4408);
   ix4411 : nor03_2x port map ( Y=>nx4410, A0=>nx5669, A1=>nx9557, A2=>
      nx10615);
   gen_11_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_11_cmp_mReg_6, QB=>
      nx5669, D=>window_11_6, CLK=>start, R=>rst);
   ix4409 : nor03_2x port map ( Y=>nx4408, A0=>gen_11_cmp_mReg_6, A1=>
      nx10065, A2=>nx10623);
   ix4445 : nand02 port map ( Y=>gen_11_cmp_BSCmp_op2_7, A0=>nx5673, A1=>
      nx5679);
   ix5674 : nor02_2x port map ( Y=>nx5673, A0=>nx4440, A1=>nx4436);
   ix4441 : nor03_2x port map ( Y=>nx4440, A0=>gen_11_cmp_mReg_6, A1=>nx9563, 
      A2=>nx10593);
   ix4437 : nor03_2x port map ( Y=>nx4436, A0=>nx5669, A1=>nx10599, A2=>
      nx10609);
   ix5680 : nor02_2x port map ( Y=>nx5679, A0=>nx4432, A1=>nx4430);
   ix4433 : nor03_2x port map ( Y=>nx4432, A0=>nx5683, A1=>nx9557, A2=>
      nx10617);
   gen_11_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_11_cmp_mReg_7, QB=>
      nx5683, D=>window_11_7, CLK=>start, R=>rst);
   ix4431 : nor03_2x port map ( Y=>nx4430, A0=>gen_11_cmp_mReg_7, A1=>
      nx10065, A2=>nx10625);
   ix4467 : nand02 port map ( Y=>gen_11_cmp_BSCmp_op2_8, A0=>nx5687, A1=>
      nx5693);
   ix5688 : nor02_2x port map ( Y=>nx5687, A0=>nx4462, A1=>nx4458);
   ix4463 : nor03_2x port map ( Y=>nx4462, A0=>gen_11_cmp_mReg_7, A1=>nx9563, 
      A2=>nx10593);
   ix4459 : nor03_2x port map ( Y=>nx4458, A0=>nx5683, A1=>nx10599, A2=>
      nx10609);
   ix5694 : nor02_2x port map ( Y=>nx5693, A0=>nx4454, A1=>nx4452);
   ix4455 : nor03_2x port map ( Y=>nx4454, A0=>nx5696, A1=>nx9557, A2=>
      nx10617);
   gen_11_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_11_cmp_mReg_8, QB=>
      nx5696, D=>window_11_8, CLK=>start, R=>rst);
   ix4453 : nor03_2x port map ( Y=>nx4452, A0=>gen_11_cmp_mReg_8, A1=>
      nx10067, A2=>nx10625);
   ix4489 : nand02 port map ( Y=>gen_11_cmp_BSCmp_op2_9, A0=>nx5703, A1=>
      nx5709);
   ix5704 : nor02_2x port map ( Y=>nx5703, A0=>nx4484, A1=>nx4480);
   ix4485 : nor03_2x port map ( Y=>nx4484, A0=>gen_11_cmp_mReg_8, A1=>nx9563, 
      A2=>nx10593);
   ix4481 : nor03_2x port map ( Y=>nx4480, A0=>nx5696, A1=>nx10599, A2=>
      nx10609);
   ix5710 : nor02_2x port map ( Y=>nx5709, A0=>nx4476, A1=>nx4474);
   ix4477 : nor03_2x port map ( Y=>nx4476, A0=>nx5713, A1=>nx9557, A2=>
      nx10617);
   gen_11_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_11_cmp_mReg_9, QB=>
      nx5713, D=>window_11_9, CLK=>start, R=>rst);
   ix4475 : nor03_2x port map ( Y=>nx4474, A0=>gen_11_cmp_mReg_9, A1=>
      nx10067, A2=>nx10625);
   ix4511 : nand02 port map ( Y=>gen_11_cmp_BSCmp_op2_10, A0=>nx5717, A1=>
      nx5723);
   ix5718 : nor02_2x port map ( Y=>nx5717, A0=>nx4506, A1=>nx4502);
   ix4507 : nor03_2x port map ( Y=>nx4506, A0=>gen_11_cmp_mReg_9, A1=>nx9563, 
      A2=>nx10593);
   ix4503 : nor03_2x port map ( Y=>nx4502, A0=>nx5713, A1=>nx10599, A2=>
      nx10609);
   ix5724 : nor02_2x port map ( Y=>nx5723, A0=>nx4498, A1=>nx4496);
   ix4499 : nor03_2x port map ( Y=>nx4498, A0=>nx5727, A1=>nx9557, A2=>
      nx10617);
   gen_11_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_11_cmp_mReg_10, QB=>
      nx5727, D=>window_11_10, CLK=>start, R=>rst);
   ix4497 : nor03_2x port map ( Y=>nx4496, A0=>gen_11_cmp_mReg_10, A1=>
      nx10067, A2=>nx10625);
   ix4533 : nand02 port map ( Y=>gen_11_cmp_BSCmp_op2_11, A0=>nx5731, A1=>
      nx5737);
   ix5732 : nor02_2x port map ( Y=>nx5731, A0=>nx4528, A1=>nx4524);
   ix4529 : nor03_2x port map ( Y=>nx4528, A0=>gen_11_cmp_mReg_10, A1=>
      nx9563, A2=>nx10593);
   ix4525 : nor03_2x port map ( Y=>nx4524, A0=>nx5727, A1=>nx10599, A2=>
      nx10609);
   ix5738 : nor02_2x port map ( Y=>nx5737, A0=>nx4520, A1=>nx4518);
   ix4521 : nor03_2x port map ( Y=>nx4520, A0=>nx5740, A1=>nx9557, A2=>
      nx10617);
   gen_11_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_11_cmp_mReg_11, QB=>
      nx5740, D=>window_11_11, CLK=>start, R=>rst);
   ix4519 : nor03_2x port map ( Y=>nx4518, A0=>gen_11_cmp_mReg_11, A1=>
      nx10067, A2=>nx10625);
   ix4555 : nand02 port map ( Y=>gen_11_cmp_BSCmp_op2_12, A0=>nx5747, A1=>
      nx5753);
   ix5748 : nor02_2x port map ( Y=>nx5747, A0=>nx4550, A1=>nx4546);
   ix4551 : nor03_2x port map ( Y=>nx4550, A0=>gen_11_cmp_mReg_11, A1=>
      nx9563, A2=>nx10593);
   ix4547 : nor03_2x port map ( Y=>nx4546, A0=>nx5740, A1=>nx10599, A2=>
      nx10609);
   ix5754 : nor02_2x port map ( Y=>nx5753, A0=>nx4542, A1=>nx4540);
   ix4543 : nor03_2x port map ( Y=>nx4542, A0=>nx5757, A1=>nx9559, A2=>
      nx10617);
   gen_11_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_11_cmp_mReg_12, QB=>
      nx5757, D=>window_11_12, CLK=>start, R=>rst);
   ix4541 : nor03_2x port map ( Y=>nx4540, A0=>gen_11_cmp_mReg_12, A1=>
      nx10067, A2=>nx10625);
   ix4577 : nand02 port map ( Y=>gen_11_cmp_BSCmp_op2_13, A0=>nx5761, A1=>
      nx5767);
   ix5762 : nor02_2x port map ( Y=>nx5761, A0=>nx4572, A1=>nx4568);
   ix4573 : nor03_2x port map ( Y=>nx4572, A0=>gen_11_cmp_mReg_12, A1=>
      nx9565, A2=>nx10595);
   ix4569 : nor03_2x port map ( Y=>nx4568, A0=>nx5757, A1=>nx10599, A2=>
      nx10611);
   ix5768 : nor02_2x port map ( Y=>nx5767, A0=>nx4564, A1=>nx4562);
   ix4565 : nor03_2x port map ( Y=>nx4564, A0=>nx5771, A1=>nx9559, A2=>
      nx10619);
   gen_11_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_11_cmp_mReg_13, QB=>
      nx5771, D=>window_11_13, CLK=>start, R=>rst);
   ix4563 : nor03_2x port map ( Y=>nx4562, A0=>gen_11_cmp_mReg_13, A1=>
      nx10067, A2=>nx10627);
   ix4599 : nand02 port map ( Y=>gen_11_cmp_BSCmp_op2_14, A0=>nx5775, A1=>
      nx5781);
   ix5776 : nor02_2x port map ( Y=>nx5775, A0=>nx4594, A1=>nx4590);
   ix4595 : nor03_2x port map ( Y=>nx4594, A0=>gen_11_cmp_mReg_13, A1=>
      nx9565, A2=>nx10595);
   ix4591 : nor03_2x port map ( Y=>nx4590, A0=>nx5771, A1=>nx10601, A2=>
      nx10611);
   ix5782 : nor02_2x port map ( Y=>nx5781, A0=>nx4586, A1=>nx4584);
   ix4587 : nor03_2x port map ( Y=>nx4586, A0=>nx5785, A1=>nx9559, A2=>
      nx10619);
   gen_11_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_11_cmp_mReg_14, QB=>
      nx5785, D=>window_11_14, CLK=>start, R=>rst);
   ix4585 : nor03_2x port map ( Y=>nx4584, A0=>gen_11_cmp_mReg_14, A1=>
      nx10067, A2=>nx10627);
   ix4621 : nand02 port map ( Y=>gen_11_cmp_BSCmp_op2_15, A0=>nx5791, A1=>
      nx5797);
   ix5792 : nor02_2x port map ( Y=>nx5791, A0=>nx4616, A1=>nx4612);
   ix4617 : nor03_2x port map ( Y=>nx4616, A0=>gen_11_cmp_mReg_14, A1=>
      nx9565, A2=>nx10595);
   ix4613 : nor03_2x port map ( Y=>nx4612, A0=>nx5785, A1=>nx10601, A2=>
      nx10611);
   ix5798 : nor02_2x port map ( Y=>nx5797, A0=>nx4608, A1=>nx4606);
   ix4609 : nor03_2x port map ( Y=>nx4608, A0=>nx5800, A1=>nx9559, A2=>
      nx10619);
   gen_11_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_11_cmp_mReg_15, QB=>
      nx5800, D=>window_11_15, CLK=>start, R=>rst);
   ix4607 : nor03_2x port map ( Y=>nx4606, A0=>gen_11_cmp_mReg_15, A1=>
      nx10069, A2=>nx10627);
   ix4631 : nand02 port map ( Y=>gen_11_cmp_BSCmp_op2_16, A0=>nx5804, A1=>
      nx5797);
   ix5805 : nor02_2x port map ( Y=>nx5804, A0=>nx4626, A1=>nx4622);
   ix4627 : nor03_2x port map ( Y=>nx4626, A0=>gen_11_cmp_mReg_15, A1=>
      nx9565, A2=>nx10595);
   ix4623 : nor03_2x port map ( Y=>nx4622, A0=>nx5800, A1=>nx10601, A2=>
      nx10611);
   ix4699 : nand02 port map ( Y=>gen_12_cmp_BSCmp_op2_1, A0=>nx5811, A1=>
      nx5831);
   ix5812 : nor02_2x port map ( Y=>nx5811, A0=>nx4694, A1=>nx4690);
   ix4695 : nor03_2x port map ( Y=>nx4694, A0=>gen_12_cmp_mReg_0, A1=>nx9549, 
      A2=>nx10631);
   gen_12_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_12_cmp_mReg_0, QB=>
      nx5817, D=>window_12_0, CLK=>start, R=>rst);
   ix5822 : inv01 port map ( Y=>nx5821, A=>gen_12_cmp_pMux_0);
   ix4691 : nor03_2x port map ( Y=>nx4690, A0=>nx5817, A1=>nx10637, A2=>
      nx10647);
   ix5830 : inv02 port map ( Y=>nx5829, A=>gen_12_cmp_pMux_2);
   ix5832 : nor02_2x port map ( Y=>nx5831, A0=>nx4680, A1=>nx4678);
   ix4681 : nor03_2x port map ( Y=>nx4680, A0=>nx5834, A1=>nx9543, A2=>
      nx10655);
   gen_12_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_12_cmp_mReg_1, QB=>
      nx5834, D=>window_12_1, CLK=>start, R=>rst);
   ix4679 : nor03_2x port map ( Y=>nx4678, A0=>gen_12_cmp_mReg_1, A1=>
      nx10071, A2=>nx10663);
   ix4639 : nor03_2x port map ( Y=>nx4638, A0=>nx9549, A1=>nx5829, A2=>
      gen_12_cmp_pMux_0);
   ix4721 : nand02 port map ( Y=>gen_12_cmp_BSCmp_op2_2, A0=>nx5847, A1=>
      nx5853);
   ix5848 : nor02_2x port map ( Y=>nx5847, A0=>nx4716, A1=>nx4712);
   ix4717 : nor03_2x port map ( Y=>nx4716, A0=>gen_12_cmp_mReg_1, A1=>nx9549, 
      A2=>nx10631);
   ix4713 : nor03_2x port map ( Y=>nx4712, A0=>nx5834, A1=>nx10637, A2=>
      nx10647);
   ix5854 : nor02_2x port map ( Y=>nx5853, A0=>nx4708, A1=>nx4706);
   ix4709 : nor03_2x port map ( Y=>nx4708, A0=>nx5857, A1=>nx9543, A2=>
      nx10655);
   gen_12_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_12_cmp_mReg_2, QB=>
      nx5857, D=>window_12_2, CLK=>start, R=>rst);
   ix4707 : nor03_2x port map ( Y=>nx4706, A0=>gen_12_cmp_mReg_2, A1=>
      nx10071, A2=>nx10663);
   ix4743 : nand02 port map ( Y=>gen_12_cmp_BSCmp_op2_3, A0=>nx5861, A1=>
      nx5867);
   ix5862 : nor02_2x port map ( Y=>nx5861, A0=>nx4738, A1=>nx4734);
   ix4739 : nor03_2x port map ( Y=>nx4738, A0=>gen_12_cmp_mReg_2, A1=>nx9549, 
      A2=>nx10631);
   ix4735 : nor03_2x port map ( Y=>nx4734, A0=>nx5857, A1=>nx10637, A2=>
      nx10647);
   ix5868 : nor02_2x port map ( Y=>nx5867, A0=>nx4730, A1=>nx4728);
   ix4731 : nor03_2x port map ( Y=>nx4730, A0=>nx5871, A1=>nx9543, A2=>
      nx10655);
   gen_12_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_12_cmp_mReg_3, QB=>
      nx5871, D=>window_12_3, CLK=>start, R=>rst);
   ix4729 : nor03_2x port map ( Y=>nx4728, A0=>gen_12_cmp_mReg_3, A1=>
      nx10071, A2=>nx10663);
   ix4765 : nand02 port map ( Y=>gen_12_cmp_BSCmp_op2_4, A0=>nx5875, A1=>
      nx5881);
   ix5876 : nor02_2x port map ( Y=>nx5875, A0=>nx4760, A1=>nx4756);
   ix4761 : nor03_2x port map ( Y=>nx4760, A0=>gen_12_cmp_mReg_3, A1=>nx9549, 
      A2=>nx10631);
   ix4757 : nor03_2x port map ( Y=>nx4756, A0=>nx5871, A1=>nx10637, A2=>
      nx10647);
   ix5882 : nor02_2x port map ( Y=>nx5881, A0=>nx4752, A1=>nx4750);
   ix4753 : nor03_2x port map ( Y=>nx4752, A0=>nx5884, A1=>nx9543, A2=>
      nx10655);
   gen_12_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_12_cmp_mReg_4, QB=>
      nx5884, D=>window_12_4, CLK=>start, R=>rst);
   ix4751 : nor03_2x port map ( Y=>nx4750, A0=>gen_12_cmp_mReg_4, A1=>
      nx10071, A2=>nx10663);
   ix4787 : nand02 port map ( Y=>gen_12_cmp_BSCmp_op2_5, A0=>nx5891, A1=>
      nx5897);
   ix5892 : nor02_2x port map ( Y=>nx5891, A0=>nx4782, A1=>nx4778);
   ix4783 : nor03_2x port map ( Y=>nx4782, A0=>gen_12_cmp_mReg_4, A1=>nx9549, 
      A2=>nx10631);
   ix4779 : nor03_2x port map ( Y=>nx4778, A0=>nx5884, A1=>nx10637, A2=>
      nx10647);
   ix5898 : nor02_2x port map ( Y=>nx5897, A0=>nx4774, A1=>nx4772);
   ix4775 : nor03_2x port map ( Y=>nx4774, A0=>nx5901, A1=>nx9545, A2=>
      nx10655);
   gen_12_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_12_cmp_mReg_5, QB=>
      nx5901, D=>window_12_5, CLK=>start, R=>rst);
   ix4773 : nor03_2x port map ( Y=>nx4772, A0=>gen_12_cmp_mReg_5, A1=>
      nx10071, A2=>nx10663);
   ix4809 : nand02 port map ( Y=>gen_12_cmp_BSCmp_op2_6, A0=>nx5905, A1=>
      nx5911);
   ix5906 : nor02_2x port map ( Y=>nx5905, A0=>nx4804, A1=>nx4800);
   ix4805 : nor03_2x port map ( Y=>nx4804, A0=>gen_12_cmp_mReg_5, A1=>nx9551, 
      A2=>nx10631);
   ix4801 : nor03_2x port map ( Y=>nx4800, A0=>nx5901, A1=>nx10637, A2=>
      nx10647);
   ix5912 : nor02_2x port map ( Y=>nx5911, A0=>nx4796, A1=>nx4794);
   ix4797 : nor03_2x port map ( Y=>nx4796, A0=>nx5915, A1=>nx9545, A2=>
      nx10655);
   gen_12_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_12_cmp_mReg_6, QB=>
      nx5915, D=>window_12_6, CLK=>start, R=>rst);
   ix4795 : nor03_2x port map ( Y=>nx4794, A0=>gen_12_cmp_mReg_6, A1=>
      nx10071, A2=>nx10663);
   ix4831 : nand02 port map ( Y=>gen_12_cmp_BSCmp_op2_7, A0=>nx5919, A1=>
      nx5925);
   ix5920 : nor02_2x port map ( Y=>nx5919, A0=>nx4826, A1=>nx4822);
   ix4827 : nor03_2x port map ( Y=>nx4826, A0=>gen_12_cmp_mReg_6, A1=>nx9551, 
      A2=>nx10633);
   ix4823 : nor03_2x port map ( Y=>nx4822, A0=>nx5915, A1=>nx10639, A2=>
      nx10649);
   ix5926 : nor02_2x port map ( Y=>nx5925, A0=>nx4818, A1=>nx4816);
   ix4819 : nor03_2x port map ( Y=>nx4818, A0=>nx5928, A1=>nx9545, A2=>
      nx10657);
   gen_12_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_12_cmp_mReg_7, QB=>
      nx5928, D=>window_12_7, CLK=>start, R=>rst);
   ix4817 : nor03_2x port map ( Y=>nx4816, A0=>gen_12_cmp_mReg_7, A1=>
      nx10071, A2=>nx10665);
   ix4853 : nand02 port map ( Y=>gen_12_cmp_BSCmp_op2_8, A0=>nx5935, A1=>
      nx5941);
   ix5936 : nor02_2x port map ( Y=>nx5935, A0=>nx4848, A1=>nx4844);
   ix4849 : nor03_2x port map ( Y=>nx4848, A0=>gen_12_cmp_mReg_7, A1=>nx9551, 
      A2=>nx10633);
   ix4845 : nor03_2x port map ( Y=>nx4844, A0=>nx5928, A1=>nx10639, A2=>
      nx10649);
   ix5942 : nor02_2x port map ( Y=>nx5941, A0=>nx4840, A1=>nx4838);
   ix4841 : nor03_2x port map ( Y=>nx4840, A0=>nx5945, A1=>nx9545, A2=>
      nx10657);
   gen_12_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_12_cmp_mReg_8, QB=>
      nx5945, D=>window_12_8, CLK=>start, R=>rst);
   ix4839 : nor03_2x port map ( Y=>nx4838, A0=>gen_12_cmp_mReg_8, A1=>
      nx10073, A2=>nx10665);
   ix4875 : nand02 port map ( Y=>gen_12_cmp_BSCmp_op2_9, A0=>nx5949, A1=>
      nx5955);
   ix5950 : nor02_2x port map ( Y=>nx5949, A0=>nx4870, A1=>nx4866);
   ix4871 : nor03_2x port map ( Y=>nx4870, A0=>gen_12_cmp_mReg_8, A1=>nx9551, 
      A2=>nx10633);
   ix4867 : nor03_2x port map ( Y=>nx4866, A0=>nx5945, A1=>nx10639, A2=>
      nx10649);
   ix5956 : nor02_2x port map ( Y=>nx5955, A0=>nx4862, A1=>nx4860);
   ix4863 : nor03_2x port map ( Y=>nx4862, A0=>nx5959, A1=>nx9545, A2=>
      nx10657);
   gen_12_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_12_cmp_mReg_9, QB=>
      nx5959, D=>window_12_9, CLK=>start, R=>rst);
   ix4861 : nor03_2x port map ( Y=>nx4860, A0=>gen_12_cmp_mReg_9, A1=>
      nx10073, A2=>nx10665);
   ix4897 : nand02 port map ( Y=>gen_12_cmp_BSCmp_op2_10, A0=>nx5963, A1=>
      nx5969);
   ix5964 : nor02_2x port map ( Y=>nx5963, A0=>nx4892, A1=>nx4888);
   ix4893 : nor03_2x port map ( Y=>nx4892, A0=>gen_12_cmp_mReg_9, A1=>nx9551, 
      A2=>nx10633);
   ix4889 : nor03_2x port map ( Y=>nx4888, A0=>nx5959, A1=>nx10639, A2=>
      nx10649);
   ix5970 : nor02_2x port map ( Y=>nx5969, A0=>nx4884, A1=>nx4882);
   ix4885 : nor03_2x port map ( Y=>nx4884, A0=>nx5972, A1=>nx9545, A2=>
      nx10657);
   gen_12_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_12_cmp_mReg_10, QB=>
      nx5972, D=>window_12_10, CLK=>start, R=>rst);
   ix4883 : nor03_2x port map ( Y=>nx4882, A0=>gen_12_cmp_mReg_10, A1=>
      nx10073, A2=>nx10665);
   ix4919 : nand02 port map ( Y=>gen_12_cmp_BSCmp_op2_11, A0=>nx5979, A1=>
      nx5985);
   ix5980 : nor02_2x port map ( Y=>nx5979, A0=>nx4914, A1=>nx4910);
   ix4915 : nor03_2x port map ( Y=>nx4914, A0=>gen_12_cmp_mReg_10, A1=>
      nx9551, A2=>nx10633);
   ix4911 : nor03_2x port map ( Y=>nx4910, A0=>nx5972, A1=>nx10639, A2=>
      nx10649);
   ix5986 : nor02_2x port map ( Y=>nx5985, A0=>nx4906, A1=>nx4904);
   ix4907 : nor03_2x port map ( Y=>nx4906, A0=>nx5989, A1=>nx9545, A2=>
      nx10657);
   gen_12_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_12_cmp_mReg_11, QB=>
      nx5989, D=>window_12_11, CLK=>start, R=>rst);
   ix4905 : nor03_2x port map ( Y=>nx4904, A0=>gen_12_cmp_mReg_11, A1=>
      nx10073, A2=>nx10665);
   ix4941 : nand02 port map ( Y=>gen_12_cmp_BSCmp_op2_12, A0=>nx5993, A1=>
      nx5999);
   ix5994 : nor02_2x port map ( Y=>nx5993, A0=>nx4936, A1=>nx4932);
   ix4937 : nor03_2x port map ( Y=>nx4936, A0=>gen_12_cmp_mReg_11, A1=>
      nx9551, A2=>nx10633);
   ix4933 : nor03_2x port map ( Y=>nx4932, A0=>nx5989, A1=>nx10639, A2=>
      nx10649);
   ix6000 : nor02_2x port map ( Y=>nx5999, A0=>nx4928, A1=>nx4926);
   ix4929 : nor03_2x port map ( Y=>nx4928, A0=>nx6003, A1=>nx9547, A2=>
      nx10657);
   gen_12_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_12_cmp_mReg_12, QB=>
      nx6003, D=>window_12_12, CLK=>start, R=>rst);
   ix4927 : nor03_2x port map ( Y=>nx4926, A0=>gen_12_cmp_mReg_12, A1=>
      nx10073, A2=>nx10665);
   ix4963 : nand02 port map ( Y=>gen_12_cmp_BSCmp_op2_13, A0=>nx6007, A1=>
      nx6013);
   ix6008 : nor02_2x port map ( Y=>nx6007, A0=>nx4958, A1=>nx4954);
   ix4959 : nor03_2x port map ( Y=>nx4958, A0=>gen_12_cmp_mReg_12, A1=>
      nx9553, A2=>nx10635);
   ix4955 : nor03_2x port map ( Y=>nx4954, A0=>nx6003, A1=>nx10639, A2=>
      nx10651);
   ix6014 : nor02_2x port map ( Y=>nx6013, A0=>nx4950, A1=>nx4948);
   ix4951 : nor03_2x port map ( Y=>nx4950, A0=>nx6016, A1=>nx9547, A2=>
      nx10659);
   gen_12_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_12_cmp_mReg_13, QB=>
      nx6016, D=>window_12_13, CLK=>start, R=>rst);
   ix4949 : nor03_2x port map ( Y=>nx4948, A0=>gen_12_cmp_mReg_13, A1=>
      nx10073, A2=>nx10667);
   ix4985 : nand02 port map ( Y=>gen_12_cmp_BSCmp_op2_14, A0=>nx6023, A1=>
      nx6029);
   ix6024 : nor02_2x port map ( Y=>nx6023, A0=>nx4980, A1=>nx4976);
   ix4981 : nor03_2x port map ( Y=>nx4980, A0=>gen_12_cmp_mReg_13, A1=>
      nx9553, A2=>nx10635);
   ix4977 : nor03_2x port map ( Y=>nx4976, A0=>nx6016, A1=>nx10641, A2=>
      nx10651);
   ix6030 : nor02_2x port map ( Y=>nx6029, A0=>nx4972, A1=>nx4970);
   ix4973 : nor03_2x port map ( Y=>nx4972, A0=>nx6033, A1=>nx9547, A2=>
      nx10659);
   gen_12_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_12_cmp_mReg_14, QB=>
      nx6033, D=>window_12_14, CLK=>start, R=>rst);
   ix4971 : nor03_2x port map ( Y=>nx4970, A0=>gen_12_cmp_mReg_14, A1=>
      nx10073, A2=>nx10667);
   ix5007 : nand02 port map ( Y=>gen_12_cmp_BSCmp_op2_15, A0=>nx6037, A1=>
      nx6043);
   ix6038 : nor02_2x port map ( Y=>nx6037, A0=>nx5002, A1=>nx4998);
   ix5003 : nor03_2x port map ( Y=>nx5002, A0=>gen_12_cmp_mReg_14, A1=>
      nx9553, A2=>nx10635);
   ix4999 : nor03_2x port map ( Y=>nx4998, A0=>nx6033, A1=>nx10641, A2=>
      nx10651);
   ix6044 : nor02_2x port map ( Y=>nx6043, A0=>nx4994, A1=>nx4992);
   ix4995 : nor03_2x port map ( Y=>nx4994, A0=>nx6047, A1=>nx9547, A2=>
      nx10659);
   gen_12_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_12_cmp_mReg_15, QB=>
      nx6047, D=>window_12_15, CLK=>start, R=>rst);
   ix4993 : nor03_2x port map ( Y=>nx4992, A0=>gen_12_cmp_mReg_15, A1=>
      nx10075, A2=>nx10667);
   ix5017 : nand02 port map ( Y=>gen_12_cmp_BSCmp_op2_16, A0=>nx6051, A1=>
      nx6043);
   ix6052 : nor02_2x port map ( Y=>nx6051, A0=>nx5012, A1=>nx5008);
   ix5013 : nor03_2x port map ( Y=>nx5012, A0=>gen_12_cmp_mReg_15, A1=>
      nx9553, A2=>nx10635);
   ix5009 : nor03_2x port map ( Y=>nx5008, A0=>nx6047, A1=>nx10641, A2=>
      nx10651);
   ix5085 : nand02 port map ( Y=>gen_13_cmp_BSCmp_op2_1, A0=>nx6058, A1=>
      nx6077);
   ix6059 : nor02_2x port map ( Y=>nx6058, A0=>nx5080, A1=>nx5076);
   ix5081 : nor03_2x port map ( Y=>nx5080, A0=>gen_13_cmp_mReg_0, A1=>nx9537, 
      A2=>nx10671);
   gen_13_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_13_cmp_mReg_0, QB=>
      nx6063, D=>window_13_0, CLK=>start, R=>rst);
   ix6068 : inv01 port map ( Y=>nx6067, A=>gen_13_cmp_pMux_0);
   ix5077 : nor03_2x port map ( Y=>nx5076, A0=>nx6063, A1=>nx10677, A2=>
      nx10687);
   ix6076 : inv02 port map ( Y=>nx6075, A=>gen_13_cmp_pMux_2);
   ix6078 : nor02_2x port map ( Y=>nx6077, A0=>nx5066, A1=>nx5064);
   ix5067 : nor03_2x port map ( Y=>nx5066, A0=>nx6080, A1=>nx9531, A2=>
      nx10695);
   gen_13_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_13_cmp_mReg_1, QB=>
      nx6080, D=>window_13_1, CLK=>start, R=>rst);
   ix5065 : nor03_2x port map ( Y=>nx5064, A0=>gen_13_cmp_mReg_1, A1=>
      nx10077, A2=>nx10703);
   ix5025 : nor03_2x port map ( Y=>nx5024, A0=>nx9537, A1=>nx6075, A2=>
      gen_13_cmp_pMux_0);
   ix5107 : nand02 port map ( Y=>gen_13_cmp_BSCmp_op2_2, A0=>nx6093, A1=>
      nx6099);
   ix6094 : nor02_2x port map ( Y=>nx6093, A0=>nx5102, A1=>nx5098);
   ix5103 : nor03_2x port map ( Y=>nx5102, A0=>gen_13_cmp_mReg_1, A1=>nx9537, 
      A2=>nx10671);
   ix5099 : nor03_2x port map ( Y=>nx5098, A0=>nx6080, A1=>nx10677, A2=>
      nx10687);
   ix6100 : nor02_2x port map ( Y=>nx6099, A0=>nx5094, A1=>nx5092);
   ix5095 : nor03_2x port map ( Y=>nx5094, A0=>nx6102, A1=>nx9531, A2=>
      nx10695);
   gen_13_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_13_cmp_mReg_2, QB=>
      nx6102, D=>window_13_2, CLK=>start, R=>rst);
   ix5093 : nor03_2x port map ( Y=>nx5092, A0=>gen_13_cmp_mReg_2, A1=>
      nx10077, A2=>nx10703);
   ix5129 : nand02 port map ( Y=>gen_13_cmp_BSCmp_op2_3, A0=>nx6107, A1=>
      nx6113);
   ix6108 : nor02_2x port map ( Y=>nx6107, A0=>nx5124, A1=>nx5120);
   ix5125 : nor03_2x port map ( Y=>nx5124, A0=>gen_13_cmp_mReg_2, A1=>nx9537, 
      A2=>nx10671);
   ix5121 : nor03_2x port map ( Y=>nx5120, A0=>nx6102, A1=>nx10677, A2=>
      nx10687);
   ix6114 : nor02_2x port map ( Y=>nx6113, A0=>nx5116, A1=>nx5114);
   ix5117 : nor03_2x port map ( Y=>nx5116, A0=>nx6117, A1=>nx9531, A2=>
      nx10695);
   gen_13_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_13_cmp_mReg_3, QB=>
      nx6117, D=>window_13_3, CLK=>start, R=>rst);
   ix5115 : nor03_2x port map ( Y=>nx5114, A0=>gen_13_cmp_mReg_3, A1=>
      nx10077, A2=>nx10703);
   ix5151 : nand02 port map ( Y=>gen_13_cmp_BSCmp_op2_4, A0=>nx6123, A1=>
      nx6127);
   ix6124 : nor02_2x port map ( Y=>nx6123, A0=>nx5146, A1=>nx5142);
   ix5147 : nor03_2x port map ( Y=>nx5146, A0=>gen_13_cmp_mReg_3, A1=>nx9537, 
      A2=>nx10671);
   ix5143 : nor03_2x port map ( Y=>nx5142, A0=>nx6117, A1=>nx10677, A2=>
      nx10687);
   ix6128 : nor02_2x port map ( Y=>nx6127, A0=>nx5138, A1=>nx5136);
   ix5139 : nor03_2x port map ( Y=>nx5138, A0=>nx6131, A1=>nx9531, A2=>
      nx10695);
   gen_13_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_13_cmp_mReg_4, QB=>
      nx6131, D=>window_13_4, CLK=>start, R=>rst);
   ix5137 : nor03_2x port map ( Y=>nx5136, A0=>gen_13_cmp_mReg_4, A1=>
      nx10077, A2=>nx10703);
   ix5173 : nand02 port map ( Y=>gen_13_cmp_BSCmp_op2_5, A0=>nx6137, A1=>
      nx6143);
   ix6138 : nor02_2x port map ( Y=>nx6137, A0=>nx5168, A1=>nx5164);
   ix5169 : nor03_2x port map ( Y=>nx5168, A0=>gen_13_cmp_mReg_4, A1=>nx9537, 
      A2=>nx10671);
   ix5165 : nor03_2x port map ( Y=>nx5164, A0=>nx6131, A1=>nx10677, A2=>
      nx10687);
   ix6144 : nor02_2x port map ( Y=>nx6143, A0=>nx5160, A1=>nx5158);
   ix5161 : nor03_2x port map ( Y=>nx5160, A0=>nx6146, A1=>nx9533, A2=>
      nx10695);
   gen_13_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_13_cmp_mReg_5, QB=>
      nx6146, D=>window_13_5, CLK=>start, R=>rst);
   ix5159 : nor03_2x port map ( Y=>nx5158, A0=>gen_13_cmp_mReg_5, A1=>
      nx10077, A2=>nx10703);
   ix5195 : nand02 port map ( Y=>gen_13_cmp_BSCmp_op2_6, A0=>nx6151, A1=>
      nx6157);
   ix6152 : nor02_2x port map ( Y=>nx6151, A0=>nx5190, A1=>nx5186);
   ix5191 : nor03_2x port map ( Y=>nx5190, A0=>gen_13_cmp_mReg_5, A1=>nx9539, 
      A2=>nx10671);
   ix5187 : nor03_2x port map ( Y=>nx5186, A0=>nx6146, A1=>nx10677, A2=>
      nx10687);
   ix6158 : nor02_2x port map ( Y=>nx6157, A0=>nx5182, A1=>nx5180);
   ix5183 : nor03_2x port map ( Y=>nx5182, A0=>nx6161, A1=>nx9533, A2=>
      nx10695);
   gen_13_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_13_cmp_mReg_6, QB=>
      nx6161, D=>window_13_6, CLK=>start, R=>rst);
   ix5181 : nor03_2x port map ( Y=>nx5180, A0=>gen_13_cmp_mReg_6, A1=>
      nx10077, A2=>nx10703);
   ix5217 : nand02 port map ( Y=>gen_13_cmp_BSCmp_op2_7, A0=>nx6167, A1=>
      nx6171);
   ix6168 : nor02_2x port map ( Y=>nx6167, A0=>nx5212, A1=>nx5208);
   ix5213 : nor03_2x port map ( Y=>nx5212, A0=>gen_13_cmp_mReg_6, A1=>nx9539, 
      A2=>nx10673);
   ix5209 : nor03_2x port map ( Y=>nx5208, A0=>nx6161, A1=>nx10679, A2=>
      nx10689);
   ix6172 : nor02_2x port map ( Y=>nx6171, A0=>nx5204, A1=>nx5202);
   ix5205 : nor03_2x port map ( Y=>nx5204, A0=>nx6175, A1=>nx9533, A2=>
      nx10697);
   gen_13_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_13_cmp_mReg_7, QB=>
      nx6175, D=>window_13_7, CLK=>start, R=>rst);
   ix5203 : nor03_2x port map ( Y=>nx5202, A0=>gen_13_cmp_mReg_7, A1=>
      nx10077, A2=>nx10705);
   ix5239 : nand02 port map ( Y=>gen_13_cmp_BSCmp_op2_8, A0=>nx6181, A1=>
      nx6186);
   ix6182 : nor02_2x port map ( Y=>nx6181, A0=>nx5234, A1=>nx5230);
   ix5235 : nor03_2x port map ( Y=>nx5234, A0=>gen_13_cmp_mReg_7, A1=>nx9539, 
      A2=>nx10673);
   ix5231 : nor03_2x port map ( Y=>nx5230, A0=>nx6175, A1=>nx10679, A2=>
      nx10689);
   ix6187 : nor02_2x port map ( Y=>nx6186, A0=>nx5226, A1=>nx5224);
   ix5227 : nor03_2x port map ( Y=>nx5226, A0=>nx6189, A1=>nx9533, A2=>
      nx10697);
   gen_13_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_13_cmp_mReg_8, QB=>
      nx6189, D=>window_13_8, CLK=>start, R=>rst);
   ix5225 : nor03_2x port map ( Y=>nx5224, A0=>gen_13_cmp_mReg_8, A1=>
      nx10079, A2=>nx10705);
   ix5261 : nand02 port map ( Y=>gen_13_cmp_BSCmp_op2_9, A0=>nx6193, A1=>
      nx6199);
   ix6194 : nor02_2x port map ( Y=>nx6193, A0=>nx5256, A1=>nx5252);
   ix5257 : nor03_2x port map ( Y=>nx5256, A0=>gen_13_cmp_mReg_8, A1=>nx9539, 
      A2=>nx10673);
   ix5253 : nor03_2x port map ( Y=>nx5252, A0=>nx6189, A1=>nx10679, A2=>
      nx10689);
   ix6200 : nor02_2x port map ( Y=>nx6199, A0=>nx5248, A1=>nx5246);
   ix5249 : nor03_2x port map ( Y=>nx5248, A0=>nx6203, A1=>nx9533, A2=>
      nx10697);
   gen_13_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_13_cmp_mReg_9, QB=>
      nx6203, D=>window_13_9, CLK=>start, R=>rst);
   ix5247 : nor03_2x port map ( Y=>nx5246, A0=>gen_13_cmp_mReg_9, A1=>
      nx10079, A2=>nx10705);
   ix5283 : nand02 port map ( Y=>gen_13_cmp_BSCmp_op2_10, A0=>nx6209, A1=>
      nx6215);
   ix6210 : nor02_2x port map ( Y=>nx6209, A0=>nx5278, A1=>nx5274);
   ix5279 : nor03_2x port map ( Y=>nx5278, A0=>gen_13_cmp_mReg_9, A1=>nx9539, 
      A2=>nx10673);
   ix5275 : nor03_2x port map ( Y=>nx5274, A0=>nx6203, A1=>nx10679, A2=>
      nx10689);
   ix6216 : nor02_2x port map ( Y=>nx6215, A0=>nx5270, A1=>nx5268);
   ix5271 : nor03_2x port map ( Y=>nx5270, A0=>nx6218, A1=>nx9533, A2=>
      nx10697);
   gen_13_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_13_cmp_mReg_10, QB=>
      nx6218, D=>window_13_10, CLK=>start, R=>rst);
   ix5269 : nor03_2x port map ( Y=>nx5268, A0=>gen_13_cmp_mReg_10, A1=>
      nx10079, A2=>nx10705);
   ix5305 : nand02 port map ( Y=>gen_13_cmp_BSCmp_op2_11, A0=>nx6223, A1=>
      nx6229);
   ix6224 : nor02_2x port map ( Y=>nx6223, A0=>nx5300, A1=>nx5296);
   ix5301 : nor03_2x port map ( Y=>nx5300, A0=>gen_13_cmp_mReg_10, A1=>
      nx9539, A2=>nx10673);
   ix5297 : nor03_2x port map ( Y=>nx5296, A0=>nx6218, A1=>nx10679, A2=>
      nx10689);
   ix6230 : nor02_2x port map ( Y=>nx6229, A0=>nx5292, A1=>nx5290);
   ix5293 : nor03_2x port map ( Y=>nx5292, A0=>nx6233, A1=>nx9533, A2=>
      nx10697);
   gen_13_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_13_cmp_mReg_11, QB=>
      nx6233, D=>window_13_11, CLK=>start, R=>rst);
   ix5291 : nor03_2x port map ( Y=>nx5290, A0=>gen_13_cmp_mReg_11, A1=>
      nx10079, A2=>nx10705);
   ix5327 : nand02 port map ( Y=>gen_13_cmp_BSCmp_op2_12, A0=>nx6239, A1=>
      nx6245);
   ix6240 : nor02_2x port map ( Y=>nx6239, A0=>nx5322, A1=>nx5318);
   ix5323 : nor03_2x port map ( Y=>nx5322, A0=>gen_13_cmp_mReg_11, A1=>
      nx9539, A2=>nx10673);
   ix5319 : nor03_2x port map ( Y=>nx5318, A0=>nx6233, A1=>nx10679, A2=>
      nx10689);
   ix6246 : nor02_2x port map ( Y=>nx6245, A0=>nx5314, A1=>nx5312);
   ix5315 : nor03_2x port map ( Y=>nx5314, A0=>nx6248, A1=>nx9535, A2=>
      nx10697);
   gen_13_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_13_cmp_mReg_12, QB=>
      nx6248, D=>window_13_12, CLK=>start, R=>rst);
   ix5313 : nor03_2x port map ( Y=>nx5312, A0=>gen_13_cmp_mReg_12, A1=>
      nx10079, A2=>nx10705);
   ix5349 : nand02 port map ( Y=>gen_13_cmp_BSCmp_op2_13, A0=>nx6255, A1=>
      nx6261);
   ix6256 : nor02_2x port map ( Y=>nx6255, A0=>nx5344, A1=>nx5340);
   ix5345 : nor03_2x port map ( Y=>nx5344, A0=>gen_13_cmp_mReg_12, A1=>
      nx9541, A2=>nx10675);
   ix5341 : nor03_2x port map ( Y=>nx5340, A0=>nx6248, A1=>nx10679, A2=>
      nx10691);
   ix6262 : nor02_2x port map ( Y=>nx6261, A0=>nx5336, A1=>nx5334);
   ix5337 : nor03_2x port map ( Y=>nx5336, A0=>nx6265, A1=>nx9535, A2=>
      nx10699);
   gen_13_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_13_cmp_mReg_13, QB=>
      nx6265, D=>window_13_13, CLK=>start, R=>rst);
   ix5335 : nor03_2x port map ( Y=>nx5334, A0=>gen_13_cmp_mReg_13, A1=>
      nx10079, A2=>nx10707);
   ix5371 : nand02 port map ( Y=>gen_13_cmp_BSCmp_op2_14, A0=>nx6269, A1=>
      nx6275);
   ix6270 : nor02_2x port map ( Y=>nx6269, A0=>nx5366, A1=>nx5362);
   ix5367 : nor03_2x port map ( Y=>nx5366, A0=>gen_13_cmp_mReg_13, A1=>
      nx9541, A2=>nx10675);
   ix5363 : nor03_2x port map ( Y=>nx5362, A0=>nx6265, A1=>nx10681, A2=>
      nx10691);
   ix6276 : nor02_2x port map ( Y=>nx6275, A0=>nx5358, A1=>nx5356);
   ix5359 : nor03_2x port map ( Y=>nx5358, A0=>nx6279, A1=>nx9535, A2=>
      nx10699);
   gen_13_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_13_cmp_mReg_14, QB=>
      nx6279, D=>window_13_14, CLK=>start, R=>rst);
   ix5357 : nor03_2x port map ( Y=>nx5356, A0=>gen_13_cmp_mReg_14, A1=>
      nx10079, A2=>nx10707);
   ix5393 : nand02 port map ( Y=>gen_13_cmp_BSCmp_op2_15, A0=>nx6283, A1=>
      nx6289);
   ix6284 : nor02_2x port map ( Y=>nx6283, A0=>nx5388, A1=>nx5384);
   ix5389 : nor03_2x port map ( Y=>nx5388, A0=>gen_13_cmp_mReg_14, A1=>
      nx9541, A2=>nx10675);
   ix5385 : nor03_2x port map ( Y=>nx5384, A0=>nx6279, A1=>nx10681, A2=>
      nx10691);
   ix6290 : nor02_2x port map ( Y=>nx6289, A0=>nx5380, A1=>nx5378);
   ix5381 : nor03_2x port map ( Y=>nx5380, A0=>nx6292, A1=>nx9535, A2=>
      nx10699);
   gen_13_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_13_cmp_mReg_15, QB=>
      nx6292, D=>window_13_15, CLK=>start, R=>rst);
   ix5379 : nor03_2x port map ( Y=>nx5378, A0=>gen_13_cmp_mReg_15, A1=>
      nx10081, A2=>nx10707);
   ix5403 : nand02 port map ( Y=>gen_13_cmp_BSCmp_op2_16, A0=>nx6299, A1=>
      nx6289);
   ix6300 : nor02_2x port map ( Y=>nx6299, A0=>nx5398, A1=>nx5394);
   ix5399 : nor03_2x port map ( Y=>nx5398, A0=>gen_13_cmp_mReg_15, A1=>
      nx9541, A2=>nx10675);
   ix5395 : nor03_2x port map ( Y=>nx5394, A0=>nx6292, A1=>nx10681, A2=>
      nx10691);
   ix5471 : nand02 port map ( Y=>gen_14_cmp_BSCmp_op2_1, A0=>nx6305, A1=>
      nx6325);
   ix6306 : nor02_2x port map ( Y=>nx6305, A0=>nx5466, A1=>nx5462);
   ix5467 : nor03_2x port map ( Y=>nx5466, A0=>gen_14_cmp_mReg_0, A1=>nx9525, 
      A2=>nx10711);
   gen_14_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_14_cmp_mReg_0, QB=>
      nx6311, D=>window_14_0, CLK=>start, R=>rst);
   ix6316 : inv01 port map ( Y=>nx6314, A=>gen_14_cmp_pMux_0);
   ix5463 : nor03_2x port map ( Y=>nx5462, A0=>nx6311, A1=>nx10717, A2=>
      nx10727);
   ix6324 : inv02 port map ( Y=>nx6323, A=>gen_14_cmp_pMux_2);
   ix6326 : nor02_2x port map ( Y=>nx6325, A0=>nx5452, A1=>nx5450);
   ix5453 : nor03_2x port map ( Y=>nx5452, A0=>nx6329, A1=>nx9519, A2=>
      nx10735);
   gen_14_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_14_cmp_mReg_1, QB=>
      nx6329, D=>window_14_1, CLK=>start, R=>rst);
   ix5451 : nor03_2x port map ( Y=>nx5450, A0=>gen_14_cmp_mReg_1, A1=>
      nx10083, A2=>nx10743);
   ix5411 : nor03_2x port map ( Y=>nx5410, A0=>nx9525, A1=>nx6323, A2=>
      gen_14_cmp_pMux_0);
   ix5493 : nand02 port map ( Y=>gen_14_cmp_BSCmp_op2_2, A0=>nx6339, A1=>
      nx6345);
   ix6340 : nor02_2x port map ( Y=>nx6339, A0=>nx5488, A1=>nx5484);
   ix5489 : nor03_2x port map ( Y=>nx5488, A0=>gen_14_cmp_mReg_1, A1=>nx9525, 
      A2=>nx10711);
   ix5485 : nor03_2x port map ( Y=>nx5484, A0=>nx6329, A1=>nx10717, A2=>
      nx10727);
   ix6346 : nor02_2x port map ( Y=>nx6345, A0=>nx5480, A1=>nx5478);
   ix5481 : nor03_2x port map ( Y=>nx5480, A0=>nx6349, A1=>nx9519, A2=>
      nx10735);
   gen_14_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_14_cmp_mReg_2, QB=>
      nx6349, D=>window_14_2, CLK=>start, R=>rst);
   ix5479 : nor03_2x port map ( Y=>nx5478, A0=>gen_14_cmp_mReg_2, A1=>
      nx10083, A2=>nx10743);
   ix5515 : nand02 port map ( Y=>gen_14_cmp_BSCmp_op2_3, A0=>nx6355, A1=>
      nx6359);
   ix6356 : nor02_2x port map ( Y=>nx6355, A0=>nx5510, A1=>nx5506);
   ix5511 : nor03_2x port map ( Y=>nx5510, A0=>gen_14_cmp_mReg_2, A1=>nx9525, 
      A2=>nx10711);
   ix5507 : nor03_2x port map ( Y=>nx5506, A0=>nx6349, A1=>nx10717, A2=>
      nx10727);
   ix6360 : nor02_2x port map ( Y=>nx6359, A0=>nx5502, A1=>nx5500);
   ix5503 : nor03_2x port map ( Y=>nx5502, A0=>nx6363, A1=>nx9519, A2=>
      nx10735);
   gen_14_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_14_cmp_mReg_3, QB=>
      nx6363, D=>window_14_3, CLK=>start, R=>rst);
   ix5501 : nor03_2x port map ( Y=>nx5500, A0=>gen_14_cmp_mReg_3, A1=>
      nx10083, A2=>nx10743);
   ix5537 : nand02 port map ( Y=>gen_14_cmp_BSCmp_op2_4, A0=>nx6369, A1=>
      nx6375);
   ix6370 : nor02_2x port map ( Y=>nx6369, A0=>nx5532, A1=>nx5528);
   ix5533 : nor03_2x port map ( Y=>nx5532, A0=>gen_14_cmp_mReg_3, A1=>nx9525, 
      A2=>nx10711);
   ix5529 : nor03_2x port map ( Y=>nx5528, A0=>nx6363, A1=>nx10717, A2=>
      nx10727);
   ix6376 : nor02_2x port map ( Y=>nx6375, A0=>nx5524, A1=>nx5522);
   ix5525 : nor03_2x port map ( Y=>nx5524, A0=>nx6378, A1=>nx9519, A2=>
      nx10735);
   gen_14_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_14_cmp_mReg_4, QB=>
      nx6378, D=>window_14_4, CLK=>start, R=>rst);
   ix5523 : nor03_2x port map ( Y=>nx5522, A0=>gen_14_cmp_mReg_4, A1=>
      nx10083, A2=>nx10743);
   ix5559 : nand02 port map ( Y=>gen_14_cmp_BSCmp_op2_5, A0=>nx6383, A1=>
      nx6389);
   ix6384 : nor02_2x port map ( Y=>nx6383, A0=>nx5554, A1=>nx5550);
   ix5555 : nor03_2x port map ( Y=>nx5554, A0=>gen_14_cmp_mReg_4, A1=>nx9525, 
      A2=>nx10711);
   ix5551 : nor03_2x port map ( Y=>nx5550, A0=>nx6378, A1=>nx10717, A2=>
      nx10727);
   ix6390 : nor02_2x port map ( Y=>nx6389, A0=>nx5546, A1=>nx5544);
   ix5547 : nor03_2x port map ( Y=>nx5546, A0=>nx6393, A1=>nx9521, A2=>
      nx10735);
   gen_14_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_14_cmp_mReg_5, QB=>
      nx6393, D=>window_14_5, CLK=>start, R=>rst);
   ix5545 : nor03_2x port map ( Y=>nx5544, A0=>gen_14_cmp_mReg_5, A1=>
      nx10083, A2=>nx10743);
   ix5581 : nand02 port map ( Y=>gen_14_cmp_BSCmp_op2_6, A0=>nx6399, A1=>
      nx6403);
   ix6400 : nor02_2x port map ( Y=>nx6399, A0=>nx5576, A1=>nx5572);
   ix5577 : nor03_2x port map ( Y=>nx5576, A0=>gen_14_cmp_mReg_5, A1=>nx9527, 
      A2=>nx10711);
   ix5573 : nor03_2x port map ( Y=>nx5572, A0=>nx6393, A1=>nx10717, A2=>
      nx10727);
   ix6404 : nor02_2x port map ( Y=>nx6403, A0=>nx5568, A1=>nx5566);
   ix5569 : nor03_2x port map ( Y=>nx5568, A0=>nx6407, A1=>nx9521, A2=>
      nx10735);
   gen_14_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_14_cmp_mReg_6, QB=>
      nx6407, D=>window_14_6, CLK=>start, R=>rst);
   ix5567 : nor03_2x port map ( Y=>nx5566, A0=>gen_14_cmp_mReg_6, A1=>
      nx10083, A2=>nx10743);
   ix5603 : nand02 port map ( Y=>gen_14_cmp_BSCmp_op2_7, A0=>nx6413, A1=>
      nx6419);
   ix6414 : nor02_2x port map ( Y=>nx6413, A0=>nx5598, A1=>nx5594);
   ix5599 : nor03_2x port map ( Y=>nx5598, A0=>gen_14_cmp_mReg_6, A1=>nx9527, 
      A2=>nx10713);
   ix5595 : nor03_2x port map ( Y=>nx5594, A0=>nx6407, A1=>nx10719, A2=>
      nx10729);
   ix6420 : nor02_2x port map ( Y=>nx6419, A0=>nx5590, A1=>nx5588);
   ix5591 : nor03_2x port map ( Y=>nx5590, A0=>nx6422, A1=>nx9521, A2=>
      nx10737);
   gen_14_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_14_cmp_mReg_7, QB=>
      nx6422, D=>window_14_7, CLK=>start, R=>rst);
   ix5589 : nor03_2x port map ( Y=>nx5588, A0=>gen_14_cmp_mReg_7, A1=>
      nx10083, A2=>nx10745);
   ix5625 : nand02 port map ( Y=>gen_14_cmp_BSCmp_op2_8, A0=>nx6427, A1=>
      nx6433);
   ix6428 : nor02_2x port map ( Y=>nx6427, A0=>nx5620, A1=>nx5616);
   ix5621 : nor03_2x port map ( Y=>nx5620, A0=>gen_14_cmp_mReg_7, A1=>nx9527, 
      A2=>nx10713);
   ix5617 : nor03_2x port map ( Y=>nx5616, A0=>nx6422, A1=>nx10719, A2=>
      nx10729);
   ix6434 : nor02_2x port map ( Y=>nx6433, A0=>nx5612, A1=>nx5610);
   ix5613 : nor03_2x port map ( Y=>nx5612, A0=>nx6437, A1=>nx9521, A2=>
      nx10737);
   gen_14_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_14_cmp_mReg_8, QB=>
      nx6437, D=>window_14_8, CLK=>start, R=>rst);
   ix5611 : nor03_2x port map ( Y=>nx5610, A0=>gen_14_cmp_mReg_8, A1=>
      nx10085, A2=>nx10745);
   ix5647 : nand02 port map ( Y=>gen_14_cmp_BSCmp_op2_9, A0=>nx6443, A1=>
      nx6447);
   ix6444 : nor02_2x port map ( Y=>nx6443, A0=>nx5642, A1=>nx5638);
   ix5643 : nor03_2x port map ( Y=>nx5642, A0=>gen_14_cmp_mReg_8, A1=>nx9527, 
      A2=>nx10713);
   ix5639 : nor03_2x port map ( Y=>nx5638, A0=>nx6437, A1=>nx10719, A2=>
      nx10729);
   ix6448 : nor02_2x port map ( Y=>nx6447, A0=>nx5634, A1=>nx5632);
   ix5635 : nor03_2x port map ( Y=>nx5634, A0=>nx6451, A1=>nx9521, A2=>
      nx10737);
   gen_14_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_14_cmp_mReg_9, QB=>
      nx6451, D=>window_14_9, CLK=>start, R=>rst);
   ix5633 : nor03_2x port map ( Y=>nx5632, A0=>gen_14_cmp_mReg_9, A1=>
      nx10085, A2=>nx10745);
   ix5669 : nand02 port map ( Y=>gen_14_cmp_BSCmp_op2_10, A0=>nx6457, A1=>
      nx6463);
   ix6458 : nor02_2x port map ( Y=>nx6457, A0=>nx5664, A1=>nx5660);
   ix5665 : nor03_2x port map ( Y=>nx5664, A0=>gen_14_cmp_mReg_9, A1=>nx9527, 
      A2=>nx10713);
   ix5661 : nor03_2x port map ( Y=>nx5660, A0=>nx6451, A1=>nx10719, A2=>
      nx10729);
   ix6464 : nor02_2x port map ( Y=>nx6463, A0=>nx5656, A1=>nx5654);
   ix5657 : nor03_2x port map ( Y=>nx5656, A0=>nx6466, A1=>nx9521, A2=>
      nx10737);
   gen_14_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_14_cmp_mReg_10, QB=>
      nx6466, D=>window_14_10, CLK=>start, R=>rst);
   ix5655 : nor03_2x port map ( Y=>nx5654, A0=>gen_14_cmp_mReg_10, A1=>
      nx10085, A2=>nx10745);
   ix5691 : nand02 port map ( Y=>gen_14_cmp_BSCmp_op2_11, A0=>nx6471, A1=>
      nx6477);
   ix6472 : nor02_2x port map ( Y=>nx6471, A0=>nx5686, A1=>nx5682);
   ix5687 : nor03_2x port map ( Y=>nx5686, A0=>gen_14_cmp_mReg_10, A1=>
      nx9527, A2=>nx10713);
   ix5683 : nor03_2x port map ( Y=>nx5682, A0=>nx6466, A1=>nx10719, A2=>
      nx10729);
   ix6478 : nor02_2x port map ( Y=>nx6477, A0=>nx5678, A1=>nx5676);
   ix5679 : nor03_2x port map ( Y=>nx5678, A0=>nx6481, A1=>nx9521, A2=>
      nx10737);
   gen_14_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_14_cmp_mReg_11, QB=>
      nx6481, D=>window_14_11, CLK=>start, R=>rst);
   ix5677 : nor03_2x port map ( Y=>nx5676, A0=>gen_14_cmp_mReg_11, A1=>
      nx10085, A2=>nx10745);
   ix5713 : nand02 port map ( Y=>gen_14_cmp_BSCmp_op2_12, A0=>nx6487, A1=>
      nx6491);
   ix6488 : nor02_2x port map ( Y=>nx6487, A0=>nx5708, A1=>nx5704);
   ix5709 : nor03_2x port map ( Y=>nx5708, A0=>gen_14_cmp_mReg_11, A1=>
      nx9527, A2=>nx10713);
   ix5705 : nor03_2x port map ( Y=>nx5704, A0=>nx6481, A1=>nx10719, A2=>
      nx10729);
   ix6492 : nor02_2x port map ( Y=>nx6491, A0=>nx5700, A1=>nx5698);
   ix5701 : nor03_2x port map ( Y=>nx5700, A0=>nx6495, A1=>nx9523, A2=>
      nx10737);
   gen_14_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_14_cmp_mReg_12, QB=>
      nx6495, D=>window_14_12, CLK=>start, R=>rst);
   ix5699 : nor03_2x port map ( Y=>nx5698, A0=>gen_14_cmp_mReg_12, A1=>
      nx10085, A2=>nx10745);
   ix5735 : nand02 port map ( Y=>gen_14_cmp_BSCmp_op2_13, A0=>nx6501, A1=>
      nx6507);
   ix6502 : nor02_2x port map ( Y=>nx6501, A0=>nx5730, A1=>nx5726);
   ix5731 : nor03_2x port map ( Y=>nx5730, A0=>gen_14_cmp_mReg_12, A1=>
      nx9529, A2=>nx10715);
   ix5727 : nor03_2x port map ( Y=>nx5726, A0=>nx6495, A1=>nx10719, A2=>
      nx10731);
   ix6508 : nor02_2x port map ( Y=>nx6507, A0=>nx5722, A1=>nx5720);
   ix5723 : nor03_2x port map ( Y=>nx5722, A0=>nx6510, A1=>nx9523, A2=>
      nx10739);
   gen_14_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_14_cmp_mReg_13, QB=>
      nx6510, D=>window_14_13, CLK=>start, R=>rst);
   ix5721 : nor03_2x port map ( Y=>nx5720, A0=>gen_14_cmp_mReg_13, A1=>
      nx10085, A2=>nx10747);
   ix5757 : nand02 port map ( Y=>gen_14_cmp_BSCmp_op2_14, A0=>nx6515, A1=>
      nx6521);
   ix6516 : nor02_2x port map ( Y=>nx6515, A0=>nx5752, A1=>nx5748);
   ix5753 : nor03_2x port map ( Y=>nx5752, A0=>gen_14_cmp_mReg_13, A1=>
      nx9529, A2=>nx10715);
   ix5749 : nor03_2x port map ( Y=>nx5748, A0=>nx6510, A1=>nx10721, A2=>
      nx10731);
   ix6522 : nor02_2x port map ( Y=>nx6521, A0=>nx5744, A1=>nx5742);
   ix5745 : nor03_2x port map ( Y=>nx5744, A0=>nx6525, A1=>nx9523, A2=>
      nx10739);
   gen_14_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_14_cmp_mReg_14, QB=>
      nx6525, D=>window_14_14, CLK=>start, R=>rst);
   ix5743 : nor03_2x port map ( Y=>nx5742, A0=>gen_14_cmp_mReg_14, A1=>
      nx10085, A2=>nx10747);
   ix5779 : nand02 port map ( Y=>gen_14_cmp_BSCmp_op2_15, A0=>nx6531, A1=>
      nx6535);
   ix6532 : nor02_2x port map ( Y=>nx6531, A0=>nx5774, A1=>nx5770);
   ix5775 : nor03_2x port map ( Y=>nx5774, A0=>gen_14_cmp_mReg_14, A1=>
      nx9529, A2=>nx10715);
   ix5771 : nor03_2x port map ( Y=>nx5770, A0=>nx6525, A1=>nx10721, A2=>
      nx10731);
   ix6536 : nor02_2x port map ( Y=>nx6535, A0=>nx5766, A1=>nx5764);
   ix5767 : nor03_2x port map ( Y=>nx5766, A0=>nx6539, A1=>nx9523, A2=>
      nx10739);
   gen_14_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_14_cmp_mReg_15, QB=>
      nx6539, D=>window_14_15, CLK=>start, R=>rst);
   ix5765 : nor03_2x port map ( Y=>nx5764, A0=>gen_14_cmp_mReg_15, A1=>
      nx10087, A2=>nx10747);
   ix5789 : nand02 port map ( Y=>gen_14_cmp_BSCmp_op2_16, A0=>nx6545, A1=>
      nx6535);
   ix6546 : nor02_2x port map ( Y=>nx6545, A0=>nx5784, A1=>nx5780);
   ix5785 : nor03_2x port map ( Y=>nx5784, A0=>gen_14_cmp_mReg_15, A1=>
      nx9529, A2=>nx10715);
   ix5781 : nor03_2x port map ( Y=>nx5780, A0=>nx6539, A1=>nx10721, A2=>
      nx10731);
   ix5857 : nand02 port map ( Y=>gen_15_cmp_BSCmp_op2_1, A0=>nx6553, A1=>
      nx6571);
   ix6554 : nor02_2x port map ( Y=>nx6553, A0=>nx5852, A1=>nx5848);
   ix5853 : nor03_2x port map ( Y=>nx5852, A0=>gen_15_cmp_mReg_0, A1=>nx9513, 
      A2=>nx10751);
   gen_15_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_15_cmp_mReg_0, QB=>
      nx6557, D=>window_15_0, CLK=>start, R=>rst);
   ix6562 : inv01 port map ( Y=>nx6561, A=>gen_15_cmp_pMux_0);
   ix5849 : nor03_2x port map ( Y=>nx5848, A0=>nx6557, A1=>nx10757, A2=>
      nx10767);
   ix6570 : inv02 port map ( Y=>nx6569, A=>gen_15_cmp_pMux_2);
   ix6572 : nor02_2x port map ( Y=>nx6571, A0=>nx5838, A1=>nx5836);
   ix5839 : nor03_2x port map ( Y=>nx5838, A0=>nx6574, A1=>nx9507, A2=>
      nx10775);
   gen_15_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_15_cmp_mReg_1, QB=>
      nx6574, D=>window_15_1, CLK=>start, R=>rst);
   ix5837 : nor03_2x port map ( Y=>nx5836, A0=>gen_15_cmp_mReg_1, A1=>
      nx10089, A2=>nx10783);
   ix5797 : nor03_2x port map ( Y=>nx5796, A0=>nx9513, A1=>nx6569, A2=>
      gen_15_cmp_pMux_0);
   ix5879 : nand02 port map ( Y=>gen_15_cmp_BSCmp_op2_2, A0=>nx6585, A1=>
      nx6591);
   ix6586 : nor02_2x port map ( Y=>nx6585, A0=>nx5874, A1=>nx5870);
   ix5875 : nor03_2x port map ( Y=>nx5874, A0=>gen_15_cmp_mReg_1, A1=>nx9513, 
      A2=>nx10751);
   ix5871 : nor03_2x port map ( Y=>nx5870, A0=>nx6574, A1=>nx10757, A2=>
      nx10767);
   ix6592 : nor02_2x port map ( Y=>nx6591, A0=>nx5866, A1=>nx5864);
   ix5867 : nor03_2x port map ( Y=>nx5866, A0=>nx6595, A1=>nx9507, A2=>
      nx10775);
   gen_15_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_15_cmp_mReg_2, QB=>
      nx6595, D=>window_15_2, CLK=>start, R=>rst);
   ix5865 : nor03_2x port map ( Y=>nx5864, A0=>gen_15_cmp_mReg_2, A1=>
      nx10089, A2=>nx10783);
   ix5901 : nand02 port map ( Y=>gen_15_cmp_BSCmp_op2_3, A0=>nx6601, A1=>
      nx6605);
   ix6602 : nor02_2x port map ( Y=>nx6601, A0=>nx5896, A1=>nx5892);
   ix5897 : nor03_2x port map ( Y=>nx5896, A0=>gen_15_cmp_mReg_2, A1=>nx9513, 
      A2=>nx10751);
   ix5893 : nor03_2x port map ( Y=>nx5892, A0=>nx6595, A1=>nx10757, A2=>
      nx10767);
   ix6606 : nor02_2x port map ( Y=>nx6605, A0=>nx5888, A1=>nx5886);
   ix5889 : nor03_2x port map ( Y=>nx5888, A0=>nx6609, A1=>nx9507, A2=>
      nx10775);
   gen_15_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_15_cmp_mReg_3, QB=>
      nx6609, D=>window_15_3, CLK=>start, R=>rst);
   ix5887 : nor03_2x port map ( Y=>nx5886, A0=>gen_15_cmp_mReg_3, A1=>
      nx10089, A2=>nx10783);
   ix5923 : nand02 port map ( Y=>gen_15_cmp_BSCmp_op2_4, A0=>nx6615, A1=>
      nx6621);
   ix6616 : nor02_2x port map ( Y=>nx6615, A0=>nx5918, A1=>nx5914);
   ix5919 : nor03_2x port map ( Y=>nx5918, A0=>gen_15_cmp_mReg_3, A1=>nx9513, 
      A2=>nx10751);
   ix5915 : nor03_2x port map ( Y=>nx5914, A0=>nx6609, A1=>nx10757, A2=>
      nx10767);
   ix6622 : nor02_2x port map ( Y=>nx6621, A0=>nx5910, A1=>nx5908);
   ix5911 : nor03_2x port map ( Y=>nx5910, A0=>nx6625, A1=>nx9507, A2=>
      nx10775);
   gen_15_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_15_cmp_mReg_4, QB=>
      nx6625, D=>window_15_4, CLK=>start, R=>rst);
   ix5909 : nor03_2x port map ( Y=>nx5908, A0=>gen_15_cmp_mReg_4, A1=>
      nx10089, A2=>nx10783);
   ix5945 : nand02 port map ( Y=>gen_15_cmp_BSCmp_op2_5, A0=>nx6631, A1=>
      nx6635);
   ix6632 : nor02_2x port map ( Y=>nx6631, A0=>nx5940, A1=>nx5936);
   ix5941 : nor03_2x port map ( Y=>nx5940, A0=>gen_15_cmp_mReg_4, A1=>nx9513, 
      A2=>nx10751);
   ix5937 : nor03_2x port map ( Y=>nx5936, A0=>nx6625, A1=>nx10757, A2=>
      nx10767);
   ix6636 : nor02_2x port map ( Y=>nx6635, A0=>nx5932, A1=>nx5930);
   ix5933 : nor03_2x port map ( Y=>nx5932, A0=>nx6639, A1=>nx9509, A2=>
      nx10775);
   gen_15_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_15_cmp_mReg_5, QB=>
      nx6639, D=>window_15_5, CLK=>start, R=>rst);
   ix5931 : nor03_2x port map ( Y=>nx5930, A0=>gen_15_cmp_mReg_5, A1=>
      nx10089, A2=>nx10783);
   ix5967 : nand02 port map ( Y=>gen_15_cmp_BSCmp_op2_6, A0=>nx6645, A1=>
      nx6651);
   ix6646 : nor02_2x port map ( Y=>nx6645, A0=>nx5962, A1=>nx5958);
   ix5963 : nor03_2x port map ( Y=>nx5962, A0=>gen_15_cmp_mReg_5, A1=>nx9515, 
      A2=>nx10751);
   ix5959 : nor03_2x port map ( Y=>nx5958, A0=>nx6639, A1=>nx10757, A2=>
      nx10767);
   ix6652 : nor02_2x port map ( Y=>nx6651, A0=>nx5954, A1=>nx5952);
   ix5955 : nor03_2x port map ( Y=>nx5954, A0=>nx6654, A1=>nx9509, A2=>
      nx10775);
   gen_15_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_15_cmp_mReg_6, QB=>
      nx6654, D=>window_15_6, CLK=>start, R=>rst);
   ix5953 : nor03_2x port map ( Y=>nx5952, A0=>gen_15_cmp_mReg_6, A1=>
      nx10089, A2=>nx10783);
   ix5989 : nand02 port map ( Y=>gen_15_cmp_BSCmp_op2_7, A0=>nx6659, A1=>
      nx6665);
   ix6660 : nor02_2x port map ( Y=>nx6659, A0=>nx5984, A1=>nx5980);
   ix5985 : nor03_2x port map ( Y=>nx5984, A0=>gen_15_cmp_mReg_6, A1=>nx9515, 
      A2=>nx10753);
   ix5981 : nor03_2x port map ( Y=>nx5980, A0=>nx6654, A1=>nx10759, A2=>
      nx10769);
   ix6666 : nor02_2x port map ( Y=>nx6665, A0=>nx5976, A1=>nx5974);
   ix5977 : nor03_2x port map ( Y=>nx5976, A0=>nx6669, A1=>nx9509, A2=>
      nx10777);
   gen_15_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_15_cmp_mReg_7, QB=>
      nx6669, D=>window_15_7, CLK=>start, R=>rst);
   ix5975 : nor03_2x port map ( Y=>nx5974, A0=>gen_15_cmp_mReg_7, A1=>
      nx10089, A2=>nx10785);
   ix6011 : nand02 port map ( Y=>gen_15_cmp_BSCmp_op2_8, A0=>nx6675, A1=>
      nx6679);
   ix6676 : nor02_2x port map ( Y=>nx6675, A0=>nx6006, A1=>nx6002);
   ix6007 : nor03_2x port map ( Y=>nx6006, A0=>gen_15_cmp_mReg_7, A1=>nx9515, 
      A2=>nx10753);
   ix6003 : nor03_2x port map ( Y=>nx6002, A0=>nx6669, A1=>nx10759, A2=>
      nx10769);
   ix6680 : nor02_2x port map ( Y=>nx6679, A0=>nx5998, A1=>nx5996);
   ix5999 : nor03_2x port map ( Y=>nx5998, A0=>nx6683, A1=>nx9509, A2=>
      nx10777);
   gen_15_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_15_cmp_mReg_8, QB=>
      nx6683, D=>window_15_8, CLK=>start, R=>rst);
   ix5997 : nor03_2x port map ( Y=>nx5996, A0=>gen_15_cmp_mReg_8, A1=>
      nx10091, A2=>nx10785);
   ix6033 : nand02 port map ( Y=>gen_15_cmp_BSCmp_op2_9, A0=>nx6689, A1=>
      nx6695);
   ix6690 : nor02_2x port map ( Y=>nx6689, A0=>nx6028, A1=>nx6024);
   ix6029 : nor03_2x port map ( Y=>nx6028, A0=>gen_15_cmp_mReg_8, A1=>nx9515, 
      A2=>nx10753);
   ix6025 : nor03_2x port map ( Y=>nx6024, A0=>nx6683, A1=>nx10759, A2=>
      nx10769);
   ix6696 : nor02_2x port map ( Y=>nx6695, A0=>nx6020, A1=>nx6018);
   ix6021 : nor03_2x port map ( Y=>nx6020, A0=>nx6698, A1=>nx9509, A2=>
      nx10777);
   gen_15_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_15_cmp_mReg_9, QB=>
      nx6698, D=>window_15_9, CLK=>start, R=>rst);
   ix6019 : nor03_2x port map ( Y=>nx6018, A0=>gen_15_cmp_mReg_9, A1=>
      nx10091, A2=>nx10785);
   ix6055 : nand02 port map ( Y=>gen_15_cmp_BSCmp_op2_10, A0=>nx6703, A1=>
      nx6709);
   ix6704 : nor02_2x port map ( Y=>nx6703, A0=>nx6050, A1=>nx6046);
   ix6051 : nor03_2x port map ( Y=>nx6050, A0=>gen_15_cmp_mReg_9, A1=>nx9515, 
      A2=>nx10753);
   ix6047 : nor03_2x port map ( Y=>nx6046, A0=>nx6698, A1=>nx10759, A2=>
      nx10769);
   ix6710 : nor02_2x port map ( Y=>nx6709, A0=>nx6042, A1=>nx6040);
   ix6043 : nor03_2x port map ( Y=>nx6042, A0=>nx6713, A1=>nx9509, A2=>
      nx10777);
   gen_15_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_15_cmp_mReg_10, QB=>
      nx6713, D=>window_15_10, CLK=>start, R=>rst);
   ix6041 : nor03_2x port map ( Y=>nx6040, A0=>gen_15_cmp_mReg_10, A1=>
      nx10091, A2=>nx10785);
   ix6077 : nand02 port map ( Y=>gen_15_cmp_BSCmp_op2_11, A0=>nx6719, A1=>
      nx6723);
   ix6720 : nor02_2x port map ( Y=>nx6719, A0=>nx6072, A1=>nx6068);
   ix6073 : nor03_2x port map ( Y=>nx6072, A0=>gen_15_cmp_mReg_10, A1=>
      nx9515, A2=>nx10753);
   ix6069 : nor03_2x port map ( Y=>nx6068, A0=>nx6713, A1=>nx10759, A2=>
      nx10769);
   ix6724 : nor02_2x port map ( Y=>nx6723, A0=>nx6064, A1=>nx6062);
   ix6065 : nor03_2x port map ( Y=>nx6064, A0=>nx6727, A1=>nx9509, A2=>
      nx10777);
   gen_15_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_15_cmp_mReg_11, QB=>
      nx6727, D=>window_15_11, CLK=>start, R=>rst);
   ix6063 : nor03_2x port map ( Y=>nx6062, A0=>gen_15_cmp_mReg_11, A1=>
      nx10091, A2=>nx10785);
   ix6099 : nand02 port map ( Y=>gen_15_cmp_BSCmp_op2_12, A0=>nx6733, A1=>
      nx6739);
   ix6734 : nor02_2x port map ( Y=>nx6733, A0=>nx6094, A1=>nx6090);
   ix6095 : nor03_2x port map ( Y=>nx6094, A0=>gen_15_cmp_mReg_11, A1=>
      nx9515, A2=>nx10753);
   ix6091 : nor03_2x port map ( Y=>nx6090, A0=>nx6727, A1=>nx10759, A2=>
      nx10769);
   ix6740 : nor02_2x port map ( Y=>nx6739, A0=>nx6086, A1=>nx6084);
   ix6087 : nor03_2x port map ( Y=>nx6086, A0=>nx6742, A1=>nx9511, A2=>
      nx10777);
   gen_15_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_15_cmp_mReg_12, QB=>
      nx6742, D=>window_15_12, CLK=>start, R=>rst);
   ix6085 : nor03_2x port map ( Y=>nx6084, A0=>gen_15_cmp_mReg_12, A1=>
      nx10091, A2=>nx10785);
   ix6121 : nand02 port map ( Y=>gen_15_cmp_BSCmp_op2_13, A0=>nx6747, A1=>
      nx6753);
   ix6748 : nor02_2x port map ( Y=>nx6747, A0=>nx6116, A1=>nx6112);
   ix6117 : nor03_2x port map ( Y=>nx6116, A0=>gen_15_cmp_mReg_12, A1=>
      nx9517, A2=>nx10755);
   ix6113 : nor03_2x port map ( Y=>nx6112, A0=>nx6742, A1=>nx10759, A2=>
      nx10771);
   ix6754 : nor02_2x port map ( Y=>nx6753, A0=>nx6108, A1=>nx6106);
   ix6109 : nor03_2x port map ( Y=>nx6108, A0=>nx6757, A1=>nx9511, A2=>
      nx10779);
   gen_15_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_15_cmp_mReg_13, QB=>
      nx6757, D=>window_15_13, CLK=>start, R=>rst);
   ix6107 : nor03_2x port map ( Y=>nx6106, A0=>gen_15_cmp_mReg_13, A1=>
      nx10091, A2=>nx10787);
   ix6143 : nand02 port map ( Y=>gen_15_cmp_BSCmp_op2_14, A0=>nx6763, A1=>
      nx6767);
   ix6764 : nor02_2x port map ( Y=>nx6763, A0=>nx6138, A1=>nx6134);
   ix6139 : nor03_2x port map ( Y=>nx6138, A0=>gen_15_cmp_mReg_13, A1=>
      nx9517, A2=>nx10755);
   ix6135 : nor03_2x port map ( Y=>nx6134, A0=>nx6757, A1=>nx10761, A2=>
      nx10771);
   ix6768 : nor02_2x port map ( Y=>nx6767, A0=>nx6130, A1=>nx6128);
   ix6131 : nor03_2x port map ( Y=>nx6130, A0=>nx6771, A1=>nx9511, A2=>
      nx10779);
   gen_15_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_15_cmp_mReg_14, QB=>
      nx6771, D=>window_15_14, CLK=>start, R=>rst);
   ix6129 : nor03_2x port map ( Y=>nx6128, A0=>gen_15_cmp_mReg_14, A1=>
      nx10091, A2=>nx10787);
   ix6165 : nand02 port map ( Y=>gen_15_cmp_BSCmp_op2_15, A0=>nx6777, A1=>
      nx6783);
   ix6778 : nor02_2x port map ( Y=>nx6777, A0=>nx6160, A1=>nx6156);
   ix6161 : nor03_2x port map ( Y=>nx6160, A0=>gen_15_cmp_mReg_14, A1=>
      nx9517, A2=>nx10755);
   ix6157 : nor03_2x port map ( Y=>nx6156, A0=>nx6771, A1=>nx10761, A2=>
      nx10771);
   ix6784 : nor02_2x port map ( Y=>nx6783, A0=>nx6152, A1=>nx6150);
   ix6153 : nor03_2x port map ( Y=>nx6152, A0=>nx6786, A1=>nx9511, A2=>
      nx10779);
   gen_15_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_15_cmp_mReg_15, QB=>
      nx6786, D=>window_15_15, CLK=>start, R=>rst);
   ix6151 : nor03_2x port map ( Y=>nx6150, A0=>gen_15_cmp_mReg_15, A1=>
      nx10093, A2=>nx10787);
   ix6175 : nand02 port map ( Y=>gen_15_cmp_BSCmp_op2_16, A0=>nx6791, A1=>
      nx6783);
   ix6792 : nor02_2x port map ( Y=>nx6791, A0=>nx6170, A1=>nx6166);
   ix6171 : nor03_2x port map ( Y=>nx6170, A0=>gen_15_cmp_mReg_15, A1=>
      nx9517, A2=>nx10755);
   ix6167 : nor03_2x port map ( Y=>nx6166, A0=>nx6786, A1=>nx10761, A2=>
      nx10771);
   ix6243 : nand02 port map ( Y=>gen_16_cmp_BSCmp_op2_1, A0=>nx6799, A1=>
      nx6817);
   ix6800 : nor02_2x port map ( Y=>nx6799, A0=>nx6238, A1=>nx6234);
   ix6239 : nor03_2x port map ( Y=>nx6238, A0=>gen_16_cmp_mReg_0, A1=>nx9501, 
      A2=>nx10791);
   gen_16_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_16_cmp_mReg_0, QB=>
      nx6805, D=>window_16_0, CLK=>start, R=>rst);
   ix6809 : inv01 port map ( Y=>nx6808, A=>gen_16_cmp_pMux_0);
   ix6235 : nor03_2x port map ( Y=>nx6234, A0=>nx6805, A1=>nx10797, A2=>
      nx10807);
   ix6816 : inv02 port map ( Y=>nx6815, A=>gen_16_cmp_pMux_2);
   ix6818 : nor02_2x port map ( Y=>nx6817, A0=>nx6224, A1=>nx6222);
   ix6225 : nor03_2x port map ( Y=>nx6224, A0=>nx6821, A1=>nx9495, A2=>
      nx10815);
   gen_16_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_16_cmp_mReg_1, QB=>
      nx6821, D=>window_16_1, CLK=>start, R=>rst);
   ix6223 : nor03_2x port map ( Y=>nx6222, A0=>gen_16_cmp_mReg_1, A1=>
      nx10095, A2=>nx10823);
   ix6183 : nor03_2x port map ( Y=>nx6182, A0=>nx9501, A1=>nx6815, A2=>
      gen_16_cmp_pMux_0);
   ix6265 : nand02 port map ( Y=>gen_16_cmp_BSCmp_op2_2, A0=>nx6832, A1=>
      nx6839);
   ix6834 : nor02_2x port map ( Y=>nx6832, A0=>nx6260, A1=>nx6256);
   ix6261 : nor03_2x port map ( Y=>nx6260, A0=>gen_16_cmp_mReg_1, A1=>nx9501, 
      A2=>nx10791);
   ix6257 : nor03_2x port map ( Y=>nx6256, A0=>nx6821, A1=>nx10797, A2=>
      nx10807);
   ix6840 : nor02_2x port map ( Y=>nx6839, A0=>nx6252, A1=>nx6250);
   ix6253 : nor03_2x port map ( Y=>nx6252, A0=>nx6843, A1=>nx9495, A2=>
      nx10815);
   gen_16_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_16_cmp_mReg_2, QB=>
      nx6843, D=>window_16_2, CLK=>start, R=>rst);
   ix6251 : nor03_2x port map ( Y=>nx6250, A0=>gen_16_cmp_mReg_2, A1=>
      nx10095, A2=>nx10823);
   ix6287 : nand02 port map ( Y=>gen_16_cmp_BSCmp_op2_3, A0=>nx6849, A1=>
      nx6853);
   ix6850 : nor02_2x port map ( Y=>nx6849, A0=>nx6282, A1=>nx6278);
   ix6283 : nor03_2x port map ( Y=>nx6282, A0=>gen_16_cmp_mReg_2, A1=>nx9501, 
      A2=>nx10791);
   ix6279 : nor03_2x port map ( Y=>nx6278, A0=>nx6843, A1=>nx10797, A2=>
      nx10807);
   ix6854 : nor02_2x port map ( Y=>nx6853, A0=>nx6274, A1=>nx6272);
   ix6275 : nor03_2x port map ( Y=>nx6274, A0=>nx6857, A1=>nx9495, A2=>
      nx10815);
   gen_16_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_16_cmp_mReg_3, QB=>
      nx6857, D=>window_16_3, CLK=>start, R=>rst);
   ix6273 : nor03_2x port map ( Y=>nx6272, A0=>gen_16_cmp_mReg_3, A1=>
      nx10095, A2=>nx10823);
   ix6309 : nand02 port map ( Y=>gen_16_cmp_BSCmp_op2_4, A0=>nx6863, A1=>
      nx6867);
   ix6864 : nor02_2x port map ( Y=>nx6863, A0=>nx6304, A1=>nx6300);
   ix6305 : nor03_2x port map ( Y=>nx6304, A0=>gen_16_cmp_mReg_3, A1=>nx9501, 
      A2=>nx10791);
   ix6301 : nor03_2x port map ( Y=>nx6300, A0=>nx6857, A1=>nx10797, A2=>
      nx10807);
   ix6868 : nor02_2x port map ( Y=>nx6867, A0=>nx6296, A1=>nx6294);
   ix6297 : nor03_2x port map ( Y=>nx6296, A0=>nx6871, A1=>nx9495, A2=>
      nx10815);
   gen_16_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_16_cmp_mReg_4, QB=>
      nx6871, D=>window_16_4, CLK=>start, R=>rst);
   ix6295 : nor03_2x port map ( Y=>nx6294, A0=>gen_16_cmp_mReg_4, A1=>
      nx10095, A2=>nx10823);
   ix6331 : nand02 port map ( Y=>gen_16_cmp_BSCmp_op2_5, A0=>nx6875, A1=>
      nx6881);
   ix6876 : nor02_2x port map ( Y=>nx6875, A0=>nx6326, A1=>nx6322);
   ix6327 : nor03_2x port map ( Y=>nx6326, A0=>gen_16_cmp_mReg_4, A1=>nx9501, 
      A2=>nx10791);
   ix6323 : nor03_2x port map ( Y=>nx6322, A0=>nx6871, A1=>nx10797, A2=>
      nx10807);
   ix6882 : nor02_2x port map ( Y=>nx6881, A0=>nx6318, A1=>nx6316);
   ix6319 : nor03_2x port map ( Y=>nx6318, A0=>nx6885, A1=>nx9497, A2=>
      nx10815);
   gen_16_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_16_cmp_mReg_5, QB=>
      nx6885, D=>window_16_5, CLK=>start, R=>rst);
   ix6317 : nor03_2x port map ( Y=>nx6316, A0=>gen_16_cmp_mReg_5, A1=>
      nx10095, A2=>nx10823);
   ix6353 : nand02 port map ( Y=>gen_16_cmp_BSCmp_op2_6, A0=>nx6889, A1=>
      nx6895);
   ix6890 : nor02_2x port map ( Y=>nx6889, A0=>nx6348, A1=>nx6344);
   ix6349 : nor03_2x port map ( Y=>nx6348, A0=>gen_16_cmp_mReg_5, A1=>nx9503, 
      A2=>nx10791);
   ix6345 : nor03_2x port map ( Y=>nx6344, A0=>nx6885, A1=>nx10797, A2=>
      nx10807);
   ix6896 : nor02_2x port map ( Y=>nx6895, A0=>nx6340, A1=>nx6338);
   ix6341 : nor03_2x port map ( Y=>nx6340, A0=>nx6898, A1=>nx9497, A2=>
      nx10815);
   gen_16_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_16_cmp_mReg_6, QB=>
      nx6898, D=>window_16_6, CLK=>start, R=>rst);
   ix6339 : nor03_2x port map ( Y=>nx6338, A0=>gen_16_cmp_mReg_6, A1=>
      nx10095, A2=>nx10823);
   ix6375 : nand02 port map ( Y=>gen_16_cmp_BSCmp_op2_7, A0=>nx6905, A1=>
      nx6911);
   ix6906 : nor02_2x port map ( Y=>nx6905, A0=>nx6370, A1=>nx6366);
   ix6371 : nor03_2x port map ( Y=>nx6370, A0=>gen_16_cmp_mReg_6, A1=>nx9503, 
      A2=>nx10793);
   ix6367 : nor03_2x port map ( Y=>nx6366, A0=>nx6898, A1=>nx10799, A2=>
      nx10809);
   ix6912 : nor02_2x port map ( Y=>nx6911, A0=>nx6362, A1=>nx6360);
   ix6363 : nor03_2x port map ( Y=>nx6362, A0=>nx6915, A1=>nx9497, A2=>
      nx10817);
   gen_16_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_16_cmp_mReg_7, QB=>
      nx6915, D=>window_16_7, CLK=>start, R=>rst);
   ix6361 : nor03_2x port map ( Y=>nx6360, A0=>gen_16_cmp_mReg_7, A1=>
      nx10095, A2=>nx10825);
   ix6397 : nand02 port map ( Y=>gen_16_cmp_BSCmp_op2_8, A0=>nx6919, A1=>
      nx6925);
   ix6920 : nor02_2x port map ( Y=>nx6919, A0=>nx6392, A1=>nx6388);
   ix6393 : nor03_2x port map ( Y=>nx6392, A0=>gen_16_cmp_mReg_7, A1=>nx9503, 
      A2=>nx10793);
   ix6389 : nor03_2x port map ( Y=>nx6388, A0=>nx6915, A1=>nx10799, A2=>
      nx10809);
   ix6926 : nor02_2x port map ( Y=>nx6925, A0=>nx6384, A1=>nx6382);
   ix6385 : nor03_2x port map ( Y=>nx6384, A0=>nx6929, A1=>nx9497, A2=>
      nx10817);
   gen_16_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_16_cmp_mReg_8, QB=>
      nx6929, D=>window_16_8, CLK=>start, R=>rst);
   ix6383 : nor03_2x port map ( Y=>nx6382, A0=>gen_16_cmp_mReg_8, A1=>
      nx10097, A2=>nx10825);
   ix6419 : nand02 port map ( Y=>gen_16_cmp_BSCmp_op2_9, A0=>nx6933, A1=>
      nx6939);
   ix6934 : nor02_2x port map ( Y=>nx6933, A0=>nx6414, A1=>nx6410);
   ix6415 : nor03_2x port map ( Y=>nx6414, A0=>gen_16_cmp_mReg_8, A1=>nx9503, 
      A2=>nx10793);
   ix6411 : nor03_2x port map ( Y=>nx6410, A0=>nx6929, A1=>nx10799, A2=>
      nx10809);
   ix6940 : nor02_2x port map ( Y=>nx6939, A0=>nx6406, A1=>nx6404);
   ix6407 : nor03_2x port map ( Y=>nx6406, A0=>nx6943, A1=>nx9497, A2=>
      nx10817);
   gen_16_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_16_cmp_mReg_9, QB=>
      nx6943, D=>window_16_9, CLK=>start, R=>rst);
   ix6405 : nor03_2x port map ( Y=>nx6404, A0=>gen_16_cmp_mReg_9, A1=>
      nx10097, A2=>nx10825);
   ix6441 : nand02 port map ( Y=>gen_16_cmp_BSCmp_op2_10, A0=>nx6949, A1=>
      nx6955);
   ix6950 : nor02_2x port map ( Y=>nx6949, A0=>nx6436, A1=>nx6432);
   ix6437 : nor03_2x port map ( Y=>nx6436, A0=>gen_16_cmp_mReg_9, A1=>nx9503, 
      A2=>nx10793);
   ix6433 : nor03_2x port map ( Y=>nx6432, A0=>nx6943, A1=>nx10799, A2=>
      nx10809);
   ix6956 : nor02_2x port map ( Y=>nx6955, A0=>nx6428, A1=>nx6426);
   ix6429 : nor03_2x port map ( Y=>nx6428, A0=>nx6958, A1=>nx9497, A2=>
      nx10817);
   gen_16_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_16_cmp_mReg_10, QB=>
      nx6958, D=>window_16_10, CLK=>start, R=>rst);
   ix6427 : nor03_2x port map ( Y=>nx6426, A0=>gen_16_cmp_mReg_10, A1=>
      nx10097, A2=>nx10825);
   ix6463 : nand02 port map ( Y=>gen_16_cmp_BSCmp_op2_11, A0=>nx6962, A1=>
      nx6967);
   ix6963 : nor02_2x port map ( Y=>nx6962, A0=>nx6458, A1=>nx6454);
   ix6459 : nor03_2x port map ( Y=>nx6458, A0=>gen_16_cmp_mReg_10, A1=>
      nx9503, A2=>nx10793);
   ix6455 : nor03_2x port map ( Y=>nx6454, A0=>nx6958, A1=>nx10799, A2=>
      nx10809);
   ix6968 : nor02_2x port map ( Y=>nx6967, A0=>nx6450, A1=>nx6448);
   ix6451 : nor03_2x port map ( Y=>nx6450, A0=>nx6971, A1=>nx9497, A2=>
      nx10817);
   gen_16_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_16_cmp_mReg_11, QB=>
      nx6971, D=>window_16_11, CLK=>start, R=>rst);
   ix6449 : nor03_2x port map ( Y=>nx6448, A0=>gen_16_cmp_mReg_11, A1=>
      nx10097, A2=>nx10825);
   ix6485 : nand02 port map ( Y=>gen_16_cmp_BSCmp_op2_12, A0=>nx6977, A1=>
      nx6983);
   ix6978 : nor02_2x port map ( Y=>nx6977, A0=>nx6480, A1=>nx6476);
   ix6481 : nor03_2x port map ( Y=>nx6480, A0=>gen_16_cmp_mReg_11, A1=>
      nx9503, A2=>nx10793);
   ix6477 : nor03_2x port map ( Y=>nx6476, A0=>nx6971, A1=>nx10799, A2=>
      nx10809);
   ix6984 : nor02_2x port map ( Y=>nx6983, A0=>nx6472, A1=>nx6470);
   ix6473 : nor03_2x port map ( Y=>nx6472, A0=>nx6987, A1=>nx9499, A2=>
      nx10817);
   gen_16_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_16_cmp_mReg_12, QB=>
      nx6987, D=>window_16_12, CLK=>start, R=>rst);
   ix6471 : nor03_2x port map ( Y=>nx6470, A0=>gen_16_cmp_mReg_12, A1=>
      nx10097, A2=>nx10825);
   ix6507 : nand02 port map ( Y=>gen_16_cmp_BSCmp_op2_13, A0=>nx6991, A1=>
      nx6997);
   ix6992 : nor02_2x port map ( Y=>nx6991, A0=>nx6502, A1=>nx6498);
   ix6503 : nor03_2x port map ( Y=>nx6502, A0=>gen_16_cmp_mReg_12, A1=>
      nx9505, A2=>nx10795);
   ix6499 : nor03_2x port map ( Y=>nx6498, A0=>nx6987, A1=>nx10799, A2=>
      nx10811);
   ix6998 : nor02_2x port map ( Y=>nx6997, A0=>nx6494, A1=>nx6492);
   ix6495 : nor03_2x port map ( Y=>nx6494, A0=>nx7001, A1=>nx9499, A2=>
      nx10819);
   gen_16_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_16_cmp_mReg_13, QB=>
      nx7001, D=>window_16_13, CLK=>start, R=>rst);
   ix6493 : nor03_2x port map ( Y=>nx6492, A0=>gen_16_cmp_mReg_13, A1=>
      nx10097, A2=>nx10827);
   ix6529 : nand02 port map ( Y=>gen_16_cmp_BSCmp_op2_14, A0=>nx7007, A1=>
      nx7011);
   ix7008 : nor02_2x port map ( Y=>nx7007, A0=>nx6524, A1=>nx6520);
   ix6525 : nor03_2x port map ( Y=>nx6524, A0=>gen_16_cmp_mReg_13, A1=>
      nx9505, A2=>nx10795);
   ix6521 : nor03_2x port map ( Y=>nx6520, A0=>nx7001, A1=>nx10801, A2=>
      nx10811);
   ix7012 : nor02_2x port map ( Y=>nx7011, A0=>nx6516, A1=>nx6514);
   ix6517 : nor03_2x port map ( Y=>nx6516, A0=>nx7015, A1=>nx9499, A2=>
      nx10819);
   gen_16_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_16_cmp_mReg_14, QB=>
      nx7015, D=>window_16_14, CLK=>start, R=>rst);
   ix6515 : nor03_2x port map ( Y=>nx6514, A0=>gen_16_cmp_mReg_14, A1=>
      nx10097, A2=>nx10827);
   ix6551 : nand02 port map ( Y=>gen_16_cmp_BSCmp_op2_15, A0=>nx7019, A1=>
      nx7025);
   ix7020 : nor02_2x port map ( Y=>nx7019, A0=>nx6546, A1=>nx6542);
   ix6547 : nor03_2x port map ( Y=>nx6546, A0=>gen_16_cmp_mReg_14, A1=>
      nx9505, A2=>nx10795);
   ix6543 : nor03_2x port map ( Y=>nx6542, A0=>nx7015, A1=>nx10801, A2=>
      nx10811);
   ix7026 : nor02_2x port map ( Y=>nx7025, A0=>nx6538, A1=>nx6536);
   ix6539 : nor03_2x port map ( Y=>nx6538, A0=>nx7029, A1=>nx9499, A2=>
      nx10819);
   gen_16_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_16_cmp_mReg_15, QB=>
      nx7029, D=>window_16_15, CLK=>start, R=>rst);
   ix6537 : nor03_2x port map ( Y=>nx6536, A0=>gen_16_cmp_mReg_15, A1=>
      nx10099, A2=>nx10827);
   ix6561 : nand02 port map ( Y=>gen_16_cmp_BSCmp_op2_16, A0=>nx7033, A1=>
      nx7025);
   ix7034 : nor02_2x port map ( Y=>nx7033, A0=>nx6556, A1=>nx6552);
   ix6557 : nor03_2x port map ( Y=>nx6556, A0=>gen_16_cmp_mReg_15, A1=>
      nx9505, A2=>nx10795);
   ix6553 : nor03_2x port map ( Y=>nx6552, A0=>nx7029, A1=>nx10801, A2=>
      nx10811);
   ix6629 : nand02 port map ( Y=>gen_17_cmp_BSCmp_op2_1, A0=>nx7040, A1=>
      nx7059);
   ix7041 : nor02_2x port map ( Y=>nx7040, A0=>nx6624, A1=>nx6620);
   ix6625 : nor03_2x port map ( Y=>nx6624, A0=>gen_17_cmp_mReg_0, A1=>nx9489, 
      A2=>nx10831);
   gen_17_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_17_cmp_mReg_0, QB=>
      nx7045, D=>window_17_0, CLK=>start, R=>rst);
   ix7050 : inv01 port map ( Y=>nx7049, A=>gen_17_cmp_pMux_0);
   ix6621 : nor03_2x port map ( Y=>nx6620, A0=>nx7045, A1=>nx10837, A2=>
      nx10847);
   ix7058 : inv02 port map ( Y=>nx7057, A=>gen_17_cmp_pMux_2);
   ix7060 : nor02_2x port map ( Y=>nx7059, A0=>nx6610, A1=>nx6608);
   ix6611 : nor03_2x port map ( Y=>nx6610, A0=>nx7062, A1=>nx9483, A2=>
      nx10855);
   gen_17_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_17_cmp_mReg_1, QB=>
      nx7062, D=>window_17_1, CLK=>start, R=>rst);
   ix6609 : nor03_2x port map ( Y=>nx6608, A0=>gen_17_cmp_mReg_1, A1=>
      nx10101, A2=>nx10863);
   ix6569 : nor03_2x port map ( Y=>nx6568, A0=>nx9489, A1=>nx7057, A2=>
      gen_17_cmp_pMux_0);
   ix6651 : nand02 port map ( Y=>gen_17_cmp_BSCmp_op2_2, A0=>nx7075, A1=>
      nx7081);
   ix7076 : nor02_2x port map ( Y=>nx7075, A0=>nx6646, A1=>nx6642);
   ix6647 : nor03_2x port map ( Y=>nx6646, A0=>gen_17_cmp_mReg_1, A1=>nx9489, 
      A2=>nx10831);
   ix6643 : nor03_2x port map ( Y=>nx6642, A0=>nx7062, A1=>nx10837, A2=>
      nx10847);
   ix7082 : nor02_2x port map ( Y=>nx7081, A0=>nx6638, A1=>nx6636);
   ix6639 : nor03_2x port map ( Y=>nx6638, A0=>nx7084, A1=>nx9483, A2=>
      nx10855);
   gen_17_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_17_cmp_mReg_2, QB=>
      nx7084, D=>window_17_2, CLK=>start, R=>rst);
   ix6637 : nor03_2x port map ( Y=>nx6636, A0=>gen_17_cmp_mReg_2, A1=>
      nx10101, A2=>nx10863);
   ix6673 : nand02 port map ( Y=>gen_17_cmp_BSCmp_op2_3, A0=>nx7089, A1=>
      nx7095);
   ix7090 : nor02_2x port map ( Y=>nx7089, A0=>nx6668, A1=>nx6664);
   ix6669 : nor03_2x port map ( Y=>nx6668, A0=>gen_17_cmp_mReg_2, A1=>nx9489, 
      A2=>nx10831);
   ix6665 : nor03_2x port map ( Y=>nx6664, A0=>nx7084, A1=>nx10837, A2=>
      nx10847);
   ix7096 : nor02_2x port map ( Y=>nx7095, A0=>nx6660, A1=>nx6658);
   ix6661 : nor03_2x port map ( Y=>nx6660, A0=>nx7099, A1=>nx9483, A2=>
      nx10855);
   gen_17_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_17_cmp_mReg_3, QB=>
      nx7099, D=>window_17_3, CLK=>start, R=>rst);
   ix6659 : nor03_2x port map ( Y=>nx6658, A0=>gen_17_cmp_mReg_3, A1=>
      nx10101, A2=>nx10863);
   ix6695 : nand02 port map ( Y=>gen_17_cmp_BSCmp_op2_4, A0=>nx7105, A1=>
      nx7109);
   ix7106 : nor02_2x port map ( Y=>nx7105, A0=>nx6690, A1=>nx6686);
   ix6691 : nor03_2x port map ( Y=>nx6690, A0=>gen_17_cmp_mReg_3, A1=>nx9489, 
      A2=>nx10831);
   ix6687 : nor03_2x port map ( Y=>nx6686, A0=>nx7099, A1=>nx10837, A2=>
      nx10847);
   ix7110 : nor02_2x port map ( Y=>nx7109, A0=>nx6682, A1=>nx6680);
   ix6683 : nor03_2x port map ( Y=>nx6682, A0=>nx7113, A1=>nx9483, A2=>
      nx10855);
   gen_17_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_17_cmp_mReg_4, QB=>
      nx7113, D=>window_17_4, CLK=>start, R=>rst);
   ix6681 : nor03_2x port map ( Y=>nx6680, A0=>gen_17_cmp_mReg_4, A1=>
      nx10101, A2=>nx10863);
   ix6717 : nand02 port map ( Y=>gen_17_cmp_BSCmp_op2_5, A0=>nx7119, A1=>
      nx7125);
   ix7120 : nor02_2x port map ( Y=>nx7119, A0=>nx6712, A1=>nx6708);
   ix6713 : nor03_2x port map ( Y=>nx6712, A0=>gen_17_cmp_mReg_4, A1=>nx9489, 
      A2=>nx10831);
   ix6709 : nor03_2x port map ( Y=>nx6708, A0=>nx7113, A1=>nx10837, A2=>
      nx10847);
   ix7126 : nor02_2x port map ( Y=>nx7125, A0=>nx6704, A1=>nx6702);
   ix6705 : nor03_2x port map ( Y=>nx6704, A0=>nx7128, A1=>nx9485, A2=>
      nx10855);
   gen_17_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_17_cmp_mReg_5, QB=>
      nx7128, D=>window_17_5, CLK=>start, R=>rst);
   ix6703 : nor03_2x port map ( Y=>nx6702, A0=>gen_17_cmp_mReg_5, A1=>
      nx10101, A2=>nx10863);
   ix6739 : nand02 port map ( Y=>gen_17_cmp_BSCmp_op2_6, A0=>nx7133, A1=>
      nx7139);
   ix7134 : nor02_2x port map ( Y=>nx7133, A0=>nx6734, A1=>nx6730);
   ix6735 : nor03_2x port map ( Y=>nx6734, A0=>gen_17_cmp_mReg_5, A1=>nx9491, 
      A2=>nx10831);
   ix6731 : nor03_2x port map ( Y=>nx6730, A0=>nx7128, A1=>nx10837, A2=>
      nx10847);
   ix7140 : nor02_2x port map ( Y=>nx7139, A0=>nx6726, A1=>nx6724);
   ix6727 : nor03_2x port map ( Y=>nx6726, A0=>nx7143, A1=>nx9485, A2=>
      nx10855);
   gen_17_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_17_cmp_mReg_6, QB=>
      nx7143, D=>window_17_6, CLK=>start, R=>rst);
   ix6725 : nor03_2x port map ( Y=>nx6724, A0=>gen_17_cmp_mReg_6, A1=>
      nx10101, A2=>nx10863);
   ix6761 : nand02 port map ( Y=>gen_17_cmp_BSCmp_op2_7, A0=>nx7149, A1=>
      nx7153);
   ix7150 : nor02_2x port map ( Y=>nx7149, A0=>nx6756, A1=>nx6752);
   ix6757 : nor03_2x port map ( Y=>nx6756, A0=>gen_17_cmp_mReg_6, A1=>nx9491, 
      A2=>nx10833);
   ix6753 : nor03_2x port map ( Y=>nx6752, A0=>nx7143, A1=>nx10839, A2=>
      nx10849);
   ix7154 : nor02_2x port map ( Y=>nx7153, A0=>nx6748, A1=>nx6746);
   ix6749 : nor03_2x port map ( Y=>nx6748, A0=>nx7157, A1=>nx9485, A2=>
      nx10857);
   gen_17_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_17_cmp_mReg_7, QB=>
      nx7157, D=>window_17_7, CLK=>start, R=>rst);
   ix6747 : nor03_2x port map ( Y=>nx6746, A0=>gen_17_cmp_mReg_7, A1=>
      nx10101, A2=>nx10865);
   ix6783 : nand02 port map ( Y=>gen_17_cmp_BSCmp_op2_8, A0=>nx7163, A1=>
      nx7169);
   ix7164 : nor02_2x port map ( Y=>nx7163, A0=>nx6778, A1=>nx6774);
   ix6779 : nor03_2x port map ( Y=>nx6778, A0=>gen_17_cmp_mReg_7, A1=>nx9491, 
      A2=>nx10833);
   ix6775 : nor03_2x port map ( Y=>nx6774, A0=>nx7157, A1=>nx10839, A2=>
      nx10849);
   ix7170 : nor02_2x port map ( Y=>nx7169, A0=>nx6770, A1=>nx6768);
   ix6771 : nor03_2x port map ( Y=>nx6770, A0=>nx7172, A1=>nx9485, A2=>
      nx10857);
   gen_17_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_17_cmp_mReg_8, QB=>
      nx7172, D=>window_17_8, CLK=>start, R=>rst);
   ix6769 : nor03_2x port map ( Y=>nx6768, A0=>gen_17_cmp_mReg_8, A1=>
      nx10103, A2=>nx10865);
   ix6805 : nand02 port map ( Y=>gen_17_cmp_BSCmp_op2_9, A0=>nx7177, A1=>
      nx7183);
   ix7178 : nor02_2x port map ( Y=>nx7177, A0=>nx6800, A1=>nx6796);
   ix6801 : nor03_2x port map ( Y=>nx6800, A0=>gen_17_cmp_mReg_8, A1=>nx9491, 
      A2=>nx10833);
   ix6797 : nor03_2x port map ( Y=>nx6796, A0=>nx7172, A1=>nx10839, A2=>
      nx10849);
   ix7184 : nor02_2x port map ( Y=>nx7183, A0=>nx6792, A1=>nx6790);
   ix6793 : nor03_2x port map ( Y=>nx6792, A0=>nx7187, A1=>nx9485, A2=>
      nx10857);
   gen_17_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_17_cmp_mReg_9, QB=>
      nx7187, D=>window_17_9, CLK=>start, R=>rst);
   ix6791 : nor03_2x port map ( Y=>nx6790, A0=>gen_17_cmp_mReg_9, A1=>
      nx10103, A2=>nx10865);
   ix6827 : nand02 port map ( Y=>gen_17_cmp_BSCmp_op2_10, A0=>nx7193, A1=>
      nx7197);
   ix7194 : nor02_2x port map ( Y=>nx7193, A0=>nx6822, A1=>nx6818);
   ix6823 : nor03_2x port map ( Y=>nx6822, A0=>gen_17_cmp_mReg_9, A1=>nx9491, 
      A2=>nx10833);
   ix6819 : nor03_2x port map ( Y=>nx6818, A0=>nx7187, A1=>nx10839, A2=>
      nx10849);
   ix7198 : nor02_2x port map ( Y=>nx7197, A0=>nx6814, A1=>nx6812);
   ix6815 : nor03_2x port map ( Y=>nx6814, A0=>nx7201, A1=>nx9485, A2=>
      nx10857);
   gen_17_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_17_cmp_mReg_10, QB=>
      nx7201, D=>window_17_10, CLK=>start, R=>rst);
   ix6813 : nor03_2x port map ( Y=>nx6812, A0=>gen_17_cmp_mReg_10, A1=>
      nx10103, A2=>nx10865);
   ix6849 : nand02 port map ( Y=>gen_17_cmp_BSCmp_op2_11, A0=>nx7207, A1=>
      nx7213);
   ix7208 : nor02_2x port map ( Y=>nx7207, A0=>nx6844, A1=>nx6840);
   ix6845 : nor03_2x port map ( Y=>nx6844, A0=>gen_17_cmp_mReg_10, A1=>
      nx9491, A2=>nx10833);
   ix6841 : nor03_2x port map ( Y=>nx6840, A0=>nx7201, A1=>nx10839, A2=>
      nx10849);
   ix7214 : nor02_2x port map ( Y=>nx7213, A0=>nx6836, A1=>nx6834);
   ix6837 : nor03_2x port map ( Y=>nx6836, A0=>nx7216, A1=>nx9485, A2=>
      nx10857);
   gen_17_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_17_cmp_mReg_11, QB=>
      nx7216, D=>window_17_11, CLK=>start, R=>rst);
   ix6835 : nor03_2x port map ( Y=>nx6834, A0=>gen_17_cmp_mReg_11, A1=>
      nx10103, A2=>nx10865);
   ix6871 : nand02 port map ( Y=>gen_17_cmp_BSCmp_op2_12, A0=>nx7221, A1=>
      nx7227);
   ix7222 : nor02_2x port map ( Y=>nx7221, A0=>nx6866, A1=>nx6862);
   ix6867 : nor03_2x port map ( Y=>nx6866, A0=>gen_17_cmp_mReg_11, A1=>
      nx9491, A2=>nx10833);
   ix6863 : nor03_2x port map ( Y=>nx6862, A0=>nx7216, A1=>nx10839, A2=>
      nx10849);
   ix7228 : nor02_2x port map ( Y=>nx7227, A0=>nx6858, A1=>nx6856);
   ix6859 : nor03_2x port map ( Y=>nx6858, A0=>nx7231, A1=>nx9487, A2=>
      nx10857);
   gen_17_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_17_cmp_mReg_12, QB=>
      nx7231, D=>window_17_12, CLK=>start, R=>rst);
   ix6857 : nor03_2x port map ( Y=>nx6856, A0=>gen_17_cmp_mReg_12, A1=>
      nx10103, A2=>nx10865);
   ix6893 : nand02 port map ( Y=>gen_17_cmp_BSCmp_op2_13, A0=>nx7237, A1=>
      nx7241);
   ix7238 : nor02_2x port map ( Y=>nx7237, A0=>nx6888, A1=>nx6884);
   ix6889 : nor03_2x port map ( Y=>nx6888, A0=>gen_17_cmp_mReg_12, A1=>
      nx9493, A2=>nx10835);
   ix6885 : nor03_2x port map ( Y=>nx6884, A0=>nx7231, A1=>nx10839, A2=>
      nx10851);
   ix7242 : nor02_2x port map ( Y=>nx7241, A0=>nx6880, A1=>nx6878);
   ix6881 : nor03_2x port map ( Y=>nx6880, A0=>nx7245, A1=>nx9487, A2=>
      nx10859);
   gen_17_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_17_cmp_mReg_13, QB=>
      nx7245, D=>window_17_13, CLK=>start, R=>rst);
   ix6879 : nor03_2x port map ( Y=>nx6878, A0=>gen_17_cmp_mReg_13, A1=>
      nx10103, A2=>nx10867);
   ix6915 : nand02 port map ( Y=>gen_17_cmp_BSCmp_op2_14, A0=>nx7251, A1=>
      nx7257);
   ix7252 : nor02_2x port map ( Y=>nx7251, A0=>nx6910, A1=>nx6906);
   ix6911 : nor03_2x port map ( Y=>nx6910, A0=>gen_17_cmp_mReg_13, A1=>
      nx9493, A2=>nx10835);
   ix6907 : nor03_2x port map ( Y=>nx6906, A0=>nx7245, A1=>nx10841, A2=>
      nx10851);
   ix7258 : nor02_2x port map ( Y=>nx7257, A0=>nx6902, A1=>nx6900);
   ix6903 : nor03_2x port map ( Y=>nx6902, A0=>nx7260, A1=>nx9487, A2=>
      nx10859);
   gen_17_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_17_cmp_mReg_14, QB=>
      nx7260, D=>window_17_14, CLK=>start, R=>rst);
   ix6901 : nor03_2x port map ( Y=>nx6900, A0=>gen_17_cmp_mReg_14, A1=>
      nx10103, A2=>nx10867);
   ix6937 : nand02 port map ( Y=>gen_17_cmp_BSCmp_op2_15, A0=>nx7265, A1=>
      nx7271);
   ix7266 : nor02_2x port map ( Y=>nx7265, A0=>nx6932, A1=>nx6928);
   ix6933 : nor03_2x port map ( Y=>nx6932, A0=>gen_17_cmp_mReg_14, A1=>
      nx9493, A2=>nx10835);
   ix6929 : nor03_2x port map ( Y=>nx6928, A0=>nx7260, A1=>nx10841, A2=>
      nx10851);
   ix7272 : nor02_2x port map ( Y=>nx7271, A0=>nx6924, A1=>nx6922);
   ix6925 : nor03_2x port map ( Y=>nx6924, A0=>nx7275, A1=>nx9487, A2=>
      nx10859);
   gen_17_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_17_cmp_mReg_15, QB=>
      nx7275, D=>window_17_15, CLK=>start, R=>rst);
   ix6923 : nor03_2x port map ( Y=>nx6922, A0=>gen_17_cmp_mReg_15, A1=>
      nx10105, A2=>nx10867);
   ix6947 : nand02 port map ( Y=>gen_17_cmp_BSCmp_op2_16, A0=>nx7281, A1=>
      nx7271);
   ix7282 : nor02_2x port map ( Y=>nx7281, A0=>nx6942, A1=>nx6938);
   ix6943 : nor03_2x port map ( Y=>nx6942, A0=>gen_17_cmp_mReg_15, A1=>
      nx9493, A2=>nx10835);
   ix6939 : nor03_2x port map ( Y=>nx6938, A0=>nx7275, A1=>nx10841, A2=>
      nx10851);
   ix7015 : nand02 port map ( Y=>gen_18_cmp_BSCmp_op2_1, A0=>nx7287, A1=>
      nx7307);
   ix7288 : nor02_2x port map ( Y=>nx7287, A0=>nx7010, A1=>nx7006);
   ix7011 : nor03_2x port map ( Y=>nx7010, A0=>gen_18_cmp_mReg_0, A1=>nx9477, 
      A2=>nx10871);
   gen_18_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_18_cmp_mReg_0, QB=>
      nx7293, D=>window_18_0, CLK=>start, R=>rst);
   ix7298 : inv01 port map ( Y=>nx7297, A=>gen_18_cmp_pMux_0);
   ix7007 : nor03_2x port map ( Y=>nx7006, A0=>nx7293, A1=>nx10877, A2=>
      nx10887);
   ix7306 : inv02 port map ( Y=>nx7305, A=>gen_18_cmp_pMux_2);
   ix7308 : nor02_2x port map ( Y=>nx7307, A0=>nx6996, A1=>nx6994);
   ix6997 : nor03_2x port map ( Y=>nx6996, A0=>nx7311, A1=>nx9471, A2=>
      nx10895);
   gen_18_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_18_cmp_mReg_1, QB=>
      nx7311, D=>window_18_1, CLK=>start, R=>rst);
   ix6995 : nor03_2x port map ( Y=>nx6994, A0=>gen_18_cmp_mReg_1, A1=>
      nx10107, A2=>nx10903);
   ix6955 : nor03_2x port map ( Y=>nx6954, A0=>nx9477, A1=>nx7305, A2=>
      gen_18_cmp_pMux_0);
   ix7037 : nand02 port map ( Y=>gen_18_cmp_BSCmp_op2_2, A0=>nx7323, A1=>
      nx7329);
   ix7324 : nor02_2x port map ( Y=>nx7323, A0=>nx7032, A1=>nx7028);
   ix7033 : nor03_2x port map ( Y=>nx7032, A0=>gen_18_cmp_mReg_1, A1=>nx9477, 
      A2=>nx10871);
   ix7029 : nor03_2x port map ( Y=>nx7028, A0=>nx7311, A1=>nx10877, A2=>
      nx10887);
   ix7330 : nor02_2x port map ( Y=>nx7329, A0=>nx7024, A1=>nx7022);
   ix7025 : nor03_2x port map ( Y=>nx7024, A0=>nx7333, A1=>nx9471, A2=>
      nx10895);
   gen_18_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_18_cmp_mReg_2, QB=>
      nx7333, D=>window_18_2, CLK=>start, R=>rst);
   ix7023 : nor03_2x port map ( Y=>nx7022, A0=>gen_18_cmp_mReg_2, A1=>
      nx10107, A2=>nx10903);
   ix7059 : nand02 port map ( Y=>gen_18_cmp_BSCmp_op2_3, A0=>nx7339, A1=>
      nx7344);
   ix7340 : nor02_2x port map ( Y=>nx7339, A0=>nx7054, A1=>nx7050);
   ix7055 : nor03_2x port map ( Y=>nx7054, A0=>gen_18_cmp_mReg_2, A1=>nx9477, 
      A2=>nx10871);
   ix7051 : nor03_2x port map ( Y=>nx7050, A0=>nx7333, A1=>nx10877, A2=>
      nx10887);
   ix7345 : nor02_2x port map ( Y=>nx7344, A0=>nx7046, A1=>nx7044);
   ix7047 : nor03_2x port map ( Y=>nx7046, A0=>nx7347, A1=>nx9471, A2=>
      nx10895);
   gen_18_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_18_cmp_mReg_3, QB=>
      nx7347, D=>window_18_3, CLK=>start, R=>rst);
   ix7045 : nor03_2x port map ( Y=>nx7044, A0=>gen_18_cmp_mReg_3, A1=>
      nx10107, A2=>nx10903);
   ix7081 : nand02 port map ( Y=>gen_18_cmp_BSCmp_op2_4, A0=>nx7351, A1=>
      nx7357);
   ix7352 : nor02_2x port map ( Y=>nx7351, A0=>nx7076, A1=>nx7072);
   ix7077 : nor03_2x port map ( Y=>nx7076, A0=>gen_18_cmp_mReg_3, A1=>nx9477, 
      A2=>nx10871);
   ix7073 : nor03_2x port map ( Y=>nx7072, A0=>nx7347, A1=>nx10877, A2=>
      nx10887);
   ix7358 : nor02_2x port map ( Y=>nx7357, A0=>nx7068, A1=>nx7066);
   ix7069 : nor03_2x port map ( Y=>nx7068, A0=>nx7361, A1=>nx9471, A2=>
      nx10895);
   gen_18_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_18_cmp_mReg_4, QB=>
      nx7361, D=>window_18_4, CLK=>start, R=>rst);
   ix7067 : nor03_2x port map ( Y=>nx7066, A0=>gen_18_cmp_mReg_4, A1=>
      nx10107, A2=>nx10903);
   ix7103 : nand02 port map ( Y=>gen_18_cmp_BSCmp_op2_5, A0=>nx7367, A1=>
      nx7373);
   ix7368 : nor02_2x port map ( Y=>nx7367, A0=>nx7098, A1=>nx7094);
   ix7099 : nor03_2x port map ( Y=>nx7098, A0=>gen_18_cmp_mReg_4, A1=>nx9477, 
      A2=>nx10871);
   ix7095 : nor03_2x port map ( Y=>nx7094, A0=>nx7361, A1=>nx10877, A2=>
      nx10887);
   ix7374 : nor02_2x port map ( Y=>nx7373, A0=>nx7090, A1=>nx7088);
   ix7091 : nor03_2x port map ( Y=>nx7090, A0=>nx7376, A1=>nx9473, A2=>
      nx10895);
   gen_18_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_18_cmp_mReg_5, QB=>
      nx7376, D=>window_18_5, CLK=>start, R=>rst);
   ix7089 : nor03_2x port map ( Y=>nx7088, A0=>gen_18_cmp_mReg_5, A1=>
      nx10107, A2=>nx10903);
   ix7125 : nand02 port map ( Y=>gen_18_cmp_BSCmp_op2_6, A0=>nx7381, A1=>
      nx7387);
   ix7382 : nor02_2x port map ( Y=>nx7381, A0=>nx7120, A1=>nx7116);
   ix7121 : nor03_2x port map ( Y=>nx7120, A0=>gen_18_cmp_mReg_5, A1=>nx9479, 
      A2=>nx10871);
   ix7117 : nor03_2x port map ( Y=>nx7116, A0=>nx7376, A1=>nx10877, A2=>
      nx10887);
   ix7388 : nor02_2x port map ( Y=>nx7387, A0=>nx7112, A1=>nx7110);
   ix7113 : nor03_2x port map ( Y=>nx7112, A0=>nx7391, A1=>nx9473, A2=>
      nx10895);
   gen_18_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_18_cmp_mReg_6, QB=>
      nx7391, D=>window_18_6, CLK=>start, R=>rst);
   ix7111 : nor03_2x port map ( Y=>nx7110, A0=>gen_18_cmp_mReg_6, A1=>
      nx10107, A2=>nx10903);
   ix7147 : nand02 port map ( Y=>gen_18_cmp_BSCmp_op2_7, A0=>nx7397, A1=>
      nx7403);
   ix7398 : nor02_2x port map ( Y=>nx7397, A0=>nx7142, A1=>nx7138);
   ix7143 : nor03_2x port map ( Y=>nx7142, A0=>gen_18_cmp_mReg_6, A1=>nx9479, 
      A2=>nx10873);
   ix7139 : nor03_2x port map ( Y=>nx7138, A0=>nx7391, A1=>nx10879, A2=>
      nx10889);
   ix7404 : nor02_2x port map ( Y=>nx7403, A0=>nx7134, A1=>nx7132);
   ix7135 : nor03_2x port map ( Y=>nx7134, A0=>nx7406, A1=>nx9473, A2=>
      nx10897);
   gen_18_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_18_cmp_mReg_7, QB=>
      nx7406, D=>window_18_7, CLK=>start, R=>rst);
   ix7133 : nor03_2x port map ( Y=>nx7132, A0=>gen_18_cmp_mReg_7, A1=>
      nx10107, A2=>nx10905);
   ix7169 : nand02 port map ( Y=>gen_18_cmp_BSCmp_op2_8, A0=>nx7413, A1=>
      nx7419);
   ix7414 : nor02_2x port map ( Y=>nx7413, A0=>nx7164, A1=>nx7160);
   ix7165 : nor03_2x port map ( Y=>nx7164, A0=>gen_18_cmp_mReg_7, A1=>nx9479, 
      A2=>nx10873);
   ix7161 : nor03_2x port map ( Y=>nx7160, A0=>nx7406, A1=>nx10879, A2=>
      nx10889);
   ix7420 : nor02_2x port map ( Y=>nx7419, A0=>nx7156, A1=>nx7154);
   ix7157 : nor03_2x port map ( Y=>nx7156, A0=>nx7423, A1=>nx9473, A2=>
      nx10897);
   gen_18_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_18_cmp_mReg_8, QB=>
      nx7423, D=>window_18_8, CLK=>start, R=>rst);
   ix7155 : nor03_2x port map ( Y=>nx7154, A0=>gen_18_cmp_mReg_8, A1=>
      nx10109, A2=>nx10905);
   ix7191 : nand02 port map ( Y=>gen_18_cmp_BSCmp_op2_9, A0=>nx7427, A1=>
      nx7433);
   ix7428 : nor02_2x port map ( Y=>nx7427, A0=>nx7186, A1=>nx7182);
   ix7187 : nor03_2x port map ( Y=>nx7186, A0=>gen_18_cmp_mReg_8, A1=>nx9479, 
      A2=>nx10873);
   ix7183 : nor03_2x port map ( Y=>nx7182, A0=>nx7423, A1=>nx10879, A2=>
      nx10889);
   ix7434 : nor02_2x port map ( Y=>nx7433, A0=>nx7178, A1=>nx7176);
   ix7179 : nor03_2x port map ( Y=>nx7178, A0=>nx7437, A1=>nx9473, A2=>
      nx10897);
   gen_18_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_18_cmp_mReg_9, QB=>
      nx7437, D=>window_18_9, CLK=>start, R=>rst);
   ix7177 : nor03_2x port map ( Y=>nx7176, A0=>gen_18_cmp_mReg_9, A1=>
      nx10109, A2=>nx10905);
   ix7213 : nand02 port map ( Y=>gen_18_cmp_BSCmp_op2_10, A0=>nx7441, A1=>
      nx7447);
   ix7442 : nor02_2x port map ( Y=>nx7441, A0=>nx7208, A1=>nx7204);
   ix7209 : nor03_2x port map ( Y=>nx7208, A0=>gen_18_cmp_mReg_9, A1=>nx9479, 
      A2=>nx10873);
   ix7205 : nor03_2x port map ( Y=>nx7204, A0=>nx7437, A1=>nx10879, A2=>
      nx10889);
   ix7448 : nor02_2x port map ( Y=>nx7447, A0=>nx7200, A1=>nx7198);
   ix7201 : nor03_2x port map ( Y=>nx7200, A0=>nx7450, A1=>nx9473, A2=>
      nx10897);
   gen_18_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_18_cmp_mReg_10, QB=>
      nx7450, D=>window_18_10, CLK=>start, R=>rst);
   ix7199 : nor03_2x port map ( Y=>nx7198, A0=>gen_18_cmp_mReg_10, A1=>
      nx10109, A2=>nx10905);
   ix7235 : nand02 port map ( Y=>gen_18_cmp_BSCmp_op2_11, A0=>nx7457, A1=>
      nx7463);
   ix7458 : nor02_2x port map ( Y=>nx7457, A0=>nx7230, A1=>nx7226);
   ix7231 : nor03_2x port map ( Y=>nx7230, A0=>gen_18_cmp_mReg_10, A1=>
      nx9479, A2=>nx10873);
   ix7227 : nor03_2x port map ( Y=>nx7226, A0=>nx7450, A1=>nx10879, A2=>
      nx10889);
   ix7464 : nor02_2x port map ( Y=>nx7463, A0=>nx7222, A1=>nx7220);
   ix7223 : nor03_2x port map ( Y=>nx7222, A0=>nx7467, A1=>nx9473, A2=>
      nx10897);
   gen_18_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_18_cmp_mReg_11, QB=>
      nx7467, D=>window_18_11, CLK=>start, R=>rst);
   ix7221 : nor03_2x port map ( Y=>nx7220, A0=>gen_18_cmp_mReg_11, A1=>
      nx10109, A2=>nx10905);
   ix7257 : nand02 port map ( Y=>gen_18_cmp_BSCmp_op2_12, A0=>nx7471, A1=>
      nx7477);
   ix7472 : nor02_2x port map ( Y=>nx7471, A0=>nx7252, A1=>nx7248);
   ix7253 : nor03_2x port map ( Y=>nx7252, A0=>gen_18_cmp_mReg_11, A1=>
      nx9479, A2=>nx10873);
   ix7249 : nor03_2x port map ( Y=>nx7248, A0=>nx7467, A1=>nx10879, A2=>
      nx10889);
   ix7478 : nor02_2x port map ( Y=>nx7477, A0=>nx7244, A1=>nx7242);
   ix7245 : nor03_2x port map ( Y=>nx7244, A0=>nx7481, A1=>nx9475, A2=>
      nx10897);
   gen_18_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_18_cmp_mReg_12, QB=>
      nx7481, D=>window_18_12, CLK=>start, R=>rst);
   ix7243 : nor03_2x port map ( Y=>nx7242, A0=>gen_18_cmp_mReg_12, A1=>
      nx10109, A2=>nx10905);
   ix7279 : nand02 port map ( Y=>gen_18_cmp_BSCmp_op2_13, A0=>nx7485, A1=>
      nx7491);
   ix7486 : nor02_2x port map ( Y=>nx7485, A0=>nx7274, A1=>nx7270);
   ix7275 : nor03_2x port map ( Y=>nx7274, A0=>gen_18_cmp_mReg_12, A1=>
      nx9481, A2=>nx10875);
   ix7271 : nor03_2x port map ( Y=>nx7270, A0=>nx7481, A1=>nx10879, A2=>
      nx10891);
   ix7492 : nor02_2x port map ( Y=>nx7491, A0=>nx7266, A1=>nx7264);
   ix7267 : nor03_2x port map ( Y=>nx7266, A0=>nx7494, A1=>nx9475, A2=>
      nx10899);
   gen_18_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_18_cmp_mReg_13, QB=>
      nx7494, D=>window_18_13, CLK=>start, R=>rst);
   ix7265 : nor03_2x port map ( Y=>nx7264, A0=>gen_18_cmp_mReg_13, A1=>
      nx10109, A2=>nx10907);
   ix7301 : nand02 port map ( Y=>gen_18_cmp_BSCmp_op2_14, A0=>nx7501, A1=>
      nx7507);
   ix7502 : nor02_2x port map ( Y=>nx7501, A0=>nx7296, A1=>nx7292);
   ix7297 : nor03_2x port map ( Y=>nx7296, A0=>gen_18_cmp_mReg_13, A1=>
      nx9481, A2=>nx10875);
   ix7293 : nor03_2x port map ( Y=>nx7292, A0=>nx7494, A1=>nx10881, A2=>
      nx10891);
   ix7508 : nor02_2x port map ( Y=>nx7507, A0=>nx7288, A1=>nx7286);
   ix7289 : nor03_2x port map ( Y=>nx7288, A0=>nx7511, A1=>nx9475, A2=>
      nx10899);
   gen_18_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_18_cmp_mReg_14, QB=>
      nx7511, D=>window_18_14, CLK=>start, R=>rst);
   ix7287 : nor03_2x port map ( Y=>nx7286, A0=>gen_18_cmp_mReg_14, A1=>
      nx10109, A2=>nx10907);
   ix7323 : nand02 port map ( Y=>gen_18_cmp_BSCmp_op2_15, A0=>nx7515, A1=>
      nx7521);
   ix7516 : nor02_2x port map ( Y=>nx7515, A0=>nx7318, A1=>nx7314);
   ix7319 : nor03_2x port map ( Y=>nx7318, A0=>gen_18_cmp_mReg_14, A1=>
      nx9481, A2=>nx10875);
   ix7315 : nor03_2x port map ( Y=>nx7314, A0=>nx7511, A1=>nx10881, A2=>
      nx10891);
   ix7522 : nor02_2x port map ( Y=>nx7521, A0=>nx7310, A1=>nx7308);
   ix7311 : nor03_2x port map ( Y=>nx7310, A0=>nx7525, A1=>nx9475, A2=>
      nx10899);
   gen_18_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_18_cmp_mReg_15, QB=>
      nx7525, D=>window_18_15, CLK=>start, R=>rst);
   ix7309 : nor03_2x port map ( Y=>nx7308, A0=>gen_18_cmp_mReg_15, A1=>
      nx10111, A2=>nx10907);
   ix7333 : nand02 port map ( Y=>gen_18_cmp_BSCmp_op2_16, A0=>nx7529, A1=>
      nx7521);
   ix7530 : nor02_2x port map ( Y=>nx7529, A0=>nx7328, A1=>nx7324);
   ix7329 : nor03_2x port map ( Y=>nx7328, A0=>gen_18_cmp_mReg_15, A1=>
      nx9481, A2=>nx10875);
   ix7325 : nor03_2x port map ( Y=>nx7324, A0=>nx7525, A1=>nx10881, A2=>
      nx10891);
   ix7401 : nand02 port map ( Y=>gen_19_cmp_BSCmp_op2_1, A0=>nx7536, A1=>
      nx7555);
   ix7537 : nor02_2x port map ( Y=>nx7536, A0=>nx7396, A1=>nx7392);
   ix7397 : nor03_2x port map ( Y=>nx7396, A0=>gen_19_cmp_mReg_0, A1=>nx9465, 
      A2=>nx10911);
   gen_19_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_19_cmp_mReg_0, QB=>
      nx7541, D=>window_19_0, CLK=>start, R=>rst);
   ix7546 : inv01 port map ( Y=>nx7545, A=>gen_19_cmp_pMux_0);
   ix7393 : nor03_2x port map ( Y=>nx7392, A0=>nx7541, A1=>nx10917, A2=>
      nx10927);
   ix7554 : inv02 port map ( Y=>nx7553, A=>gen_19_cmp_pMux_2);
   ix7556 : nor02_2x port map ( Y=>nx7555, A0=>nx7382, A1=>nx7380);
   ix7383 : nor03_2x port map ( Y=>nx7382, A0=>nx7558, A1=>nx9459, A2=>
      nx10935);
   gen_19_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_19_cmp_mReg_1, QB=>
      nx7558, D=>window_19_1, CLK=>start, R=>rst);
   ix7381 : nor03_2x port map ( Y=>nx7380, A0=>gen_19_cmp_mReg_1, A1=>
      nx10113, A2=>nx10943);
   ix7341 : nor03_2x port map ( Y=>nx7340, A0=>nx9465, A1=>nx7553, A2=>
      gen_19_cmp_pMux_0);
   ix7423 : nand02 port map ( Y=>gen_19_cmp_BSCmp_op2_2, A0=>nx7571, A1=>
      nx7577);
   ix7572 : nor02_2x port map ( Y=>nx7571, A0=>nx7418, A1=>nx7414);
   ix7419 : nor03_2x port map ( Y=>nx7418, A0=>gen_19_cmp_mReg_1, A1=>nx9465, 
      A2=>nx10911);
   ix7415 : nor03_2x port map ( Y=>nx7414, A0=>nx7558, A1=>nx10917, A2=>
      nx10927);
   ix7578 : nor02_2x port map ( Y=>nx7577, A0=>nx7410, A1=>nx7408);
   ix7411 : nor03_2x port map ( Y=>nx7410, A0=>nx7580, A1=>nx9459, A2=>
      nx10935);
   gen_19_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_19_cmp_mReg_2, QB=>
      nx7580, D=>window_19_2, CLK=>start, R=>rst);
   ix7409 : nor03_2x port map ( Y=>nx7408, A0=>gen_19_cmp_mReg_2, A1=>
      nx10113, A2=>nx10943);
   ix7445 : nand02 port map ( Y=>gen_19_cmp_BSCmp_op2_3, A0=>nx7585, A1=>
      nx7591);
   ix7586 : nor02_2x port map ( Y=>nx7585, A0=>nx7440, A1=>nx7436);
   ix7441 : nor03_2x port map ( Y=>nx7440, A0=>gen_19_cmp_mReg_2, A1=>nx9465, 
      A2=>nx10911);
   ix7437 : nor03_2x port map ( Y=>nx7436, A0=>nx7580, A1=>nx10917, A2=>
      nx10927);
   ix7592 : nor02_2x port map ( Y=>nx7591, A0=>nx7432, A1=>nx7430);
   ix7433 : nor03_2x port map ( Y=>nx7432, A0=>nx7595, A1=>nx9459, A2=>
      nx10935);
   gen_19_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_19_cmp_mReg_3, QB=>
      nx7595, D=>window_19_3, CLK=>start, R=>rst);
   ix7431 : nor03_2x port map ( Y=>nx7430, A0=>gen_19_cmp_mReg_3, A1=>
      nx10113, A2=>nx10943);
   ix7467 : nand02 port map ( Y=>gen_19_cmp_BSCmp_op2_4, A0=>nx7601, A1=>
      nx7605);
   ix7602 : nor02_2x port map ( Y=>nx7601, A0=>nx7462, A1=>nx7458);
   ix7463 : nor03_2x port map ( Y=>nx7462, A0=>gen_19_cmp_mReg_3, A1=>nx9465, 
      A2=>nx10911);
   ix7459 : nor03_2x port map ( Y=>nx7458, A0=>nx7595, A1=>nx10917, A2=>
      nx10927);
   ix7606 : nor02_2x port map ( Y=>nx7605, A0=>nx7454, A1=>nx7452);
   ix7455 : nor03_2x port map ( Y=>nx7454, A0=>nx7609, A1=>nx9459, A2=>
      nx10935);
   gen_19_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_19_cmp_mReg_4, QB=>
      nx7609, D=>window_19_4, CLK=>start, R=>rst);
   ix7453 : nor03_2x port map ( Y=>nx7452, A0=>gen_19_cmp_mReg_4, A1=>
      nx10113, A2=>nx10943);
   ix7489 : nand02 port map ( Y=>gen_19_cmp_BSCmp_op2_5, A0=>nx7615, A1=>
      nx7621);
   ix7616 : nor02_2x port map ( Y=>nx7615, A0=>nx7484, A1=>nx7480);
   ix7485 : nor03_2x port map ( Y=>nx7484, A0=>gen_19_cmp_mReg_4, A1=>nx9465, 
      A2=>nx10911);
   ix7481 : nor03_2x port map ( Y=>nx7480, A0=>nx7609, A1=>nx10917, A2=>
      nx10927);
   ix7622 : nor02_2x port map ( Y=>nx7621, A0=>nx7476, A1=>nx7474);
   ix7477 : nor03_2x port map ( Y=>nx7476, A0=>nx7624, A1=>nx9461, A2=>
      nx10935);
   gen_19_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_19_cmp_mReg_5, QB=>
      nx7624, D=>window_19_5, CLK=>start, R=>rst);
   ix7475 : nor03_2x port map ( Y=>nx7474, A0=>gen_19_cmp_mReg_5, A1=>
      nx10113, A2=>nx10943);
   ix7511 : nand02 port map ( Y=>gen_19_cmp_BSCmp_op2_6, A0=>nx7629, A1=>
      nx7635);
   ix7630 : nor02_2x port map ( Y=>nx7629, A0=>nx7506, A1=>nx7502);
   ix7507 : nor03_2x port map ( Y=>nx7506, A0=>gen_19_cmp_mReg_5, A1=>nx9467, 
      A2=>nx10911);
   ix7503 : nor03_2x port map ( Y=>nx7502, A0=>nx7624, A1=>nx10917, A2=>
      nx10927);
   ix7636 : nor02_2x port map ( Y=>nx7635, A0=>nx7498, A1=>nx7496);
   ix7499 : nor03_2x port map ( Y=>nx7498, A0=>nx7639, A1=>nx9461, A2=>
      nx10935);
   gen_19_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_19_cmp_mReg_6, QB=>
      nx7639, D=>window_19_6, CLK=>start, R=>rst);
   ix7497 : nor03_2x port map ( Y=>nx7496, A0=>gen_19_cmp_mReg_6, A1=>
      nx10113, A2=>nx10943);
   ix7533 : nand02 port map ( Y=>gen_19_cmp_BSCmp_op2_7, A0=>nx7645, A1=>
      nx7649);
   ix7646 : nor02_2x port map ( Y=>nx7645, A0=>nx7528, A1=>nx7524);
   ix7529 : nor03_2x port map ( Y=>nx7528, A0=>gen_19_cmp_mReg_6, A1=>nx9467, 
      A2=>nx10913);
   ix7525 : nor03_2x port map ( Y=>nx7524, A0=>nx7639, A1=>nx10919, A2=>
      nx10929);
   ix7650 : nor02_2x port map ( Y=>nx7649, A0=>nx7520, A1=>nx7518);
   ix7521 : nor03_2x port map ( Y=>nx7520, A0=>nx7653, A1=>nx9461, A2=>
      nx10937);
   gen_19_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_19_cmp_mReg_7, QB=>
      nx7653, D=>window_19_7, CLK=>start, R=>rst);
   ix7519 : nor03_2x port map ( Y=>nx7518, A0=>gen_19_cmp_mReg_7, A1=>
      nx10113, A2=>nx10945);
   ix7555 : nand02 port map ( Y=>gen_19_cmp_BSCmp_op2_8, A0=>nx7659, A1=>
      nx7665);
   ix7660 : nor02_2x port map ( Y=>nx7659, A0=>nx7550, A1=>nx7546);
   ix7551 : nor03_2x port map ( Y=>nx7550, A0=>gen_19_cmp_mReg_7, A1=>nx9467, 
      A2=>nx10913);
   ix7547 : nor03_2x port map ( Y=>nx7546, A0=>nx7653, A1=>nx10919, A2=>
      nx10929);
   ix7666 : nor02_2x port map ( Y=>nx7665, A0=>nx7542, A1=>nx7540);
   ix7543 : nor03_2x port map ( Y=>nx7542, A0=>nx7668, A1=>nx9461, A2=>
      nx10937);
   gen_19_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_19_cmp_mReg_8, QB=>
      nx7668, D=>window_19_8, CLK=>start, R=>rst);
   ix7541 : nor03_2x port map ( Y=>nx7540, A0=>gen_19_cmp_mReg_8, A1=>
      nx10115, A2=>nx10945);
   ix7577 : nand02 port map ( Y=>gen_19_cmp_BSCmp_op2_9, A0=>nx7673, A1=>
      nx7679);
   ix7674 : nor02_2x port map ( Y=>nx7673, A0=>nx7572, A1=>nx7568);
   ix7573 : nor03_2x port map ( Y=>nx7572, A0=>gen_19_cmp_mReg_8, A1=>nx9467, 
      A2=>nx10913);
   ix7569 : nor03_2x port map ( Y=>nx7568, A0=>nx7668, A1=>nx10919, A2=>
      nx10929);
   ix7680 : nor02_2x port map ( Y=>nx7679, A0=>nx7564, A1=>nx7562);
   ix7565 : nor03_2x port map ( Y=>nx7564, A0=>nx7683, A1=>nx9461, A2=>
      nx10937);
   gen_19_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_19_cmp_mReg_9, QB=>
      nx7683, D=>window_19_9, CLK=>start, R=>rst);
   ix7563 : nor03_2x port map ( Y=>nx7562, A0=>gen_19_cmp_mReg_9, A1=>
      nx10115, A2=>nx10945);
   ix7599 : nand02 port map ( Y=>gen_19_cmp_BSCmp_op2_10, A0=>nx7689, A1=>
      nx7693);
   ix7690 : nor02_2x port map ( Y=>nx7689, A0=>nx7594, A1=>nx7590);
   ix7595 : nor03_2x port map ( Y=>nx7594, A0=>gen_19_cmp_mReg_9, A1=>nx9467, 
      A2=>nx10913);
   ix7591 : nor03_2x port map ( Y=>nx7590, A0=>nx7683, A1=>nx10919, A2=>
      nx10929);
   ix7694 : nor02_2x port map ( Y=>nx7693, A0=>nx7586, A1=>nx7584);
   ix7587 : nor03_2x port map ( Y=>nx7586, A0=>nx7697, A1=>nx9461, A2=>
      nx10937);
   gen_19_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_19_cmp_mReg_10, QB=>
      nx7697, D=>window_19_10, CLK=>start, R=>rst);
   ix7585 : nor03_2x port map ( Y=>nx7584, A0=>gen_19_cmp_mReg_10, A1=>
      nx10115, A2=>nx10945);
   ix7621 : nand02 port map ( Y=>gen_19_cmp_BSCmp_op2_11, A0=>nx7703, A1=>
      nx7709);
   ix7704 : nor02_2x port map ( Y=>nx7703, A0=>nx7616, A1=>nx7612);
   ix7617 : nor03_2x port map ( Y=>nx7616, A0=>gen_19_cmp_mReg_10, A1=>
      nx9467, A2=>nx10913);
   ix7613 : nor03_2x port map ( Y=>nx7612, A0=>nx7697, A1=>nx10919, A2=>
      nx10929);
   ix7710 : nor02_2x port map ( Y=>nx7709, A0=>nx7608, A1=>nx7606);
   ix7609 : nor03_2x port map ( Y=>nx7608, A0=>nx7713, A1=>nx9461, A2=>
      nx10937);
   gen_19_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_19_cmp_mReg_11, QB=>
      nx7713, D=>window_19_11, CLK=>start, R=>rst);
   ix7607 : nor03_2x port map ( Y=>nx7606, A0=>gen_19_cmp_mReg_11, A1=>
      nx10115, A2=>nx10945);
   ix7643 : nand02 port map ( Y=>gen_19_cmp_BSCmp_op2_12, A0=>nx7719, A1=>
      nx7725);
   ix7720 : nor02_2x port map ( Y=>nx7719, A0=>nx7638, A1=>nx7634);
   ix7639 : nor03_2x port map ( Y=>nx7638, A0=>gen_19_cmp_mReg_11, A1=>
      nx9467, A2=>nx10913);
   ix7635 : nor03_2x port map ( Y=>nx7634, A0=>nx7713, A1=>nx10919, A2=>
      nx10929);
   ix7726 : nor02_2x port map ( Y=>nx7725, A0=>nx7630, A1=>nx7628);
   ix7631 : nor03_2x port map ( Y=>nx7630, A0=>nx7729, A1=>nx9463, A2=>
      nx10937);
   gen_19_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_19_cmp_mReg_12, QB=>
      nx7729, D=>window_19_12, CLK=>start, R=>rst);
   ix7629 : nor03_2x port map ( Y=>nx7628, A0=>gen_19_cmp_mReg_12, A1=>
      nx10115, A2=>nx10945);
   ix7665 : nand02 port map ( Y=>gen_19_cmp_BSCmp_op2_13, A0=>nx7733, A1=>
      nx7737);
   ix7734 : nor02_2x port map ( Y=>nx7733, A0=>nx7660, A1=>nx7656);
   ix7661 : nor03_2x port map ( Y=>nx7660, A0=>gen_19_cmp_mReg_12, A1=>
      nx9469, A2=>nx10915);
   ix7657 : nor03_2x port map ( Y=>nx7656, A0=>nx7729, A1=>nx10919, A2=>
      nx10931);
   ix7738 : nor02_2x port map ( Y=>nx7737, A0=>nx7652, A1=>nx7650);
   ix7653 : nor03_2x port map ( Y=>nx7652, A0=>nx7741, A1=>nx9463, A2=>
      nx10939);
   gen_19_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_19_cmp_mReg_13, QB=>
      nx7741, D=>window_19_13, CLK=>start, R=>rst);
   ix7651 : nor03_2x port map ( Y=>nx7650, A0=>gen_19_cmp_mReg_13, A1=>
      nx10115, A2=>nx10947);
   ix7687 : nand02 port map ( Y=>gen_19_cmp_BSCmp_op2_14, A0=>nx7747, A1=>
      nx7753);
   ix7748 : nor02_2x port map ( Y=>nx7747, A0=>nx7682, A1=>nx7678);
   ix7683 : nor03_2x port map ( Y=>nx7682, A0=>gen_19_cmp_mReg_13, A1=>
      nx9469, A2=>nx10915);
   ix7679 : nor03_2x port map ( Y=>nx7678, A0=>nx7741, A1=>nx10921, A2=>
      nx10931);
   ix7754 : nor02_2x port map ( Y=>nx7753, A0=>nx7674, A1=>nx7672);
   ix7675 : nor03_2x port map ( Y=>nx7674, A0=>nx7757, A1=>nx9463, A2=>
      nx10939);
   gen_19_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_19_cmp_mReg_14, QB=>
      nx7757, D=>window_19_14, CLK=>start, R=>rst);
   ix7673 : nor03_2x port map ( Y=>nx7672, A0=>gen_19_cmp_mReg_14, A1=>
      nx10115, A2=>nx10947);
   ix7709 : nand02 port map ( Y=>gen_19_cmp_BSCmp_op2_15, A0=>nx7762, A1=>
      nx7767);
   ix7763 : nor02_2x port map ( Y=>nx7762, A0=>nx7704, A1=>nx7700);
   ix7705 : nor03_2x port map ( Y=>nx7704, A0=>gen_19_cmp_mReg_14, A1=>
      nx9469, A2=>nx10915);
   ix7701 : nor03_2x port map ( Y=>nx7700, A0=>nx7757, A1=>nx10921, A2=>
      nx10931);
   ix7768 : nor02_2x port map ( Y=>nx7767, A0=>nx7696, A1=>nx7694);
   ix7697 : nor03_2x port map ( Y=>nx7696, A0=>nx7771, A1=>nx9463, A2=>
      nx10939);
   gen_19_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_19_cmp_mReg_15, QB=>
      nx7771, D=>window_19_15, CLK=>start, R=>rst);
   ix7695 : nor03_2x port map ( Y=>nx7694, A0=>gen_19_cmp_mReg_15, A1=>
      nx10117, A2=>nx10947);
   ix7719 : nand02 port map ( Y=>gen_19_cmp_BSCmp_op2_16, A0=>nx7775, A1=>
      nx7767);
   ix7776 : nor02_2x port map ( Y=>nx7775, A0=>nx7714, A1=>nx7710);
   ix7715 : nor03_2x port map ( Y=>nx7714, A0=>gen_19_cmp_mReg_15, A1=>
      nx9469, A2=>nx10915);
   ix7711 : nor03_2x port map ( Y=>nx7710, A0=>nx7771, A1=>nx10921, A2=>
      nx10931);
   ix7787 : nand02 port map ( Y=>gen_20_cmp_BSCmp_op2_1, A0=>nx7783, A1=>
      nx7803);
   ix7784 : nor02_2x port map ( Y=>nx7783, A0=>nx7782, A1=>nx7778);
   ix7783 : nor03_2x port map ( Y=>nx7782, A0=>gen_20_cmp_mReg_0, A1=>nx9453, 
      A2=>nx10951);
   gen_20_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_20_cmp_mReg_0, QB=>
      nx7789, D=>window_20_0, CLK=>start, R=>rst);
   ix7794 : inv01 port map ( Y=>nx7792, A=>gen_20_cmp_pMux_0);
   ix7779 : nor03_2x port map ( Y=>nx7778, A0=>nx7789, A1=>nx10957, A2=>
      nx10967);
   ix7802 : inv02 port map ( Y=>nx7801, A=>gen_20_cmp_pMux_2);
   ix7804 : nor02_2x port map ( Y=>nx7803, A0=>nx7768, A1=>nx7766);
   ix7769 : nor03_2x port map ( Y=>nx7768, A0=>nx7807, A1=>nx9447, A2=>
      nx10975);
   gen_20_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_20_cmp_mReg_1, QB=>
      nx7807, D=>window_20_1, CLK=>start, R=>rst);
   ix7767 : nor03_2x port map ( Y=>nx7766, A0=>gen_20_cmp_mReg_1, A1=>
      nx10119, A2=>nx10983);
   ix7727 : nor03_2x port map ( Y=>nx7726, A0=>nx9453, A1=>nx7801, A2=>
      gen_20_cmp_pMux_0);
   ix7809 : nand02 port map ( Y=>gen_20_cmp_BSCmp_op2_2, A0=>nx7817, A1=>
      nx7823);
   ix7818 : nor02_2x port map ( Y=>nx7817, A0=>nx7804, A1=>nx7800);
   ix7805 : nor03_2x port map ( Y=>nx7804, A0=>gen_20_cmp_mReg_1, A1=>nx9453, 
      A2=>nx10951);
   ix7801 : nor03_2x port map ( Y=>nx7800, A0=>nx7807, A1=>nx10957, A2=>
      nx10967);
   ix7824 : nor02_2x port map ( Y=>nx7823, A0=>nx7796, A1=>nx7794);
   ix7797 : nor03_2x port map ( Y=>nx7796, A0=>nx7827, A1=>nx9447, A2=>
      nx10975);
   gen_20_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_20_cmp_mReg_2, QB=>
      nx7827, D=>window_20_2, CLK=>start, R=>rst);
   ix7795 : nor03_2x port map ( Y=>nx7794, A0=>gen_20_cmp_mReg_2, A1=>
      nx10119, A2=>nx10983);
   ix7831 : nand02 port map ( Y=>gen_20_cmp_BSCmp_op2_3, A0=>nx7833, A1=>
      nx7837);
   ix7834 : nor02_2x port map ( Y=>nx7833, A0=>nx7826, A1=>nx7822);
   ix7827 : nor03_2x port map ( Y=>nx7826, A0=>gen_20_cmp_mReg_2, A1=>nx9453, 
      A2=>nx10951);
   ix7823 : nor03_2x port map ( Y=>nx7822, A0=>nx7827, A1=>nx10957, A2=>
      nx10967);
   ix7838 : nor02_2x port map ( Y=>nx7837, A0=>nx7818, A1=>nx7816);
   ix7819 : nor03_2x port map ( Y=>nx7818, A0=>nx7841, A1=>nx9447, A2=>
      nx10975);
   gen_20_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_20_cmp_mReg_3, QB=>
      nx7841, D=>window_20_3, CLK=>start, R=>rst);
   ix7817 : nor03_2x port map ( Y=>nx7816, A0=>gen_20_cmp_mReg_3, A1=>
      nx10119, A2=>nx10983);
   ix7853 : nand02 port map ( Y=>gen_20_cmp_BSCmp_op2_4, A0=>nx7847, A1=>
      nx7853);
   ix7848 : nor02_2x port map ( Y=>nx7847, A0=>nx7848, A1=>nx7844);
   ix7849 : nor03_2x port map ( Y=>nx7848, A0=>gen_20_cmp_mReg_3, A1=>nx9453, 
      A2=>nx10951);
   ix7845 : nor03_2x port map ( Y=>nx7844, A0=>nx7841, A1=>nx10957, A2=>
      nx10967);
   ix7854 : nor02_2x port map ( Y=>nx7853, A0=>nx7840, A1=>nx7838);
   ix7841 : nor03_2x port map ( Y=>nx7840, A0=>nx7856, A1=>nx9447, A2=>
      nx10975);
   gen_20_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_20_cmp_mReg_4, QB=>
      nx7856, D=>window_20_4, CLK=>start, R=>rst);
   ix7839 : nor03_2x port map ( Y=>nx7838, A0=>gen_20_cmp_mReg_4, A1=>
      nx10119, A2=>nx10983);
   ix7875 : nand02 port map ( Y=>gen_20_cmp_BSCmp_op2_5, A0=>nx7861, A1=>
      nx7867);
   ix7862 : nor02_2x port map ( Y=>nx7861, A0=>nx7870, A1=>nx7866);
   ix7871 : nor03_2x port map ( Y=>nx7870, A0=>gen_20_cmp_mReg_4, A1=>nx9453, 
      A2=>nx10951);
   ix7867 : nor03_2x port map ( Y=>nx7866, A0=>nx7856, A1=>nx10957, A2=>
      nx10967);
   ix7868 : nor02_2x port map ( Y=>nx7867, A0=>nx7862, A1=>nx7860);
   ix7863 : nor03_2x port map ( Y=>nx7862, A0=>nx7871, A1=>nx9449, A2=>
      nx10975);
   gen_20_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_20_cmp_mReg_5, QB=>
      nx7871, D=>window_20_5, CLK=>start, R=>rst);
   ix7861 : nor03_2x port map ( Y=>nx7860, A0=>gen_20_cmp_mReg_5, A1=>
      nx10119, A2=>nx10983);
   ix7897 : nand02 port map ( Y=>gen_20_cmp_BSCmp_op2_6, A0=>nx7877, A1=>
      nx7881);
   ix7878 : nor02_2x port map ( Y=>nx7877, A0=>nx7892, A1=>nx7888);
   ix7893 : nor03_2x port map ( Y=>nx7892, A0=>gen_20_cmp_mReg_5, A1=>nx9455, 
      A2=>nx10951);
   ix7889 : nor03_2x port map ( Y=>nx7888, A0=>nx7871, A1=>nx10957, A2=>
      nx10967);
   ix7882 : nor02_2x port map ( Y=>nx7881, A0=>nx7884, A1=>nx7882);
   ix7885 : nor03_2x port map ( Y=>nx7884, A0=>nx7885, A1=>nx9449, A2=>
      nx10975);
   gen_20_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_20_cmp_mReg_6, QB=>
      nx7885, D=>window_20_6, CLK=>start, R=>rst);
   ix7883 : nor03_2x port map ( Y=>nx7882, A0=>gen_20_cmp_mReg_6, A1=>
      nx10119, A2=>nx10983);
   ix7919 : nand02 port map ( Y=>gen_20_cmp_BSCmp_op2_7, A0=>nx7891, A1=>
      nx7897);
   ix7892 : nor02_2x port map ( Y=>nx7891, A0=>nx7914, A1=>nx7910);
   ix7915 : nor03_2x port map ( Y=>nx7914, A0=>gen_20_cmp_mReg_6, A1=>nx9455, 
      A2=>nx10953);
   ix7911 : nor03_2x port map ( Y=>nx7910, A0=>nx7885, A1=>nx10959, A2=>
      nx10969);
   ix7898 : nor02_2x port map ( Y=>nx7897, A0=>nx7906, A1=>nx7904);
   ix7907 : nor03_2x port map ( Y=>nx7906, A0=>nx7900, A1=>nx9449, A2=>
      nx10977);
   gen_20_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_20_cmp_mReg_7, QB=>
      nx7900, D=>window_20_7, CLK=>start, R=>rst);
   ix7905 : nor03_2x port map ( Y=>nx7904, A0=>gen_20_cmp_mReg_7, A1=>
      nx10119, A2=>nx10985);
   ix7941 : nand02 port map ( Y=>gen_20_cmp_BSCmp_op2_8, A0=>nx7905, A1=>
      nx7911);
   ix7906 : nor02_2x port map ( Y=>nx7905, A0=>nx7936, A1=>nx7932);
   ix7937 : nor03_2x port map ( Y=>nx7936, A0=>gen_20_cmp_mReg_7, A1=>nx9455, 
      A2=>nx10953);
   ix7933 : nor03_2x port map ( Y=>nx7932, A0=>nx7900, A1=>nx10959, A2=>
      nx10969);
   ix7912 : nor02_2x port map ( Y=>nx7911, A0=>nx7928, A1=>nx7926);
   ix7929 : nor03_2x port map ( Y=>nx7928, A0=>nx7915, A1=>nx9449, A2=>
      nx10977);
   gen_20_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_20_cmp_mReg_8, QB=>
      nx7915, D=>window_20_8, CLK=>start, R=>rst);
   ix7927 : nor03_2x port map ( Y=>nx7926, A0=>gen_20_cmp_mReg_8, A1=>
      nx10121, A2=>nx10985);
   ix7963 : nand02 port map ( Y=>gen_20_cmp_BSCmp_op2_9, A0=>nx7921, A1=>
      nx7925);
   ix7922 : nor02_2x port map ( Y=>nx7921, A0=>nx7958, A1=>nx7954);
   ix7959 : nor03_2x port map ( Y=>nx7958, A0=>gen_20_cmp_mReg_8, A1=>nx9455, 
      A2=>nx10953);
   ix7955 : nor03_2x port map ( Y=>nx7954, A0=>nx7915, A1=>nx10959, A2=>
      nx10969);
   ix7926 : nor02_2x port map ( Y=>nx7925, A0=>nx7950, A1=>nx7948);
   ix7951 : nor03_2x port map ( Y=>nx7950, A0=>nx7929, A1=>nx9449, A2=>
      nx10977);
   gen_20_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_20_cmp_mReg_9, QB=>
      nx7929, D=>window_20_9, CLK=>start, R=>rst);
   ix7949 : nor03_2x port map ( Y=>nx7948, A0=>gen_20_cmp_mReg_9, A1=>
      nx10121, A2=>nx10985);
   ix7985 : nand02 port map ( Y=>gen_20_cmp_BSCmp_op2_10, A0=>nx7935, A1=>
      nx7941);
   ix7936 : nor02_2x port map ( Y=>nx7935, A0=>nx7980, A1=>nx7976);
   ix7981 : nor03_2x port map ( Y=>nx7980, A0=>gen_20_cmp_mReg_9, A1=>nx9455, 
      A2=>nx10953);
   ix7977 : nor03_2x port map ( Y=>nx7976, A0=>nx7929, A1=>nx10959, A2=>
      nx10969);
   ix7942 : nor02_2x port map ( Y=>nx7941, A0=>nx7972, A1=>nx7970);
   ix7973 : nor03_2x port map ( Y=>nx7972, A0=>nx7944, A1=>nx9449, A2=>
      nx10977);
   gen_20_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_20_cmp_mReg_10, QB=>
      nx7944, D=>window_20_10, CLK=>start, R=>rst);
   ix7971 : nor03_2x port map ( Y=>nx7970, A0=>gen_20_cmp_mReg_10, A1=>
      nx10121, A2=>nx10985);
   ix8007 : nand02 port map ( Y=>gen_20_cmp_BSCmp_op2_11, A0=>nx7949, A1=>
      nx7955);
   ix7950 : nor02_2x port map ( Y=>nx7949, A0=>nx8002, A1=>nx7998);
   ix8003 : nor03_2x port map ( Y=>nx8002, A0=>gen_20_cmp_mReg_10, A1=>
      nx9455, A2=>nx10953);
   ix7999 : nor03_2x port map ( Y=>nx7998, A0=>nx7944, A1=>nx10959, A2=>
      nx10969);
   ix7956 : nor02_2x port map ( Y=>nx7955, A0=>nx7994, A1=>nx7992);
   ix7995 : nor03_2x port map ( Y=>nx7994, A0=>nx7959, A1=>nx9449, A2=>
      nx10977);
   gen_20_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_20_cmp_mReg_11, QB=>
      nx7959, D=>window_20_11, CLK=>start, R=>rst);
   ix7993 : nor03_2x port map ( Y=>nx7992, A0=>gen_20_cmp_mReg_11, A1=>
      nx10121, A2=>nx10985);
   ix8029 : nand02 port map ( Y=>gen_20_cmp_BSCmp_op2_12, A0=>nx7965, A1=>
      nx7969);
   ix7966 : nor02_2x port map ( Y=>nx7965, A0=>nx8024, A1=>nx8020);
   ix8025 : nor03_2x port map ( Y=>nx8024, A0=>gen_20_cmp_mReg_11, A1=>
      nx9455, A2=>nx10953);
   ix8021 : nor03_2x port map ( Y=>nx8020, A0=>nx7959, A1=>nx10959, A2=>
      nx10969);
   ix7970 : nor02_2x port map ( Y=>nx7969, A0=>nx8016, A1=>nx8014);
   ix8017 : nor03_2x port map ( Y=>nx8016, A0=>nx7973, A1=>nx9451, A2=>
      nx10977);
   gen_20_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_20_cmp_mReg_12, QB=>
      nx7973, D=>window_20_12, CLK=>start, R=>rst);
   ix8015 : nor03_2x port map ( Y=>nx8014, A0=>gen_20_cmp_mReg_12, A1=>
      nx10121, A2=>nx10985);
   ix8051 : nand02 port map ( Y=>gen_20_cmp_BSCmp_op2_13, A0=>nx7979, A1=>
      nx7985);
   ix7980 : nor02_2x port map ( Y=>nx7979, A0=>nx8046, A1=>nx8042);
   ix8047 : nor03_2x port map ( Y=>nx8046, A0=>gen_20_cmp_mReg_12, A1=>
      nx9457, A2=>nx10955);
   ix8043 : nor03_2x port map ( Y=>nx8042, A0=>nx7973, A1=>nx10959, A2=>
      nx10971);
   ix7986 : nor02_2x port map ( Y=>nx7985, A0=>nx8038, A1=>nx8036);
   ix8039 : nor03_2x port map ( Y=>nx8038, A0=>nx7988, A1=>nx9451, A2=>
      nx10979);
   gen_20_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_20_cmp_mReg_13, QB=>
      nx7988, D=>window_20_13, CLK=>start, R=>rst);
   ix8037 : nor03_2x port map ( Y=>nx8036, A0=>gen_20_cmp_mReg_13, A1=>
      nx10121, A2=>nx10987);
   ix8073 : nand02 port map ( Y=>gen_20_cmp_BSCmp_op2_14, A0=>nx7993, A1=>
      nx7999);
   ix7994 : nor02_2x port map ( Y=>nx7993, A0=>nx8068, A1=>nx8064);
   ix8069 : nor03_2x port map ( Y=>nx8068, A0=>gen_20_cmp_mReg_13, A1=>
      nx9457, A2=>nx10955);
   ix8065 : nor03_2x port map ( Y=>nx8064, A0=>nx7988, A1=>nx10961, A2=>
      nx10971);
   ix8000 : nor02_2x port map ( Y=>nx7999, A0=>nx8060, A1=>nx8058);
   ix8061 : nor03_2x port map ( Y=>nx8060, A0=>nx8003, A1=>nx9451, A2=>
      nx10979);
   gen_20_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_20_cmp_mReg_14, QB=>
      nx8003, D=>window_20_14, CLK=>start, R=>rst);
   ix8059 : nor03_2x port map ( Y=>nx8058, A0=>gen_20_cmp_mReg_14, A1=>
      nx10121, A2=>nx10987);
   ix8095 : nand02 port map ( Y=>gen_20_cmp_BSCmp_op2_15, A0=>nx8009, A1=>
      nx8013);
   ix8010 : nor02_2x port map ( Y=>nx8009, A0=>nx8090, A1=>nx8086);
   ix8091 : nor03_2x port map ( Y=>nx8090, A0=>gen_20_cmp_mReg_14, A1=>
      nx9457, A2=>nx10955);
   ix8087 : nor03_2x port map ( Y=>nx8086, A0=>nx8003, A1=>nx10961, A2=>
      nx10971);
   ix8014 : nor02_2x port map ( Y=>nx8013, A0=>nx8082, A1=>nx8080);
   ix8083 : nor03_2x port map ( Y=>nx8082, A0=>nx8017, A1=>nx9451, A2=>
      nx10979);
   gen_20_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_20_cmp_mReg_15, QB=>
      nx8017, D=>window_20_15, CLK=>start, R=>rst);
   ix8081 : nor03_2x port map ( Y=>nx8080, A0=>gen_20_cmp_mReg_15, A1=>
      nx10123, A2=>nx10987);
   ix8105 : nand02 port map ( Y=>gen_20_cmp_BSCmp_op2_16, A0=>nx8023, A1=>
      nx8013);
   ix8024 : nor02_2x port map ( Y=>nx8023, A0=>nx8100, A1=>nx8096);
   ix8101 : nor03_2x port map ( Y=>nx8100, A0=>gen_20_cmp_mReg_15, A1=>
      nx9457, A2=>nx10955);
   ix8097 : nor03_2x port map ( Y=>nx8096, A0=>nx8017, A1=>nx10961, A2=>
      nx10971);
   ix8173 : nand02 port map ( Y=>gen_21_cmp_BSCmp_op2_1, A0=>nx8031, A1=>
      nx8049);
   ix8032 : nor02_2x port map ( Y=>nx8031, A0=>nx8168, A1=>nx8164);
   ix8169 : nor03_2x port map ( Y=>nx8168, A0=>gen_21_cmp_mReg_0, A1=>nx9441, 
      A2=>nx10991);
   gen_21_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_21_cmp_mReg_0, QB=>
      nx8035, D=>window_21_0, CLK=>start, R=>rst);
   ix8040 : inv01 port map ( Y=>nx8039, A=>gen_21_cmp_pMux_0);
   ix8165 : nor03_2x port map ( Y=>nx8164, A0=>nx8035, A1=>nx10997, A2=>
      nx11007);
   ix8048 : inv02 port map ( Y=>nx8047, A=>gen_21_cmp_pMux_2);
   ix8050 : nor02_2x port map ( Y=>nx8049, A0=>nx8154, A1=>nx8152);
   ix8155 : nor03_2x port map ( Y=>nx8154, A0=>nx8053, A1=>nx9435, A2=>
      nx11015);
   gen_21_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_21_cmp_mReg_1, QB=>
      nx8053, D=>window_21_1, CLK=>start, R=>rst);
   ix8153 : nor03_2x port map ( Y=>nx8152, A0=>gen_21_cmp_mReg_1, A1=>
      nx10125, A2=>nx11023);
   ix8113 : nor03_2x port map ( Y=>nx8112, A0=>nx9441, A1=>nx8047, A2=>
      gen_21_cmp_pMux_0);
   ix8195 : nand02 port map ( Y=>gen_21_cmp_BSCmp_op2_2, A0=>nx8065, A1=>
      nx8069);
   ix8066 : nor02_2x port map ( Y=>nx8065, A0=>nx8190, A1=>nx8186);
   ix8191 : nor03_2x port map ( Y=>nx8190, A0=>gen_21_cmp_mReg_1, A1=>nx9441, 
      A2=>nx10991);
   ix8187 : nor03_2x port map ( Y=>nx8186, A0=>nx8053, A1=>nx10997, A2=>
      nx11007);
   ix8070 : nor02_2x port map ( Y=>nx8069, A0=>nx8182, A1=>nx8180);
   ix8183 : nor03_2x port map ( Y=>nx8182, A0=>nx8073, A1=>nx9435, A2=>
      nx11015);
   gen_21_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_21_cmp_mReg_2, QB=>
      nx8073, D=>window_21_2, CLK=>start, R=>rst);
   ix8181 : nor03_2x port map ( Y=>nx8180, A0=>gen_21_cmp_mReg_2, A1=>
      nx10125, A2=>nx11023);
   ix8217 : nand02 port map ( Y=>gen_21_cmp_BSCmp_op2_3, A0=>nx8077, A1=>
      nx8083);
   ix8078 : nor02_2x port map ( Y=>nx8077, A0=>nx8212, A1=>nx8208);
   ix8213 : nor03_2x port map ( Y=>nx8212, A0=>gen_21_cmp_mReg_2, A1=>nx9441, 
      A2=>nx10991);
   ix8209 : nor03_2x port map ( Y=>nx8208, A0=>nx8073, A1=>nx10997, A2=>
      nx11007);
   ix8084 : nor02_2x port map ( Y=>nx8083, A0=>nx8204, A1=>nx8202);
   ix8205 : nor03_2x port map ( Y=>nx8204, A0=>nx8087, A1=>nx9435, A2=>
      nx11015);
   gen_21_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_21_cmp_mReg_3, QB=>
      nx8087, D=>window_21_3, CLK=>start, R=>rst);
   ix8203 : nor03_2x port map ( Y=>nx8202, A0=>gen_21_cmp_mReg_3, A1=>
      nx10125, A2=>nx11023);
   ix8239 : nand02 port map ( Y=>gen_21_cmp_BSCmp_op2_4, A0=>nx8091, A1=>
      nx8097);
   ix8092 : nor02_2x port map ( Y=>nx8091, A0=>nx8234, A1=>nx8230);
   ix8235 : nor03_2x port map ( Y=>nx8234, A0=>gen_21_cmp_mReg_3, A1=>nx9441, 
      A2=>nx10991);
   ix8231 : nor03_2x port map ( Y=>nx8230, A0=>nx8087, A1=>nx10997, A2=>
      nx11007);
   ix8098 : nor02_2x port map ( Y=>nx8097, A0=>nx8226, A1=>nx8224);
   ix8227 : nor03_2x port map ( Y=>nx8226, A0=>nx8101, A1=>nx9435, A2=>
      nx11015);
   gen_21_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_21_cmp_mReg_4, QB=>
      nx8101, D=>window_21_4, CLK=>start, R=>rst);
   ix8225 : nor03_2x port map ( Y=>nx8224, A0=>gen_21_cmp_mReg_4, A1=>
      nx10125, A2=>nx11023);
   ix8261 : nand02 port map ( Y=>gen_21_cmp_BSCmp_op2_5, A0=>nx8107, A1=>
      nx8113);
   ix8108 : nor02_2x port map ( Y=>nx8107, A0=>nx8256, A1=>nx8252);
   ix8257 : nor03_2x port map ( Y=>nx8256, A0=>gen_21_cmp_mReg_4, A1=>nx9441, 
      A2=>nx10991);
   ix8253 : nor03_2x port map ( Y=>nx8252, A0=>nx8101, A1=>nx10997, A2=>
      nx11007);
   ix8114 : nor02_2x port map ( Y=>nx8113, A0=>nx8248, A1=>nx8246);
   ix8249 : nor03_2x port map ( Y=>nx8248, A0=>nx8116, A1=>nx9437, A2=>
      nx11015);
   gen_21_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_21_cmp_mReg_5, QB=>
      nx8116, D=>window_21_5, CLK=>start, R=>rst);
   ix8247 : nor03_2x port map ( Y=>nx8246, A0=>gen_21_cmp_mReg_5, A1=>
      nx10125, A2=>nx11023);
   ix8283 : nand02 port map ( Y=>gen_21_cmp_BSCmp_op2_6, A0=>nx8120, A1=>
      nx8125);
   ix8121 : nor02_2x port map ( Y=>nx8120, A0=>nx8278, A1=>nx8274);
   ix8279 : nor03_2x port map ( Y=>nx8278, A0=>gen_21_cmp_mReg_5, A1=>nx9443, 
      A2=>nx10991);
   ix8275 : nor03_2x port map ( Y=>nx8274, A0=>nx8116, A1=>nx10997, A2=>
      nx11007);
   ix8126 : nor02_2x port map ( Y=>nx8125, A0=>nx8270, A1=>nx8268);
   ix8271 : nor03_2x port map ( Y=>nx8270, A0=>nx8129, A1=>nx9437, A2=>
      nx11015);
   gen_21_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_21_cmp_mReg_6, QB=>
      nx8129, D=>window_21_6, CLK=>start, R=>rst);
   ix8269 : nor03_2x port map ( Y=>nx8268, A0=>gen_21_cmp_mReg_6, A1=>
      nx10125, A2=>nx11023);
   ix8305 : nand02 port map ( Y=>gen_21_cmp_BSCmp_op2_7, A0=>nx8135, A1=>
      nx8141);
   ix8136 : nor02_2x port map ( Y=>nx8135, A0=>nx8300, A1=>nx8296);
   ix8301 : nor03_2x port map ( Y=>nx8300, A0=>gen_21_cmp_mReg_6, A1=>nx9443, 
      A2=>nx10993);
   ix8297 : nor03_2x port map ( Y=>nx8296, A0=>nx8129, A1=>nx10999, A2=>
      nx11009);
   ix8142 : nor02_2x port map ( Y=>nx8141, A0=>nx8292, A1=>nx8290);
   ix8293 : nor03_2x port map ( Y=>nx8292, A0=>nx8145, A1=>nx9437, A2=>
      nx11017);
   gen_21_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_21_cmp_mReg_7, QB=>
      nx8145, D=>window_21_7, CLK=>start, R=>rst);
   ix8291 : nor03_2x port map ( Y=>nx8290, A0=>gen_21_cmp_mReg_7, A1=>
      nx10125, A2=>nx11025);
   ix8327 : nand02 port map ( Y=>gen_21_cmp_BSCmp_op2_8, A0=>nx8149, A1=>
      nx8155);
   ix8150 : nor02_2x port map ( Y=>nx8149, A0=>nx8322, A1=>nx8318);
   ix8323 : nor03_2x port map ( Y=>nx8322, A0=>gen_21_cmp_mReg_7, A1=>nx9443, 
      A2=>nx10993);
   ix8319 : nor03_2x port map ( Y=>nx8318, A0=>nx8145, A1=>nx10999, A2=>
      nx11009);
   ix8156 : nor02_2x port map ( Y=>nx8155, A0=>nx8314, A1=>nx8312);
   ix8315 : nor03_2x port map ( Y=>nx8314, A0=>nx8159, A1=>nx9437, A2=>
      nx11017);
   gen_21_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_21_cmp_mReg_8, QB=>
      nx8159, D=>window_21_8, CLK=>start, R=>rst);
   ix8313 : nor03_2x port map ( Y=>nx8312, A0=>gen_21_cmp_mReg_8, A1=>
      nx10127, A2=>nx11025);
   ix8349 : nand02 port map ( Y=>gen_21_cmp_BSCmp_op2_9, A0=>nx8165, A1=>
      nx8169);
   ix8166 : nor02_2x port map ( Y=>nx8165, A0=>nx8344, A1=>nx8340);
   ix8345 : nor03_2x port map ( Y=>nx8344, A0=>gen_21_cmp_mReg_8, A1=>nx9443, 
      A2=>nx10993);
   ix8341 : nor03_2x port map ( Y=>nx8340, A0=>nx8159, A1=>nx10999, A2=>
      nx11009);
   ix8170 : nor02_2x port map ( Y=>nx8169, A0=>nx8336, A1=>nx8334);
   ix8337 : nor03_2x port map ( Y=>nx8336, A0=>nx8173, A1=>nx9437, A2=>
      nx11017);
   gen_21_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_21_cmp_mReg_9, QB=>
      nx8173, D=>window_21_9, CLK=>start, R=>rst);
   ix8335 : nor03_2x port map ( Y=>nx8334, A0=>gen_21_cmp_mReg_9, A1=>
      nx10127, A2=>nx11025);
   ix8371 : nand02 port map ( Y=>gen_21_cmp_BSCmp_op2_10, A0=>nx8177, A1=>
      nx8183);
   ix8178 : nor02_2x port map ( Y=>nx8177, A0=>nx8366, A1=>nx8362);
   ix8367 : nor03_2x port map ( Y=>nx8366, A0=>gen_21_cmp_mReg_9, A1=>nx9443, 
      A2=>nx10993);
   ix8363 : nor03_2x port map ( Y=>nx8362, A0=>nx8173, A1=>nx10999, A2=>
      nx11009);
   ix8184 : nor02_2x port map ( Y=>nx8183, A0=>nx8358, A1=>nx8356);
   ix8359 : nor03_2x port map ( Y=>nx8358, A0=>nx8187, A1=>nx9437, A2=>
      nx11017);
   gen_21_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_21_cmp_mReg_10, QB=>
      nx8187, D=>window_21_10, CLK=>start, R=>rst);
   ix8357 : nor03_2x port map ( Y=>nx8356, A0=>gen_21_cmp_mReg_10, A1=>
      nx10127, A2=>nx11025);
   ix8393 : nand02 port map ( Y=>gen_21_cmp_BSCmp_op2_11, A0=>nx8191, A1=>
      nx8197);
   ix8192 : nor02_2x port map ( Y=>nx8191, A0=>nx8388, A1=>nx8384);
   ix8389 : nor03_2x port map ( Y=>nx8388, A0=>gen_21_cmp_mReg_10, A1=>
      nx9443, A2=>nx10993);
   ix8385 : nor03_2x port map ( Y=>nx8384, A0=>nx8187, A1=>nx10999, A2=>
      nx11009);
   ix8198 : nor02_2x port map ( Y=>nx8197, A0=>nx8380, A1=>nx8378);
   ix8381 : nor03_2x port map ( Y=>nx8380, A0=>nx8200, A1=>nx9437, A2=>
      nx11017);
   gen_21_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_21_cmp_mReg_11, QB=>
      nx8200, D=>window_21_11, CLK=>start, R=>rst);
   ix8379 : nor03_2x port map ( Y=>nx8378, A0=>gen_21_cmp_mReg_11, A1=>
      nx10127, A2=>nx11025);
   ix8415 : nand02 port map ( Y=>gen_21_cmp_BSCmp_op2_12, A0=>nx8207, A1=>
      nx8213);
   ix8208 : nor02_2x port map ( Y=>nx8207, A0=>nx8410, A1=>nx8406);
   ix8411 : nor03_2x port map ( Y=>nx8410, A0=>gen_21_cmp_mReg_11, A1=>
      nx9443, A2=>nx10993);
   ix8407 : nor03_2x port map ( Y=>nx8406, A0=>nx8200, A1=>nx10999, A2=>
      nx11009);
   ix8214 : nor02_2x port map ( Y=>nx8213, A0=>nx8402, A1=>nx8400);
   ix8403 : nor03_2x port map ( Y=>nx8402, A0=>nx8217, A1=>nx9439, A2=>
      nx11017);
   gen_21_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_21_cmp_mReg_12, QB=>
      nx8217, D=>window_21_12, CLK=>start, R=>rst);
   ix8401 : nor03_2x port map ( Y=>nx8400, A0=>gen_21_cmp_mReg_12, A1=>
      nx10127, A2=>nx11025);
   ix8437 : nand02 port map ( Y=>gen_21_cmp_BSCmp_op2_13, A0=>nx8221, A1=>
      nx8227);
   ix8222 : nor02_2x port map ( Y=>nx8221, A0=>nx8432, A1=>nx8428);
   ix8433 : nor03_2x port map ( Y=>nx8432, A0=>gen_21_cmp_mReg_12, A1=>
      nx9445, A2=>nx10995);
   ix8429 : nor03_2x port map ( Y=>nx8428, A0=>nx8217, A1=>nx10999, A2=>
      nx11011);
   ix8228 : nor02_2x port map ( Y=>nx8227, A0=>nx8424, A1=>nx8422);
   ix8425 : nor03_2x port map ( Y=>nx8424, A0=>nx8231, A1=>nx9439, A2=>
      nx11019);
   gen_21_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_21_cmp_mReg_13, QB=>
      nx8231, D=>window_21_13, CLK=>start, R=>rst);
   ix8423 : nor03_2x port map ( Y=>nx8422, A0=>gen_21_cmp_mReg_13, A1=>
      nx10127, A2=>nx11027);
   ix8459 : nand02 port map ( Y=>gen_21_cmp_BSCmp_op2_14, A0=>nx8235, A1=>
      nx8241);
   ix8236 : nor02_2x port map ( Y=>nx8235, A0=>nx8454, A1=>nx8450);
   ix8455 : nor03_2x port map ( Y=>nx8454, A0=>gen_21_cmp_mReg_13, A1=>
      nx9445, A2=>nx10995);
   ix8451 : nor03_2x port map ( Y=>nx8450, A0=>nx8231, A1=>nx11001, A2=>
      nx11011);
   ix8242 : nor02_2x port map ( Y=>nx8241, A0=>nx8446, A1=>nx8444);
   ix8447 : nor03_2x port map ( Y=>nx8446, A0=>nx8244, A1=>nx9439, A2=>
      nx11019);
   gen_21_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_21_cmp_mReg_14, QB=>
      nx8244, D=>window_21_14, CLK=>start, R=>rst);
   ix8445 : nor03_2x port map ( Y=>nx8444, A0=>gen_21_cmp_mReg_14, A1=>
      nx10127, A2=>nx11027);
   ix8481 : nand02 port map ( Y=>gen_21_cmp_BSCmp_op2_15, A0=>nx8251, A1=>
      nx8257);
   ix8252 : nor02_2x port map ( Y=>nx8251, A0=>nx8476, A1=>nx8472);
   ix8477 : nor03_2x port map ( Y=>nx8476, A0=>gen_21_cmp_mReg_14, A1=>
      nx9445, A2=>nx10995);
   ix8473 : nor03_2x port map ( Y=>nx8472, A0=>nx8244, A1=>nx11001, A2=>
      nx11011);
   ix8258 : nor02_2x port map ( Y=>nx8257, A0=>nx8468, A1=>nx8466);
   ix8469 : nor03_2x port map ( Y=>nx8468, A0=>nx8261, A1=>nx9439, A2=>
      nx11019);
   gen_21_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_21_cmp_mReg_15, QB=>
      nx8261, D=>window_21_15, CLK=>start, R=>rst);
   ix8467 : nor03_2x port map ( Y=>nx8466, A0=>gen_21_cmp_mReg_15, A1=>
      nx10129, A2=>nx11027);
   ix8491 : nand02 port map ( Y=>gen_21_cmp_BSCmp_op2_16, A0=>nx8265, A1=>
      nx8257);
   ix8266 : nor02_2x port map ( Y=>nx8265, A0=>nx8486, A1=>nx8482);
   ix8487 : nor03_2x port map ( Y=>nx8486, A0=>gen_21_cmp_mReg_15, A1=>
      nx9445, A2=>nx10995);
   ix8483 : nor03_2x port map ( Y=>nx8482, A0=>nx8261, A1=>nx11001, A2=>
      nx11011);
   ix8559 : nand02 port map ( Y=>gen_22_cmp_BSCmp_op2_1, A0=>nx8273, A1=>
      nx8293);
   ix8274 : nor02_2x port map ( Y=>nx8273, A0=>nx8554, A1=>nx8550);
   ix8555 : nor03_2x port map ( Y=>nx8554, A0=>gen_22_cmp_mReg_0, A1=>nx9429, 
      A2=>nx11031);
   gen_22_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_22_cmp_mReg_0, QB=>
      nx8279, D=>window_22_0, CLK=>start, R=>rst);
   ix8284 : inv01 port map ( Y=>nx8283, A=>gen_22_cmp_pMux_0);
   ix8551 : nor03_2x port map ( Y=>nx8550, A0=>nx8279, A1=>nx11037, A2=>
      nx11047);
   ix8292 : inv02 port map ( Y=>nx8291, A=>gen_22_cmp_pMux_2);
   ix8294 : nor02_2x port map ( Y=>nx8293, A0=>nx8540, A1=>nx8538);
   ix8541 : nor03_2x port map ( Y=>nx8540, A0=>nx8297, A1=>nx9423, A2=>
      nx11055);
   gen_22_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_22_cmp_mReg_1, QB=>
      nx8297, D=>window_22_1, CLK=>start, R=>rst);
   ix8539 : nor03_2x port map ( Y=>nx8538, A0=>gen_22_cmp_mReg_1, A1=>
      nx10131, A2=>nx11063);
   ix8499 : nor03_2x port map ( Y=>nx8498, A0=>nx9429, A1=>nx8291, A2=>
      gen_22_cmp_pMux_0);
   ix8581 : nand02 port map ( Y=>gen_22_cmp_BSCmp_op2_2, A0=>nx8308, A1=>
      nx8313);
   ix8309 : nor02_2x port map ( Y=>nx8308, A0=>nx8576, A1=>nx8572);
   ix8577 : nor03_2x port map ( Y=>nx8576, A0=>gen_22_cmp_mReg_1, A1=>nx9429, 
      A2=>nx11031);
   ix8573 : nor03_2x port map ( Y=>nx8572, A0=>nx8297, A1=>nx11037, A2=>
      nx11047);
   ix8314 : nor02_2x port map ( Y=>nx8313, A0=>nx8568, A1=>nx8566);
   ix8569 : nor03_2x port map ( Y=>nx8568, A0=>nx8317, A1=>nx9423, A2=>
      nx11055);
   gen_22_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_22_cmp_mReg_2, QB=>
      nx8317, D=>window_22_2, CLK=>start, R=>rst);
   ix8567 : nor03_2x port map ( Y=>nx8566, A0=>gen_22_cmp_mReg_2, A1=>
      nx10131, A2=>nx11063);
   ix8603 : nand02 port map ( Y=>gen_22_cmp_BSCmp_op2_3, A0=>nx8323, A1=>
      nx8329);
   ix8324 : nor02_2x port map ( Y=>nx8323, A0=>nx8598, A1=>nx8594);
   ix8599 : nor03_2x port map ( Y=>nx8598, A0=>gen_22_cmp_mReg_2, A1=>nx9429, 
      A2=>nx11031);
   ix8595 : nor03_2x port map ( Y=>nx8594, A0=>nx8317, A1=>nx11037, A2=>
      nx11047);
   ix8330 : nor02_2x port map ( Y=>nx8329, A0=>nx8590, A1=>nx8588);
   ix8591 : nor03_2x port map ( Y=>nx8590, A0=>nx8332, A1=>nx9423, A2=>
      nx11055);
   gen_22_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_22_cmp_mReg_3, QB=>
      nx8332, D=>window_22_3, CLK=>start, R=>rst);
   ix8589 : nor03_2x port map ( Y=>nx8588, A0=>gen_22_cmp_mReg_3, A1=>
      nx10131, A2=>nx11063);
   ix8625 : nand02 port map ( Y=>gen_22_cmp_BSCmp_op2_4, A0=>nx8339, A1=>
      nx8345);
   ix8340 : nor02_2x port map ( Y=>nx8339, A0=>nx8620, A1=>nx8616);
   ix8621 : nor03_2x port map ( Y=>nx8620, A0=>gen_22_cmp_mReg_3, A1=>nx9429, 
      A2=>nx11031);
   ix8617 : nor03_2x port map ( Y=>nx8616, A0=>nx8332, A1=>nx11037, A2=>
      nx11047);
   ix8346 : nor02_2x port map ( Y=>nx8345, A0=>nx8612, A1=>nx8610);
   ix8613 : nor03_2x port map ( Y=>nx8612, A0=>nx8349, A1=>nx9423, A2=>
      nx11055);
   gen_22_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_22_cmp_mReg_4, QB=>
      nx8349, D=>window_22_4, CLK=>start, R=>rst);
   ix8611 : nor03_2x port map ( Y=>nx8610, A0=>gen_22_cmp_mReg_4, A1=>
      nx10131, A2=>nx11063);
   ix8647 : nand02 port map ( Y=>gen_22_cmp_BSCmp_op2_5, A0=>nx8353, A1=>
      nx8359);
   ix8354 : nor02_2x port map ( Y=>nx8353, A0=>nx8642, A1=>nx8638);
   ix8643 : nor03_2x port map ( Y=>nx8642, A0=>gen_22_cmp_mReg_4, A1=>nx9429, 
      A2=>nx11031);
   ix8639 : nor03_2x port map ( Y=>nx8638, A0=>nx8349, A1=>nx11037, A2=>
      nx11047);
   ix8360 : nor02_2x port map ( Y=>nx8359, A0=>nx8634, A1=>nx8632);
   ix8635 : nor03_2x port map ( Y=>nx8634, A0=>nx8363, A1=>nx9425, A2=>
      nx11055);
   gen_22_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_22_cmp_mReg_5, QB=>
      nx8363, D=>window_22_5, CLK=>start, R=>rst);
   ix8633 : nor03_2x port map ( Y=>nx8632, A0=>gen_22_cmp_mReg_5, A1=>
      nx10131, A2=>nx11063);
   ix8669 : nand02 port map ( Y=>gen_22_cmp_BSCmp_op2_6, A0=>nx8367, A1=>
      nx8373);
   ix8368 : nor02_2x port map ( Y=>nx8367, A0=>nx8664, A1=>nx8660);
   ix8665 : nor03_2x port map ( Y=>nx8664, A0=>gen_22_cmp_mReg_5, A1=>nx9431, 
      A2=>nx11031);
   ix8661 : nor03_2x port map ( Y=>nx8660, A0=>nx8363, A1=>nx11037, A2=>
      nx11047);
   ix8374 : nor02_2x port map ( Y=>nx8373, A0=>nx8656, A1=>nx8654);
   ix8657 : nor03_2x port map ( Y=>nx8656, A0=>nx8376, A1=>nx9425, A2=>
      nx11055);
   gen_22_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_22_cmp_mReg_6, QB=>
      nx8376, D=>window_22_6, CLK=>start, R=>rst);
   ix8655 : nor03_2x port map ( Y=>nx8654, A0=>gen_22_cmp_mReg_6, A1=>
      nx10131, A2=>nx11063);
   ix8691 : nand02 port map ( Y=>gen_22_cmp_BSCmp_op2_7, A0=>nx8383, A1=>
      nx8389);
   ix8384 : nor02_2x port map ( Y=>nx8383, A0=>nx8686, A1=>nx8682);
   ix8687 : nor03_2x port map ( Y=>nx8686, A0=>gen_22_cmp_mReg_6, A1=>nx9431, 
      A2=>nx11033);
   ix8683 : nor03_2x port map ( Y=>nx8682, A0=>nx8376, A1=>nx11039, A2=>
      nx11049);
   ix8390 : nor02_2x port map ( Y=>nx8389, A0=>nx8678, A1=>nx8676);
   ix8679 : nor03_2x port map ( Y=>nx8678, A0=>nx8393, A1=>nx9425, A2=>
      nx11057);
   gen_22_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_22_cmp_mReg_7, QB=>
      nx8393, D=>window_22_7, CLK=>start, R=>rst);
   ix8677 : nor03_2x port map ( Y=>nx8676, A0=>gen_22_cmp_mReg_7, A1=>
      nx10131, A2=>nx11065);
   ix8713 : nand02 port map ( Y=>gen_22_cmp_BSCmp_op2_8, A0=>nx8397, A1=>
      nx8403);
   ix8398 : nor02_2x port map ( Y=>nx8397, A0=>nx8708, A1=>nx8704);
   ix8709 : nor03_2x port map ( Y=>nx8708, A0=>gen_22_cmp_mReg_7, A1=>nx9431, 
      A2=>nx11033);
   ix8705 : nor03_2x port map ( Y=>nx8704, A0=>nx8393, A1=>nx11039, A2=>
      nx11049);
   ix8404 : nor02_2x port map ( Y=>nx8403, A0=>nx8700, A1=>nx8698);
   ix8701 : nor03_2x port map ( Y=>nx8700, A0=>nx8407, A1=>nx9425, A2=>
      nx11057);
   gen_22_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_22_cmp_mReg_8, QB=>
      nx8407, D=>window_22_8, CLK=>start, R=>rst);
   ix8699 : nor03_2x port map ( Y=>nx8698, A0=>gen_22_cmp_mReg_8, A1=>
      nx10133, A2=>nx11065);
   ix8735 : nand02 port map ( Y=>gen_22_cmp_BSCmp_op2_9, A0=>nx8411, A1=>
      nx8417);
   ix8412 : nor02_2x port map ( Y=>nx8411, A0=>nx8730, A1=>nx8726);
   ix8731 : nor03_2x port map ( Y=>nx8730, A0=>gen_22_cmp_mReg_8, A1=>nx9431, 
      A2=>nx11033);
   ix8727 : nor03_2x port map ( Y=>nx8726, A0=>nx8407, A1=>nx11039, A2=>
      nx11049);
   ix8418 : nor02_2x port map ( Y=>nx8417, A0=>nx8722, A1=>nx8720);
   ix8723 : nor03_2x port map ( Y=>nx8722, A0=>nx8420, A1=>nx9425, A2=>
      nx11057);
   gen_22_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_22_cmp_mReg_9, QB=>
      nx8420, D=>window_22_9, CLK=>start, R=>rst);
   ix8721 : nor03_2x port map ( Y=>nx8720, A0=>gen_22_cmp_mReg_9, A1=>
      nx10133, A2=>nx11065);
   ix8757 : nand02 port map ( Y=>gen_22_cmp_BSCmp_op2_10, A0=>nx8427, A1=>
      nx8433);
   ix8428 : nor02_2x port map ( Y=>nx8427, A0=>nx8752, A1=>nx8748);
   ix8753 : nor03_2x port map ( Y=>nx8752, A0=>gen_22_cmp_mReg_9, A1=>nx9431, 
      A2=>nx11033);
   ix8749 : nor03_2x port map ( Y=>nx8748, A0=>nx8420, A1=>nx11039, A2=>
      nx11049);
   ix8434 : nor02_2x port map ( Y=>nx8433, A0=>nx8744, A1=>nx8742);
   ix8745 : nor03_2x port map ( Y=>nx8744, A0=>nx8437, A1=>nx9425, A2=>
      nx11057);
   gen_22_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_22_cmp_mReg_10, QB=>
      nx8437, D=>window_22_10, CLK=>start, R=>rst);
   ix8743 : nor03_2x port map ( Y=>nx8742, A0=>gen_22_cmp_mReg_10, A1=>
      nx10133, A2=>nx11065);
   ix8779 : nand02 port map ( Y=>gen_22_cmp_BSCmp_op2_11, A0=>nx8441, A1=>
      nx8447);
   ix8442 : nor02_2x port map ( Y=>nx8441, A0=>nx8774, A1=>nx8770);
   ix8775 : nor03_2x port map ( Y=>nx8774, A0=>gen_22_cmp_mReg_10, A1=>
      nx9431, A2=>nx11033);
   ix8771 : nor03_2x port map ( Y=>nx8770, A0=>nx8437, A1=>nx11039, A2=>
      nx11049);
   ix8448 : nor02_2x port map ( Y=>nx8447, A0=>nx8766, A1=>nx8764);
   ix8767 : nor03_2x port map ( Y=>nx8766, A0=>nx8451, A1=>nx9425, A2=>
      nx11057);
   gen_22_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_22_cmp_mReg_11, QB=>
      nx8451, D=>window_22_11, CLK=>start, R=>rst);
   ix8765 : nor03_2x port map ( Y=>nx8764, A0=>gen_22_cmp_mReg_11, A1=>
      nx10133, A2=>nx11065);
   ix8801 : nand02 port map ( Y=>gen_22_cmp_BSCmp_op2_12, A0=>nx8455, A1=>
      nx8461);
   ix8456 : nor02_2x port map ( Y=>nx8455, A0=>nx8796, A1=>nx8792);
   ix8797 : nor03_2x port map ( Y=>nx8796, A0=>gen_22_cmp_mReg_11, A1=>
      nx9431, A2=>nx11033);
   ix8793 : nor03_2x port map ( Y=>nx8792, A0=>nx8451, A1=>nx11039, A2=>
      nx11049);
   ix8462 : nor02_2x port map ( Y=>nx8461, A0=>nx8788, A1=>nx8786);
   ix8789 : nor03_2x port map ( Y=>nx8788, A0=>nx8464, A1=>nx9427, A2=>
      nx11057);
   gen_22_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_22_cmp_mReg_12, QB=>
      nx8464, D=>window_22_12, CLK=>start, R=>rst);
   ix8787 : nor03_2x port map ( Y=>nx8786, A0=>gen_22_cmp_mReg_12, A1=>
      nx10133, A2=>nx11065);
   ix8823 : nand02 port map ( Y=>gen_22_cmp_BSCmp_op2_13, A0=>nx8471, A1=>
      nx8477);
   ix8472 : nor02_2x port map ( Y=>nx8471, A0=>nx8818, A1=>nx8814);
   ix8819 : nor03_2x port map ( Y=>nx8818, A0=>gen_22_cmp_mReg_12, A1=>
      nx9433, A2=>nx11035);
   ix8815 : nor03_2x port map ( Y=>nx8814, A0=>nx8464, A1=>nx11039, A2=>
      nx11051);
   ix8478 : nor02_2x port map ( Y=>nx8477, A0=>nx8810, A1=>nx8808);
   ix8811 : nor03_2x port map ( Y=>nx8810, A0=>nx8481, A1=>nx9427, A2=>
      nx11059);
   gen_22_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_22_cmp_mReg_13, QB=>
      nx8481, D=>window_22_13, CLK=>start, R=>rst);
   ix8809 : nor03_2x port map ( Y=>nx8808, A0=>gen_22_cmp_mReg_13, A1=>
      nx10133, A2=>nx11067);
   ix8845 : nand02 port map ( Y=>gen_22_cmp_BSCmp_op2_14, A0=>nx8487, A1=>
      nx8493);
   ix8488 : nor02_2x port map ( Y=>nx8487, A0=>nx8840, A1=>nx8836);
   ix8841 : nor03_2x port map ( Y=>nx8840, A0=>gen_22_cmp_mReg_13, A1=>
      nx9433, A2=>nx11035);
   ix8837 : nor03_2x port map ( Y=>nx8836, A0=>nx8481, A1=>nx11041, A2=>
      nx11051);
   ix8494 : nor02_2x port map ( Y=>nx8493, A0=>nx8832, A1=>nx8830);
   ix8833 : nor03_2x port map ( Y=>nx8832, A0=>nx8497, A1=>nx9427, A2=>
      nx11059);
   gen_22_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_22_cmp_mReg_14, QB=>
      nx8497, D=>window_22_14, CLK=>start, R=>rst);
   ix8831 : nor03_2x port map ( Y=>nx8830, A0=>gen_22_cmp_mReg_14, A1=>
      nx10133, A2=>nx11067);
   ix8867 : nand02 port map ( Y=>gen_22_cmp_BSCmp_op2_15, A0=>nx8502, A1=>
      nx8506);
   ix8503 : nor02_2x port map ( Y=>nx8502, A0=>nx8862, A1=>nx8858);
   ix8863 : nor03_2x port map ( Y=>nx8862, A0=>gen_22_cmp_mReg_14, A1=>
      nx9433, A2=>nx11035);
   ix8859 : nor03_2x port map ( Y=>nx8858, A0=>nx8497, A1=>nx11041, A2=>
      nx11051);
   ix8507 : nor02_2x port map ( Y=>nx8506, A0=>nx8854, A1=>nx8852);
   ix8855 : nor03_2x port map ( Y=>nx8854, A0=>nx8509, A1=>nx9427, A2=>
      nx11059);
   gen_22_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_22_cmp_mReg_15, QB=>
      nx8509, D=>window_22_15, CLK=>start, R=>rst);
   ix8853 : nor03_2x port map ( Y=>nx8852, A0=>gen_22_cmp_mReg_15, A1=>
      nx10135, A2=>nx11067);
   ix8877 : nand02 port map ( Y=>gen_22_cmp_BSCmp_op2_16, A0=>nx8515, A1=>
      nx8506);
   ix8516 : nor02_2x port map ( Y=>nx8515, A0=>nx8872, A1=>nx8868);
   ix8873 : nor03_2x port map ( Y=>nx8872, A0=>gen_22_cmp_mReg_15, A1=>
      nx9433, A2=>nx11035);
   ix8869 : nor03_2x port map ( Y=>nx8868, A0=>nx8509, A1=>nx11041, A2=>
      nx11051);
   ix8945 : nand02 port map ( Y=>gen_23_cmp_BSCmp_op2_1, A0=>nx8523, A1=>
      nx8543);
   ix8524 : nor02_2x port map ( Y=>nx8523, A0=>nx8940, A1=>nx8936);
   ix8941 : nor03_2x port map ( Y=>nx8940, A0=>gen_23_cmp_mReg_0, A1=>nx9417, 
      A2=>nx11071);
   gen_23_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_23_cmp_mReg_0, QB=>
      nx8529, D=>window_23_0, CLK=>start, R=>rst);
   ix8534 : inv01 port map ( Y=>nx8533, A=>gen_23_cmp_pMux_0);
   ix8937 : nor03_2x port map ( Y=>nx8936, A0=>nx8529, A1=>nx11077, A2=>
      nx11087);
   ix8542 : inv02 port map ( Y=>nx8541, A=>gen_23_cmp_pMux_2);
   ix8544 : nor02_2x port map ( Y=>nx8543, A0=>nx8926, A1=>nx8924);
   ix8927 : nor03_2x port map ( Y=>nx8926, A0=>nx8547, A1=>nx9411, A2=>
      nx11095);
   gen_23_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_23_cmp_mReg_1, QB=>
      nx8547, D=>window_23_1, CLK=>start, R=>rst);
   ix8925 : nor03_2x port map ( Y=>nx8924, A0=>gen_23_cmp_mReg_1, A1=>
      nx10137, A2=>nx11103);
   ix8885 : nor03_2x port map ( Y=>nx8884, A0=>nx9417, A1=>nx8541, A2=>
      gen_23_cmp_pMux_0);
   ix8967 : nand02 port map ( Y=>gen_23_cmp_BSCmp_op2_2, A0=>nx8559, A1=>
      nx8563);
   ix8560 : nor02_2x port map ( Y=>nx8559, A0=>nx8962, A1=>nx8958);
   ix8963 : nor03_2x port map ( Y=>nx8962, A0=>gen_23_cmp_mReg_1, A1=>nx9417, 
      A2=>nx11071);
   ix8959 : nor03_2x port map ( Y=>nx8958, A0=>nx8547, A1=>nx11077, A2=>
      nx11087);
   ix8564 : nor02_2x port map ( Y=>nx8563, A0=>nx8954, A1=>nx8952);
   ix8955 : nor03_2x port map ( Y=>nx8954, A0=>nx8567, A1=>nx9411, A2=>
      nx11095);
   gen_23_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_23_cmp_mReg_2, QB=>
      nx8567, D=>window_23_2, CLK=>start, R=>rst);
   ix8953 : nor03_2x port map ( Y=>nx8952, A0=>gen_23_cmp_mReg_2, A1=>
      nx10137, A2=>nx11103);
   ix8989 : nand02 port map ( Y=>gen_23_cmp_BSCmp_op2_3, A0=>nx8573, A1=>
      nx8577);
   ix8574 : nor02_2x port map ( Y=>nx8573, A0=>nx8984, A1=>nx8980);
   ix8985 : nor03_2x port map ( Y=>nx8984, A0=>gen_23_cmp_mReg_2, A1=>nx9417, 
      A2=>nx11071);
   ix8981 : nor03_2x port map ( Y=>nx8980, A0=>nx8567, A1=>nx11077, A2=>
      nx11087);
   ix8578 : nor02_2x port map ( Y=>nx8577, A0=>nx8976, A1=>nx8974);
   ix8977 : nor03_2x port map ( Y=>nx8976, A0=>nx8581, A1=>nx9411, A2=>
      nx11095);
   gen_23_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_23_cmp_mReg_3, QB=>
      nx8581, D=>window_23_3, CLK=>start, R=>rst);
   ix8975 : nor03_2x port map ( Y=>nx8974, A0=>gen_23_cmp_mReg_3, A1=>
      nx10137, A2=>nx11103);
   ix9011 : nand02 port map ( Y=>gen_23_cmp_BSCmp_op2_4, A0=>nx8585, A1=>
      nx8591);
   ix8586 : nor02_2x port map ( Y=>nx8585, A0=>nx9006, A1=>nx9002);
   ix9007 : nor03_2x port map ( Y=>nx9006, A0=>gen_23_cmp_mReg_3, A1=>nx9417, 
      A2=>nx11071);
   ix9003 : nor03_2x port map ( Y=>nx9002, A0=>nx8581, A1=>nx11077, A2=>
      nx11087);
   ix8592 : nor02_2x port map ( Y=>nx8591, A0=>nx8998, A1=>nx8996);
   ix8999 : nor03_2x port map ( Y=>nx8998, A0=>nx8595, A1=>nx9411, A2=>
      nx11095);
   gen_23_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_23_cmp_mReg_4, QB=>
      nx8595, D=>window_23_4, CLK=>start, R=>rst);
   ix8997 : nor03_2x port map ( Y=>nx8996, A0=>gen_23_cmp_mReg_4, A1=>
      nx10137, A2=>nx11103);
   ix9033 : nand02 port map ( Y=>gen_23_cmp_BSCmp_op2_5, A0=>nx8599, A1=>
      nx8605);
   ix8600 : nor02_2x port map ( Y=>nx8599, A0=>nx9028, A1=>nx9024);
   ix9029 : nor03_2x port map ( Y=>nx9028, A0=>gen_23_cmp_mReg_4, A1=>nx9417, 
      A2=>nx11071);
   ix9025 : nor03_2x port map ( Y=>nx9024, A0=>nx8595, A1=>nx11077, A2=>
      nx11087);
   ix8606 : nor02_2x port map ( Y=>nx8605, A0=>nx9020, A1=>nx9018);
   ix9021 : nor03_2x port map ( Y=>nx9020, A0=>nx8608, A1=>nx9413, A2=>
      nx11095);
   gen_23_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_23_cmp_mReg_5, QB=>
      nx8608, D=>window_23_5, CLK=>start, R=>rst);
   ix9019 : nor03_2x port map ( Y=>nx9018, A0=>gen_23_cmp_mReg_5, A1=>
      nx10137, A2=>nx11103);
   ix9055 : nand02 port map ( Y=>gen_23_cmp_BSCmp_op2_6, A0=>nx8615, A1=>
      nx8621);
   ix8616 : nor02_2x port map ( Y=>nx8615, A0=>nx9050, A1=>nx9046);
   ix9051 : nor03_2x port map ( Y=>nx9050, A0=>gen_23_cmp_mReg_5, A1=>nx9419, 
      A2=>nx11071);
   ix9047 : nor03_2x port map ( Y=>nx9046, A0=>nx8608, A1=>nx11077, A2=>
      nx11087);
   ix8622 : nor02_2x port map ( Y=>nx8621, A0=>nx9042, A1=>nx9040);
   ix9043 : nor03_2x port map ( Y=>nx9042, A0=>nx8625, A1=>nx9413, A2=>
      nx11095);
   gen_23_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_23_cmp_mReg_6, QB=>
      nx8625, D=>window_23_6, CLK=>start, R=>rst);
   ix9041 : nor03_2x port map ( Y=>nx9040, A0=>gen_23_cmp_mReg_6, A1=>
      nx10137, A2=>nx11103);
   ix9077 : nand02 port map ( Y=>gen_23_cmp_BSCmp_op2_7, A0=>nx8629, A1=>
      nx8635);
   ix8630 : nor02_2x port map ( Y=>nx8629, A0=>nx9072, A1=>nx9068);
   ix9073 : nor03_2x port map ( Y=>nx9072, A0=>gen_23_cmp_mReg_6, A1=>nx9419, 
      A2=>nx11073);
   ix9069 : nor03_2x port map ( Y=>nx9068, A0=>nx8625, A1=>nx11079, A2=>
      nx11089);
   ix8636 : nor02_2x port map ( Y=>nx8635, A0=>nx9064, A1=>nx9062);
   ix9065 : nor03_2x port map ( Y=>nx9064, A0=>nx8639, A1=>nx9413, A2=>
      nx11097);
   gen_23_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_23_cmp_mReg_7, QB=>
      nx8639, D=>window_23_7, CLK=>start, R=>rst);
   ix9063 : nor03_2x port map ( Y=>nx9062, A0=>gen_23_cmp_mReg_7, A1=>
      nx10137, A2=>nx11105);
   ix9099 : nand02 port map ( Y=>gen_23_cmp_BSCmp_op2_8, A0=>nx8643, A1=>
      nx8649);
   ix8644 : nor02_2x port map ( Y=>nx8643, A0=>nx9094, A1=>nx9090);
   ix9095 : nor03_2x port map ( Y=>nx9094, A0=>gen_23_cmp_mReg_7, A1=>nx9419, 
      A2=>nx11073);
   ix9091 : nor03_2x port map ( Y=>nx9090, A0=>nx8639, A1=>nx11079, A2=>
      nx11089);
   ix8650 : nor02_2x port map ( Y=>nx8649, A0=>nx9086, A1=>nx9084);
   ix9087 : nor03_2x port map ( Y=>nx9086, A0=>nx8652, A1=>nx9413, A2=>
      nx11097);
   gen_23_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_23_cmp_mReg_8, QB=>
      nx8652, D=>window_23_8, CLK=>start, R=>rst);
   ix9085 : nor03_2x port map ( Y=>nx9084, A0=>gen_23_cmp_mReg_8, A1=>
      nx10139, A2=>nx11105);
   ix9121 : nand02 port map ( Y=>gen_23_cmp_BSCmp_op2_9, A0=>nx8659, A1=>
      nx8665);
   ix8660 : nor02_2x port map ( Y=>nx8659, A0=>nx9116, A1=>nx9112);
   ix9117 : nor03_2x port map ( Y=>nx9116, A0=>gen_23_cmp_mReg_8, A1=>nx9419, 
      A2=>nx11073);
   ix9113 : nor03_2x port map ( Y=>nx9112, A0=>nx8652, A1=>nx11079, A2=>
      nx11089);
   ix8666 : nor02_2x port map ( Y=>nx8665, A0=>nx9108, A1=>nx9106);
   ix9109 : nor03_2x port map ( Y=>nx9108, A0=>nx8669, A1=>nx9413, A2=>
      nx11097);
   gen_23_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_23_cmp_mReg_9, QB=>
      nx8669, D=>window_23_9, CLK=>start, R=>rst);
   ix9107 : nor03_2x port map ( Y=>nx9106, A0=>gen_23_cmp_mReg_9, A1=>
      nx10139, A2=>nx11105);
   ix9143 : nand02 port map ( Y=>gen_23_cmp_BSCmp_op2_10, A0=>nx8673, A1=>
      nx8679);
   ix8674 : nor02_2x port map ( Y=>nx8673, A0=>nx9138, A1=>nx9134);
   ix9139 : nor03_2x port map ( Y=>nx9138, A0=>gen_23_cmp_mReg_9, A1=>nx9419, 
      A2=>nx11073);
   ix9135 : nor03_2x port map ( Y=>nx9134, A0=>nx8669, A1=>nx11079, A2=>
      nx11089);
   ix8680 : nor02_2x port map ( Y=>nx8679, A0=>nx9130, A1=>nx9128);
   ix9131 : nor03_2x port map ( Y=>nx9130, A0=>nx8683, A1=>nx9413, A2=>
      nx11097);
   gen_23_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_23_cmp_mReg_10, QB=>
      nx8683, D=>window_23_10, CLK=>start, R=>rst);
   ix9129 : nor03_2x port map ( Y=>nx9128, A0=>gen_23_cmp_mReg_10, A1=>
      nx10139, A2=>nx11105);
   ix9165 : nand02 port map ( Y=>gen_23_cmp_BSCmp_op2_11, A0=>nx8687, A1=>
      nx8693);
   ix8688 : nor02_2x port map ( Y=>nx8687, A0=>nx9160, A1=>nx9156);
   ix9161 : nor03_2x port map ( Y=>nx9160, A0=>gen_23_cmp_mReg_10, A1=>
      nx9419, A2=>nx11073);
   ix9157 : nor03_2x port map ( Y=>nx9156, A0=>nx8683, A1=>nx11079, A2=>
      nx11089);
   ix8694 : nor02_2x port map ( Y=>nx8693, A0=>nx9152, A1=>nx9150);
   ix9153 : nor03_2x port map ( Y=>nx9152, A0=>nx8696, A1=>nx9413, A2=>
      nx11097);
   gen_23_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_23_cmp_mReg_11, QB=>
      nx8696, D=>window_23_11, CLK=>start, R=>rst);
   ix9151 : nor03_2x port map ( Y=>nx9150, A0=>gen_23_cmp_mReg_11, A1=>
      nx10139, A2=>nx11105);
   ix9187 : nand02 port map ( Y=>gen_23_cmp_BSCmp_op2_12, A0=>nx8703, A1=>
      nx8709);
   ix8704 : nor02_2x port map ( Y=>nx8703, A0=>nx9182, A1=>nx9178);
   ix9183 : nor03_2x port map ( Y=>nx9182, A0=>gen_23_cmp_mReg_11, A1=>
      nx9419, A2=>nx11073);
   ix9179 : nor03_2x port map ( Y=>nx9178, A0=>nx8696, A1=>nx11079, A2=>
      nx11089);
   ix8710 : nor02_2x port map ( Y=>nx8709, A0=>nx9174, A1=>nx9172);
   ix9175 : nor03_2x port map ( Y=>nx9174, A0=>nx8713, A1=>nx9415, A2=>
      nx11097);
   gen_23_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_23_cmp_mReg_12, QB=>
      nx8713, D=>window_23_12, CLK=>start, R=>rst);
   ix9173 : nor03_2x port map ( Y=>nx9172, A0=>gen_23_cmp_mReg_12, A1=>
      nx10139, A2=>nx11105);
   ix9209 : nand02 port map ( Y=>gen_23_cmp_BSCmp_op2_13, A0=>nx8717, A1=>
      nx8723);
   ix8718 : nor02_2x port map ( Y=>nx8717, A0=>nx9204, A1=>nx9200);
   ix9205 : nor03_2x port map ( Y=>nx9204, A0=>gen_23_cmp_mReg_12, A1=>
      nx9421, A2=>nx11075);
   ix9201 : nor03_2x port map ( Y=>nx9200, A0=>nx8713, A1=>nx11079, A2=>
      nx11091);
   ix8724 : nor02_2x port map ( Y=>nx8723, A0=>nx9196, A1=>nx9194);
   ix9197 : nor03_2x port map ( Y=>nx9196, A0=>nx8727, A1=>nx9415, A2=>
      nx11099);
   gen_23_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_23_cmp_mReg_13, QB=>
      nx8727, D=>window_23_13, CLK=>start, R=>rst);
   ix9195 : nor03_2x port map ( Y=>nx9194, A0=>gen_23_cmp_mReg_13, A1=>
      nx10139, A2=>nx11107);
   ix9231 : nand02 port map ( Y=>gen_23_cmp_BSCmp_op2_14, A0=>nx8731, A1=>
      nx8737);
   ix8732 : nor02_2x port map ( Y=>nx8731, A0=>nx9226, A1=>nx9222);
   ix9227 : nor03_2x port map ( Y=>nx9226, A0=>gen_23_cmp_mReg_13, A1=>
      nx9421, A2=>nx11075);
   ix9223 : nor03_2x port map ( Y=>nx9222, A0=>nx8727, A1=>nx11081, A2=>
      nx11091);
   ix8738 : nor02_2x port map ( Y=>nx8737, A0=>nx9218, A1=>nx9216);
   ix9219 : nor03_2x port map ( Y=>nx9218, A0=>nx8740, A1=>nx9415, A2=>
      nx11099);
   gen_23_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_23_cmp_mReg_14, QB=>
      nx8740, D=>window_23_14, CLK=>start, R=>rst);
   ix9217 : nor03_2x port map ( Y=>nx9216, A0=>gen_23_cmp_mReg_14, A1=>
      nx10139, A2=>nx11107);
   ix9253 : nand02 port map ( Y=>gen_23_cmp_BSCmp_op2_15, A0=>nx8747, A1=>
      nx8753);
   ix8748 : nor02_2x port map ( Y=>nx8747, A0=>nx9248, A1=>nx9244);
   ix9249 : nor03_2x port map ( Y=>nx9248, A0=>gen_23_cmp_mReg_14, A1=>
      nx9421, A2=>nx11075);
   ix9245 : nor03_2x port map ( Y=>nx9244, A0=>nx8740, A1=>nx11081, A2=>
      nx11091);
   ix8754 : nor02_2x port map ( Y=>nx8753, A0=>nx9240, A1=>nx9238);
   ix9241 : nor03_2x port map ( Y=>nx9240, A0=>nx8757, A1=>nx9415, A2=>
      nx11099);
   gen_23_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_23_cmp_mReg_15, QB=>
      nx8757, D=>window_23_15, CLK=>start, R=>rst);
   ix9239 : nor03_2x port map ( Y=>nx9238, A0=>gen_23_cmp_mReg_15, A1=>
      nx10141, A2=>nx11107);
   ix9263 : nand02 port map ( Y=>gen_23_cmp_BSCmp_op2_16, A0=>nx8761, A1=>
      nx8753);
   ix8762 : nor02_2x port map ( Y=>nx8761, A0=>nx9258, A1=>nx9254);
   ix9259 : nor03_2x port map ( Y=>nx9258, A0=>gen_23_cmp_mReg_15, A1=>
      nx9421, A2=>nx11075);
   ix9255 : nor03_2x port map ( Y=>nx9254, A0=>nx8757, A1=>nx11081, A2=>
      nx11091);
   ix9331 : nand02 port map ( Y=>gen_24_cmp_BSCmp_op2_1, A0=>nx8769, A1=>
      nx8789);
   ix8770 : nor02_2x port map ( Y=>nx8769, A0=>nx9326, A1=>nx9322);
   ix9327 : nor03_2x port map ( Y=>nx9326, A0=>gen_24_cmp_mReg_0, A1=>nx9405, 
      A2=>nx11111);
   gen_24_cmp_mRegCmp_reg_Q_0 : dffr port map ( Q=>gen_24_cmp_mReg_0, QB=>
      nx8775, D=>window_24_0, CLK=>start, R=>rst);
   ix8780 : inv01 port map ( Y=>nx8779, A=>gen_24_cmp_pMux_0);
   ix9323 : nor03_2x port map ( Y=>nx9322, A0=>nx8775, A1=>nx11117, A2=>
      nx11127);
   ix8788 : inv02 port map ( Y=>nx8787, A=>gen_24_cmp_pMux_2);
   ix8790 : nor02_2x port map ( Y=>nx8789, A0=>nx9312, A1=>nx9310);
   ix9313 : nor03_2x port map ( Y=>nx9312, A0=>nx8793, A1=>nx9399, A2=>
      nx11135);
   gen_24_cmp_mRegCmp_reg_Q_1 : dffr port map ( Q=>gen_24_cmp_mReg_1, QB=>
      nx8793, D=>window_24_1, CLK=>start, R=>rst);
   ix9311 : nor03_2x port map ( Y=>nx9310, A0=>gen_24_cmp_mReg_1, A1=>
      nx10143, A2=>nx11143);
   ix9271 : nor03_2x port map ( Y=>nx9270, A0=>nx9405, A1=>nx8787, A2=>
      gen_24_cmp_pMux_0);
   ix9353 : nand02 port map ( Y=>gen_24_cmp_BSCmp_op2_2, A0=>nx8804, A1=>
      nx8809);
   ix8805 : nor02_2x port map ( Y=>nx8804, A0=>nx9348, A1=>nx9344);
   ix9349 : nor03_2x port map ( Y=>nx9348, A0=>gen_24_cmp_mReg_1, A1=>nx9405, 
      A2=>nx11111);
   ix9345 : nor03_2x port map ( Y=>nx9344, A0=>nx8793, A1=>nx11117, A2=>
      nx11127);
   ix8810 : nor02_2x port map ( Y=>nx8809, A0=>nx9340, A1=>nx9338);
   ix9341 : nor03_2x port map ( Y=>nx9340, A0=>nx8813, A1=>nx9399, A2=>
      nx11135);
   gen_24_cmp_mRegCmp_reg_Q_2 : dffr port map ( Q=>gen_24_cmp_mReg_2, QB=>
      nx8813, D=>window_24_2, CLK=>start, R=>rst);
   ix9339 : nor03_2x port map ( Y=>nx9338, A0=>gen_24_cmp_mReg_2, A1=>
      nx10143, A2=>nx11143);
   ix9375 : nand02 port map ( Y=>gen_24_cmp_BSCmp_op2_3, A0=>nx8819, A1=>
      nx8825);
   ix8820 : nor02_2x port map ( Y=>nx8819, A0=>nx9370, A1=>nx9366);
   ix9371 : nor03_2x port map ( Y=>nx9370, A0=>gen_24_cmp_mReg_2, A1=>nx9405, 
      A2=>nx11111);
   ix9367 : nor03_2x port map ( Y=>nx9366, A0=>nx8813, A1=>nx11117, A2=>
      nx11127);
   ix8826 : nor02_2x port map ( Y=>nx8825, A0=>nx9362, A1=>nx9360);
   ix9363 : nor03_2x port map ( Y=>nx9362, A0=>nx8828, A1=>nx9399, A2=>
      nx11135);
   gen_24_cmp_mRegCmp_reg_Q_3 : dffr port map ( Q=>gen_24_cmp_mReg_3, QB=>
      nx8828, D=>window_24_3, CLK=>start, R=>rst);
   ix9361 : nor03_2x port map ( Y=>nx9360, A0=>gen_24_cmp_mReg_3, A1=>
      nx10143, A2=>nx11143);
   ix9397 : nand02 port map ( Y=>gen_24_cmp_BSCmp_op2_4, A0=>nx8835, A1=>
      nx8841);
   ix8836 : nor02_2x port map ( Y=>nx8835, A0=>nx9392, A1=>nx9388);
   ix9393 : nor03_2x port map ( Y=>nx9392, A0=>gen_24_cmp_mReg_3, A1=>nx9405, 
      A2=>nx11111);
   ix9389 : nor03_2x port map ( Y=>nx9388, A0=>nx8828, A1=>nx11117, A2=>
      nx11127);
   ix8842 : nor02_2x port map ( Y=>nx8841, A0=>nx9384, A1=>nx9382);
   ix9385 : nor03_2x port map ( Y=>nx9384, A0=>nx8845, A1=>nx9399, A2=>
      nx11135);
   gen_24_cmp_mRegCmp_reg_Q_4 : dffr port map ( Q=>gen_24_cmp_mReg_4, QB=>
      nx8845, D=>window_24_4, CLK=>start, R=>rst);
   ix9383 : nor03_2x port map ( Y=>nx9382, A0=>gen_24_cmp_mReg_4, A1=>
      nx10143, A2=>nx11143);
   ix9419 : nand02 port map ( Y=>gen_24_cmp_BSCmp_op2_5, A0=>nx8849, A1=>
      nx8855);
   ix8850 : nor02_2x port map ( Y=>nx8849, A0=>nx9414, A1=>nx9410);
   ix9415 : nor03_2x port map ( Y=>nx9414, A0=>gen_24_cmp_mReg_4, A1=>nx9405, 
      A2=>nx11111);
   ix9411 : nor03_2x port map ( Y=>nx9410, A0=>nx8845, A1=>nx11117, A2=>
      nx11127);
   ix8856 : nor02_2x port map ( Y=>nx8855, A0=>nx9406, A1=>nx9404);
   ix9407 : nor03_2x port map ( Y=>nx9406, A0=>nx8859, A1=>nx9401, A2=>
      nx11135);
   gen_24_cmp_mRegCmp_reg_Q_5 : dffr port map ( Q=>gen_24_cmp_mReg_5, QB=>
      nx8859, D=>window_24_5, CLK=>start, R=>rst);
   ix9405 : nor03_2x port map ( Y=>nx9404, A0=>gen_24_cmp_mReg_5, A1=>
      nx10143, A2=>nx11143);
   ix9441 : nand02 port map ( Y=>gen_24_cmp_BSCmp_op2_6, A0=>nx8863, A1=>
      nx8869);
   ix8864 : nor02_2x port map ( Y=>nx8863, A0=>nx9436, A1=>nx9432);
   ix9437 : nor03_2x port map ( Y=>nx9436, A0=>gen_24_cmp_mReg_5, A1=>nx9407, 
      A2=>nx11111);
   ix9433 : nor03_2x port map ( Y=>nx9432, A0=>nx8859, A1=>nx11117, A2=>
      nx11127);
   ix8870 : nor02_2x port map ( Y=>nx8869, A0=>nx9428, A1=>nx9426);
   ix9429 : nor03_2x port map ( Y=>nx9428, A0=>nx8873, A1=>nx9401, A2=>
      nx11135);
   gen_24_cmp_mRegCmp_reg_Q_6 : dffr port map ( Q=>gen_24_cmp_mReg_6, QB=>
      nx8873, D=>window_24_6, CLK=>start, R=>rst);
   ix9427 : nor03_2x port map ( Y=>nx9426, A0=>gen_24_cmp_mReg_6, A1=>
      nx10143, A2=>nx11143);
   ix9463 : nand02 port map ( Y=>gen_24_cmp_BSCmp_op2_7, A0=>nx8879, A1=>
      nx8885);
   ix8880 : nor02_2x port map ( Y=>nx8879, A0=>nx9458, A1=>nx9454);
   ix9459 : nor03_2x port map ( Y=>nx9458, A0=>gen_24_cmp_mReg_6, A1=>nx9407, 
      A2=>nx11113);
   ix9455 : nor03_2x port map ( Y=>nx9454, A0=>nx8873, A1=>nx11119, A2=>
      nx11129);
   ix8886 : nor02_2x port map ( Y=>nx8885, A0=>nx9450, A1=>nx9448);
   ix9451 : nor03_2x port map ( Y=>nx9450, A0=>nx8888, A1=>nx9401, A2=>
      nx11137);
   gen_24_cmp_mRegCmp_reg_Q_7 : dffr port map ( Q=>gen_24_cmp_mReg_7, QB=>
      nx8888, D=>window_24_7, CLK=>start, R=>rst);
   ix9449 : nor03_2x port map ( Y=>nx9448, A0=>gen_24_cmp_mReg_7, A1=>
      nx10143, A2=>nx11145);
   ix9485 : nand02 port map ( Y=>gen_24_cmp_BSCmp_op2_8, A0=>nx8892, A1=>
      nx8897);
   ix8893 : nor02_2x port map ( Y=>nx8892, A0=>nx9480, A1=>nx9476);
   ix9481 : nor03_2x port map ( Y=>nx9480, A0=>gen_24_cmp_mReg_7, A1=>nx9407, 
      A2=>nx11113);
   ix9477 : nor03_2x port map ( Y=>nx9476, A0=>nx8888, A1=>nx11119, A2=>
      nx11129);
   ix8898 : nor02_2x port map ( Y=>nx8897, A0=>nx9472, A1=>nx9470);
   ix9473 : nor03_2x port map ( Y=>nx9472, A0=>nx8901, A1=>nx9401, A2=>
      nx11137);
   gen_24_cmp_mRegCmp_reg_Q_8 : dffr port map ( Q=>gen_24_cmp_mReg_8, QB=>
      nx8901, D=>window_24_8, CLK=>start, R=>rst);
   ix9471 : nor03_2x port map ( Y=>nx9470, A0=>gen_24_cmp_mReg_8, A1=>
      nx10145, A2=>nx11145);
   ix9507 : nand02 port map ( Y=>gen_24_cmp_BSCmp_op2_9, A0=>nx8907, A1=>
      nx8913);
   ix8908 : nor02_2x port map ( Y=>nx8907, A0=>nx9502, A1=>nx9498);
   ix9503 : nor03_2x port map ( Y=>nx9502, A0=>gen_24_cmp_mReg_8, A1=>nx9407, 
      A2=>nx11113);
   ix9499 : nor03_2x port map ( Y=>nx9498, A0=>nx8901, A1=>nx11119, A2=>
      nx11129);
   ix8914 : nor02_2x port map ( Y=>nx8913, A0=>nx9494, A1=>nx9492);
   ix9495 : nor03_2x port map ( Y=>nx9494, A0=>nx8917, A1=>nx9401, A2=>
      nx11137);
   gen_24_cmp_mRegCmp_reg_Q_9 : dffr port map ( Q=>gen_24_cmp_mReg_9, QB=>
      nx8917, D=>window_24_9, CLK=>start, R=>rst);
   ix9493 : nor03_2x port map ( Y=>nx9492, A0=>gen_24_cmp_mReg_9, A1=>
      nx10145, A2=>nx11145);
   ix9529 : nand02 port map ( Y=>gen_24_cmp_BSCmp_op2_10, A0=>nx8921, A1=>
      nx8927);
   ix8922 : nor02_2x port map ( Y=>nx8921, A0=>nx9524, A1=>nx9520);
   ix9525 : nor03_2x port map ( Y=>nx9524, A0=>gen_24_cmp_mReg_9, A1=>nx9407, 
      A2=>nx11113);
   ix9521 : nor03_2x port map ( Y=>nx9520, A0=>nx8917, A1=>nx11119, A2=>
      nx11129);
   ix8928 : nor02_2x port map ( Y=>nx8927, A0=>nx9516, A1=>nx9514);
   ix9517 : nor03_2x port map ( Y=>nx9516, A0=>nx8931, A1=>nx9401, A2=>
      nx11137);
   gen_24_cmp_mRegCmp_reg_Q_10 : dffr port map ( Q=>gen_24_cmp_mReg_10, QB=>
      nx8931, D=>window_24_10, CLK=>start, R=>rst);
   ix9515 : nor03_2x port map ( Y=>nx9514, A0=>gen_24_cmp_mReg_10, A1=>
      nx10145, A2=>nx11145);
   ix9551 : nand02 port map ( Y=>gen_24_cmp_BSCmp_op2_11, A0=>nx8937, A1=>
      nx8941);
   ix8938 : nor02_2x port map ( Y=>nx8937, A0=>nx9546, A1=>nx9542);
   ix9547 : nor03_2x port map ( Y=>nx9546, A0=>gen_24_cmp_mReg_10, A1=>
      nx9407, A2=>nx11113);
   ix9543 : nor03_2x port map ( Y=>nx9542, A0=>nx8931, A1=>nx11119, A2=>
      nx11129);
   ix8942 : nor02_2x port map ( Y=>nx8941, A0=>nx9538, A1=>nx9536);
   ix9539 : nor03_2x port map ( Y=>nx9538, A0=>nx8945, A1=>nx9401, A2=>
      nx11137);
   gen_24_cmp_mRegCmp_reg_Q_11 : dffr port map ( Q=>gen_24_cmp_mReg_11, QB=>
      nx8945, D=>window_24_11, CLK=>start, R=>rst);
   ix9537 : nor03_2x port map ( Y=>nx9536, A0=>gen_24_cmp_mReg_11, A1=>
      nx10145, A2=>nx11145);
   ix9573 : nand02 port map ( Y=>gen_24_cmp_BSCmp_op2_12, A0=>nx8949, A1=>
      nx8955);
   ix8950 : nor02_2x port map ( Y=>nx8949, A0=>nx9568, A1=>nx9564);
   ix9569 : nor03_2x port map ( Y=>nx9568, A0=>gen_24_cmp_mReg_11, A1=>
      nx9407, A2=>nx11113);
   ix9565 : nor03_2x port map ( Y=>nx9564, A0=>nx8945, A1=>nx11119, A2=>
      nx11129);
   ix8956 : nor02_2x port map ( Y=>nx8955, A0=>nx9560, A1=>nx9558);
   ix9561 : nor03_2x port map ( Y=>nx9560, A0=>nx8959, A1=>nx9403, A2=>
      nx11137);
   gen_24_cmp_mRegCmp_reg_Q_12 : dffr port map ( Q=>gen_24_cmp_mReg_12, QB=>
      nx8959, D=>window_24_12, CLK=>start, R=>rst);
   ix9559 : nor03_2x port map ( Y=>nx9558, A0=>gen_24_cmp_mReg_12, A1=>
      nx10145, A2=>nx11145);
   ix9595 : nand02 port map ( Y=>gen_24_cmp_BSCmp_op2_13, A0=>nx8963, A1=>
      nx8969);
   ix8964 : nor02_2x port map ( Y=>nx8963, A0=>nx9590, A1=>nx9586);
   ix9591 : nor03_2x port map ( Y=>nx9590, A0=>gen_24_cmp_mReg_12, A1=>
      nx9409, A2=>nx11115);
   ix9587 : nor03_2x port map ( Y=>nx9586, A0=>nx8959, A1=>nx11119, A2=>
      nx11131);
   ix8970 : nor02_2x port map ( Y=>nx8969, A0=>nx9582, A1=>nx9580);
   ix9583 : nor03_2x port map ( Y=>nx9582, A0=>nx8972, A1=>nx9403, A2=>
      nx11139);
   gen_24_cmp_mRegCmp_reg_Q_13 : dffr port map ( Q=>gen_24_cmp_mReg_13, QB=>
      nx8972, D=>window_24_13, CLK=>start, R=>rst);
   ix9581 : nor03_2x port map ( Y=>nx9580, A0=>gen_24_cmp_mReg_13, A1=>
      nx10145, A2=>nx11147);
   ix9617 : nand02 port map ( Y=>gen_24_cmp_BSCmp_op2_14, A0=>nx8979, A1=>
      nx8985);
   ix8980 : nor02_2x port map ( Y=>nx8979, A0=>nx9612, A1=>nx9608);
   ix9613 : nor03_2x port map ( Y=>nx9612, A0=>gen_24_cmp_mReg_13, A1=>
      nx9409, A2=>nx11115);
   ix9609 : nor03_2x port map ( Y=>nx9608, A0=>nx8972, A1=>nx11121, A2=>
      nx11131);
   ix8986 : nor02_2x port map ( Y=>nx8985, A0=>nx9604, A1=>nx9602);
   ix9605 : nor03_2x port map ( Y=>nx9604, A0=>nx8989, A1=>nx9403, A2=>
      nx11139);
   gen_24_cmp_mRegCmp_reg_Q_14 : dffr port map ( Q=>gen_24_cmp_mReg_14, QB=>
      nx8989, D=>window_24_14, CLK=>start, R=>rst);
   ix9603 : nor03_2x port map ( Y=>nx9602, A0=>gen_24_cmp_mReg_14, A1=>
      nx10145, A2=>nx11147);
   ix9639 : nand02 port map ( Y=>gen_24_cmp_BSCmp_op2_15, A0=>nx8993, A1=>
      nx8999);
   ix8994 : nor02_2x port map ( Y=>nx8993, A0=>nx9634, A1=>nx9630);
   ix9635 : nor03_2x port map ( Y=>nx9634, A0=>gen_24_cmp_mReg_14, A1=>
      nx9409, A2=>nx11115);
   ix9631 : nor03_2x port map ( Y=>nx9630, A0=>nx8989, A1=>nx11121, A2=>
      nx11131);
   ix9000 : nor02_2x port map ( Y=>nx8999, A0=>nx9626, A1=>nx9624);
   ix9627 : nor03_2x port map ( Y=>nx9626, A0=>nx9003, A1=>nx9403, A2=>
      nx11139);
   gen_24_cmp_mRegCmp_reg_Q_15 : dffr port map ( Q=>gen_24_cmp_mReg_15, QB=>
      nx9003, D=>window_24_15, CLK=>start, R=>rst);
   ix9625 : nor03_2x port map ( Y=>nx9624, A0=>gen_24_cmp_mReg_15, A1=>
      nx10147, A2=>nx11147);
   ix9649 : nand02 port map ( Y=>gen_24_cmp_BSCmp_op2_16, A0=>nx9007, A1=>
      nx8999);
   ix9008 : nor02_2x port map ( Y=>nx9007, A0=>nx9644, A1=>nx9640);
   ix9645 : nor03_2x port map ( Y=>nx9644, A0=>gen_24_cmp_mReg_15, A1=>
      nx9409, A2=>nx11115);
   ix9641 : nor03_2x port map ( Y=>nx9640, A0=>nx9003, A1=>nx11121, A2=>
      nx11131);
   ix19 : nor02_2x port map ( Y=>gen_0_cmp_BSCmp_carryIn, A0=>nx2871, A1=>
      nx9014);
   ix9015 : nor02_2x port map ( Y=>nx9014, A0=>nx10161, A1=>nx2862);
   ix39 : nand02 port map ( Y=>gen_0_cmp_BSCmp_op2_0, A0=>nx9017, A1=>nx9023
   );
   ix9018 : nor02_2x port map ( Y=>nx9017, A0=>nx34, A1=>nx26);
   ix35 : nor03_2x port map ( Y=>nx34, A0=>nx2859, A1=>nx9691, A2=>nx10179);
   ix27 : nor03_2x port map ( Y=>nx26, A0=>gen_0_cmp_mReg_0, A1=>nx10003, A2
      =>nx10187);
   ix9024 : nand03 port map ( Y=>nx9023, A0=>nx10161, A1=>nx9691, A2=>nx2862
   );
   ix405 : nor02_2x port map ( Y=>gen_1_cmp_BSCmp_carryIn, A0=>nx3115, A1=>
      nx9027);
   ix9028 : nor02_2x port map ( Y=>nx9027, A0=>nx10201, A1=>nx3107);
   ix425 : nand02 port map ( Y=>gen_1_cmp_BSCmp_op2_0, A0=>nx9031, A1=>
      nx9036);
   ix9032 : nor02_2x port map ( Y=>nx9031, A0=>nx420, A1=>nx412);
   ix421 : nor03_2x port map ( Y=>nx420, A0=>nx3103, A1=>nx9679, A2=>nx10219
   );
   ix413 : nor03_2x port map ( Y=>nx412, A0=>gen_1_cmp_mReg_0, A1=>nx10009, 
      A2=>nx10227);
   ix9037 : nand03 port map ( Y=>nx9036, A0=>nx10201, A1=>nx9679, A2=>nx3107
   );
   ix791 : nor02_2x port map ( Y=>gen_2_cmp_BSCmp_carryIn, A0=>nx3363, A1=>
      nx9039);
   ix9040 : nor02_2x port map ( Y=>nx9039, A0=>nx10241, A1=>nx3356);
   ix811 : nand02 port map ( Y=>gen_2_cmp_BSCmp_op2_0, A0=>nx9043, A1=>
      nx9049);
   ix9044 : nor02_2x port map ( Y=>nx9043, A0=>nx806, A1=>nx798);
   ix807 : nor03_2x port map ( Y=>nx806, A0=>nx3353, A1=>nx9667, A2=>nx10259
   );
   ix799 : nor03_2x port map ( Y=>nx798, A0=>gen_2_cmp_mReg_0, A1=>nx10015, 
      A2=>nx10267);
   ix9050 : nand03 port map ( Y=>nx9049, A0=>nx10241, A1=>nx9667, A2=>nx3356
   );
   ix1177 : nor02_2x port map ( Y=>gen_3_cmp_BSCmp_carryIn, A0=>nx3611, A1=>
      nx9053);
   ix9054 : nor02_2x port map ( Y=>nx9053, A0=>nx10281, A1=>nx3603);
   ix1197 : nand02 port map ( Y=>gen_3_cmp_BSCmp_op2_0, A0=>nx9057, A1=>
      nx9061);
   ix9058 : nor02_2x port map ( Y=>nx9057, A0=>nx1192, A1=>nx1184);
   ix1193 : nor03_2x port map ( Y=>nx1192, A0=>nx3599, A1=>nx9655, A2=>
      nx10299);
   ix1185 : nor03_2x port map ( Y=>nx1184, A0=>gen_3_cmp_mReg_0, A1=>nx10021, 
      A2=>nx10307);
   ix9062 : nand03 port map ( Y=>nx9061, A0=>nx10281, A1=>nx9655, A2=>nx3603
   );
   ix1563 : nor02_2x port map ( Y=>gen_4_cmp_BSCmp_carryIn, A0=>nx3857, A1=>
      nx9065);
   ix9066 : nor02_2x port map ( Y=>nx9065, A0=>nx10321, A1=>nx3849);
   ix1583 : nand02 port map ( Y=>gen_4_cmp_BSCmp_op2_0, A0=>nx9069, A1=>
      nx9073);
   ix9070 : nor02_2x port map ( Y=>nx9069, A0=>nx1578, A1=>nx1570);
   ix1579 : nor03_2x port map ( Y=>nx1578, A0=>nx3845, A1=>nx9643, A2=>
      nx10339);
   ix1571 : nor03_2x port map ( Y=>nx1570, A0=>gen_4_cmp_mReg_0, A1=>nx10027, 
      A2=>nx10347);
   ix9074 : nand03 port map ( Y=>nx9073, A0=>nx10321, A1=>nx9643, A2=>nx3849
   );
   ix1949 : nor02_2x port map ( Y=>gen_5_cmp_BSCmp_carryIn, A0=>nx4101, A1=>
      nx9077);
   ix9078 : nor02_2x port map ( Y=>nx9077, A0=>nx10361, A1=>nx4093);
   ix1969 : nand02 port map ( Y=>gen_5_cmp_BSCmp_op2_0, A0=>nx9080, A1=>
      nx9085);
   ix9081 : nor02_2x port map ( Y=>nx9080, A0=>nx1964, A1=>nx1956);
   ix1965 : nor03_2x port map ( Y=>nx1964, A0=>nx4089, A1=>nx9631, A2=>
      nx10379);
   ix1957 : nor03_2x port map ( Y=>nx1956, A0=>gen_5_cmp_mReg_0, A1=>nx10033, 
      A2=>nx10387);
   ix9086 : nand03 port map ( Y=>nx9085, A0=>nx10361, A1=>nx9631, A2=>nx4093
   );
   ix2335 : nor02_2x port map ( Y=>gen_6_cmp_BSCmp_carryIn, A0=>nx4349, A1=>
      nx9089);
   ix9090 : nor02_2x port map ( Y=>nx9089, A0=>nx10401, A1=>nx4340);
   ix2355 : nand02 port map ( Y=>gen_6_cmp_BSCmp_op2_0, A0=>nx9093, A1=>
      nx9099);
   ix9094 : nor02_2x port map ( Y=>nx9093, A0=>nx2350, A1=>nx2342);
   ix2351 : nor03_2x port map ( Y=>nx2350, A0=>nx4337, A1=>nx9619, A2=>
      nx10419);
   ix2343 : nor03_2x port map ( Y=>nx2342, A0=>gen_6_cmp_mReg_0, A1=>nx10039, 
      A2=>nx10427);
   ix9100 : nand03 port map ( Y=>nx9099, A0=>nx10401, A1=>nx9619, A2=>nx4340
   );
   ix2721 : nor02_2x port map ( Y=>gen_7_cmp_BSCmp_carryIn, A0=>nx4595, A1=>
      nx9102);
   ix9103 : nor02_2x port map ( Y=>nx9102, A0=>nx10441, A1=>nx4587);
   ix2741 : nand02 port map ( Y=>gen_7_cmp_BSCmp_op2_0, A0=>nx9105, A1=>
      nx9111);
   ix9106 : nor02_2x port map ( Y=>nx9105, A0=>nx2736, A1=>nx2728);
   ix2737 : nor03_2x port map ( Y=>nx2736, A0=>nx4583, A1=>nx9607, A2=>
      nx10459);
   ix2729 : nor03_2x port map ( Y=>nx2728, A0=>gen_7_cmp_mReg_0, A1=>nx10045, 
      A2=>nx10467);
   ix9112 : nand03 port map ( Y=>nx9111, A0=>nx10441, A1=>nx9607, A2=>nx4587
   );
   ix3107 : nor02_2x port map ( Y=>gen_8_cmp_BSCmp_carryIn, A0=>nx4841, A1=>
      nx9115);
   ix9116 : nor02_2x port map ( Y=>nx9115, A0=>nx10481, A1=>nx4834);
   ix3127 : nand02 port map ( Y=>gen_8_cmp_BSCmp_op2_0, A0=>nx9119, A1=>
      nx9124);
   ix9120 : nor02_2x port map ( Y=>nx9119, A0=>nx3122, A1=>nx3114);
   ix3123 : nor03_2x port map ( Y=>nx3122, A0=>nx4831, A1=>nx9595, A2=>
      nx10499);
   ix3115 : nor03_2x port map ( Y=>nx3114, A0=>gen_8_cmp_mReg_0, A1=>nx10051, 
      A2=>nx10507);
   ix9125 : nand03 port map ( Y=>nx9124, A0=>nx10481, A1=>nx9595, A2=>nx4834
   );
   ix3493 : nor02_2x port map ( Y=>gen_9_cmp_BSCmp_carryIn, A0=>nx5085, A1=>
      nx9127);
   ix9128 : nor02_2x port map ( Y=>nx9127, A0=>nx10521, A1=>nx5077);
   ix3513 : nand02 port map ( Y=>gen_9_cmp_BSCmp_op2_0, A0=>nx9131, A1=>
      nx9137);
   ix9132 : nor02_2x port map ( Y=>nx9131, A0=>nx3508, A1=>nx3500);
   ix3509 : nor03_2x port map ( Y=>nx3508, A0=>nx5073, A1=>nx9583, A2=>
      nx10539);
   ix3501 : nor03_2x port map ( Y=>nx3500, A0=>gen_9_cmp_mReg_0, A1=>nx10057, 
      A2=>nx10547);
   ix9138 : nand03 port map ( Y=>nx9137, A0=>nx10521, A1=>nx9583, A2=>nx5077
   );
   ix3879 : nor02_2x port map ( Y=>gen_10_cmp_BSCmp_carryIn, A0=>nx5335, A1
      =>nx9141);
   ix9142 : nor02_2x port map ( Y=>nx9141, A0=>nx10561, A1=>nx5327);
   ix3899 : nand02 port map ( Y=>gen_10_cmp_BSCmp_op2_0, A0=>nx9145, A1=>
      nx9149);
   ix9146 : nor02_2x port map ( Y=>nx9145, A0=>nx3894, A1=>nx3886);
   ix3895 : nor03_2x port map ( Y=>nx3894, A0=>nx5323, A1=>nx9571, A2=>
      nx10579);
   ix3887 : nor03_2x port map ( Y=>nx3886, A0=>gen_10_cmp_mReg_0, A1=>
      nx10063, A2=>nx10587);
   ix9150 : nand03 port map ( Y=>nx9149, A0=>nx10561, A1=>nx9571, A2=>nx5327
   );
   ix4265 : nor02_2x port map ( Y=>gen_11_cmp_BSCmp_carryIn, A0=>nx5585, A1
      =>nx9153);
   ix9154 : nor02_2x port map ( Y=>nx9153, A0=>nx10601, A1=>nx5577);
   ix4285 : nand02 port map ( Y=>gen_11_cmp_BSCmp_op2_0, A0=>nx9157, A1=>
      nx9161);
   ix9158 : nor02_2x port map ( Y=>nx9157, A0=>nx4280, A1=>nx4272);
   ix4281 : nor03_2x port map ( Y=>nx4280, A0=>nx5573, A1=>nx9559, A2=>
      nx10619);
   ix4273 : nor03_2x port map ( Y=>nx4272, A0=>gen_11_cmp_mReg_0, A1=>
      nx10069, A2=>nx10627);
   ix9162 : nand03 port map ( Y=>nx9161, A0=>nx10601, A1=>nx9559, A2=>nx5577
   );
   ix4651 : nor02_2x port map ( Y=>gen_12_cmp_BSCmp_carryIn, A0=>nx5829, A1
      =>nx9165);
   ix9166 : nor02_2x port map ( Y=>nx9165, A0=>nx10641, A1=>nx5821);
   ix4671 : nand02 port map ( Y=>gen_12_cmp_BSCmp_op2_0, A0=>nx9168, A1=>
      nx9173);
   ix9169 : nor02_2x port map ( Y=>nx9168, A0=>nx4666, A1=>nx4658);
   ix4667 : nor03_2x port map ( Y=>nx4666, A0=>nx5817, A1=>nx9547, A2=>
      nx10659);
   ix4659 : nor03_2x port map ( Y=>nx4658, A0=>gen_12_cmp_mReg_0, A1=>
      nx10075, A2=>nx10667);
   ix9174 : nand03 port map ( Y=>nx9173, A0=>nx10641, A1=>nx9547, A2=>nx5821
   );
   ix5037 : nor02_2x port map ( Y=>gen_13_cmp_BSCmp_carryIn, A0=>nx6075, A1
      =>nx9177);
   ix9178 : nor02_2x port map ( Y=>nx9177, A0=>nx10681, A1=>nx6067);
   ix5057 : nand02 port map ( Y=>gen_13_cmp_BSCmp_op2_0, A0=>nx9181, A1=>
      nx9187);
   ix9182 : nor02_2x port map ( Y=>nx9181, A0=>nx5052, A1=>nx5044);
   ix5053 : nor03_2x port map ( Y=>nx5052, A0=>nx6063, A1=>nx9535, A2=>
      nx10699);
   ix5045 : nor03_2x port map ( Y=>nx5044, A0=>gen_13_cmp_mReg_0, A1=>
      nx10081, A2=>nx10707);
   ix9188 : nand03 port map ( Y=>nx9187, A0=>nx10681, A1=>nx9535, A2=>nx6067
   );
   ix5423 : nor02_2x port map ( Y=>gen_14_cmp_BSCmp_carryIn, A0=>nx6323, A1
      =>nx9190);
   ix9191 : nor02_2x port map ( Y=>nx9190, A0=>nx10721, A1=>nx6314);
   ix5443 : nand02 port map ( Y=>gen_14_cmp_BSCmp_op2_0, A0=>nx9193, A1=>
      nx9199);
   ix9194 : nor02_2x port map ( Y=>nx9193, A0=>nx5438, A1=>nx5430);
   ix5439 : nor03_2x port map ( Y=>nx5438, A0=>nx6311, A1=>nx9523, A2=>
      nx10739);
   ix5431 : nor03_2x port map ( Y=>nx5430, A0=>gen_14_cmp_mReg_0, A1=>
      nx10087, A2=>nx10747);
   ix9200 : nand03 port map ( Y=>nx9199, A0=>nx10721, A1=>nx9523, A2=>nx6314
   );
   ix5809 : nor02_2x port map ( Y=>gen_15_cmp_BSCmp_carryIn, A0=>nx6569, A1
      =>nx9203);
   ix9204 : nor02_2x port map ( Y=>nx9203, A0=>nx10761, A1=>nx6561);
   ix5829 : nand02 port map ( Y=>gen_15_cmp_BSCmp_op2_0, A0=>nx9207, A1=>
      nx9212);
   ix9208 : nor02_2x port map ( Y=>nx9207, A0=>nx5824, A1=>nx5816);
   ix5825 : nor03_2x port map ( Y=>nx5824, A0=>nx6557, A1=>nx9511, A2=>
      nx10779);
   ix5817 : nor03_2x port map ( Y=>nx5816, A0=>gen_15_cmp_mReg_0, A1=>
      nx10093, A2=>nx10787);
   ix9213 : nand03 port map ( Y=>nx9212, A0=>nx10761, A1=>nx9511, A2=>nx6561
   );
   ix6195 : nor02_2x port map ( Y=>gen_16_cmp_BSCmp_carryIn, A0=>nx6815, A1
      =>nx9215);
   ix9216 : nor02_2x port map ( Y=>nx9215, A0=>nx10801, A1=>nx6808);
   ix6215 : nand02 port map ( Y=>gen_16_cmp_BSCmp_op2_0, A0=>nx9219, A1=>
      nx9225);
   ix9220 : nor02_2x port map ( Y=>nx9219, A0=>nx6210, A1=>nx6202);
   ix6211 : nor03_2x port map ( Y=>nx6210, A0=>nx6805, A1=>nx9499, A2=>
      nx10819);
   ix6203 : nor03_2x port map ( Y=>nx6202, A0=>gen_16_cmp_mReg_0, A1=>
      nx10099, A2=>nx10827);
   ix9226 : nand03 port map ( Y=>nx9225, A0=>nx10801, A1=>nx9499, A2=>nx6808
   );
   ix6581 : nor02_2x port map ( Y=>gen_17_cmp_BSCmp_carryIn, A0=>nx7057, A1
      =>nx9229);
   ix9230 : nor02_2x port map ( Y=>nx9229, A0=>nx10841, A1=>nx7049);
   ix6601 : nand02 port map ( Y=>gen_17_cmp_BSCmp_op2_0, A0=>nx9233, A1=>
      nx9237);
   ix9234 : nor02_2x port map ( Y=>nx9233, A0=>nx6596, A1=>nx6588);
   ix6597 : nor03_2x port map ( Y=>nx6596, A0=>nx7045, A1=>nx9487, A2=>
      nx10859);
   ix6589 : nor03_2x port map ( Y=>nx6588, A0=>gen_17_cmp_mReg_0, A1=>
      nx10105, A2=>nx10867);
   ix9238 : nand03 port map ( Y=>nx9237, A0=>nx10841, A1=>nx9487, A2=>nx7049
   );
   ix6967 : nor02_2x port map ( Y=>gen_18_cmp_BSCmp_carryIn, A0=>nx7305, A1
      =>nx9241);
   ix9242 : nor02_2x port map ( Y=>nx9241, A0=>nx10881, A1=>nx7297);
   ix6987 : nand02 port map ( Y=>gen_18_cmp_BSCmp_op2_0, A0=>nx9245, A1=>
      nx9249);
   ix9246 : nor02_2x port map ( Y=>nx9245, A0=>nx6982, A1=>nx6974);
   ix6983 : nor03_2x port map ( Y=>nx6982, A0=>nx7293, A1=>nx9475, A2=>
      nx10899);
   ix6975 : nor03_2x port map ( Y=>nx6974, A0=>gen_18_cmp_mReg_0, A1=>
      nx10111, A2=>nx10907);
   ix9250 : nand03 port map ( Y=>nx9249, A0=>nx10881, A1=>nx9475, A2=>nx7297
   );
   ix7353 : nor02_2x port map ( Y=>gen_19_cmp_BSCmp_carryIn, A0=>nx7553, A1
      =>nx9253);
   ix9254 : nor02_2x port map ( Y=>nx9253, A0=>nx10921, A1=>nx7545);
   ix7373 : nand02 port map ( Y=>gen_19_cmp_BSCmp_op2_0, A0=>nx9257, A1=>
      nx9263);
   ix9258 : nor02_2x port map ( Y=>nx9257, A0=>nx7368, A1=>nx7360);
   ix7369 : nor03_2x port map ( Y=>nx7368, A0=>nx7541, A1=>nx9463, A2=>
      nx10939);
   ix7361 : nor03_2x port map ( Y=>nx7360, A0=>gen_19_cmp_mReg_0, A1=>
      nx10117, A2=>nx10947);
   ix9264 : nand03 port map ( Y=>nx9263, A0=>nx10921, A1=>nx9463, A2=>nx7545
   );
   ix7739 : nor02_2x port map ( Y=>gen_20_cmp_BSCmp_carryIn, A0=>nx7801, A1
      =>nx9267);
   ix9268 : nor02_2x port map ( Y=>nx9267, A0=>nx10961, A1=>nx7792);
   ix7759 : nand02 port map ( Y=>gen_20_cmp_BSCmp_op2_0, A0=>nx9271, A1=>
      nx9275);
   ix9272 : nor02_2x port map ( Y=>nx9271, A0=>nx7754, A1=>nx7746);
   ix7755 : nor03_2x port map ( Y=>nx7754, A0=>nx7789, A1=>nx9451, A2=>
      nx10979);
   ix7747 : nor03_2x port map ( Y=>nx7746, A0=>gen_20_cmp_mReg_0, A1=>
      nx10123, A2=>nx10987);
   ix9276 : nand03 port map ( Y=>nx9275, A0=>nx10961, A1=>nx9451, A2=>nx7792
   );
   ix8125 : nor02_2x port map ( Y=>gen_21_cmp_BSCmp_carryIn, A0=>nx8047, A1
      =>nx9278);
   ix9279 : nor02_2x port map ( Y=>nx9278, A0=>nx11001, A1=>nx8039);
   ix8145 : nand02 port map ( Y=>gen_21_cmp_BSCmp_op2_0, A0=>nx9281, A1=>
      nx9287);
   ix9282 : nor02_2x port map ( Y=>nx9281, A0=>nx8140, A1=>nx8132);
   ix8141 : nor03_2x port map ( Y=>nx8140, A0=>nx8035, A1=>nx9439, A2=>
      nx11019);
   ix8133 : nor03_2x port map ( Y=>nx8132, A0=>gen_21_cmp_mReg_0, A1=>
      nx10129, A2=>nx11027);
   ix9288 : nand03 port map ( Y=>nx9287, A0=>nx11001, A1=>nx9439, A2=>nx8039
   );
   ix8511 : nor02_2x port map ( Y=>gen_22_cmp_BSCmp_carryIn, A0=>nx8291, A1
      =>nx9291);
   ix9292 : nor02_2x port map ( Y=>nx9291, A0=>nx11041, A1=>nx8283);
   ix8531 : nand02 port map ( Y=>gen_22_cmp_BSCmp_op2_0, A0=>nx9295, A1=>
      nx9301);
   ix9296 : nor02_2x port map ( Y=>nx9295, A0=>nx8526, A1=>nx8518);
   ix8527 : nor03_2x port map ( Y=>nx8526, A0=>nx8279, A1=>nx9427, A2=>
      nx11059);
   ix8519 : nor03_2x port map ( Y=>nx8518, A0=>gen_22_cmp_mReg_0, A1=>
      nx10135, A2=>nx11067);
   ix9302 : nand03 port map ( Y=>nx9301, A0=>nx11041, A1=>nx9427, A2=>nx8283
   );
   ix8897 : nor02_2x port map ( Y=>gen_23_cmp_BSCmp_carryIn, A0=>nx8541, A1
      =>nx9305);
   ix9306 : nor02_2x port map ( Y=>nx9305, A0=>nx11081, A1=>nx8533);
   ix8917 : nand02 port map ( Y=>gen_23_cmp_BSCmp_op2_0, A0=>nx9308, A1=>
      nx9315);
   ix9310 : nor02_2x port map ( Y=>nx9308, A0=>nx8912, A1=>nx8904);
   ix8913 : nor03_2x port map ( Y=>nx8912, A0=>nx8529, A1=>nx9415, A2=>
      nx11099);
   ix8905 : nor03_2x port map ( Y=>nx8904, A0=>gen_23_cmp_mReg_0, A1=>
      nx10141, A2=>nx11107);
   ix9316 : nand03 port map ( Y=>nx9315, A0=>nx11081, A1=>nx9415, A2=>nx8533
   );
   ix9283 : nor02_2x port map ( Y=>gen_24_cmp_BSCmp_carryIn, A0=>nx8787, A1
      =>nx9319);
   ix9320 : nor02_2x port map ( Y=>nx9319, A0=>nx11121, A1=>nx8779);
   ix9303 : nand02 port map ( Y=>gen_24_cmp_BSCmp_op2_0, A0=>nx9323, A1=>
      nx9327);
   ix9324 : nor02_2x port map ( Y=>nx9323, A0=>nx9298, A1=>nx9290);
   ix9299 : nor03_2x port map ( Y=>nx9298, A0=>nx8775, A1=>nx9403, A2=>
      nx11139);
   ix9291 : nor03_2x port map ( Y=>nx9290, A0=>gen_24_cmp_mReg_0, A1=>
      nx10147, A2=>nx11147);
   ix9328 : nand03 port map ( Y=>nx9327, A0=>nx11121, A1=>nx9403, A2=>nx8779
   );
   ix2840 : nor02_2x port map ( Y=>nx2839, A0=>nx11197, A1=>nx11171);
   CounterCmp_reg_outp_0 : dffs_ni port map ( Q=>OPEN, QB=>nx9333, D=>nx2839, 
      CLK=>clk, S=>nx9670);
   ix9671 : inv01 port map ( Y=>nx9670, A=>nx9336);
   ix9338 : nor02_2x port map ( Y=>nx9336, A0=>restartDetection, A1=>rst);
   StartCaptuerCmp_reg_f : dffr port map ( Q=>restartDetection, QB=>OPEN, D
      =>nx9650, CLK=>start, R=>nx9664);
   ix9665 : inv01 port map ( Y=>nx9664, A=>nx9343);
   ix9344 : nor02_2x port map ( Y=>nx9343, A0=>StartCaptuerCmp_d, A1=>rst);
   StartCaptuerCmp_reg_d : dff port map ( Q=>StartCaptuerCmp_d, QB=>OPEN, D
      =>restartDetection, CLK=>nx9397);
   firtStartLachCmp_reg_Q_0 : dffr port map ( Q=>OPEN, QB=>nx9353, D=>nx9650, 
      CLK=>start, R=>rst);
   ix2834 : oai21 port map ( Y=>nx2833, A0=>nx9357, A1=>nx9353, B0=>nx9365);
   CounterCmp_reg_outp_2 : dffr port map ( Q=>OPEN, QB=>nx9357, D=>nx2823, 
      CLK=>clk, R=>nx9670);
   CounterCmp_reg_outp_1 : dffr port map ( Q=>OPEN, QB=>nx9361, D=>nx2813, 
      CLK=>clk, R=>nx9670);
   CounterCmp_reg_outp_3 : dffr port map ( Q=>done, QB=>nx9365, D=>nx2833, 
      CLK=>clk, R=>nx9670);
   ix9374 : inv02 port map ( Y=>nx9375, A=>nx9373);
   ix9376 : inv02 port map ( Y=>nx9377, A=>nx11201);
   ix9378 : inv02 port map ( Y=>nx9379, A=>nx11201);
   ix9380 : inv02 port map ( Y=>nx9381, A=>nx11201);
   ix9388 : inv01 port map ( Y=>nx9389, A=>nx9333);
   ix9390 : inv01 port map ( Y=>nx9391, A=>clk);
   ix9392 : inv01 port map ( Y=>nx9393, A=>clk);
   ix9394 : inv01 port map ( Y=>nx9395, A=>clk);
   ix9396 : inv01 port map ( Y=>nx9397, A=>clk);
   ix9398 : inv04 port map ( Y=>nx9399, A=>nx8787);
   ix9400 : inv04 port map ( Y=>nx9401, A=>nx8787);
   ix9402 : inv04 port map ( Y=>nx9403, A=>nx8787);
   ix9404 : inv04 port map ( Y=>nx9405, A=>nx11121);
   ix9406 : inv04 port map ( Y=>nx9407, A=>nx11121);
   ix9408 : inv04 port map ( Y=>nx9409, A=>nx11123);
   ix9410 : inv04 port map ( Y=>nx9411, A=>nx8541);
   ix9412 : inv04 port map ( Y=>nx9413, A=>nx8541);
   ix9414 : inv04 port map ( Y=>nx9415, A=>nx8541);
   ix9416 : inv04 port map ( Y=>nx9417, A=>nx11081);
   ix9418 : inv04 port map ( Y=>nx9419, A=>nx11081);
   ix9420 : inv04 port map ( Y=>nx9421, A=>nx11083);
   ix9422 : inv04 port map ( Y=>nx9423, A=>nx8291);
   ix9424 : inv04 port map ( Y=>nx9425, A=>nx8291);
   ix9426 : inv04 port map ( Y=>nx9427, A=>nx8291);
   ix9428 : inv04 port map ( Y=>nx9429, A=>nx11041);
   ix9430 : inv04 port map ( Y=>nx9431, A=>nx11041);
   ix9432 : inv04 port map ( Y=>nx9433, A=>nx11043);
   ix9434 : inv04 port map ( Y=>nx9435, A=>nx8047);
   ix9436 : inv04 port map ( Y=>nx9437, A=>nx8047);
   ix9438 : inv04 port map ( Y=>nx9439, A=>nx8047);
   ix9440 : inv04 port map ( Y=>nx9441, A=>nx11001);
   ix9442 : inv04 port map ( Y=>nx9443, A=>nx11001);
   ix9444 : inv04 port map ( Y=>nx9445, A=>nx11003);
   ix9446 : inv04 port map ( Y=>nx9447, A=>nx7801);
   ix9448 : inv04 port map ( Y=>nx9449, A=>nx7801);
   ix9450 : inv04 port map ( Y=>nx9451, A=>nx7801);
   ix9452 : inv04 port map ( Y=>nx9453, A=>nx10961);
   ix9454 : inv04 port map ( Y=>nx9455, A=>nx10961);
   ix9456 : inv04 port map ( Y=>nx9457, A=>nx10963);
   ix9458 : inv04 port map ( Y=>nx9459, A=>nx7553);
   ix9460 : inv04 port map ( Y=>nx9461, A=>nx7553);
   ix9462 : inv04 port map ( Y=>nx9463, A=>nx7553);
   ix9464 : inv04 port map ( Y=>nx9465, A=>nx10921);
   ix9466 : inv04 port map ( Y=>nx9467, A=>nx10921);
   ix9468 : inv04 port map ( Y=>nx9469, A=>nx10923);
   ix9470 : inv04 port map ( Y=>nx9471, A=>nx7305);
   ix9472 : inv04 port map ( Y=>nx9473, A=>nx7305);
   ix9474 : inv04 port map ( Y=>nx9475, A=>nx7305);
   ix9476 : inv04 port map ( Y=>nx9477, A=>nx10881);
   ix9478 : inv04 port map ( Y=>nx9479, A=>nx10881);
   ix9480 : inv04 port map ( Y=>nx9481, A=>nx10883);
   ix9482 : inv04 port map ( Y=>nx9483, A=>nx7057);
   ix9484 : inv04 port map ( Y=>nx9485, A=>nx7057);
   ix9486 : inv04 port map ( Y=>nx9487, A=>nx7057);
   ix9488 : inv04 port map ( Y=>nx9489, A=>nx10841);
   ix9490 : inv04 port map ( Y=>nx9491, A=>nx10841);
   ix9492 : inv04 port map ( Y=>nx9493, A=>nx10843);
   ix9494 : inv04 port map ( Y=>nx9495, A=>nx6815);
   ix9496 : inv04 port map ( Y=>nx9497, A=>nx6815);
   ix9498 : inv04 port map ( Y=>nx9499, A=>nx6815);
   ix9500 : inv04 port map ( Y=>nx9501, A=>nx10801);
   ix9502 : inv04 port map ( Y=>nx9503, A=>nx10801);
   ix9504 : inv04 port map ( Y=>nx9505, A=>nx10803);
   ix9506 : inv04 port map ( Y=>nx9507, A=>nx6569);
   ix9508 : inv04 port map ( Y=>nx9509, A=>nx6569);
   ix9510 : inv04 port map ( Y=>nx9511, A=>nx6569);
   ix9512 : inv04 port map ( Y=>nx9513, A=>nx10761);
   ix9514 : inv04 port map ( Y=>nx9515, A=>nx10761);
   ix9516 : inv04 port map ( Y=>nx9517, A=>nx10763);
   ix9518 : inv04 port map ( Y=>nx9519, A=>nx6323);
   ix9520 : inv04 port map ( Y=>nx9521, A=>nx6323);
   ix9522 : inv04 port map ( Y=>nx9523, A=>nx6323);
   ix9524 : inv04 port map ( Y=>nx9525, A=>nx10721);
   ix9526 : inv04 port map ( Y=>nx9527, A=>nx10721);
   ix9528 : inv04 port map ( Y=>nx9529, A=>nx10723);
   ix9530 : inv04 port map ( Y=>nx9531, A=>nx6075);
   ix9532 : inv04 port map ( Y=>nx9533, A=>nx6075);
   ix9534 : inv04 port map ( Y=>nx9535, A=>nx6075);
   ix9536 : inv04 port map ( Y=>nx9537, A=>nx10681);
   ix9538 : inv04 port map ( Y=>nx9539, A=>nx10681);
   ix9540 : inv04 port map ( Y=>nx9541, A=>nx10683);
   ix9542 : inv04 port map ( Y=>nx9543, A=>nx5829);
   ix9544 : inv04 port map ( Y=>nx9545, A=>nx5829);
   ix9546 : inv04 port map ( Y=>nx9547, A=>nx5829);
   ix9548 : inv04 port map ( Y=>nx9549, A=>nx10641);
   ix9550 : inv04 port map ( Y=>nx9551, A=>nx10641);
   ix9552 : inv04 port map ( Y=>nx9553, A=>nx10643);
   ix9554 : inv04 port map ( Y=>nx9555, A=>nx5585);
   ix9556 : inv04 port map ( Y=>nx9557, A=>nx5585);
   ix9558 : inv04 port map ( Y=>nx9559, A=>nx5585);
   ix9560 : inv04 port map ( Y=>nx9561, A=>nx10601);
   ix9562 : inv04 port map ( Y=>nx9563, A=>nx10601);
   ix9564 : inv04 port map ( Y=>nx9565, A=>nx10603);
   ix9566 : inv04 port map ( Y=>nx9567, A=>nx5335);
   ix9568 : inv04 port map ( Y=>nx9569, A=>nx5335);
   ix9570 : inv04 port map ( Y=>nx9571, A=>nx5335);
   ix9572 : inv04 port map ( Y=>nx9573, A=>nx10561);
   ix9574 : inv04 port map ( Y=>nx9575, A=>nx10561);
   ix9576 : inv04 port map ( Y=>nx9577, A=>nx10563);
   ix9578 : inv04 port map ( Y=>nx9579, A=>nx5085);
   ix9580 : inv04 port map ( Y=>nx9581, A=>nx5085);
   ix9582 : inv04 port map ( Y=>nx9583, A=>nx5085);
   ix9584 : inv04 port map ( Y=>nx9585, A=>nx10521);
   ix9586 : inv04 port map ( Y=>nx9587, A=>nx10521);
   ix9588 : inv04 port map ( Y=>nx9589, A=>nx10523);
   ix9590 : inv04 port map ( Y=>nx9591, A=>nx4841);
   ix9592 : inv04 port map ( Y=>nx9593, A=>nx4841);
   ix9594 : inv04 port map ( Y=>nx9595, A=>nx4841);
   ix9596 : inv04 port map ( Y=>nx9597, A=>nx10481);
   ix9598 : inv04 port map ( Y=>nx9599, A=>nx10481);
   ix9600 : inv04 port map ( Y=>nx9601, A=>nx10483);
   ix9602 : inv04 port map ( Y=>nx9603, A=>nx4595);
   ix9604 : inv04 port map ( Y=>nx9605, A=>nx4595);
   ix9606 : inv04 port map ( Y=>nx9607, A=>nx4595);
   ix9608 : inv04 port map ( Y=>nx9609, A=>nx10441);
   ix9610 : inv04 port map ( Y=>nx9611, A=>nx10441);
   ix9612 : inv04 port map ( Y=>nx9613, A=>nx10443);
   ix9614 : inv04 port map ( Y=>nx9615, A=>nx4349);
   ix9616 : inv04 port map ( Y=>nx9617, A=>nx4349);
   ix9618 : inv04 port map ( Y=>nx9619, A=>nx4349);
   ix9620 : inv04 port map ( Y=>nx9621, A=>nx10401);
   ix9622 : inv04 port map ( Y=>nx9623, A=>nx10401);
   ix9624 : inv04 port map ( Y=>nx9625, A=>nx10403);
   ix9626 : inv04 port map ( Y=>nx9627, A=>nx4101);
   ix9628 : inv04 port map ( Y=>nx9629, A=>nx4101);
   ix9630 : inv04 port map ( Y=>nx9631, A=>nx4101);
   ix9632 : inv04 port map ( Y=>nx9633, A=>nx10361);
   ix9634 : inv04 port map ( Y=>nx9635, A=>nx10361);
   ix9636 : inv04 port map ( Y=>nx9637, A=>nx10363);
   ix9638 : inv04 port map ( Y=>nx9639, A=>nx3857);
   ix9640 : inv04 port map ( Y=>nx9641, A=>nx3857);
   ix9642 : inv04 port map ( Y=>nx9643, A=>nx3857);
   ix9644 : inv04 port map ( Y=>nx9645, A=>nx10321);
   ix9646 : inv04 port map ( Y=>nx9647, A=>nx10321);
   ix9648 : inv04 port map ( Y=>nx9649, A=>nx10323);
   ix9650 : inv04 port map ( Y=>nx9651, A=>nx3611);
   ix9652 : inv04 port map ( Y=>nx9653, A=>nx3611);
   ix9654 : inv04 port map ( Y=>nx9655, A=>nx3611);
   ix9656 : inv04 port map ( Y=>nx9657, A=>nx10281);
   ix9658 : inv04 port map ( Y=>nx9659, A=>nx10281);
   ix9660 : inv04 port map ( Y=>nx9661, A=>nx10283);
   ix9662 : inv04 port map ( Y=>nx9663, A=>nx3363);
   ix9664 : inv04 port map ( Y=>nx9665, A=>nx3363);
   ix9666 : inv04 port map ( Y=>nx9667, A=>nx3363);
   ix9668 : inv04 port map ( Y=>nx9669, A=>nx10241);
   ix9670 : inv04 port map ( Y=>nx9671, A=>nx10241);
   ix9672 : inv04 port map ( Y=>nx9673, A=>nx10243);
   ix9674 : inv04 port map ( Y=>nx9675, A=>nx3115);
   ix9676 : inv04 port map ( Y=>nx9677, A=>nx3115);
   ix9678 : inv04 port map ( Y=>nx9679, A=>nx3115);
   ix9680 : inv04 port map ( Y=>nx9681, A=>nx10201);
   ix9682 : inv04 port map ( Y=>nx9683, A=>nx10201);
   ix9684 : inv04 port map ( Y=>nx9685, A=>nx10203);
   ix9686 : inv04 port map ( Y=>nx9687, A=>nx2871);
   ix9688 : inv04 port map ( Y=>nx9689, A=>nx2871);
   ix9690 : inv04 port map ( Y=>nx9691, A=>nx2871);
   ix9692 : inv04 port map ( Y=>nx9693, A=>nx10161);
   ix9694 : inv04 port map ( Y=>nx9695, A=>nx10161);
   ix9696 : inv04 port map ( Y=>nx9697, A=>nx10163);
   ix9698 : inv01 port map ( Y=>nx9699, A=>gen_24_cmp_BSCmp_op2_16);
   ix9700 : inv02 port map ( Y=>nx9701, A=>nx9699);
   ix9702 : inv02 port map ( Y=>nx9703, A=>nx9699);
   ix9704 : inv02 port map ( Y=>nx9705, A=>nx9699);
   ix9706 : inv02 port map ( Y=>nx9707, A=>nx9699);
   ix9708 : inv02 port map ( Y=>nx9709, A=>nx9699);
   ix9710 : inv01 port map ( Y=>nx9711, A=>gen_23_cmp_BSCmp_op2_16);
   ix9712 : inv02 port map ( Y=>nx9713, A=>nx9711);
   ix9714 : inv02 port map ( Y=>nx9715, A=>nx9711);
   ix9716 : inv02 port map ( Y=>nx9717, A=>nx9711);
   ix9718 : inv02 port map ( Y=>nx9719, A=>nx9711);
   ix9720 : inv02 port map ( Y=>nx9721, A=>nx9711);
   ix9722 : inv01 port map ( Y=>nx9723, A=>gen_22_cmp_BSCmp_op2_16);
   ix9724 : inv02 port map ( Y=>nx9725, A=>nx9723);
   ix9726 : inv02 port map ( Y=>nx9727, A=>nx9723);
   ix9728 : inv02 port map ( Y=>nx9729, A=>nx9723);
   ix9730 : inv02 port map ( Y=>nx9731, A=>nx9723);
   ix9732 : inv02 port map ( Y=>nx9733, A=>nx9723);
   ix9734 : inv01 port map ( Y=>nx9735, A=>gen_21_cmp_BSCmp_op2_16);
   ix9736 : inv02 port map ( Y=>nx9737, A=>nx9735);
   ix9738 : inv02 port map ( Y=>nx9739, A=>nx9735);
   ix9740 : inv02 port map ( Y=>nx9741, A=>nx9735);
   ix9742 : inv02 port map ( Y=>nx9743, A=>nx9735);
   ix9744 : inv02 port map ( Y=>nx9745, A=>nx9735);
   ix9746 : inv01 port map ( Y=>nx9747, A=>gen_20_cmp_BSCmp_op2_16);
   ix9748 : inv02 port map ( Y=>nx9749, A=>nx9747);
   ix9750 : inv02 port map ( Y=>nx9751, A=>nx9747);
   ix9752 : inv02 port map ( Y=>nx9753, A=>nx9747);
   ix9754 : inv02 port map ( Y=>nx9755, A=>nx9747);
   ix9756 : inv02 port map ( Y=>nx9757, A=>nx9747);
   ix9758 : inv01 port map ( Y=>nx9759, A=>gen_19_cmp_BSCmp_op2_16);
   ix9760 : inv02 port map ( Y=>nx9761, A=>nx9759);
   ix9762 : inv02 port map ( Y=>nx9763, A=>nx9759);
   ix9764 : inv02 port map ( Y=>nx9765, A=>nx9759);
   ix9766 : inv02 port map ( Y=>nx9767, A=>nx9759);
   ix9768 : inv02 port map ( Y=>nx9769, A=>nx9759);
   ix9770 : inv01 port map ( Y=>nx9771, A=>gen_18_cmp_BSCmp_op2_16);
   ix9772 : inv02 port map ( Y=>nx9773, A=>nx9771);
   ix9774 : inv02 port map ( Y=>nx9775, A=>nx9771);
   ix9776 : inv02 port map ( Y=>nx9777, A=>nx9771);
   ix9778 : inv02 port map ( Y=>nx9779, A=>nx9771);
   ix9780 : inv02 port map ( Y=>nx9781, A=>nx9771);
   ix9782 : inv01 port map ( Y=>nx9783, A=>gen_17_cmp_BSCmp_op2_16);
   ix9784 : inv02 port map ( Y=>nx9785, A=>nx9783);
   ix9786 : inv02 port map ( Y=>nx9787, A=>nx9783);
   ix9788 : inv02 port map ( Y=>nx9789, A=>nx9783);
   ix9790 : inv02 port map ( Y=>nx9791, A=>nx9783);
   ix9792 : inv02 port map ( Y=>nx9793, A=>nx9783);
   ix9794 : inv01 port map ( Y=>nx9795, A=>gen_16_cmp_BSCmp_op2_16);
   ix9796 : inv02 port map ( Y=>nx9797, A=>nx9795);
   ix9798 : inv02 port map ( Y=>nx9799, A=>nx9795);
   ix9800 : inv02 port map ( Y=>nx9801, A=>nx9795);
   ix9802 : inv02 port map ( Y=>nx9803, A=>nx9795);
   ix9804 : inv02 port map ( Y=>nx9805, A=>nx9795);
   ix9806 : inv01 port map ( Y=>nx9807, A=>gen_15_cmp_BSCmp_op2_16);
   ix9808 : inv02 port map ( Y=>nx9809, A=>nx9807);
   ix9810 : inv02 port map ( Y=>nx9811, A=>nx9807);
   ix9812 : inv02 port map ( Y=>nx9813, A=>nx9807);
   ix9814 : inv02 port map ( Y=>nx9815, A=>nx9807);
   ix9816 : inv02 port map ( Y=>nx9817, A=>nx9807);
   ix9818 : inv01 port map ( Y=>nx9819, A=>gen_14_cmp_BSCmp_op2_16);
   ix9820 : inv02 port map ( Y=>nx9821, A=>nx9819);
   ix9822 : inv02 port map ( Y=>nx9823, A=>nx9819);
   ix9824 : inv02 port map ( Y=>nx9825, A=>nx9819);
   ix9826 : inv02 port map ( Y=>nx9827, A=>nx9819);
   ix9828 : inv02 port map ( Y=>nx9829, A=>nx9819);
   ix9830 : inv01 port map ( Y=>nx9831, A=>gen_13_cmp_BSCmp_op2_16);
   ix9832 : inv02 port map ( Y=>nx9833, A=>nx9831);
   ix9834 : inv02 port map ( Y=>nx9835, A=>nx9831);
   ix9836 : inv02 port map ( Y=>nx9837, A=>nx9831);
   ix9838 : inv02 port map ( Y=>nx9839, A=>nx9831);
   ix9840 : inv02 port map ( Y=>nx9841, A=>nx9831);
   ix9842 : inv01 port map ( Y=>nx9843, A=>gen_12_cmp_BSCmp_op2_16);
   ix9844 : inv02 port map ( Y=>nx9845, A=>nx9843);
   ix9846 : inv02 port map ( Y=>nx9847, A=>nx9843);
   ix9848 : inv02 port map ( Y=>nx9849, A=>nx9843);
   ix9850 : inv02 port map ( Y=>nx9851, A=>nx9843);
   ix9852 : inv02 port map ( Y=>nx9853, A=>nx9843);
   ix9854 : inv01 port map ( Y=>nx9855, A=>gen_11_cmp_BSCmp_op2_16);
   ix9856 : inv02 port map ( Y=>nx9857, A=>nx9855);
   ix9858 : inv02 port map ( Y=>nx9859, A=>nx9855);
   ix9860 : inv02 port map ( Y=>nx9861, A=>nx9855);
   ix9862 : inv02 port map ( Y=>nx9863, A=>nx9855);
   ix9864 : inv02 port map ( Y=>nx9865, A=>nx9855);
   ix9866 : inv01 port map ( Y=>nx9867, A=>gen_10_cmp_BSCmp_op2_16);
   ix9868 : inv02 port map ( Y=>nx9869, A=>nx9867);
   ix9870 : inv02 port map ( Y=>nx9871, A=>nx9867);
   ix9872 : inv02 port map ( Y=>nx9873, A=>nx9867);
   ix9874 : inv02 port map ( Y=>nx9875, A=>nx9867);
   ix9876 : inv02 port map ( Y=>nx9877, A=>nx9867);
   ix9878 : inv01 port map ( Y=>nx9879, A=>gen_9_cmp_BSCmp_op2_16);
   ix9880 : inv02 port map ( Y=>nx9881, A=>nx9879);
   ix9882 : inv02 port map ( Y=>nx9883, A=>nx9879);
   ix9884 : inv02 port map ( Y=>nx9885, A=>nx9879);
   ix9886 : inv02 port map ( Y=>nx9887, A=>nx9879);
   ix9888 : inv02 port map ( Y=>nx9889, A=>nx9879);
   ix9890 : inv01 port map ( Y=>nx9891, A=>gen_8_cmp_BSCmp_op2_16);
   ix9892 : inv02 port map ( Y=>nx9893, A=>nx9891);
   ix9894 : inv02 port map ( Y=>nx9895, A=>nx9891);
   ix9896 : inv02 port map ( Y=>nx9897, A=>nx9891);
   ix9898 : inv02 port map ( Y=>nx9899, A=>nx9891);
   ix9900 : inv02 port map ( Y=>nx9901, A=>nx9891);
   ix9902 : inv01 port map ( Y=>nx9903, A=>gen_7_cmp_BSCmp_op2_16);
   ix9904 : inv02 port map ( Y=>nx9905, A=>nx9903);
   ix9906 : inv02 port map ( Y=>nx9907, A=>nx9903);
   ix9908 : inv02 port map ( Y=>nx9909, A=>nx9903);
   ix9910 : inv02 port map ( Y=>nx9911, A=>nx9903);
   ix9912 : inv02 port map ( Y=>nx9913, A=>nx9903);
   ix9914 : inv01 port map ( Y=>nx9915, A=>gen_6_cmp_BSCmp_op2_16);
   ix9916 : inv02 port map ( Y=>nx9917, A=>nx9915);
   ix9918 : inv02 port map ( Y=>nx9919, A=>nx9915);
   ix9920 : inv02 port map ( Y=>nx9921, A=>nx9915);
   ix9922 : inv02 port map ( Y=>nx9923, A=>nx9915);
   ix9924 : inv02 port map ( Y=>nx9925, A=>nx9915);
   ix9926 : inv01 port map ( Y=>nx9927, A=>gen_5_cmp_BSCmp_op2_16);
   ix9928 : inv02 port map ( Y=>nx9929, A=>nx9927);
   ix9930 : inv02 port map ( Y=>nx9931, A=>nx9927);
   ix9932 : inv02 port map ( Y=>nx9933, A=>nx9927);
   ix9934 : inv02 port map ( Y=>nx9935, A=>nx9927);
   ix9936 : inv02 port map ( Y=>nx9937, A=>nx9927);
   ix9938 : inv01 port map ( Y=>nx9939, A=>gen_4_cmp_BSCmp_op2_16);
   ix9940 : inv02 port map ( Y=>nx9941, A=>nx9939);
   ix9942 : inv02 port map ( Y=>nx9943, A=>nx9939);
   ix9944 : inv02 port map ( Y=>nx9945, A=>nx9939);
   ix9946 : inv02 port map ( Y=>nx9947, A=>nx9939);
   ix9948 : inv02 port map ( Y=>nx9949, A=>nx9939);
   ix9950 : inv01 port map ( Y=>nx9951, A=>gen_3_cmp_BSCmp_op2_16);
   ix9952 : inv02 port map ( Y=>nx9953, A=>nx9951);
   ix9954 : inv02 port map ( Y=>nx9955, A=>nx9951);
   ix9956 : inv02 port map ( Y=>nx9957, A=>nx9951);
   ix9958 : inv02 port map ( Y=>nx9959, A=>nx9951);
   ix9960 : inv02 port map ( Y=>nx9961, A=>nx9951);
   ix9962 : inv01 port map ( Y=>nx9963, A=>gen_2_cmp_BSCmp_op2_16);
   ix9964 : inv02 port map ( Y=>nx9965, A=>nx9963);
   ix9966 : inv02 port map ( Y=>nx9967, A=>nx9963);
   ix9968 : inv02 port map ( Y=>nx9969, A=>nx9963);
   ix9970 : inv02 port map ( Y=>nx9971, A=>nx9963);
   ix9972 : inv02 port map ( Y=>nx9973, A=>nx9963);
   ix9974 : inv01 port map ( Y=>nx9975, A=>gen_1_cmp_BSCmp_op2_16);
   ix9976 : inv02 port map ( Y=>nx9977, A=>nx9975);
   ix9978 : inv02 port map ( Y=>nx9979, A=>nx9975);
   ix9980 : inv02 port map ( Y=>nx9981, A=>nx9975);
   ix9982 : inv02 port map ( Y=>nx9983, A=>nx9975);
   ix9984 : inv02 port map ( Y=>nx9985, A=>nx9975);
   ix9986 : inv01 port map ( Y=>nx9987, A=>gen_0_cmp_BSCmp_op2_16);
   ix9988 : inv02 port map ( Y=>nx9989, A=>nx9987);
   ix9990 : inv02 port map ( Y=>nx9991, A=>nx9987);
   ix9992 : inv02 port map ( Y=>nx9993, A=>nx9987);
   ix9994 : inv02 port map ( Y=>nx9995, A=>nx9987);
   ix9996 : inv02 port map ( Y=>nx9997, A=>nx9987);
   ix9998 : buf02 port map ( Y=>nx9999, A=>nx6);
   ix10000 : buf02 port map ( Y=>nx10001, A=>nx6);
   ix10002 : buf02 port map ( Y=>nx10003, A=>nx6);
   ix10004 : buf02 port map ( Y=>nx10005, A=>nx392);
   ix10006 : buf02 port map ( Y=>nx10007, A=>nx392);
   ix10008 : buf02 port map ( Y=>nx10009, A=>nx392);
   ix10010 : buf02 port map ( Y=>nx10011, A=>nx778);
   ix10012 : buf02 port map ( Y=>nx10013, A=>nx778);
   ix10014 : buf02 port map ( Y=>nx10015, A=>nx778);
   ix10016 : buf02 port map ( Y=>nx10017, A=>nx1164);
   ix10018 : buf02 port map ( Y=>nx10019, A=>nx1164);
   ix10020 : buf02 port map ( Y=>nx10021, A=>nx1164);
   ix10022 : buf02 port map ( Y=>nx10023, A=>nx1550);
   ix10024 : buf02 port map ( Y=>nx10025, A=>nx1550);
   ix10026 : buf02 port map ( Y=>nx10027, A=>nx1550);
   ix10028 : buf02 port map ( Y=>nx10029, A=>nx1936);
   ix10030 : buf02 port map ( Y=>nx10031, A=>nx1936);
   ix10032 : buf02 port map ( Y=>nx10033, A=>nx1936);
   ix10034 : buf02 port map ( Y=>nx10035, A=>nx2322);
   ix10036 : buf02 port map ( Y=>nx10037, A=>nx2322);
   ix10038 : buf02 port map ( Y=>nx10039, A=>nx2322);
   ix10040 : buf02 port map ( Y=>nx10041, A=>nx2708);
   ix10042 : buf02 port map ( Y=>nx10043, A=>nx2708);
   ix10044 : buf02 port map ( Y=>nx10045, A=>nx2708);
   ix10046 : buf02 port map ( Y=>nx10047, A=>nx3094);
   ix10048 : buf02 port map ( Y=>nx10049, A=>nx3094);
   ix10050 : buf02 port map ( Y=>nx10051, A=>nx3094);
   ix10052 : buf02 port map ( Y=>nx10053, A=>nx3480);
   ix10054 : buf02 port map ( Y=>nx10055, A=>nx3480);
   ix10056 : buf02 port map ( Y=>nx10057, A=>nx3480);
   ix10058 : buf02 port map ( Y=>nx10059, A=>nx3866);
   ix10060 : buf02 port map ( Y=>nx10061, A=>nx3866);
   ix10062 : buf02 port map ( Y=>nx10063, A=>nx3866);
   ix10064 : buf02 port map ( Y=>nx10065, A=>nx4252);
   ix10066 : buf02 port map ( Y=>nx10067, A=>nx4252);
   ix10068 : buf02 port map ( Y=>nx10069, A=>nx4252);
   ix10070 : buf02 port map ( Y=>nx10071, A=>nx4638);
   ix10072 : buf02 port map ( Y=>nx10073, A=>nx4638);
   ix10074 : buf02 port map ( Y=>nx10075, A=>nx4638);
   ix10076 : buf02 port map ( Y=>nx10077, A=>nx5024);
   ix10078 : buf02 port map ( Y=>nx10079, A=>nx5024);
   ix10080 : buf02 port map ( Y=>nx10081, A=>nx5024);
   ix10082 : buf02 port map ( Y=>nx10083, A=>nx5410);
   ix10084 : buf02 port map ( Y=>nx10085, A=>nx5410);
   ix10086 : buf02 port map ( Y=>nx10087, A=>nx5410);
   ix10088 : buf02 port map ( Y=>nx10089, A=>nx5796);
   ix10090 : buf02 port map ( Y=>nx10091, A=>nx5796);
   ix10092 : buf02 port map ( Y=>nx10093, A=>nx5796);
   ix10094 : buf02 port map ( Y=>nx10095, A=>nx6182);
   ix10096 : buf02 port map ( Y=>nx10097, A=>nx6182);
   ix10098 : buf02 port map ( Y=>nx10099, A=>nx6182);
   ix10100 : buf02 port map ( Y=>nx10101, A=>nx6568);
   ix10102 : buf02 port map ( Y=>nx10103, A=>nx6568);
   ix10104 : buf02 port map ( Y=>nx10105, A=>nx6568);
   ix10106 : buf02 port map ( Y=>nx10107, A=>nx6954);
   ix10108 : buf02 port map ( Y=>nx10109, A=>nx6954);
   ix10110 : buf02 port map ( Y=>nx10111, A=>nx6954);
   ix10112 : buf02 port map ( Y=>nx10113, A=>nx7340);
   ix10114 : buf02 port map ( Y=>nx10115, A=>nx7340);
   ix10116 : buf02 port map ( Y=>nx10117, A=>nx7340);
   ix10118 : buf02 port map ( Y=>nx10119, A=>nx7726);
   ix10120 : buf02 port map ( Y=>nx10121, A=>nx7726);
   ix10122 : buf02 port map ( Y=>nx10123, A=>nx7726);
   ix10124 : buf02 port map ( Y=>nx10125, A=>nx8112);
   ix10126 : buf02 port map ( Y=>nx10127, A=>nx8112);
   ix10128 : buf02 port map ( Y=>nx10129, A=>nx8112);
   ix10130 : buf02 port map ( Y=>nx10131, A=>nx8498);
   ix10132 : buf02 port map ( Y=>nx10133, A=>nx8498);
   ix10134 : buf02 port map ( Y=>nx10135, A=>nx8498);
   ix10136 : buf02 port map ( Y=>nx10137, A=>nx8884);
   ix10138 : buf02 port map ( Y=>nx10139, A=>nx8884);
   ix10140 : buf02 port map ( Y=>nx10141, A=>nx8884);
   ix10142 : buf02 port map ( Y=>nx10143, A=>nx9270);
   ix10144 : buf02 port map ( Y=>nx10145, A=>nx9270);
   ix10146 : buf02 port map ( Y=>nx10147, A=>nx9270);
   ix10150 : inv02 port map ( Y=>nx10151, A=>nx10149);
   ix10152 : inv02 port map ( Y=>nx10153, A=>nx10149);
   ix10154 : inv02 port map ( Y=>nx10155, A=>nx10149);
   ix10156 : inv04 port map ( Y=>nx10157, A=>gen_0_cmp_pMux_1);
   ix10158 : inv04 port map ( Y=>nx10159, A=>gen_0_cmp_pMux_1);
   ix10160 : inv04 port map ( Y=>nx10161, A=>gen_0_cmp_pMux_1);
   ix10162 : inv04 port map ( Y=>nx10163, A=>gen_0_cmp_pMux_1);
   ix10166 : inv02 port map ( Y=>nx10167, A=>nx10165);
   ix10168 : inv02 port map ( Y=>nx10169, A=>nx10165);
   ix10170 : inv02 port map ( Y=>nx10171, A=>nx10165);
   ix10174 : inv02 port map ( Y=>nx10175, A=>nx10173);
   ix10176 : inv02 port map ( Y=>nx10177, A=>nx10173);
   ix10178 : inv02 port map ( Y=>nx10179, A=>nx10173);
   ix10182 : inv02 port map ( Y=>nx10183, A=>nx10181);
   ix10184 : inv02 port map ( Y=>nx10185, A=>nx10181);
   ix10186 : inv02 port map ( Y=>nx10187, A=>nx10181);
   ix10190 : inv02 port map ( Y=>nx10191, A=>nx10189);
   ix10192 : inv02 port map ( Y=>nx10193, A=>nx10189);
   ix10194 : inv02 port map ( Y=>nx10195, A=>nx10189);
   ix10196 : inv04 port map ( Y=>nx10197, A=>gen_1_cmp_pMux_1);
   ix10198 : inv04 port map ( Y=>nx10199, A=>gen_1_cmp_pMux_1);
   ix10200 : inv04 port map ( Y=>nx10201, A=>gen_1_cmp_pMux_1);
   ix10202 : inv04 port map ( Y=>nx10203, A=>gen_1_cmp_pMux_1);
   ix10206 : inv02 port map ( Y=>nx10207, A=>nx10205);
   ix10208 : inv02 port map ( Y=>nx10209, A=>nx10205);
   ix10210 : inv02 port map ( Y=>nx10211, A=>nx10205);
   ix10214 : inv02 port map ( Y=>nx10215, A=>nx10213);
   ix10216 : inv02 port map ( Y=>nx10217, A=>nx10213);
   ix10218 : inv02 port map ( Y=>nx10219, A=>nx10213);
   ix10222 : inv02 port map ( Y=>nx10223, A=>nx10221);
   ix10224 : inv02 port map ( Y=>nx10225, A=>nx10221);
   ix10226 : inv02 port map ( Y=>nx10227, A=>nx10221);
   ix10230 : inv02 port map ( Y=>nx10231, A=>nx10229);
   ix10232 : inv02 port map ( Y=>nx10233, A=>nx10229);
   ix10234 : inv02 port map ( Y=>nx10235, A=>nx10229);
   ix10236 : inv04 port map ( Y=>nx10237, A=>gen_2_cmp_pMux_1);
   ix10238 : inv04 port map ( Y=>nx10239, A=>gen_2_cmp_pMux_1);
   ix10240 : inv04 port map ( Y=>nx10241, A=>gen_2_cmp_pMux_1);
   ix10242 : inv04 port map ( Y=>nx10243, A=>gen_2_cmp_pMux_1);
   ix10246 : inv02 port map ( Y=>nx10247, A=>nx10245);
   ix10248 : inv02 port map ( Y=>nx10249, A=>nx10245);
   ix10250 : inv02 port map ( Y=>nx10251, A=>nx10245);
   ix10254 : inv02 port map ( Y=>nx10255, A=>nx10253);
   ix10256 : inv02 port map ( Y=>nx10257, A=>nx10253);
   ix10258 : inv02 port map ( Y=>nx10259, A=>nx10253);
   ix10262 : inv02 port map ( Y=>nx10263, A=>nx10261);
   ix10264 : inv02 port map ( Y=>nx10265, A=>nx10261);
   ix10266 : inv02 port map ( Y=>nx10267, A=>nx10261);
   ix10270 : inv02 port map ( Y=>nx10271, A=>nx10269);
   ix10272 : inv02 port map ( Y=>nx10273, A=>nx10269);
   ix10274 : inv02 port map ( Y=>nx10275, A=>nx10269);
   ix10276 : inv04 port map ( Y=>nx10277, A=>gen_3_cmp_pMux_1);
   ix10278 : inv04 port map ( Y=>nx10279, A=>gen_3_cmp_pMux_1);
   ix10280 : inv04 port map ( Y=>nx10281, A=>gen_3_cmp_pMux_1);
   ix10282 : inv04 port map ( Y=>nx10283, A=>gen_3_cmp_pMux_1);
   ix10286 : inv02 port map ( Y=>nx10287, A=>nx10285);
   ix10288 : inv02 port map ( Y=>nx10289, A=>nx10285);
   ix10290 : inv02 port map ( Y=>nx10291, A=>nx10285);
   ix10294 : inv02 port map ( Y=>nx10295, A=>nx10293);
   ix10296 : inv02 port map ( Y=>nx10297, A=>nx10293);
   ix10298 : inv02 port map ( Y=>nx10299, A=>nx10293);
   ix10302 : inv02 port map ( Y=>nx10303, A=>nx10301);
   ix10304 : inv02 port map ( Y=>nx10305, A=>nx10301);
   ix10306 : inv02 port map ( Y=>nx10307, A=>nx10301);
   ix10310 : inv02 port map ( Y=>nx10311, A=>nx10309);
   ix10312 : inv02 port map ( Y=>nx10313, A=>nx10309);
   ix10314 : inv02 port map ( Y=>nx10315, A=>nx10309);
   ix10316 : inv04 port map ( Y=>nx10317, A=>gen_4_cmp_pMux_1);
   ix10318 : inv04 port map ( Y=>nx10319, A=>gen_4_cmp_pMux_1);
   ix10320 : inv04 port map ( Y=>nx10321, A=>gen_4_cmp_pMux_1);
   ix10322 : inv04 port map ( Y=>nx10323, A=>gen_4_cmp_pMux_1);
   ix10326 : inv02 port map ( Y=>nx10327, A=>nx10325);
   ix10328 : inv02 port map ( Y=>nx10329, A=>nx10325);
   ix10330 : inv02 port map ( Y=>nx10331, A=>nx10325);
   ix10334 : inv02 port map ( Y=>nx10335, A=>nx10333);
   ix10336 : inv02 port map ( Y=>nx10337, A=>nx10333);
   ix10338 : inv02 port map ( Y=>nx10339, A=>nx10333);
   ix10342 : inv02 port map ( Y=>nx10343, A=>nx10341);
   ix10344 : inv02 port map ( Y=>nx10345, A=>nx10341);
   ix10346 : inv02 port map ( Y=>nx10347, A=>nx10341);
   ix10350 : inv02 port map ( Y=>nx10351, A=>nx10349);
   ix10352 : inv02 port map ( Y=>nx10353, A=>nx10349);
   ix10354 : inv02 port map ( Y=>nx10355, A=>nx10349);
   ix10356 : inv04 port map ( Y=>nx10357, A=>gen_5_cmp_pMux_1);
   ix10358 : inv04 port map ( Y=>nx10359, A=>gen_5_cmp_pMux_1);
   ix10360 : inv04 port map ( Y=>nx10361, A=>gen_5_cmp_pMux_1);
   ix10362 : inv04 port map ( Y=>nx10363, A=>gen_5_cmp_pMux_1);
   ix10366 : inv02 port map ( Y=>nx10367, A=>nx10365);
   ix10368 : inv02 port map ( Y=>nx10369, A=>nx10365);
   ix10370 : inv02 port map ( Y=>nx10371, A=>nx10365);
   ix10374 : inv02 port map ( Y=>nx10375, A=>nx10373);
   ix10376 : inv02 port map ( Y=>nx10377, A=>nx10373);
   ix10378 : inv02 port map ( Y=>nx10379, A=>nx10373);
   ix10382 : inv02 port map ( Y=>nx10383, A=>nx10381);
   ix10384 : inv02 port map ( Y=>nx10385, A=>nx10381);
   ix10386 : inv02 port map ( Y=>nx10387, A=>nx10381);
   ix10390 : inv02 port map ( Y=>nx10391, A=>nx10389);
   ix10392 : inv02 port map ( Y=>nx10393, A=>nx10389);
   ix10394 : inv02 port map ( Y=>nx10395, A=>nx10389);
   ix10396 : inv04 port map ( Y=>nx10397, A=>gen_6_cmp_pMux_1);
   ix10398 : inv04 port map ( Y=>nx10399, A=>gen_6_cmp_pMux_1);
   ix10400 : inv04 port map ( Y=>nx10401, A=>gen_6_cmp_pMux_1);
   ix10402 : inv04 port map ( Y=>nx10403, A=>gen_6_cmp_pMux_1);
   ix10406 : inv02 port map ( Y=>nx10407, A=>nx10405);
   ix10408 : inv02 port map ( Y=>nx10409, A=>nx10405);
   ix10410 : inv02 port map ( Y=>nx10411, A=>nx10405);
   ix10414 : inv02 port map ( Y=>nx10415, A=>nx10413);
   ix10416 : inv02 port map ( Y=>nx10417, A=>nx10413);
   ix10418 : inv02 port map ( Y=>nx10419, A=>nx10413);
   ix10422 : inv02 port map ( Y=>nx10423, A=>nx10421);
   ix10424 : inv02 port map ( Y=>nx10425, A=>nx10421);
   ix10426 : inv02 port map ( Y=>nx10427, A=>nx10421);
   ix10430 : inv02 port map ( Y=>nx10431, A=>nx10429);
   ix10432 : inv02 port map ( Y=>nx10433, A=>nx10429);
   ix10434 : inv02 port map ( Y=>nx10435, A=>nx10429);
   ix10436 : inv04 port map ( Y=>nx10437, A=>gen_7_cmp_pMux_1);
   ix10438 : inv04 port map ( Y=>nx10439, A=>gen_7_cmp_pMux_1);
   ix10440 : inv04 port map ( Y=>nx10441, A=>gen_7_cmp_pMux_1);
   ix10442 : inv04 port map ( Y=>nx10443, A=>gen_7_cmp_pMux_1);
   ix10446 : inv02 port map ( Y=>nx10447, A=>nx10445);
   ix10448 : inv02 port map ( Y=>nx10449, A=>nx10445);
   ix10450 : inv02 port map ( Y=>nx10451, A=>nx10445);
   ix10454 : inv02 port map ( Y=>nx10455, A=>nx10453);
   ix10456 : inv02 port map ( Y=>nx10457, A=>nx10453);
   ix10458 : inv02 port map ( Y=>nx10459, A=>nx10453);
   ix10462 : inv02 port map ( Y=>nx10463, A=>nx10461);
   ix10464 : inv02 port map ( Y=>nx10465, A=>nx10461);
   ix10466 : inv02 port map ( Y=>nx10467, A=>nx10461);
   ix10470 : inv02 port map ( Y=>nx10471, A=>nx10469);
   ix10472 : inv02 port map ( Y=>nx10473, A=>nx10469);
   ix10474 : inv02 port map ( Y=>nx10475, A=>nx10469);
   ix10476 : inv04 port map ( Y=>nx10477, A=>gen_8_cmp_pMux_1);
   ix10478 : inv04 port map ( Y=>nx10479, A=>gen_8_cmp_pMux_1);
   ix10480 : inv04 port map ( Y=>nx10481, A=>gen_8_cmp_pMux_1);
   ix10482 : inv04 port map ( Y=>nx10483, A=>gen_8_cmp_pMux_1);
   ix10486 : inv02 port map ( Y=>nx10487, A=>nx10485);
   ix10488 : inv02 port map ( Y=>nx10489, A=>nx10485);
   ix10490 : inv02 port map ( Y=>nx10491, A=>nx10485);
   ix10494 : inv02 port map ( Y=>nx10495, A=>nx10493);
   ix10496 : inv02 port map ( Y=>nx10497, A=>nx10493);
   ix10498 : inv02 port map ( Y=>nx10499, A=>nx10493);
   ix10502 : inv02 port map ( Y=>nx10503, A=>nx10501);
   ix10504 : inv02 port map ( Y=>nx10505, A=>nx10501);
   ix10506 : inv02 port map ( Y=>nx10507, A=>nx10501);
   ix10510 : inv02 port map ( Y=>nx10511, A=>nx10509);
   ix10512 : inv02 port map ( Y=>nx10513, A=>nx10509);
   ix10514 : inv02 port map ( Y=>nx10515, A=>nx10509);
   ix10516 : inv04 port map ( Y=>nx10517, A=>gen_9_cmp_pMux_1);
   ix10518 : inv04 port map ( Y=>nx10519, A=>gen_9_cmp_pMux_1);
   ix10520 : inv04 port map ( Y=>nx10521, A=>gen_9_cmp_pMux_1);
   ix10522 : inv04 port map ( Y=>nx10523, A=>gen_9_cmp_pMux_1);
   ix10526 : inv02 port map ( Y=>nx10527, A=>nx10525);
   ix10528 : inv02 port map ( Y=>nx10529, A=>nx10525);
   ix10530 : inv02 port map ( Y=>nx10531, A=>nx10525);
   ix10534 : inv02 port map ( Y=>nx10535, A=>nx10533);
   ix10536 : inv02 port map ( Y=>nx10537, A=>nx10533);
   ix10538 : inv02 port map ( Y=>nx10539, A=>nx10533);
   ix10542 : inv02 port map ( Y=>nx10543, A=>nx10541);
   ix10544 : inv02 port map ( Y=>nx10545, A=>nx10541);
   ix10546 : inv02 port map ( Y=>nx10547, A=>nx10541);
   ix10550 : inv02 port map ( Y=>nx10551, A=>nx10549);
   ix10552 : inv02 port map ( Y=>nx10553, A=>nx10549);
   ix10554 : inv02 port map ( Y=>nx10555, A=>nx10549);
   ix10556 : inv04 port map ( Y=>nx10557, A=>gen_10_cmp_pMux_1);
   ix10558 : inv04 port map ( Y=>nx10559, A=>gen_10_cmp_pMux_1);
   ix10560 : inv04 port map ( Y=>nx10561, A=>gen_10_cmp_pMux_1);
   ix10562 : inv04 port map ( Y=>nx10563, A=>gen_10_cmp_pMux_1);
   ix10566 : inv02 port map ( Y=>nx10567, A=>nx10565);
   ix10568 : inv02 port map ( Y=>nx10569, A=>nx10565);
   ix10570 : inv02 port map ( Y=>nx10571, A=>nx10565);
   ix10574 : inv02 port map ( Y=>nx10575, A=>nx10573);
   ix10576 : inv02 port map ( Y=>nx10577, A=>nx10573);
   ix10578 : inv02 port map ( Y=>nx10579, A=>nx10573);
   ix10582 : inv02 port map ( Y=>nx10583, A=>nx10581);
   ix10584 : inv02 port map ( Y=>nx10585, A=>nx10581);
   ix10586 : inv02 port map ( Y=>nx10587, A=>nx10581);
   ix10590 : inv02 port map ( Y=>nx10591, A=>nx10589);
   ix10592 : inv02 port map ( Y=>nx10593, A=>nx10589);
   ix10594 : inv02 port map ( Y=>nx10595, A=>nx10589);
   ix10596 : inv04 port map ( Y=>nx10597, A=>gen_11_cmp_pMux_1);
   ix10598 : inv04 port map ( Y=>nx10599, A=>gen_11_cmp_pMux_1);
   ix10600 : inv04 port map ( Y=>nx10601, A=>gen_11_cmp_pMux_1);
   ix10602 : inv04 port map ( Y=>nx10603, A=>gen_11_cmp_pMux_1);
   ix10606 : inv02 port map ( Y=>nx10607, A=>nx10605);
   ix10608 : inv02 port map ( Y=>nx10609, A=>nx10605);
   ix10610 : inv02 port map ( Y=>nx10611, A=>nx10605);
   ix10614 : inv02 port map ( Y=>nx10615, A=>nx10613);
   ix10616 : inv02 port map ( Y=>nx10617, A=>nx10613);
   ix10618 : inv02 port map ( Y=>nx10619, A=>nx10613);
   ix10622 : inv02 port map ( Y=>nx10623, A=>nx10621);
   ix10624 : inv02 port map ( Y=>nx10625, A=>nx10621);
   ix10626 : inv02 port map ( Y=>nx10627, A=>nx10621);
   ix10630 : inv02 port map ( Y=>nx10631, A=>nx10629);
   ix10632 : inv02 port map ( Y=>nx10633, A=>nx10629);
   ix10634 : inv02 port map ( Y=>nx10635, A=>nx10629);
   ix10636 : inv04 port map ( Y=>nx10637, A=>gen_12_cmp_pMux_1);
   ix10638 : inv04 port map ( Y=>nx10639, A=>gen_12_cmp_pMux_1);
   ix10640 : inv04 port map ( Y=>nx10641, A=>gen_12_cmp_pMux_1);
   ix10642 : inv04 port map ( Y=>nx10643, A=>gen_12_cmp_pMux_1);
   ix10646 : inv02 port map ( Y=>nx10647, A=>nx10645);
   ix10648 : inv02 port map ( Y=>nx10649, A=>nx10645);
   ix10650 : inv02 port map ( Y=>nx10651, A=>nx10645);
   ix10654 : inv02 port map ( Y=>nx10655, A=>nx10653);
   ix10656 : inv02 port map ( Y=>nx10657, A=>nx10653);
   ix10658 : inv02 port map ( Y=>nx10659, A=>nx10653);
   ix10662 : inv02 port map ( Y=>nx10663, A=>nx10661);
   ix10664 : inv02 port map ( Y=>nx10665, A=>nx10661);
   ix10666 : inv02 port map ( Y=>nx10667, A=>nx10661);
   ix10670 : inv02 port map ( Y=>nx10671, A=>nx10669);
   ix10672 : inv02 port map ( Y=>nx10673, A=>nx10669);
   ix10674 : inv02 port map ( Y=>nx10675, A=>nx10669);
   ix10676 : inv04 port map ( Y=>nx10677, A=>gen_13_cmp_pMux_1);
   ix10678 : inv04 port map ( Y=>nx10679, A=>gen_13_cmp_pMux_1);
   ix10680 : inv04 port map ( Y=>nx10681, A=>gen_13_cmp_pMux_1);
   ix10682 : inv04 port map ( Y=>nx10683, A=>gen_13_cmp_pMux_1);
   ix10686 : inv02 port map ( Y=>nx10687, A=>nx10685);
   ix10688 : inv02 port map ( Y=>nx10689, A=>nx10685);
   ix10690 : inv02 port map ( Y=>nx10691, A=>nx10685);
   ix10694 : inv02 port map ( Y=>nx10695, A=>nx10693);
   ix10696 : inv02 port map ( Y=>nx10697, A=>nx10693);
   ix10698 : inv02 port map ( Y=>nx10699, A=>nx10693);
   ix10702 : inv02 port map ( Y=>nx10703, A=>nx10701);
   ix10704 : inv02 port map ( Y=>nx10705, A=>nx10701);
   ix10706 : inv02 port map ( Y=>nx10707, A=>nx10701);
   ix10710 : inv02 port map ( Y=>nx10711, A=>nx10709);
   ix10712 : inv02 port map ( Y=>nx10713, A=>nx10709);
   ix10714 : inv02 port map ( Y=>nx10715, A=>nx10709);
   ix10716 : inv04 port map ( Y=>nx10717, A=>gen_14_cmp_pMux_1);
   ix10718 : inv04 port map ( Y=>nx10719, A=>gen_14_cmp_pMux_1);
   ix10720 : inv04 port map ( Y=>nx10721, A=>gen_14_cmp_pMux_1);
   ix10722 : inv04 port map ( Y=>nx10723, A=>gen_14_cmp_pMux_1);
   ix10726 : inv02 port map ( Y=>nx10727, A=>nx10725);
   ix10728 : inv02 port map ( Y=>nx10729, A=>nx10725);
   ix10730 : inv02 port map ( Y=>nx10731, A=>nx10725);
   ix10734 : inv02 port map ( Y=>nx10735, A=>nx10733);
   ix10736 : inv02 port map ( Y=>nx10737, A=>nx10733);
   ix10738 : inv02 port map ( Y=>nx10739, A=>nx10733);
   ix10742 : inv02 port map ( Y=>nx10743, A=>nx10741);
   ix10744 : inv02 port map ( Y=>nx10745, A=>nx10741);
   ix10746 : inv02 port map ( Y=>nx10747, A=>nx10741);
   ix10750 : inv02 port map ( Y=>nx10751, A=>nx10749);
   ix10752 : inv02 port map ( Y=>nx10753, A=>nx10749);
   ix10754 : inv02 port map ( Y=>nx10755, A=>nx10749);
   ix10756 : inv04 port map ( Y=>nx10757, A=>gen_15_cmp_pMux_1);
   ix10758 : inv04 port map ( Y=>nx10759, A=>gen_15_cmp_pMux_1);
   ix10760 : inv04 port map ( Y=>nx10761, A=>gen_15_cmp_pMux_1);
   ix10762 : inv04 port map ( Y=>nx10763, A=>gen_15_cmp_pMux_1);
   ix10766 : inv02 port map ( Y=>nx10767, A=>nx10765);
   ix10768 : inv02 port map ( Y=>nx10769, A=>nx10765);
   ix10770 : inv02 port map ( Y=>nx10771, A=>nx10765);
   ix10774 : inv02 port map ( Y=>nx10775, A=>nx10773);
   ix10776 : inv02 port map ( Y=>nx10777, A=>nx10773);
   ix10778 : inv02 port map ( Y=>nx10779, A=>nx10773);
   ix10782 : inv02 port map ( Y=>nx10783, A=>nx10781);
   ix10784 : inv02 port map ( Y=>nx10785, A=>nx10781);
   ix10786 : inv02 port map ( Y=>nx10787, A=>nx10781);
   ix10790 : inv02 port map ( Y=>nx10791, A=>nx10789);
   ix10792 : inv02 port map ( Y=>nx10793, A=>nx10789);
   ix10794 : inv02 port map ( Y=>nx10795, A=>nx10789);
   ix10796 : inv04 port map ( Y=>nx10797, A=>gen_16_cmp_pMux_1);
   ix10798 : inv04 port map ( Y=>nx10799, A=>gen_16_cmp_pMux_1);
   ix10800 : inv04 port map ( Y=>nx10801, A=>gen_16_cmp_pMux_1);
   ix10802 : inv04 port map ( Y=>nx10803, A=>gen_16_cmp_pMux_1);
   ix10806 : inv02 port map ( Y=>nx10807, A=>nx10805);
   ix10808 : inv02 port map ( Y=>nx10809, A=>nx10805);
   ix10810 : inv02 port map ( Y=>nx10811, A=>nx10805);
   ix10814 : inv02 port map ( Y=>nx10815, A=>nx10813);
   ix10816 : inv02 port map ( Y=>nx10817, A=>nx10813);
   ix10818 : inv02 port map ( Y=>nx10819, A=>nx10813);
   ix10822 : inv02 port map ( Y=>nx10823, A=>nx10821);
   ix10824 : inv02 port map ( Y=>nx10825, A=>nx10821);
   ix10826 : inv02 port map ( Y=>nx10827, A=>nx10821);
   ix10830 : inv02 port map ( Y=>nx10831, A=>nx10829);
   ix10832 : inv02 port map ( Y=>nx10833, A=>nx10829);
   ix10834 : inv02 port map ( Y=>nx10835, A=>nx10829);
   ix10836 : inv04 port map ( Y=>nx10837, A=>gen_17_cmp_pMux_1);
   ix10838 : inv04 port map ( Y=>nx10839, A=>gen_17_cmp_pMux_1);
   ix10840 : inv04 port map ( Y=>nx10841, A=>gen_17_cmp_pMux_1);
   ix10842 : inv04 port map ( Y=>nx10843, A=>gen_17_cmp_pMux_1);
   ix10846 : inv02 port map ( Y=>nx10847, A=>nx10845);
   ix10848 : inv02 port map ( Y=>nx10849, A=>nx10845);
   ix10850 : inv02 port map ( Y=>nx10851, A=>nx10845);
   ix10854 : inv02 port map ( Y=>nx10855, A=>nx10853);
   ix10856 : inv02 port map ( Y=>nx10857, A=>nx10853);
   ix10858 : inv02 port map ( Y=>nx10859, A=>nx10853);
   ix10862 : inv02 port map ( Y=>nx10863, A=>nx10861);
   ix10864 : inv02 port map ( Y=>nx10865, A=>nx10861);
   ix10866 : inv02 port map ( Y=>nx10867, A=>nx10861);
   ix10870 : inv02 port map ( Y=>nx10871, A=>nx10869);
   ix10872 : inv02 port map ( Y=>nx10873, A=>nx10869);
   ix10874 : inv02 port map ( Y=>nx10875, A=>nx10869);
   ix10876 : inv04 port map ( Y=>nx10877, A=>gen_18_cmp_pMux_1);
   ix10878 : inv04 port map ( Y=>nx10879, A=>gen_18_cmp_pMux_1);
   ix10880 : inv04 port map ( Y=>nx10881, A=>gen_18_cmp_pMux_1);
   ix10882 : inv04 port map ( Y=>nx10883, A=>gen_18_cmp_pMux_1);
   ix10886 : inv02 port map ( Y=>nx10887, A=>nx10885);
   ix10888 : inv02 port map ( Y=>nx10889, A=>nx10885);
   ix10890 : inv02 port map ( Y=>nx10891, A=>nx10885);
   ix10894 : inv02 port map ( Y=>nx10895, A=>nx10893);
   ix10896 : inv02 port map ( Y=>nx10897, A=>nx10893);
   ix10898 : inv02 port map ( Y=>nx10899, A=>nx10893);
   ix10902 : inv02 port map ( Y=>nx10903, A=>nx10901);
   ix10904 : inv02 port map ( Y=>nx10905, A=>nx10901);
   ix10906 : inv02 port map ( Y=>nx10907, A=>nx10901);
   ix10910 : inv02 port map ( Y=>nx10911, A=>nx10909);
   ix10912 : inv02 port map ( Y=>nx10913, A=>nx10909);
   ix10914 : inv02 port map ( Y=>nx10915, A=>nx10909);
   ix10916 : inv04 port map ( Y=>nx10917, A=>gen_19_cmp_pMux_1);
   ix10918 : inv04 port map ( Y=>nx10919, A=>gen_19_cmp_pMux_1);
   ix10920 : inv04 port map ( Y=>nx10921, A=>gen_19_cmp_pMux_1);
   ix10922 : inv04 port map ( Y=>nx10923, A=>gen_19_cmp_pMux_1);
   ix10926 : inv02 port map ( Y=>nx10927, A=>nx10925);
   ix10928 : inv02 port map ( Y=>nx10929, A=>nx10925);
   ix10930 : inv02 port map ( Y=>nx10931, A=>nx10925);
   ix10934 : inv02 port map ( Y=>nx10935, A=>nx10933);
   ix10936 : inv02 port map ( Y=>nx10937, A=>nx10933);
   ix10938 : inv02 port map ( Y=>nx10939, A=>nx10933);
   ix10942 : inv02 port map ( Y=>nx10943, A=>nx10941);
   ix10944 : inv02 port map ( Y=>nx10945, A=>nx10941);
   ix10946 : inv02 port map ( Y=>nx10947, A=>nx10941);
   ix10950 : inv02 port map ( Y=>nx10951, A=>nx10949);
   ix10952 : inv02 port map ( Y=>nx10953, A=>nx10949);
   ix10954 : inv02 port map ( Y=>nx10955, A=>nx10949);
   ix10956 : inv04 port map ( Y=>nx10957, A=>gen_20_cmp_pMux_1);
   ix10958 : inv04 port map ( Y=>nx10959, A=>gen_20_cmp_pMux_1);
   ix10960 : inv04 port map ( Y=>nx10961, A=>gen_20_cmp_pMux_1);
   ix10962 : inv04 port map ( Y=>nx10963, A=>gen_20_cmp_pMux_1);
   ix10966 : inv02 port map ( Y=>nx10967, A=>nx10965);
   ix10968 : inv02 port map ( Y=>nx10969, A=>nx10965);
   ix10970 : inv02 port map ( Y=>nx10971, A=>nx10965);
   ix10974 : inv02 port map ( Y=>nx10975, A=>nx10973);
   ix10976 : inv02 port map ( Y=>nx10977, A=>nx10973);
   ix10978 : inv02 port map ( Y=>nx10979, A=>nx10973);
   ix10982 : inv02 port map ( Y=>nx10983, A=>nx10981);
   ix10984 : inv02 port map ( Y=>nx10985, A=>nx10981);
   ix10986 : inv02 port map ( Y=>nx10987, A=>nx10981);
   ix10990 : inv02 port map ( Y=>nx10991, A=>nx10989);
   ix10992 : inv02 port map ( Y=>nx10993, A=>nx10989);
   ix10994 : inv02 port map ( Y=>nx10995, A=>nx10989);
   ix10996 : inv04 port map ( Y=>nx10997, A=>gen_21_cmp_pMux_1);
   ix10998 : inv04 port map ( Y=>nx10999, A=>gen_21_cmp_pMux_1);
   ix11000 : inv04 port map ( Y=>nx11001, A=>gen_21_cmp_pMux_1);
   ix11002 : inv04 port map ( Y=>nx11003, A=>gen_21_cmp_pMux_1);
   ix11006 : inv02 port map ( Y=>nx11007, A=>nx11005);
   ix11008 : inv02 port map ( Y=>nx11009, A=>nx11005);
   ix11010 : inv02 port map ( Y=>nx11011, A=>nx11005);
   ix11014 : inv02 port map ( Y=>nx11015, A=>nx11013);
   ix11016 : inv02 port map ( Y=>nx11017, A=>nx11013);
   ix11018 : inv02 port map ( Y=>nx11019, A=>nx11013);
   ix11022 : inv02 port map ( Y=>nx11023, A=>nx11021);
   ix11024 : inv02 port map ( Y=>nx11025, A=>nx11021);
   ix11026 : inv02 port map ( Y=>nx11027, A=>nx11021);
   ix11030 : inv02 port map ( Y=>nx11031, A=>nx11029);
   ix11032 : inv02 port map ( Y=>nx11033, A=>nx11029);
   ix11034 : inv02 port map ( Y=>nx11035, A=>nx11029);
   ix11036 : inv04 port map ( Y=>nx11037, A=>gen_22_cmp_pMux_1);
   ix11038 : inv04 port map ( Y=>nx11039, A=>gen_22_cmp_pMux_1);
   ix11040 : inv04 port map ( Y=>nx11041, A=>gen_22_cmp_pMux_1);
   ix11042 : inv04 port map ( Y=>nx11043, A=>gen_22_cmp_pMux_1);
   ix11046 : inv02 port map ( Y=>nx11047, A=>nx11045);
   ix11048 : inv02 port map ( Y=>nx11049, A=>nx11045);
   ix11050 : inv02 port map ( Y=>nx11051, A=>nx11045);
   ix11054 : inv02 port map ( Y=>nx11055, A=>nx11053);
   ix11056 : inv02 port map ( Y=>nx11057, A=>nx11053);
   ix11058 : inv02 port map ( Y=>nx11059, A=>nx11053);
   ix11062 : inv02 port map ( Y=>nx11063, A=>nx11061);
   ix11064 : inv02 port map ( Y=>nx11065, A=>nx11061);
   ix11066 : inv02 port map ( Y=>nx11067, A=>nx11061);
   ix11070 : inv02 port map ( Y=>nx11071, A=>nx11069);
   ix11072 : inv02 port map ( Y=>nx11073, A=>nx11069);
   ix11074 : inv02 port map ( Y=>nx11075, A=>nx11069);
   ix11076 : inv04 port map ( Y=>nx11077, A=>gen_23_cmp_pMux_1);
   ix11078 : inv04 port map ( Y=>nx11079, A=>gen_23_cmp_pMux_1);
   ix11080 : inv04 port map ( Y=>nx11081, A=>gen_23_cmp_pMux_1);
   ix11082 : inv04 port map ( Y=>nx11083, A=>gen_23_cmp_pMux_1);
   ix11086 : inv02 port map ( Y=>nx11087, A=>nx11085);
   ix11088 : inv02 port map ( Y=>nx11089, A=>nx11085);
   ix11090 : inv02 port map ( Y=>nx11091, A=>nx11085);
   ix11094 : inv02 port map ( Y=>nx11095, A=>nx11093);
   ix11096 : inv02 port map ( Y=>nx11097, A=>nx11093);
   ix11098 : inv02 port map ( Y=>nx11099, A=>nx11093);
   ix11102 : inv02 port map ( Y=>nx11103, A=>nx11101);
   ix11104 : inv02 port map ( Y=>nx11105, A=>nx11101);
   ix11106 : inv02 port map ( Y=>nx11107, A=>nx11101);
   ix11110 : inv02 port map ( Y=>nx11111, A=>nx11109);
   ix11112 : inv02 port map ( Y=>nx11113, A=>nx11109);
   ix11114 : inv02 port map ( Y=>nx11115, A=>nx11109);
   ix11116 : inv04 port map ( Y=>nx11117, A=>gen_24_cmp_pMux_1);
   ix11118 : inv04 port map ( Y=>nx11119, A=>gen_24_cmp_pMux_1);
   ix11120 : inv04 port map ( Y=>nx11121, A=>gen_24_cmp_pMux_1);
   ix11122 : inv04 port map ( Y=>nx11123, A=>gen_24_cmp_pMux_1);
   ix11126 : inv02 port map ( Y=>nx11127, A=>nx11125);
   ix11128 : inv02 port map ( Y=>nx11129, A=>nx11125);
   ix11130 : inv02 port map ( Y=>nx11131, A=>nx11125);
   ix11134 : inv02 port map ( Y=>nx11135, A=>nx11133);
   ix11136 : inv02 port map ( Y=>nx11137, A=>nx11133);
   ix11138 : inv02 port map ( Y=>nx11139, A=>nx11133);
   ix11142 : inv02 port map ( Y=>nx11143, A=>nx11141);
   ix11144 : inv02 port map ( Y=>nx11145, A=>nx11141);
   ix11146 : inv02 port map ( Y=>nx11147, A=>nx11141);
   ix2861 : nor02_2x port map ( Y=>nx10149, A0=>nx2871, A1=>gen_0_cmp_pMux_0
   );
   ix2870 : nor02_2x port map ( Y=>nx10165, A0=>gen_0_cmp_pMux_2, A1=>nx2862
   );
   ix2880 : xnor2 port map ( Y=>nx10173, A0=>gen_0_cmp_pMux_0, A1=>nx10161);
   ix2884 : aoi21 port map ( Y=>nx10181, A0=>gen_0_cmp_pMux_1, A1=>
      gen_0_cmp_pMux_0, B0=>nx2871);
   ix3106 : nor02_2x port map ( Y=>nx10189, A0=>nx3115, A1=>gen_1_cmp_pMux_0
   );
   ix3114 : nor02_2x port map ( Y=>nx10205, A0=>gen_1_cmp_pMux_2, A1=>nx3107
   );
   ix3124 : xnor2 port map ( Y=>nx10213, A0=>gen_1_cmp_pMux_0, A1=>nx10201);
   ix3130 : aoi21 port map ( Y=>nx10221, A0=>gen_1_cmp_pMux_1, A1=>
      gen_1_cmp_pMux_0, B0=>nx3115);
   ix3355 : nor02_2x port map ( Y=>nx10229, A0=>nx3363, A1=>gen_2_cmp_pMux_0
   );
   ix3362 : nor02_2x port map ( Y=>nx10245, A0=>gen_2_cmp_pMux_2, A1=>nx3356
   );
   ix3372 : xnor2 port map ( Y=>nx10253, A0=>gen_2_cmp_pMux_0, A1=>nx10241);
   ix3378 : aoi21 port map ( Y=>nx10261, A0=>gen_2_cmp_pMux_1, A1=>
      gen_2_cmp_pMux_0, B0=>nx3363);
   ix3601 : nor02_2x port map ( Y=>nx10269, A0=>nx3611, A1=>gen_3_cmp_pMux_0
   );
   ix3610 : nor02_2x port map ( Y=>nx10285, A0=>gen_3_cmp_pMux_2, A1=>nx3603
   );
   ix3620 : xnor2 port map ( Y=>nx10293, A0=>gen_3_cmp_pMux_0, A1=>nx10281);
   ix3626 : aoi21 port map ( Y=>nx10301, A0=>gen_3_cmp_pMux_1, A1=>
      gen_3_cmp_pMux_0, B0=>nx3611);
   ix3848 : nor02_2x port map ( Y=>nx10309, A0=>nx3857, A1=>gen_4_cmp_pMux_0
   );
   ix3856 : nor02_2x port map ( Y=>nx10325, A0=>gen_4_cmp_pMux_2, A1=>nx3849
   );
   ix3866 : xnor2 port map ( Y=>nx10333, A0=>gen_4_cmp_pMux_0, A1=>nx10321);
   ix3871 : aoi21 port map ( Y=>nx10341, A0=>gen_4_cmp_pMux_1, A1=>
      gen_4_cmp_pMux_0, B0=>nx3857);
   ix4092 : nor02_2x port map ( Y=>nx10349, A0=>nx4101, A1=>gen_5_cmp_pMux_0
   );
   ix4100 : nor02_2x port map ( Y=>nx10365, A0=>gen_5_cmp_pMux_2, A1=>nx4093
   );
   ix4110 : xnor2 port map ( Y=>nx10373, A0=>gen_5_cmp_pMux_0, A1=>nx10361);
   ix4116 : aoi21 port map ( Y=>nx10381, A0=>gen_5_cmp_pMux_1, A1=>
      gen_5_cmp_pMux_0, B0=>nx4101);
   ix4339 : nor02_2x port map ( Y=>nx10389, A0=>nx4349, A1=>gen_6_cmp_pMux_0
   );
   ix4348 : nor02_2x port map ( Y=>nx10405, A0=>gen_6_cmp_pMux_2, A1=>nx4340
   );
   ix4358 : xnor2 port map ( Y=>nx10413, A0=>gen_6_cmp_pMux_0, A1=>nx10401);
   ix4362 : aoi21 port map ( Y=>nx10421, A0=>gen_6_cmp_pMux_1, A1=>
      gen_6_cmp_pMux_0, B0=>nx4349);
   ix4586 : nor02_2x port map ( Y=>nx10429, A0=>nx4595, A1=>gen_7_cmp_pMux_0
   );
   ix4594 : nor02_2x port map ( Y=>nx10445, A0=>gen_7_cmp_pMux_2, A1=>nx4587
   );
   ix4604 : xnor2 port map ( Y=>nx10453, A0=>gen_7_cmp_pMux_0, A1=>nx10441);
   ix4610 : aoi21 port map ( Y=>nx10461, A0=>gen_7_cmp_pMux_1, A1=>
      gen_7_cmp_pMux_0, B0=>nx4595);
   ix4833 : nor02_2x port map ( Y=>nx10469, A0=>nx4841, A1=>gen_8_cmp_pMux_0
   );
   ix4840 : nor02_2x port map ( Y=>nx10485, A0=>gen_8_cmp_pMux_2, A1=>nx4834
   );
   ix4850 : xnor2 port map ( Y=>nx10493, A0=>gen_8_cmp_pMux_0, A1=>nx10481);
   ix4856 : aoi21 port map ( Y=>nx10501, A0=>gen_8_cmp_pMux_1, A1=>
      gen_8_cmp_pMux_0, B0=>nx4841);
   ix5076 : nor02_2x port map ( Y=>nx10509, A0=>nx5085, A1=>gen_9_cmp_pMux_0
   );
   ix5084 : nor02_2x port map ( Y=>nx10525, A0=>gen_9_cmp_pMux_2, A1=>nx5077
   );
   ix5094 : xnor2 port map ( Y=>nx10533, A0=>gen_9_cmp_pMux_0, A1=>nx10521);
   ix5100 : aoi21 port map ( Y=>nx10541, A0=>gen_9_cmp_pMux_1, A1=>
      gen_9_cmp_pMux_0, B0=>nx5085);
   ix5326 : nor02_2x port map ( Y=>nx10549, A0=>nx5335, A1=>
      gen_10_cmp_pMux_0);
   ix5334 : nor02_2x port map ( Y=>nx10565, A0=>gen_10_cmp_pMux_2, A1=>
      nx5327);
   ix5344 : xnor2 port map ( Y=>nx10573, A0=>gen_10_cmp_pMux_0, A1=>nx10561
   );
   ix5350 : aoi21 port map ( Y=>nx10581, A0=>gen_10_cmp_pMux_1, A1=>
      gen_10_cmp_pMux_0, B0=>nx5335);
   ix5575 : nor02_2x port map ( Y=>nx10589, A0=>nx5585, A1=>
      gen_11_cmp_pMux_0);
   ix5584 : nor02_2x port map ( Y=>nx10605, A0=>gen_11_cmp_pMux_2, A1=>
      nx5577);
   ix5594 : xnor2 port map ( Y=>nx10613, A0=>gen_11_cmp_pMux_0, A1=>nx10601
   );
   ix5600 : aoi21 port map ( Y=>nx10621, A0=>gen_11_cmp_pMux_1, A1=>
      gen_11_cmp_pMux_0, B0=>nx5585);
   ix5820 : nor02_2x port map ( Y=>nx10629, A0=>nx5829, A1=>
      gen_12_cmp_pMux_0);
   ix5828 : nor02_2x port map ( Y=>nx10645, A0=>gen_12_cmp_pMux_2, A1=>
      nx5821);
   ix5838 : xnor2 port map ( Y=>nx10653, A0=>gen_12_cmp_pMux_0, A1=>nx10641
   );
   ix5844 : aoi21 port map ( Y=>nx10661, A0=>gen_12_cmp_pMux_1, A1=>
      gen_12_cmp_pMux_0, B0=>nx5829);
   ix6066 : nor02_2x port map ( Y=>nx10669, A0=>nx6075, A1=>
      gen_13_cmp_pMux_0);
   ix6074 : nor02_2x port map ( Y=>nx10685, A0=>gen_13_cmp_pMux_2, A1=>
      nx6067);
   ix6084 : xnor2 port map ( Y=>nx10693, A0=>gen_13_cmp_pMux_0, A1=>nx10681
   );
   ix6090 : aoi21 port map ( Y=>nx10701, A0=>gen_13_cmp_pMux_1, A1=>
      gen_13_cmp_pMux_0, B0=>nx6075);
   ix6313 : nor02_2x port map ( Y=>nx10709, A0=>nx6323, A1=>
      gen_14_cmp_pMux_0);
   ix6322 : nor02_2x port map ( Y=>nx10725, A0=>gen_14_cmp_pMux_2, A1=>
      nx6314);
   ix6332 : xnor2 port map ( Y=>nx10733, A0=>gen_14_cmp_pMux_0, A1=>nx10721
   );
   ix6336 : aoi21 port map ( Y=>nx10741, A0=>gen_14_cmp_pMux_1, A1=>
      gen_14_cmp_pMux_0, B0=>nx6323);
   ix6560 : nor02_2x port map ( Y=>nx10749, A0=>nx6569, A1=>
      gen_15_cmp_pMux_0);
   ix6568 : nor02_2x port map ( Y=>nx10765, A0=>gen_15_cmp_pMux_2, A1=>
      nx6561);
   ix6577 : xnor2 port map ( Y=>nx10773, A0=>gen_15_cmp_pMux_0, A1=>nx10761
   );
   ix6582 : aoi21 port map ( Y=>nx10781, A0=>gen_15_cmp_pMux_1, A1=>
      gen_15_cmp_pMux_0, B0=>nx6569);
   ix6807 : nor02_2x port map ( Y=>nx10789, A0=>nx6815, A1=>
      gen_16_cmp_pMux_0);
   ix6814 : nor02_2x port map ( Y=>nx10805, A0=>gen_16_cmp_pMux_2, A1=>
      nx6808);
   ix6824 : xnor2 port map ( Y=>nx10813, A0=>gen_16_cmp_pMux_0, A1=>nx10801
   );
   ix6830 : aoi21 port map ( Y=>nx10821, A0=>gen_16_cmp_pMux_1, A1=>
      gen_16_cmp_pMux_0, B0=>nx6815);
   ix7048 : nor02_2x port map ( Y=>nx10829, A0=>nx7057, A1=>
      gen_17_cmp_pMux_0);
   ix7056 : nor02_2x port map ( Y=>nx10845, A0=>gen_17_cmp_pMux_2, A1=>
      nx7049);
   ix7066 : xnor2 port map ( Y=>nx10853, A0=>gen_17_cmp_pMux_0, A1=>nx10841
   );
   ix7072 : aoi21 port map ( Y=>nx10861, A0=>gen_17_cmp_pMux_1, A1=>
      gen_17_cmp_pMux_0, B0=>nx7057);
   ix7295 : nor02_2x port map ( Y=>nx10869, A0=>nx7305, A1=>
      gen_18_cmp_pMux_0);
   ix7304 : nor02_2x port map ( Y=>nx10885, A0=>gen_18_cmp_pMux_2, A1=>
      nx7297);
   ix7314 : xnor2 port map ( Y=>nx10893, A0=>gen_18_cmp_pMux_0, A1=>nx10881
   );
   ix7320 : aoi21 port map ( Y=>nx10901, A0=>gen_18_cmp_pMux_1, A1=>
      gen_18_cmp_pMux_0, B0=>nx7305);
   ix7544 : nor02_2x port map ( Y=>nx10909, A0=>nx7553, A1=>
      gen_19_cmp_pMux_0);
   ix7552 : nor02_2x port map ( Y=>nx10925, A0=>gen_19_cmp_pMux_2, A1=>
      nx7545);
   ix7562 : xnor2 port map ( Y=>nx10933, A0=>gen_19_cmp_pMux_0, A1=>nx10921
   );
   ix7568 : aoi21 port map ( Y=>nx10941, A0=>gen_19_cmp_pMux_1, A1=>
      gen_19_cmp_pMux_0, B0=>nx7553);
   ix7791 : nor02_2x port map ( Y=>nx10949, A0=>nx7801, A1=>
      gen_20_cmp_pMux_0);
   ix7800 : nor02_2x port map ( Y=>nx10965, A0=>gen_20_cmp_pMux_2, A1=>
      nx7792);
   ix7810 : xnor2 port map ( Y=>nx10973, A0=>gen_20_cmp_pMux_0, A1=>nx10961
   );
   ix7814 : aoi21 port map ( Y=>nx10981, A0=>gen_20_cmp_pMux_1, A1=>
      gen_20_cmp_pMux_0, B0=>nx7801);
   ix8038 : nor02_2x port map ( Y=>nx10989, A0=>nx8047, A1=>
      gen_21_cmp_pMux_0);
   ix8046 : nor02_2x port map ( Y=>nx11005, A0=>gen_21_cmp_pMux_2, A1=>
      nx8039);
   ix8056 : xnor2 port map ( Y=>nx11013, A0=>gen_21_cmp_pMux_0, A1=>nx11001
   );
   ix8062 : aoi21 port map ( Y=>nx11021, A0=>gen_21_cmp_pMux_1, A1=>
      gen_21_cmp_pMux_0, B0=>nx8047);
   ix8282 : nor02_2x port map ( Y=>nx11029, A0=>nx8291, A1=>
      gen_22_cmp_pMux_0);
   ix8290 : nor02_2x port map ( Y=>nx11045, A0=>gen_22_cmp_pMux_2, A1=>
      nx8283);
   ix8300 : xnor2 port map ( Y=>nx11053, A0=>gen_22_cmp_pMux_0, A1=>nx11041
   );
   ix8306 : aoi21 port map ( Y=>nx11061, A0=>gen_22_cmp_pMux_1, A1=>
      gen_22_cmp_pMux_0, B0=>nx8291);
   ix8532 : nor02_2x port map ( Y=>nx11069, A0=>nx8541, A1=>
      gen_23_cmp_pMux_0);
   ix8540 : nor02_2x port map ( Y=>nx11085, A0=>gen_23_cmp_pMux_2, A1=>
      nx8533);
   ix8550 : xnor2 port map ( Y=>nx11093, A0=>gen_23_cmp_pMux_0, A1=>nx11081
   );
   ix8556 : aoi21 port map ( Y=>nx11101, A0=>gen_23_cmp_pMux_1, A1=>
      gen_23_cmp_pMux_0, B0=>nx8541);
   ix8778 : nor02_2x port map ( Y=>nx11109, A0=>nx8787, A1=>
      gen_24_cmp_pMux_0);
   ix8786 : nor02_2x port map ( Y=>nx11125, A0=>gen_24_cmp_pMux_2, A1=>
      nx8779);
   ix8796 : xnor2 port map ( Y=>nx11133, A0=>gen_24_cmp_pMux_0, A1=>nx11121
   );
   ix8802 : aoi21 port map ( Y=>nx11141, A0=>gen_24_cmp_pMux_1, A1=>
      gen_24_cmp_pMux_0, B0=>nx8787);
   ix9687 : nand02 port map ( Y=>nx9373, A0=>nx11157, A1=>nx9365);
   ix11156 : inv01 port map ( Y=>nx11157, A=>nx9353);
   ix2824 : mux21 port map ( Y=>nx2823, A0=>nx9361, A1=>nx9357, S0=>nx11201
   );
   ix2814 : mux21 port map ( Y=>nx2813, A0=>nx11197, A1=>nx9361, S0=>nx11201
   );
   ix11158 : inv02 port map ( Y=>nx11159, A=>nx11201);
   ix11160 : inv02 port map ( Y=>nx11161, A=>nx11201);
   ix11162 : inv02 port map ( Y=>nx11163, A=>nx11203);
   ix11164 : inv02 port map ( Y=>nx11165, A=>nx11203);
   ix11166 : inv02 port map ( Y=>nx11167, A=>nx11203);
   ix11168 : inv02 port map ( Y=>nx11169, A=>nx11203);
   ix11170 : inv02 port map ( Y=>nx11171, A=>nx11203);
   ix11172 : inv02 port map ( Y=>nx11173, A=>nx11197);
   ix11174 : inv02 port map ( Y=>nx11175, A=>nx11197);
   ix11176 : inv02 port map ( Y=>nx11177, A=>nx11197);
   ix11178 : inv02 port map ( Y=>nx11179, A=>nx11197);
   ix11180 : inv02 port map ( Y=>nx11181, A=>nx11197);
   ix11182 : inv02 port map ( Y=>nx11183, A=>nx11199);
   ix11184 : inv02 port map ( Y=>nx11185, A=>nx11199);
   ix11186 : inv02 port map ( Y=>nx11187, A=>nx11199);
   ix11188 : inv02 port map ( Y=>nx11189, A=>nx11199);
   ix11190 : inv01 port map ( Y=>nx11191, A=>nx11199);
   ix11196 : inv02 port map ( Y=>nx11197, A=>nx9389);
   ix11198 : inv02 port map ( Y=>nx11199, A=>nx9389);
   ix11200 : inv02 port map ( Y=>nx11201, A=>nx9375);
   ix11202 : inv02 port map ( Y=>nx11203, A=>nx9375);
end CNNMulsArch_unfold_1782 ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity RegUnit_8_16 is
   port (
      filterBus : IN std_logic_vector (7 DOWNTO 0) ;
      windowBus : IN std_logic_vector (15 DOWNTO 0) ;
      regPage1NextUnit : IN std_logic_vector (15 DOWNTO 0) ;
      regPage2NextUnit : IN std_logic_vector (15 DOWNTO 0) ;
      clk : IN std_logic ;
      rst : IN std_logic ;
      enableRegPage1 : IN std_logic ;
      enableRegPage2 : IN std_logic ;
      enableRegFilter : IN std_logic ;
      page1ReadBusOrPage2 : IN std_logic ;
      page2ReadBusOrPage1 : IN std_logic ;
      pageTurn : IN std_logic ;
      outRegPage : OUT std_logic_vector (15 DOWNTO 0) ;
      outputRegPage1 : OUT std_logic_vector (15 DOWNTO 0) ;
      outputRegPage2 : OUT std_logic_vector (15 DOWNTO 0) ;
      outFilter : OUT std_logic_vector (7 DOWNTO 0)) ;
end RegUnit_8_16 ;

architecture RegUnitArch_unfold_2792 of RegUnit_8_16 is
   signal outFilter_7_EXMPLR, outFilter_6_EXMPLR, outFilter_5_EXMPLR, 
      outFilter_4_EXMPLR, outFilter_3_EXMPLR, outFilter_2_EXMPLR, 
      outFilter_1_EXMPLR, outFilter_0_EXMPLR, regPage1Map_GND0, 
      outputRegPage1_0_EXMPLR, outputRegPage2_0_EXMPLR, 
      outputRegPage1_1_EXMPLR, outputRegPage2_1_EXMPLR, 
      outputRegPage1_2_EXMPLR, outputRegPage2_2_EXMPLR, 
      outputRegPage1_3_EXMPLR, outputRegPage2_3_EXMPLR, 
      outputRegPage1_4_EXMPLR, outputRegPage2_4_EXMPLR, 
      outputRegPage1_5_EXMPLR, outputRegPage2_5_EXMPLR, 
      outputRegPage1_6_EXMPLR, outputRegPage2_6_EXMPLR, 
      outputRegPage1_7_EXMPLR, outputRegPage2_7_EXMPLR, 
      outputRegPage1_8_EXMPLR, outputRegPage2_8_EXMPLR, 
      outputRegPage1_9_EXMPLR, outputRegPage2_9_EXMPLR, 
      outputRegPage1_10_EXMPLR, outputRegPage2_10_EXMPLR, 
      outputRegPage1_11_EXMPLR, outputRegPage2_11_EXMPLR, 
      outputRegPage1_12_EXMPLR, outputRegPage2_12_EXMPLR, 
      outputRegPage1_13_EXMPLR, outputRegPage2_13_EXMPLR, 
      outputRegPage1_14_EXMPLR, outputRegPage2_14_EXMPLR, 
      outputRegPage1_15_EXMPLR, outputRegPage2_15_EXMPLR, nx133, nx143, 
      nx153, nx163, nx173, nx183, nx193, nx203, nx213, nx223, nx233, nx243, 
      nx253, nx263, nx273, nx283, nx293, nx303, nx313, nx323, nx333, nx343, 
      nx353, nx363, nx373, nx383, nx393, nx403, nx413, nx423, nx433, nx443, 
      nx453, nx463, nx473, nx483, nx493, nx503, nx513, nx523, nx535, nx539, 
      nx544, nx546, nx551, nx553, nx558, nx560, nx565, nx567, nx572, nx574, 
      nx579, nx581, nx586, nx588, nx592, nx595, nx597, nx599, nx602, nx605, 
      nx607, nx609, nx613, nx616, nx618, nx621, nx624, nx626, nx630, nx633, 
      nx635, nx638, nx641, nx643, nx647, nx650, nx652, nx655, nx658, nx660, 
      nx664, nx667, nx669, nx672, nx675, nx677, nx681, nx684, nx686, nx689, 
      nx692, nx694, nx698, nx701, nx703, nx706, nx709, nx711, nx715, nx718, 
      nx720, nx723, nx726, nx728, nx732, nx735, nx737, nx740, nx743, nx745, 
      nx749, nx752, nx754, nx757, nx760, nx762, nx766, nx769, nx771, nx774, 
      nx777, nx779, nx783, nx786, nx788, nx791, nx794, nx796, nx800, nx803, 
      nx805, nx808, nx811, nx813, nx817, nx820, nx822, nx825, nx828, nx830, 
      nx834, nx837, nx839, nx842, nx845, nx847, nx851, nx854, nx856, nx859, 
      nx862, nx864, nx874, nx876, nx878, nx880, nx882, nx884, nx886, nx888, 
      nx890, nx892, nx894, nx896, nx898, nx904, nx906, nx908, nx910: 
   std_logic ;

begin
   outputRegPage1(15) <= regPage1Map_GND0 ;
   outputRegPage1(14) <= regPage1Map_GND0 ;
   outputRegPage1(13) <= regPage1Map_GND0 ;
   outputRegPage1(12) <= regPage1Map_GND0 ;
   outputRegPage1(11) <= regPage1Map_GND0 ;
   outputRegPage1(10) <= regPage1Map_GND0 ;
   outputRegPage1(9) <= regPage1Map_GND0 ;
   outputRegPage1(8) <= regPage1Map_GND0 ;
   outputRegPage1(7) <= regPage1Map_GND0 ;
   outputRegPage1(6) <= regPage1Map_GND0 ;
   outputRegPage1(5) <= regPage1Map_GND0 ;
   outputRegPage1(4) <= regPage1Map_GND0 ;
   outputRegPage1(3) <= regPage1Map_GND0 ;
   outputRegPage1(2) <= regPage1Map_GND0 ;
   outputRegPage1(1) <= regPage1Map_GND0 ;
   outputRegPage1(0) <= regPage1Map_GND0 ;
   outputRegPage2(15) <= regPage1Map_GND0 ;
   outputRegPage2(14) <= regPage1Map_GND0 ;
   outputRegPage2(13) <= regPage1Map_GND0 ;
   outputRegPage2(12) <= regPage1Map_GND0 ;
   outputRegPage2(11) <= regPage1Map_GND0 ;
   outputRegPage2(10) <= regPage1Map_GND0 ;
   outputRegPage2(9) <= regPage1Map_GND0 ;
   outputRegPage2(8) <= regPage1Map_GND0 ;
   outputRegPage2(7) <= regPage1Map_GND0 ;
   outputRegPage2(6) <= regPage1Map_GND0 ;
   outputRegPage2(5) <= regPage1Map_GND0 ;
   outputRegPage2(4) <= regPage1Map_GND0 ;
   outputRegPage2(3) <= regPage1Map_GND0 ;
   outputRegPage2(2) <= regPage1Map_GND0 ;
   outputRegPage2(1) <= regPage1Map_GND0 ;
   outputRegPage2(0) <= regPage1Map_GND0 ;
   outFilter(7) <= outFilter_7_EXMPLR ;
   outFilter(6) <= outFilter_6_EXMPLR ;
   outFilter(5) <= outFilter_5_EXMPLR ;
   outFilter(4) <= outFilter_4_EXMPLR ;
   outFilter(3) <= outFilter_3_EXMPLR ;
   outFilter(2) <= outFilter_2_EXMPLR ;
   outFilter(1) <= outFilter_1_EXMPLR ;
   outFilter(0) <= outFilter_0_EXMPLR ;
   ix54 : fake_gnd port map ( Y=>regPage1Map_GND0);
   regFilterMap_reg_Q_0 : dffr port map ( Q=>outFilter_0_EXMPLR, QB=>OPEN, D
      =>nx453, CLK=>clk, R=>rst);
   ix454 : nand02 port map ( Y=>nx453, A0=>nx535, A1=>nx539);
   ix536 : nand02 port map ( Y=>nx535, A0=>outFilter_0_EXMPLR, A1=>nx908);
   ix540 : nand02 port map ( Y=>nx539, A0=>filterBus(0), A1=>nx904);
   regFilterMap_reg_Q_1 : dffr port map ( Q=>outFilter_1_EXMPLR, QB=>OPEN, D
      =>nx463, CLK=>clk, R=>rst);
   ix464 : nand02 port map ( Y=>nx463, A0=>nx544, A1=>nx546);
   ix545 : nand02 port map ( Y=>nx544, A0=>outFilter_1_EXMPLR, A1=>nx908);
   ix547 : nand02 port map ( Y=>nx546, A0=>filterBus(1), A1=>nx904);
   regFilterMap_reg_Q_2 : dffr port map ( Q=>outFilter_2_EXMPLR, QB=>OPEN, D
      =>nx473, CLK=>clk, R=>rst);
   ix474 : nand02 port map ( Y=>nx473, A0=>nx551, A1=>nx553);
   ix552 : nand02 port map ( Y=>nx551, A0=>outFilter_2_EXMPLR, A1=>nx908);
   ix554 : nand02 port map ( Y=>nx553, A0=>filterBus(2), A1=>nx904);
   regFilterMap_reg_Q_3 : dffr port map ( Q=>outFilter_3_EXMPLR, QB=>OPEN, D
      =>nx483, CLK=>clk, R=>rst);
   ix484 : nand02 port map ( Y=>nx483, A0=>nx558, A1=>nx560);
   ix559 : nand02 port map ( Y=>nx558, A0=>outFilter_3_EXMPLR, A1=>nx908);
   ix561 : nand02 port map ( Y=>nx560, A0=>filterBus(3), A1=>nx904);
   regFilterMap_reg_Q_4 : dffr port map ( Q=>outFilter_4_EXMPLR, QB=>OPEN, D
      =>nx493, CLK=>clk, R=>rst);
   ix494 : nand02 port map ( Y=>nx493, A0=>nx565, A1=>nx567);
   ix566 : nand02 port map ( Y=>nx565, A0=>outFilter_4_EXMPLR, A1=>nx908);
   ix568 : nand02 port map ( Y=>nx567, A0=>filterBus(4), A1=>nx904);
   regFilterMap_reg_Q_5 : dffr port map ( Q=>outFilter_5_EXMPLR, QB=>OPEN, D
      =>nx503, CLK=>clk, R=>rst);
   ix504 : nand02 port map ( Y=>nx503, A0=>nx572, A1=>nx574);
   ix573 : nand02 port map ( Y=>nx572, A0=>outFilter_5_EXMPLR, A1=>nx908);
   ix575 : nand02 port map ( Y=>nx574, A0=>filterBus(5), A1=>nx904);
   regFilterMap_reg_Q_6 : dffr port map ( Q=>outFilter_6_EXMPLR, QB=>OPEN, D
      =>nx513, CLK=>clk, R=>rst);
   ix514 : nand02 port map ( Y=>nx513, A0=>nx579, A1=>nx581);
   ix580 : nand02 port map ( Y=>nx579, A0=>outFilter_6_EXMPLR, A1=>nx908);
   ix582 : nand02 port map ( Y=>nx581, A0=>filterBus(6), A1=>nx904);
   regFilterMap_reg_Q_7 : dffr port map ( Q=>outFilter_7_EXMPLR, QB=>OPEN, D
      =>nx523, CLK=>clk, R=>rst);
   ix524 : nand02 port map ( Y=>nx523, A0=>nx586, A1=>nx588);
   ix587 : nand02 port map ( Y=>nx586, A0=>outFilter_7_EXMPLR, A1=>nx874);
   ix589 : nand02 port map ( Y=>nx588, A0=>filterBus(7), A1=>nx906);
   ix33 : mux21 port map ( Y=>outRegPage(0), A0=>nx592, A1=>nx602, S0=>
      pageTurn);
   ix134 : oai21 port map ( Y=>nx133, A0=>nx595, A1=>nx878, B0=>nx599);
   ix596 : mux21 port map ( Y=>nx595, A0=>windowBus(0), A1=>
      regPage2NextUnit(0), S0=>page1ReadBusOrPage2);
   ix598 : nor02_2x port map ( Y=>nx597, A0=>enableRegPage1, A1=>
      page1ReadBusOrPage2);
   ix600 : nand02 port map ( Y=>nx599, A0=>outputRegPage1_0_EXMPLR, A1=>
      nx878);
   regPage1Map_reg_Q_0 : dffr port map ( Q=>outputRegPage1_0_EXMPLR, QB=>
      nx592, D=>nx133, CLK=>clk, R=>rst);
   ix144 : oai21 port map ( Y=>nx143, A0=>nx605, A1=>nx890, B0=>nx609);
   ix606 : mux21 port map ( Y=>nx605, A0=>windowBus(0), A1=>
      regPage1NextUnit(0), S0=>page2ReadBusOrPage1);
   ix608 : nor02_2x port map ( Y=>nx607, A0=>enableRegPage2, A1=>
      page2ReadBusOrPage1);
   ix610 : nand02 port map ( Y=>nx609, A0=>outputRegPage2_0_EXMPLR, A1=>
      nx890);
   regPage2Map_reg_Q_0 : dffr port map ( Q=>outputRegPage2_0_EXMPLR, QB=>
      nx602, D=>nx143, CLK=>clk, R=>rst);
   ix61 : mux21 port map ( Y=>outRegPage(1), A0=>nx613, A1=>nx621, S0=>
      pageTurn);
   ix154 : oai21 port map ( Y=>nx153, A0=>nx616, A1=>nx878, B0=>nx618);
   ix617 : mux21 port map ( Y=>nx616, A0=>windowBus(1), A1=>
      regPage2NextUnit(1), S0=>page1ReadBusOrPage2);
   ix619 : nand02 port map ( Y=>nx618, A0=>outputRegPage1_1_EXMPLR, A1=>
      nx878);
   regPage1Map_reg_Q_1 : dffr port map ( Q=>outputRegPage1_1_EXMPLR, QB=>
      nx613, D=>nx153, CLK=>clk, R=>rst);
   ix164 : oai21 port map ( Y=>nx163, A0=>nx624, A1=>nx890, B0=>nx626);
   ix625 : mux21 port map ( Y=>nx624, A0=>windowBus(1), A1=>
      regPage1NextUnit(1), S0=>page2ReadBusOrPage1);
   ix627 : nand02 port map ( Y=>nx626, A0=>outputRegPage2_1_EXMPLR, A1=>
      nx890);
   regPage2Map_reg_Q_1 : dffr port map ( Q=>outputRegPage2_1_EXMPLR, QB=>
      nx621, D=>nx163, CLK=>clk, R=>rst);
   ix89 : mux21 port map ( Y=>outRegPage(2), A0=>nx630, A1=>nx638, S0=>
      pageTurn);
   ix174 : oai21 port map ( Y=>nx173, A0=>nx633, A1=>nx878, B0=>nx635);
   ix634 : mux21 port map ( Y=>nx633, A0=>windowBus(2), A1=>
      regPage2NextUnit(2), S0=>page1ReadBusOrPage2);
   ix636 : nand02 port map ( Y=>nx635, A0=>outputRegPage1_2_EXMPLR, A1=>
      nx878);
   regPage1Map_reg_Q_2 : dffr port map ( Q=>outputRegPage1_2_EXMPLR, QB=>
      nx630, D=>nx173, CLK=>clk, R=>rst);
   ix184 : oai21 port map ( Y=>nx183, A0=>nx641, A1=>nx890, B0=>nx643);
   ix642 : mux21 port map ( Y=>nx641, A0=>windowBus(2), A1=>
      regPage1NextUnit(2), S0=>page2ReadBusOrPage1);
   ix644 : nand02 port map ( Y=>nx643, A0=>outputRegPage2_2_EXMPLR, A1=>
      nx890);
   regPage2Map_reg_Q_2 : dffr port map ( Q=>outputRegPage2_2_EXMPLR, QB=>
      nx638, D=>nx183, CLK=>clk, R=>rst);
   ix117 : mux21 port map ( Y=>outRegPage(3), A0=>nx647, A1=>nx655, S0=>
      pageTurn);
   ix194 : oai21 port map ( Y=>nx193, A0=>nx650, A1=>nx878, B0=>nx652);
   ix651 : mux21 port map ( Y=>nx650, A0=>windowBus(3), A1=>
      regPage2NextUnit(3), S0=>page1ReadBusOrPage2);
   ix653 : nand02 port map ( Y=>nx652, A0=>outputRegPage1_3_EXMPLR, A1=>
      nx880);
   regPage1Map_reg_Q_3 : dffr port map ( Q=>outputRegPage1_3_EXMPLR, QB=>
      nx647, D=>nx193, CLK=>clk, R=>rst);
   ix204 : oai21 port map ( Y=>nx203, A0=>nx658, A1=>nx890, B0=>nx660);
   ix659 : mux21 port map ( Y=>nx658, A0=>windowBus(3), A1=>
      regPage1NextUnit(3), S0=>page2ReadBusOrPage1);
   ix661 : nand02 port map ( Y=>nx660, A0=>outputRegPage2_3_EXMPLR, A1=>
      nx892);
   regPage2Map_reg_Q_3 : dffr port map ( Q=>outputRegPage2_3_EXMPLR, QB=>
      nx655, D=>nx203, CLK=>clk, R=>rst);
   ix145 : mux21 port map ( Y=>outRegPage(4), A0=>nx664, A1=>nx672, S0=>
      pageTurn);
   ix214 : oai21 port map ( Y=>nx213, A0=>nx667, A1=>nx880, B0=>nx669);
   ix668 : mux21 port map ( Y=>nx667, A0=>windowBus(4), A1=>
      regPage2NextUnit(4), S0=>page1ReadBusOrPage2);
   ix670 : nand02 port map ( Y=>nx669, A0=>outputRegPage1_4_EXMPLR, A1=>
      nx880);
   regPage1Map_reg_Q_4 : dffr port map ( Q=>outputRegPage1_4_EXMPLR, QB=>
      nx664, D=>nx213, CLK=>clk, R=>rst);
   ix224 : oai21 port map ( Y=>nx223, A0=>nx675, A1=>nx892, B0=>nx677);
   ix676 : mux21 port map ( Y=>nx675, A0=>windowBus(4), A1=>
      regPage1NextUnit(4), S0=>page2ReadBusOrPage1);
   ix678 : nand02 port map ( Y=>nx677, A0=>outputRegPage2_4_EXMPLR, A1=>
      nx892);
   regPage2Map_reg_Q_4 : dffr port map ( Q=>outputRegPage2_4_EXMPLR, QB=>
      nx672, D=>nx223, CLK=>clk, R=>rst);
   ix173 : mux21 port map ( Y=>outRegPage(5), A0=>nx681, A1=>nx689, S0=>
      pageTurn);
   ix234 : oai21 port map ( Y=>nx233, A0=>nx684, A1=>nx880, B0=>nx686);
   ix685 : mux21 port map ( Y=>nx684, A0=>windowBus(5), A1=>
      regPage2NextUnit(5), S0=>page1ReadBusOrPage2);
   ix687 : nand02 port map ( Y=>nx686, A0=>outputRegPage1_5_EXMPLR, A1=>
      nx880);
   regPage1Map_reg_Q_5 : dffr port map ( Q=>outputRegPage1_5_EXMPLR, QB=>
      nx681, D=>nx233, CLK=>clk, R=>rst);
   ix244 : oai21 port map ( Y=>nx243, A0=>nx692, A1=>nx892, B0=>nx694);
   ix693 : mux21 port map ( Y=>nx692, A0=>windowBus(5), A1=>
      regPage1NextUnit(5), S0=>page2ReadBusOrPage1);
   ix695 : nand02 port map ( Y=>nx694, A0=>outputRegPage2_5_EXMPLR, A1=>
      nx892);
   regPage2Map_reg_Q_5 : dffr port map ( Q=>outputRegPage2_5_EXMPLR, QB=>
      nx689, D=>nx243, CLK=>clk, R=>rst);
   ix201 : mux21 port map ( Y=>outRegPage(6), A0=>nx698, A1=>nx706, S0=>
      pageTurn);
   ix254 : oai21 port map ( Y=>nx253, A0=>nx701, A1=>nx880, B0=>nx703);
   ix702 : mux21 port map ( Y=>nx701, A0=>windowBus(6), A1=>
      regPage2NextUnit(6), S0=>page1ReadBusOrPage2);
   ix704 : nand02 port map ( Y=>nx703, A0=>outputRegPage1_6_EXMPLR, A1=>
      nx880);
   regPage1Map_reg_Q_6 : dffr port map ( Q=>outputRegPage1_6_EXMPLR, QB=>
      nx698, D=>nx253, CLK=>clk, R=>rst);
   ix264 : oai21 port map ( Y=>nx263, A0=>nx709, A1=>nx892, B0=>nx711);
   ix710 : mux21 port map ( Y=>nx709, A0=>windowBus(6), A1=>
      regPage1NextUnit(6), S0=>page2ReadBusOrPage1);
   ix712 : nand02 port map ( Y=>nx711, A0=>outputRegPage2_6_EXMPLR, A1=>
      nx892);
   regPage2Map_reg_Q_6 : dffr port map ( Q=>outputRegPage2_6_EXMPLR, QB=>
      nx706, D=>nx263, CLK=>clk, R=>rst);
   ix229 : mux21 port map ( Y=>outRegPage(7), A0=>nx715, A1=>nx723, S0=>
      pageTurn);
   ix274 : oai21 port map ( Y=>nx273, A0=>nx718, A1=>nx882, B0=>nx720);
   ix719 : mux21 port map ( Y=>nx718, A0=>windowBus(7), A1=>
      regPage2NextUnit(7), S0=>page1ReadBusOrPage2);
   ix721 : nand02 port map ( Y=>nx720, A0=>outputRegPage1_7_EXMPLR, A1=>
      nx882);
   regPage1Map_reg_Q_7 : dffr port map ( Q=>outputRegPage1_7_EXMPLR, QB=>
      nx715, D=>nx273, CLK=>clk, R=>rst);
   ix284 : oai21 port map ( Y=>nx283, A0=>nx726, A1=>nx894, B0=>nx728);
   ix727 : mux21 port map ( Y=>nx726, A0=>windowBus(7), A1=>
      regPage1NextUnit(7), S0=>page2ReadBusOrPage1);
   ix729 : nand02 port map ( Y=>nx728, A0=>outputRegPage2_7_EXMPLR, A1=>
      nx894);
   regPage2Map_reg_Q_7 : dffr port map ( Q=>outputRegPage2_7_EXMPLR, QB=>
      nx723, D=>nx283, CLK=>clk, R=>rst);
   ix257 : mux21 port map ( Y=>outRegPage(8), A0=>nx732, A1=>nx740, S0=>
      pageTurn);
   ix294 : oai21 port map ( Y=>nx293, A0=>nx735, A1=>nx882, B0=>nx737);
   ix736 : mux21 port map ( Y=>nx735, A0=>windowBus(8), A1=>
      regPage2NextUnit(8), S0=>page1ReadBusOrPage2);
   ix738 : nand02 port map ( Y=>nx737, A0=>outputRegPage1_8_EXMPLR, A1=>
      nx882);
   regPage1Map_reg_Q_8 : dffr port map ( Q=>outputRegPage1_8_EXMPLR, QB=>
      nx732, D=>nx293, CLK=>clk, R=>rst);
   ix304 : oai21 port map ( Y=>nx303, A0=>nx743, A1=>nx894, B0=>nx745);
   ix744 : mux21 port map ( Y=>nx743, A0=>windowBus(8), A1=>
      regPage1NextUnit(8), S0=>page2ReadBusOrPage1);
   ix746 : nand02 port map ( Y=>nx745, A0=>outputRegPage2_8_EXMPLR, A1=>
      nx894);
   regPage2Map_reg_Q_8 : dffr port map ( Q=>outputRegPage2_8_EXMPLR, QB=>
      nx740, D=>nx303, CLK=>clk, R=>rst);
   ix285 : mux21 port map ( Y=>outRegPage(9), A0=>nx749, A1=>nx757, S0=>
      pageTurn);
   ix314 : oai21 port map ( Y=>nx313, A0=>nx752, A1=>nx882, B0=>nx754);
   ix753 : mux21 port map ( Y=>nx752, A0=>windowBus(9), A1=>
      regPage2NextUnit(9), S0=>page1ReadBusOrPage2);
   ix755 : nand02 port map ( Y=>nx754, A0=>outputRegPage1_9_EXMPLR, A1=>
      nx882);
   regPage1Map_reg_Q_9 : dffr port map ( Q=>outputRegPage1_9_EXMPLR, QB=>
      nx749, D=>nx313, CLK=>clk, R=>rst);
   ix324 : oai21 port map ( Y=>nx323, A0=>nx760, A1=>nx894, B0=>nx762);
   ix761 : mux21 port map ( Y=>nx760, A0=>windowBus(9), A1=>
      regPage1NextUnit(9), S0=>page2ReadBusOrPage1);
   ix763 : nand02 port map ( Y=>nx762, A0=>outputRegPage2_9_EXMPLR, A1=>
      nx894);
   regPage2Map_reg_Q_9 : dffr port map ( Q=>outputRegPage2_9_EXMPLR, QB=>
      nx757, D=>nx323, CLK=>clk, R=>rst);
   ix313 : mux21 port map ( Y=>outRegPage(10), A0=>nx766, A1=>nx774, S0=>
      pageTurn);
   ix334 : oai21 port map ( Y=>nx333, A0=>nx769, A1=>nx882, B0=>nx771);
   ix770 : mux21 port map ( Y=>nx769, A0=>windowBus(10), A1=>
      regPage2NextUnit(10), S0=>page1ReadBusOrPage2);
   ix772 : nand02 port map ( Y=>nx771, A0=>outputRegPage1_10_EXMPLR, A1=>
      nx884);
   regPage1Map_reg_Q_10 : dffr port map ( Q=>outputRegPage1_10_EXMPLR, QB=>
      nx766, D=>nx333, CLK=>clk, R=>rst);
   ix344 : oai21 port map ( Y=>nx343, A0=>nx777, A1=>nx894, B0=>nx779);
   ix778 : mux21 port map ( Y=>nx777, A0=>windowBus(10), A1=>
      regPage1NextUnit(10), S0=>page2ReadBusOrPage1);
   ix780 : nand02 port map ( Y=>nx779, A0=>outputRegPage2_10_EXMPLR, A1=>
      nx896);
   regPage2Map_reg_Q_10 : dffr port map ( Q=>outputRegPage2_10_EXMPLR, QB=>
      nx774, D=>nx343, CLK=>clk, R=>rst);
   ix341 : mux21 port map ( Y=>outRegPage(11), A0=>nx783, A1=>nx791, S0=>
      pageTurn);
   ix354 : oai21 port map ( Y=>nx353, A0=>nx786, A1=>nx884, B0=>nx788);
   ix787 : mux21 port map ( Y=>nx786, A0=>windowBus(11), A1=>
      regPage2NextUnit(11), S0=>page1ReadBusOrPage2);
   ix789 : nand02 port map ( Y=>nx788, A0=>outputRegPage1_11_EXMPLR, A1=>
      nx884);
   regPage1Map_reg_Q_11 : dffr port map ( Q=>outputRegPage1_11_EXMPLR, QB=>
      nx783, D=>nx353, CLK=>clk, R=>rst);
   ix364 : oai21 port map ( Y=>nx363, A0=>nx794, A1=>nx896, B0=>nx796);
   ix795 : mux21 port map ( Y=>nx794, A0=>windowBus(11), A1=>
      regPage1NextUnit(11), S0=>page2ReadBusOrPage1);
   ix797 : nand02 port map ( Y=>nx796, A0=>outputRegPage2_11_EXMPLR, A1=>
      nx896);
   regPage2Map_reg_Q_11 : dffr port map ( Q=>outputRegPage2_11_EXMPLR, QB=>
      nx791, D=>nx363, CLK=>clk, R=>rst);
   ix369 : mux21 port map ( Y=>outRegPage(12), A0=>nx800, A1=>nx808, S0=>
      pageTurn);
   ix374 : oai21 port map ( Y=>nx373, A0=>nx803, A1=>nx884, B0=>nx805);
   ix804 : mux21 port map ( Y=>nx803, A0=>windowBus(12), A1=>
      regPage2NextUnit(12), S0=>page1ReadBusOrPage2);
   ix806 : nand02 port map ( Y=>nx805, A0=>outputRegPage1_12_EXMPLR, A1=>
      nx884);
   regPage1Map_reg_Q_12 : dffr port map ( Q=>outputRegPage1_12_EXMPLR, QB=>
      nx800, D=>nx373, CLK=>clk, R=>rst);
   ix384 : oai21 port map ( Y=>nx383, A0=>nx811, A1=>nx896, B0=>nx813);
   ix812 : mux21 port map ( Y=>nx811, A0=>windowBus(12), A1=>
      regPage1NextUnit(12), S0=>page2ReadBusOrPage1);
   ix814 : nand02 port map ( Y=>nx813, A0=>outputRegPage2_12_EXMPLR, A1=>
      nx896);
   regPage2Map_reg_Q_12 : dffr port map ( Q=>outputRegPage2_12_EXMPLR, QB=>
      nx808, D=>nx383, CLK=>clk, R=>rst);
   ix397 : mux21 port map ( Y=>outRegPage(13), A0=>nx817, A1=>nx825, S0=>
      pageTurn);
   ix394 : oai21 port map ( Y=>nx393, A0=>nx820, A1=>nx884, B0=>nx822);
   ix821 : mux21 port map ( Y=>nx820, A0=>windowBus(13), A1=>
      regPage2NextUnit(13), S0=>page1ReadBusOrPage2);
   ix823 : nand02 port map ( Y=>nx822, A0=>outputRegPage1_13_EXMPLR, A1=>
      nx884);
   regPage1Map_reg_Q_13 : dffr port map ( Q=>outputRegPage1_13_EXMPLR, QB=>
      nx817, D=>nx393, CLK=>clk, R=>rst);
   ix404 : oai21 port map ( Y=>nx403, A0=>nx828, A1=>nx896, B0=>nx830);
   ix829 : mux21 port map ( Y=>nx828, A0=>windowBus(13), A1=>
      regPage1NextUnit(13), S0=>page2ReadBusOrPage1);
   ix831 : nand02 port map ( Y=>nx830, A0=>outputRegPage2_13_EXMPLR, A1=>
      nx896);
   regPage2Map_reg_Q_13 : dffr port map ( Q=>outputRegPage2_13_EXMPLR, QB=>
      nx825, D=>nx403, CLK=>clk, R=>rst);
   ix425 : mux21 port map ( Y=>outRegPage(14), A0=>nx834, A1=>nx842, S0=>
      pageTurn);
   ix414 : oai21 port map ( Y=>nx413, A0=>nx837, A1=>nx886, B0=>nx839);
   ix838 : mux21 port map ( Y=>nx837, A0=>windowBus(14), A1=>
      regPage2NextUnit(14), S0=>page1ReadBusOrPage2);
   ix840 : nand02 port map ( Y=>nx839, A0=>outputRegPage1_14_EXMPLR, A1=>
      nx886);
   regPage1Map_reg_Q_14 : dffr port map ( Q=>outputRegPage1_14_EXMPLR, QB=>
      nx834, D=>nx413, CLK=>clk, R=>rst);
   ix424 : oai21 port map ( Y=>nx423, A0=>nx845, A1=>nx898, B0=>nx847);
   ix846 : mux21 port map ( Y=>nx845, A0=>windowBus(14), A1=>
      regPage1NextUnit(14), S0=>page2ReadBusOrPage1);
   ix848 : nand02 port map ( Y=>nx847, A0=>outputRegPage2_14_EXMPLR, A1=>
      nx898);
   regPage2Map_reg_Q_14 : dffr port map ( Q=>outputRegPage2_14_EXMPLR, QB=>
      nx842, D=>nx423, CLK=>clk, R=>rst);
   ix453 : mux21 port map ( Y=>outRegPage(15), A0=>nx851, A1=>nx859, S0=>
      pageTurn);
   ix434 : oai21 port map ( Y=>nx433, A0=>nx854, A1=>nx886, B0=>nx856);
   ix855 : mux21 port map ( Y=>nx854, A0=>windowBus(15), A1=>
      regPage2NextUnit(15), S0=>page1ReadBusOrPage2);
   ix857 : nand02 port map ( Y=>nx856, A0=>outputRegPage1_15_EXMPLR, A1=>
      nx886);
   regPage1Map_reg_Q_15 : dffr port map ( Q=>outputRegPage1_15_EXMPLR, QB=>
      nx851, D=>nx433, CLK=>clk, R=>rst);
   ix444 : oai21 port map ( Y=>nx443, A0=>nx862, A1=>nx898, B0=>nx864);
   ix863 : mux21 port map ( Y=>nx862, A0=>windowBus(15), A1=>
      regPage1NextUnit(15), S0=>page2ReadBusOrPage1);
   ix865 : nand02 port map ( Y=>nx864, A0=>outputRegPage2_15_EXMPLR, A1=>
      nx898);
   regPage2Map_reg_Q_15 : dffr port map ( Q=>outputRegPage2_15_EXMPLR, QB=>
      nx859, D=>nx443, CLK=>clk, R=>rst);
   ix873 : inv01 port map ( Y=>nx874, A=>nx906);
   ix875 : inv01 port map ( Y=>nx876, A=>nx597);
   ix877 : inv02 port map ( Y=>nx878, A=>nx876);
   ix879 : inv02 port map ( Y=>nx880, A=>nx876);
   ix881 : inv02 port map ( Y=>nx882, A=>nx876);
   ix883 : inv02 port map ( Y=>nx884, A=>nx876);
   ix885 : inv02 port map ( Y=>nx886, A=>nx876);
   ix887 : inv01 port map ( Y=>nx888, A=>nx607);
   ix889 : inv02 port map ( Y=>nx890, A=>nx888);
   ix891 : inv02 port map ( Y=>nx892, A=>nx888);
   ix893 : inv02 port map ( Y=>nx894, A=>nx888);
   ix895 : inv02 port map ( Y=>nx896, A=>nx888);
   ix897 : inv02 port map ( Y=>nx898, A=>nx888);
   ix903 : inv02 port map ( Y=>nx904, A=>nx910);
   ix905 : inv02 port map ( Y=>nx906, A=>nx910);
   ix907 : inv02 port map ( Y=>nx908, A=>enableRegFilter);
   ix909 : inv02 port map ( Y=>nx910, A=>enableRegFilter);
end RegUnitArch_unfold_2792 ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity RegUnit_8_16_unfolded2 is
   port (
      filterBus : IN std_logic_vector (7 DOWNTO 0) ;
      windowBus : IN std_logic_vector (15 DOWNTO 0) ;
      regPage1NextUnit : IN std_logic_vector (15 DOWNTO 0) ;
      regPage2NextUnit : IN std_logic_vector (15 DOWNTO 0) ;
      clk : IN std_logic ;
      rst : IN std_logic ;
      enableRegPage1 : IN std_logic ;
      enableRegPage2 : IN std_logic ;
      enableRegFilter : IN std_logic ;
      page1ReadBusOrPage2 : IN std_logic ;
      page2ReadBusOrPage1 : IN std_logic ;
      pageTurn : IN std_logic ;
      outRegPage : OUT std_logic_vector (15 DOWNTO 0) ;
      outputRegPage1 : OUT std_logic_vector (15 DOWNTO 0) ;
      outputRegPage2 : OUT std_logic_vector (15 DOWNTO 0) ;
      outFilter : OUT std_logic_vector (7 DOWNTO 0)) ;
end RegUnit_8_16_unfolded2 ;

architecture RegUnitArch_xmplrcopy of RegUnit_8_16_unfolded2 is
   signal outputRegPage1_15_EXMPLR, outputRegPage1_14_EXMPLR, 
      outputRegPage1_13_EXMPLR, outputRegPage1_12_EXMPLR, 
      outputRegPage1_11_EXMPLR, outputRegPage1_10_EXMPLR, 
      outputRegPage1_9_EXMPLR, outputRegPage1_8_EXMPLR, 
      outputRegPage1_7_EXMPLR, outputRegPage1_6_EXMPLR, 
      outputRegPage1_5_EXMPLR, outputRegPage1_4_EXMPLR, 
      outputRegPage1_3_EXMPLR, outputRegPage1_2_EXMPLR, 
      outputRegPage1_1_EXMPLR, outputRegPage1_0_EXMPLR, 
      outputRegPage2_15_EXMPLR, outputRegPage2_14_EXMPLR, 
      outputRegPage2_13_EXMPLR, outputRegPage2_12_EXMPLR, 
      outputRegPage2_11_EXMPLR, outputRegPage2_10_EXMPLR, 
      outputRegPage2_9_EXMPLR, outputRegPage2_8_EXMPLR, 
      outputRegPage2_7_EXMPLR, outputRegPage2_6_EXMPLR, 
      outputRegPage2_5_EXMPLR, outputRegPage2_4_EXMPLR, 
      outputRegPage2_3_EXMPLR, outputRegPage2_2_EXMPLR, 
      outputRegPage2_1_EXMPLR, outputRegPage2_0_EXMPLR, outFilter_7_EXMPLR, 
      outFilter_6_EXMPLR, outFilter_5_EXMPLR, outFilter_4_EXMPLR, 
      outFilter_3_EXMPLR, outFilter_2_EXMPLR, outFilter_1_EXMPLR, 
      outFilter_0_EXMPLR, nx345, nx355, nx365, nx375, nx385, nx395, nx405, 
      nx415, nx425, nx435, nx445, nx455, nx465, nx475, nx485, nx495, nx505, 
      nx515, nx525, nx535, nx545, nx555, nx565, nx575, nx585, nx595, nx605, 
      nx615, nx625, nx635, nx645, nx655, nx665, nx675, nx685, nx695, nx705, 
      nx715, nx725, nx735, nx747, nx751, nx756, nx758, nx763, nx765, nx770, 
      nx772, nx777, nx779, nx784, nx786, nx791, nx793, nx798, nx800, nx805, 
      nx807, nx809, nx811, nx814, nx816, nx818, nx821, nx823, nx825, nx828, 
      nx830, nx832, nx835, nx837, nx839, nx842, nx844, nx846, nx849, nx851, 
      nx853, nx856, nx858, nx860, nx863, nx865, nx867, nx870, nx872, nx874, 
      nx877, nx879, nx881, nx884, nx886, nx888, nx891, nx893, nx895, nx898, 
      nx900, nx902, nx905, nx907, nx909, nx912, nx914, nx916, nx919, nx921, 
      nx923, nx925, nx928, nx930, nx932, nx935, nx937, nx939, nx942, nx944, 
      nx946, nx949, nx951, nx953, nx956, nx958, nx960, nx963, nx965, nx967, 
      nx970, nx972, nx974, nx977, nx979, nx981, nx984, nx986, nx988, nx991, 
      nx993, nx995, nx998, nx1000, nx1002, nx1005, nx1007, nx1009, nx1012, 
      nx1014, nx1016, nx1019, nx1021, nx1023, nx1026, nx1028, nx1030, nx1054, 
      nx1056, nx1058, nx1060, nx1062, nx1064, nx1066, nx1068, nx1070, nx1072, 
      nx1074, nx1076, nx1078, nx1084, nx1086, nx1088, nx1090: std_logic ;

begin
   outputRegPage1(15) <= outputRegPage1_15_EXMPLR ;
   outputRegPage1(14) <= outputRegPage1_14_EXMPLR ;
   outputRegPage1(13) <= outputRegPage1_13_EXMPLR ;
   outputRegPage1(12) <= outputRegPage1_12_EXMPLR ;
   outputRegPage1(11) <= outputRegPage1_11_EXMPLR ;
   outputRegPage1(10) <= outputRegPage1_10_EXMPLR ;
   outputRegPage1(9) <= outputRegPage1_9_EXMPLR ;
   outputRegPage1(8) <= outputRegPage1_8_EXMPLR ;
   outputRegPage1(7) <= outputRegPage1_7_EXMPLR ;
   outputRegPage1(6) <= outputRegPage1_6_EXMPLR ;
   outputRegPage1(5) <= outputRegPage1_5_EXMPLR ;
   outputRegPage1(4) <= outputRegPage1_4_EXMPLR ;
   outputRegPage1(3) <= outputRegPage1_3_EXMPLR ;
   outputRegPage1(2) <= outputRegPage1_2_EXMPLR ;
   outputRegPage1(1) <= outputRegPage1_1_EXMPLR ;
   outputRegPage1(0) <= outputRegPage1_0_EXMPLR ;
   outputRegPage2(15) <= outputRegPage2_15_EXMPLR ;
   outputRegPage2(14) <= outputRegPage2_14_EXMPLR ;
   outputRegPage2(13) <= outputRegPage2_13_EXMPLR ;
   outputRegPage2(12) <= outputRegPage2_12_EXMPLR ;
   outputRegPage2(11) <= outputRegPage2_11_EXMPLR ;
   outputRegPage2(10) <= outputRegPage2_10_EXMPLR ;
   outputRegPage2(9) <= outputRegPage2_9_EXMPLR ;
   outputRegPage2(8) <= outputRegPage2_8_EXMPLR ;
   outputRegPage2(7) <= outputRegPage2_7_EXMPLR ;
   outputRegPage2(6) <= outputRegPage2_6_EXMPLR ;
   outputRegPage2(5) <= outputRegPage2_5_EXMPLR ;
   outputRegPage2(4) <= outputRegPage2_4_EXMPLR ;
   outputRegPage2(3) <= outputRegPage2_3_EXMPLR ;
   outputRegPage2(2) <= outputRegPage2_2_EXMPLR ;
   outputRegPage2(1) <= outputRegPage2_1_EXMPLR ;
   outputRegPage2(0) <= outputRegPage2_0_EXMPLR ;
   outFilter(7) <= outFilter_7_EXMPLR ;
   outFilter(6) <= outFilter_6_EXMPLR ;
   outFilter(5) <= outFilter_5_EXMPLR ;
   outFilter(4) <= outFilter_4_EXMPLR ;
   outFilter(3) <= outFilter_3_EXMPLR ;
   outFilter(2) <= outFilter_2_EXMPLR ;
   outFilter(1) <= outFilter_1_EXMPLR ;
   outFilter(0) <= outFilter_0_EXMPLR ;
   regFilterMap_reg_Q_0 : dffr port map ( Q=>outFilter_0_EXMPLR, QB=>OPEN, D
      =>nx665, CLK=>clk, R=>rst);
   ix666 : nand02 port map ( Y=>nx665, A0=>nx747, A1=>nx751);
   ix748 : nand02 port map ( Y=>nx747, A0=>outFilter_0_EXMPLR, A1=>nx1088);
   ix752 : nand02 port map ( Y=>nx751, A0=>filterBus(0), A1=>nx1084);
   regFilterMap_reg_Q_1 : dffr port map ( Q=>outFilter_1_EXMPLR, QB=>OPEN, D
      =>nx675, CLK=>clk, R=>rst);
   ix676 : nand02 port map ( Y=>nx675, A0=>nx756, A1=>nx758);
   ix757 : nand02 port map ( Y=>nx756, A0=>outFilter_1_EXMPLR, A1=>nx1088);
   ix759 : nand02 port map ( Y=>nx758, A0=>filterBus(1), A1=>nx1084);
   regFilterMap_reg_Q_2 : dffr port map ( Q=>outFilter_2_EXMPLR, QB=>OPEN, D
      =>nx685, CLK=>clk, R=>rst);
   ix686 : nand02 port map ( Y=>nx685, A0=>nx763, A1=>nx765);
   ix764 : nand02 port map ( Y=>nx763, A0=>outFilter_2_EXMPLR, A1=>nx1088);
   ix766 : nand02 port map ( Y=>nx765, A0=>filterBus(2), A1=>nx1084);
   regFilterMap_reg_Q_3 : dffr port map ( Q=>outFilter_3_EXMPLR, QB=>OPEN, D
      =>nx695, CLK=>clk, R=>rst);
   ix696 : nand02 port map ( Y=>nx695, A0=>nx770, A1=>nx772);
   ix771 : nand02 port map ( Y=>nx770, A0=>outFilter_3_EXMPLR, A1=>nx1088);
   ix773 : nand02 port map ( Y=>nx772, A0=>filterBus(3), A1=>nx1084);
   regFilterMap_reg_Q_4 : dffr port map ( Q=>outFilter_4_EXMPLR, QB=>OPEN, D
      =>nx705, CLK=>clk, R=>rst);
   ix706 : nand02 port map ( Y=>nx705, A0=>nx777, A1=>nx779);
   ix778 : nand02 port map ( Y=>nx777, A0=>outFilter_4_EXMPLR, A1=>nx1088);
   ix780 : nand02 port map ( Y=>nx779, A0=>filterBus(4), A1=>nx1084);
   regFilterMap_reg_Q_5 : dffr port map ( Q=>outFilter_5_EXMPLR, QB=>OPEN, D
      =>nx715, CLK=>clk, R=>rst);
   ix716 : nand02 port map ( Y=>nx715, A0=>nx784, A1=>nx786);
   ix785 : nand02 port map ( Y=>nx784, A0=>outFilter_5_EXMPLR, A1=>nx1088);
   ix787 : nand02 port map ( Y=>nx786, A0=>filterBus(5), A1=>nx1084);
   regFilterMap_reg_Q_6 : dffr port map ( Q=>outFilter_6_EXMPLR, QB=>OPEN, D
      =>nx725, CLK=>clk, R=>rst);
   ix726 : nand02 port map ( Y=>nx725, A0=>nx791, A1=>nx793);
   ix792 : nand02 port map ( Y=>nx791, A0=>outFilter_6_EXMPLR, A1=>nx1088);
   ix794 : nand02 port map ( Y=>nx793, A0=>filterBus(6), A1=>nx1084);
   regFilterMap_reg_Q_7 : dffr port map ( Q=>outFilter_7_EXMPLR, QB=>OPEN, D
      =>nx735, CLK=>clk, R=>rst);
   ix736 : nand02 port map ( Y=>nx735, A0=>nx798, A1=>nx800);
   ix799 : nand02 port map ( Y=>nx798, A0=>outFilter_7_EXMPLR, A1=>nx1054);
   ix801 : nand02 port map ( Y=>nx800, A0=>filterBus(7), A1=>nx1086);
   regPage2Map_reg_Q_0 : dffr port map ( Q=>outputRegPage2_0_EXMPLR, QB=>
      nx811, D=>nx355, CLK=>clk, R=>rst);
   ix356 : oai21 port map ( Y=>nx355, A0=>nx805, A1=>nx1058, B0=>nx809);
   ix806 : mux21 port map ( Y=>nx805, A0=>windowBus(0), A1=>
      regPage1NextUnit(0), S0=>page2ReadBusOrPage1);
   ix808 : nor02_2x port map ( Y=>nx807, A0=>enableRegPage2, A1=>
      page2ReadBusOrPage1);
   ix810 : nand02 port map ( Y=>nx809, A0=>outputRegPage2_0_EXMPLR, A1=>
      nx1058);
   regPage2Map_reg_Q_1 : dffr port map ( Q=>outputRegPage2_1_EXMPLR, QB=>
      nx818, D=>nx375, CLK=>clk, R=>rst);
   ix376 : oai21 port map ( Y=>nx375, A0=>nx814, A1=>nx1058, B0=>nx816);
   ix815 : mux21 port map ( Y=>nx814, A0=>windowBus(1), A1=>
      regPage1NextUnit(1), S0=>page2ReadBusOrPage1);
   ix817 : nand02 port map ( Y=>nx816, A0=>outputRegPage2_1_EXMPLR, A1=>
      nx1058);
   regPage2Map_reg_Q_2 : dffr port map ( Q=>outputRegPage2_2_EXMPLR, QB=>
      nx825, D=>nx395, CLK=>clk, R=>rst);
   ix396 : oai21 port map ( Y=>nx395, A0=>nx821, A1=>nx1058, B0=>nx823);
   ix822 : mux21 port map ( Y=>nx821, A0=>windowBus(2), A1=>
      regPage1NextUnit(2), S0=>page2ReadBusOrPage1);
   ix824 : nand02 port map ( Y=>nx823, A0=>outputRegPage2_2_EXMPLR, A1=>
      nx1058);
   regPage2Map_reg_Q_3 : dffr port map ( Q=>outputRegPage2_3_EXMPLR, QB=>
      nx832, D=>nx415, CLK=>clk, R=>rst);
   ix416 : oai21 port map ( Y=>nx415, A0=>nx828, A1=>nx1058, B0=>nx830);
   ix829 : mux21 port map ( Y=>nx828, A0=>windowBus(3), A1=>
      regPage1NextUnit(3), S0=>page2ReadBusOrPage1);
   ix831 : nand02 port map ( Y=>nx830, A0=>outputRegPage2_3_EXMPLR, A1=>
      nx1060);
   regPage2Map_reg_Q_4 : dffr port map ( Q=>outputRegPage2_4_EXMPLR, QB=>
      nx839, D=>nx435, CLK=>clk, R=>rst);
   ix436 : oai21 port map ( Y=>nx435, A0=>nx835, A1=>nx1060, B0=>nx837);
   ix836 : mux21 port map ( Y=>nx835, A0=>windowBus(4), A1=>
      regPage1NextUnit(4), S0=>page2ReadBusOrPage1);
   ix838 : nand02 port map ( Y=>nx837, A0=>outputRegPage2_4_EXMPLR, A1=>
      nx1060);
   regPage2Map_reg_Q_5 : dffr port map ( Q=>outputRegPage2_5_EXMPLR, QB=>
      nx846, D=>nx455, CLK=>clk, R=>rst);
   ix456 : oai21 port map ( Y=>nx455, A0=>nx842, A1=>nx1060, B0=>nx844);
   ix843 : mux21 port map ( Y=>nx842, A0=>windowBus(5), A1=>
      regPage1NextUnit(5), S0=>page2ReadBusOrPage1);
   ix845 : nand02 port map ( Y=>nx844, A0=>outputRegPage2_5_EXMPLR, A1=>
      nx1060);
   regPage2Map_reg_Q_6 : dffr port map ( Q=>outputRegPage2_6_EXMPLR, QB=>
      nx853, D=>nx475, CLK=>clk, R=>rst);
   ix476 : oai21 port map ( Y=>nx475, A0=>nx849, A1=>nx1060, B0=>nx851);
   ix850 : mux21 port map ( Y=>nx849, A0=>windowBus(6), A1=>
      regPage1NextUnit(6), S0=>page2ReadBusOrPage1);
   ix852 : nand02 port map ( Y=>nx851, A0=>outputRegPage2_6_EXMPLR, A1=>
      nx1060);
   regPage2Map_reg_Q_7 : dffr port map ( Q=>outputRegPage2_7_EXMPLR, QB=>
      nx860, D=>nx495, CLK=>clk, R=>rst);
   ix496 : oai21 port map ( Y=>nx495, A0=>nx856, A1=>nx1062, B0=>nx858);
   ix857 : mux21 port map ( Y=>nx856, A0=>windowBus(7), A1=>
      regPage1NextUnit(7), S0=>page2ReadBusOrPage1);
   ix859 : nand02 port map ( Y=>nx858, A0=>outputRegPage2_7_EXMPLR, A1=>
      nx1062);
   regPage2Map_reg_Q_8 : dffr port map ( Q=>outputRegPage2_8_EXMPLR, QB=>
      nx867, D=>nx515, CLK=>clk, R=>rst);
   ix516 : oai21 port map ( Y=>nx515, A0=>nx863, A1=>nx1062, B0=>nx865);
   ix864 : mux21 port map ( Y=>nx863, A0=>windowBus(8), A1=>
      regPage1NextUnit(8), S0=>page2ReadBusOrPage1);
   ix866 : nand02 port map ( Y=>nx865, A0=>outputRegPage2_8_EXMPLR, A1=>
      nx1062);
   regPage2Map_reg_Q_9 : dffr port map ( Q=>outputRegPage2_9_EXMPLR, QB=>
      nx874, D=>nx535, CLK=>clk, R=>rst);
   ix536 : oai21 port map ( Y=>nx535, A0=>nx870, A1=>nx1062, B0=>nx872);
   ix871 : mux21 port map ( Y=>nx870, A0=>windowBus(9), A1=>
      regPage1NextUnit(9), S0=>page2ReadBusOrPage1);
   ix873 : nand02 port map ( Y=>nx872, A0=>outputRegPage2_9_EXMPLR, A1=>
      nx1062);
   regPage2Map_reg_Q_10 : dffr port map ( Q=>outputRegPage2_10_EXMPLR, QB=>
      nx881, D=>nx555, CLK=>clk, R=>rst);
   ix556 : oai21 port map ( Y=>nx555, A0=>nx877, A1=>nx1062, B0=>nx879);
   ix878 : mux21 port map ( Y=>nx877, A0=>windowBus(10), A1=>
      regPage1NextUnit(10), S0=>page2ReadBusOrPage1);
   ix880 : nand02 port map ( Y=>nx879, A0=>outputRegPage2_10_EXMPLR, A1=>
      nx1064);
   regPage2Map_reg_Q_11 : dffr port map ( Q=>outputRegPage2_11_EXMPLR, QB=>
      nx888, D=>nx575, CLK=>clk, R=>rst);
   ix576 : oai21 port map ( Y=>nx575, A0=>nx884, A1=>nx1064, B0=>nx886);
   ix885 : mux21 port map ( Y=>nx884, A0=>windowBus(11), A1=>
      regPage1NextUnit(11), S0=>page2ReadBusOrPage1);
   ix887 : nand02 port map ( Y=>nx886, A0=>outputRegPage2_11_EXMPLR, A1=>
      nx1064);
   regPage2Map_reg_Q_12 : dffr port map ( Q=>outputRegPage2_12_EXMPLR, QB=>
      nx895, D=>nx595, CLK=>clk, R=>rst);
   ix596 : oai21 port map ( Y=>nx595, A0=>nx891, A1=>nx1064, B0=>nx893);
   ix892 : mux21 port map ( Y=>nx891, A0=>windowBus(12), A1=>
      regPage1NextUnit(12), S0=>page2ReadBusOrPage1);
   ix894 : nand02 port map ( Y=>nx893, A0=>outputRegPage2_12_EXMPLR, A1=>
      nx1064);
   regPage2Map_reg_Q_13 : dffr port map ( Q=>outputRegPage2_13_EXMPLR, QB=>
      nx902, D=>nx615, CLK=>clk, R=>rst);
   ix616 : oai21 port map ( Y=>nx615, A0=>nx898, A1=>nx1064, B0=>nx900);
   ix899 : mux21 port map ( Y=>nx898, A0=>windowBus(13), A1=>
      regPage1NextUnit(13), S0=>page2ReadBusOrPage1);
   ix901 : nand02 port map ( Y=>nx900, A0=>outputRegPage2_13_EXMPLR, A1=>
      nx1064);
   regPage2Map_reg_Q_14 : dffr port map ( Q=>outputRegPage2_14_EXMPLR, QB=>
      nx909, D=>nx635, CLK=>clk, R=>rst);
   ix636 : oai21 port map ( Y=>nx635, A0=>nx905, A1=>nx1066, B0=>nx907);
   ix906 : mux21 port map ( Y=>nx905, A0=>windowBus(14), A1=>
      regPage1NextUnit(14), S0=>page2ReadBusOrPage1);
   ix908 : nand02 port map ( Y=>nx907, A0=>outputRegPage2_14_EXMPLR, A1=>
      nx1066);
   regPage2Map_reg_Q_15 : dffr port map ( Q=>outputRegPage2_15_EXMPLR, QB=>
      nx916, D=>nx655, CLK=>clk, R=>rst);
   ix656 : oai21 port map ( Y=>nx655, A0=>nx912, A1=>nx1066, B0=>nx914);
   ix913 : mux21 port map ( Y=>nx912, A0=>windowBus(15), A1=>
      regPage1NextUnit(15), S0=>page2ReadBusOrPage1);
   ix915 : nand02 port map ( Y=>nx914, A0=>outputRegPage2_15_EXMPLR, A1=>
      nx1066);
   regPage1Map_reg_Q_0 : dffr port map ( Q=>outputRegPage1_0_EXMPLR, QB=>
      nx925, D=>nx345, CLK=>clk, R=>rst);
   ix346 : oai21 port map ( Y=>nx345, A0=>nx919, A1=>nx1070, B0=>nx923);
   ix920 : mux21 port map ( Y=>nx919, A0=>windowBus(0), A1=>
      regPage2NextUnit(0), S0=>page1ReadBusOrPage2);
   ix922 : nor02_2x port map ( Y=>nx921, A0=>enableRegPage1, A1=>
      page1ReadBusOrPage2);
   ix924 : nand02 port map ( Y=>nx923, A0=>outputRegPage1_0_EXMPLR, A1=>
      nx1070);
   regPage1Map_reg_Q_1 : dffr port map ( Q=>outputRegPage1_1_EXMPLR, QB=>
      nx932, D=>nx365, CLK=>clk, R=>rst);
   ix366 : oai21 port map ( Y=>nx365, A0=>nx928, A1=>nx1070, B0=>nx930);
   ix929 : mux21 port map ( Y=>nx928, A0=>windowBus(1), A1=>
      regPage2NextUnit(1), S0=>page1ReadBusOrPage2);
   ix931 : nand02 port map ( Y=>nx930, A0=>outputRegPage1_1_EXMPLR, A1=>
      nx1070);
   regPage1Map_reg_Q_2 : dffr port map ( Q=>outputRegPage1_2_EXMPLR, QB=>
      nx939, D=>nx385, CLK=>clk, R=>rst);
   ix386 : oai21 port map ( Y=>nx385, A0=>nx935, A1=>nx1070, B0=>nx937);
   ix936 : mux21 port map ( Y=>nx935, A0=>windowBus(2), A1=>
      regPage2NextUnit(2), S0=>page1ReadBusOrPage2);
   ix938 : nand02 port map ( Y=>nx937, A0=>outputRegPage1_2_EXMPLR, A1=>
      nx1070);
   regPage1Map_reg_Q_3 : dffr port map ( Q=>outputRegPage1_3_EXMPLR, QB=>
      nx946, D=>nx405, CLK=>clk, R=>rst);
   ix406 : oai21 port map ( Y=>nx405, A0=>nx942, A1=>nx1070, B0=>nx944);
   ix943 : mux21 port map ( Y=>nx942, A0=>windowBus(3), A1=>
      regPage2NextUnit(3), S0=>page1ReadBusOrPage2);
   ix945 : nand02 port map ( Y=>nx944, A0=>outputRegPage1_3_EXMPLR, A1=>
      nx1072);
   regPage1Map_reg_Q_4 : dffr port map ( Q=>outputRegPage1_4_EXMPLR, QB=>
      nx953, D=>nx425, CLK=>clk, R=>rst);
   ix426 : oai21 port map ( Y=>nx425, A0=>nx949, A1=>nx1072, B0=>nx951);
   ix950 : mux21 port map ( Y=>nx949, A0=>windowBus(4), A1=>
      regPage2NextUnit(4), S0=>page1ReadBusOrPage2);
   ix952 : nand02 port map ( Y=>nx951, A0=>outputRegPage1_4_EXMPLR, A1=>
      nx1072);
   regPage1Map_reg_Q_5 : dffr port map ( Q=>outputRegPage1_5_EXMPLR, QB=>
      nx960, D=>nx445, CLK=>clk, R=>rst);
   ix446 : oai21 port map ( Y=>nx445, A0=>nx956, A1=>nx1072, B0=>nx958);
   ix957 : mux21 port map ( Y=>nx956, A0=>windowBus(5), A1=>
      regPage2NextUnit(5), S0=>page1ReadBusOrPage2);
   ix959 : nand02 port map ( Y=>nx958, A0=>outputRegPage1_5_EXMPLR, A1=>
      nx1072);
   regPage1Map_reg_Q_6 : dffr port map ( Q=>outputRegPage1_6_EXMPLR, QB=>
      nx967, D=>nx465, CLK=>clk, R=>rst);
   ix466 : oai21 port map ( Y=>nx465, A0=>nx963, A1=>nx1072, B0=>nx965);
   ix964 : mux21 port map ( Y=>nx963, A0=>windowBus(6), A1=>
      regPage2NextUnit(6), S0=>page1ReadBusOrPage2);
   ix966 : nand02 port map ( Y=>nx965, A0=>outputRegPage1_6_EXMPLR, A1=>
      nx1072);
   regPage1Map_reg_Q_7 : dffr port map ( Q=>outputRegPage1_7_EXMPLR, QB=>
      nx974, D=>nx485, CLK=>clk, R=>rst);
   ix486 : oai21 port map ( Y=>nx485, A0=>nx970, A1=>nx1074, B0=>nx972);
   ix971 : mux21 port map ( Y=>nx970, A0=>windowBus(7), A1=>
      regPage2NextUnit(7), S0=>page1ReadBusOrPage2);
   ix973 : nand02 port map ( Y=>nx972, A0=>outputRegPage1_7_EXMPLR, A1=>
      nx1074);
   regPage1Map_reg_Q_8 : dffr port map ( Q=>outputRegPage1_8_EXMPLR, QB=>
      nx981, D=>nx505, CLK=>clk, R=>rst);
   ix506 : oai21 port map ( Y=>nx505, A0=>nx977, A1=>nx1074, B0=>nx979);
   ix978 : mux21 port map ( Y=>nx977, A0=>windowBus(8), A1=>
      regPage2NextUnit(8), S0=>page1ReadBusOrPage2);
   ix980 : nand02 port map ( Y=>nx979, A0=>outputRegPage1_8_EXMPLR, A1=>
      nx1074);
   regPage1Map_reg_Q_9 : dffr port map ( Q=>outputRegPage1_9_EXMPLR, QB=>
      nx988, D=>nx525, CLK=>clk, R=>rst);
   ix526 : oai21 port map ( Y=>nx525, A0=>nx984, A1=>nx1074, B0=>nx986);
   ix985 : mux21 port map ( Y=>nx984, A0=>windowBus(9), A1=>
      regPage2NextUnit(9), S0=>page1ReadBusOrPage2);
   ix987 : nand02 port map ( Y=>nx986, A0=>outputRegPage1_9_EXMPLR, A1=>
      nx1074);
   regPage1Map_reg_Q_10 : dffr port map ( Q=>outputRegPage1_10_EXMPLR, QB=>
      nx995, D=>nx545, CLK=>clk, R=>rst);
   ix546 : oai21 port map ( Y=>nx545, A0=>nx991, A1=>nx1074, B0=>nx993);
   ix992 : mux21 port map ( Y=>nx991, A0=>windowBus(10), A1=>
      regPage2NextUnit(10), S0=>page1ReadBusOrPage2);
   ix994 : nand02 port map ( Y=>nx993, A0=>outputRegPage1_10_EXMPLR, A1=>
      nx1076);
   regPage1Map_reg_Q_11 : dffr port map ( Q=>outputRegPage1_11_EXMPLR, QB=>
      nx1002, D=>nx565, CLK=>clk, R=>rst);
   ix566 : oai21 port map ( Y=>nx565, A0=>nx998, A1=>nx1076, B0=>nx1000);
   ix999 : mux21 port map ( Y=>nx998, A0=>windowBus(11), A1=>
      regPage2NextUnit(11), S0=>page1ReadBusOrPage2);
   ix1001 : nand02 port map ( Y=>nx1000, A0=>outputRegPage1_11_EXMPLR, A1=>
      nx1076);
   regPage1Map_reg_Q_12 : dffr port map ( Q=>outputRegPage1_12_EXMPLR, QB=>
      nx1009, D=>nx585, CLK=>clk, R=>rst);
   ix586 : oai21 port map ( Y=>nx585, A0=>nx1005, A1=>nx1076, B0=>nx1007);
   ix1006 : mux21 port map ( Y=>nx1005, A0=>windowBus(12), A1=>
      regPage2NextUnit(12), S0=>page1ReadBusOrPage2);
   ix1008 : nand02 port map ( Y=>nx1007, A0=>outputRegPage1_12_EXMPLR, A1=>
      nx1076);
   regPage1Map_reg_Q_13 : dffr port map ( Q=>outputRegPage1_13_EXMPLR, QB=>
      nx1016, D=>nx605, CLK=>clk, R=>rst);
   ix606 : oai21 port map ( Y=>nx605, A0=>nx1012, A1=>nx1076, B0=>nx1014);
   ix1013 : mux21 port map ( Y=>nx1012, A0=>windowBus(13), A1=>
      regPage2NextUnit(13), S0=>page1ReadBusOrPage2);
   ix1015 : nand02 port map ( Y=>nx1014, A0=>outputRegPage1_13_EXMPLR, A1=>
      nx1076);
   regPage1Map_reg_Q_14 : dffr port map ( Q=>outputRegPage1_14_EXMPLR, QB=>
      nx1023, D=>nx625, CLK=>clk, R=>rst);
   ix626 : oai21 port map ( Y=>nx625, A0=>nx1019, A1=>nx1078, B0=>nx1021);
   ix1020 : mux21 port map ( Y=>nx1019, A0=>windowBus(14), A1=>
      regPage2NextUnit(14), S0=>page1ReadBusOrPage2);
   ix1022 : nand02 port map ( Y=>nx1021, A0=>outputRegPage1_14_EXMPLR, A1=>
      nx1078);
   regPage1Map_reg_Q_15 : dffr port map ( Q=>outputRegPage1_15_EXMPLR, QB=>
      nx1030, D=>nx645, CLK=>clk, R=>rst);
   ix646 : oai21 port map ( Y=>nx645, A0=>nx1026, A1=>nx1078, B0=>nx1028);
   ix1027 : mux21 port map ( Y=>nx1026, A0=>windowBus(15), A1=>
      regPage2NextUnit(15), S0=>page1ReadBusOrPage2);
   ix1029 : nand02 port map ( Y=>nx1028, A0=>outputRegPage1_15_EXMPLR, A1=>
      nx1078);
   ix33 : mux21 port map ( Y=>outRegPage(0), A0=>nx925, A1=>nx811, S0=>
      pageTurn);
   ix61 : mux21 port map ( Y=>outRegPage(1), A0=>nx932, A1=>nx818, S0=>
      pageTurn);
   ix89 : mux21 port map ( Y=>outRegPage(2), A0=>nx939, A1=>nx825, S0=>
      pageTurn);
   ix117 : mux21 port map ( Y=>outRegPage(3), A0=>nx946, A1=>nx832, S0=>
      pageTurn);
   ix145 : mux21 port map ( Y=>outRegPage(4), A0=>nx953, A1=>nx839, S0=>
      pageTurn);
   ix173 : mux21 port map ( Y=>outRegPage(5), A0=>nx960, A1=>nx846, S0=>
      pageTurn);
   ix201 : mux21 port map ( Y=>outRegPage(6), A0=>nx967, A1=>nx853, S0=>
      pageTurn);
   ix229 : mux21 port map ( Y=>outRegPage(7), A0=>nx974, A1=>nx860, S0=>
      pageTurn);
   ix257 : mux21 port map ( Y=>outRegPage(8), A0=>nx981, A1=>nx867, S0=>
      pageTurn);
   ix285 : mux21 port map ( Y=>outRegPage(9), A0=>nx988, A1=>nx874, S0=>
      pageTurn);
   ix313 : mux21 port map ( Y=>outRegPage(10), A0=>nx995, A1=>nx881, S0=>
      pageTurn);
   ix341 : mux21 port map ( Y=>outRegPage(11), A0=>nx1002, A1=>nx888, S0=>
      pageTurn);
   ix369 : mux21 port map ( Y=>outRegPage(12), A0=>nx1009, A1=>nx895, S0=>
      pageTurn);
   ix397 : mux21 port map ( Y=>outRegPage(13), A0=>nx1016, A1=>nx902, S0=>
      pageTurn);
   ix425 : mux21 port map ( Y=>outRegPage(14), A0=>nx1023, A1=>nx909, S0=>
      pageTurn);
   ix453 : mux21 port map ( Y=>outRegPage(15), A0=>nx1030, A1=>nx916, S0=>
      pageTurn);
   ix1053 : inv01 port map ( Y=>nx1054, A=>nx1086);
   ix1055 : inv01 port map ( Y=>nx1056, A=>nx807);
   ix1057 : inv02 port map ( Y=>nx1058, A=>nx1056);
   ix1059 : inv02 port map ( Y=>nx1060, A=>nx1056);
   ix1061 : inv02 port map ( Y=>nx1062, A=>nx1056);
   ix1063 : inv02 port map ( Y=>nx1064, A=>nx1056);
   ix1065 : inv02 port map ( Y=>nx1066, A=>nx1056);
   ix1067 : inv01 port map ( Y=>nx1068, A=>nx921);
   ix1069 : inv02 port map ( Y=>nx1070, A=>nx1068);
   ix1071 : inv02 port map ( Y=>nx1072, A=>nx1068);
   ix1073 : inv02 port map ( Y=>nx1074, A=>nx1068);
   ix1075 : inv02 port map ( Y=>nx1076, A=>nx1068);
   ix1077 : inv02 port map ( Y=>nx1078, A=>nx1068);
   ix1083 : inv02 port map ( Y=>nx1084, A=>nx1090);
   ix1085 : inv02 port map ( Y=>nx1086, A=>nx1090);
   ix1087 : inv02 port map ( Y=>nx1088, A=>enableRegFilter);
   ix1089 : inv02 port map ( Y=>nx1090, A=>enableRegFilter);
end RegUnitArch_xmplrcopy ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity RegUnit_8_16_unfolded3 is
   port (
      filterBus : IN std_logic_vector (7 DOWNTO 0) ;
      windowBus : IN std_logic_vector (15 DOWNTO 0) ;
      regPage1NextUnit : IN std_logic_vector (15 DOWNTO 0) ;
      regPage2NextUnit : IN std_logic_vector (15 DOWNTO 0) ;
      clk : IN std_logic ;
      rst : IN std_logic ;
      enableRegPage1 : IN std_logic ;
      enableRegPage2 : IN std_logic ;
      enableRegFilter : IN std_logic ;
      page1ReadBusOrPage2 : IN std_logic ;
      page2ReadBusOrPage1 : IN std_logic ;
      pageTurn : IN std_logic ;
      outRegPage : OUT std_logic_vector (15 DOWNTO 0) ;
      outputRegPage1 : OUT std_logic_vector (15 DOWNTO 0) ;
      outputRegPage2 : OUT std_logic_vector (15 DOWNTO 0) ;
      outFilter : OUT std_logic_vector (7 DOWNTO 0)) ;
end RegUnit_8_16_unfolded3 ;

architecture RegUnitArch_unfold_2792_2_xmplrcopy of RegUnit_8_16_unfolded3
    is
   signal outputRegPage1_15_EXMPLR, outputRegPage1_14_EXMPLR, 
      outputRegPage1_13_EXMPLR, outputRegPage1_12_EXMPLR, 
      outputRegPage1_11_EXMPLR, outputRegPage1_10_EXMPLR, 
      outputRegPage1_9_EXMPLR, outputRegPage1_8_EXMPLR, 
      outputRegPage1_7_EXMPLR, outputRegPage1_6_EXMPLR, 
      outputRegPage1_5_EXMPLR, outputRegPage1_4_EXMPLR, 
      outputRegPage1_3_EXMPLR, outputRegPage1_2_EXMPLR, 
      outputRegPage1_1_EXMPLR, outputRegPage1_0_EXMPLR, 
      outputRegPage2_15_EXMPLR, outputRegPage2_14_EXMPLR, 
      outputRegPage2_13_EXMPLR, outputRegPage2_12_EXMPLR, 
      outputRegPage2_11_EXMPLR, outputRegPage2_10_EXMPLR, 
      outputRegPage2_9_EXMPLR, outputRegPage2_8_EXMPLR, 
      outputRegPage2_7_EXMPLR, outputRegPage2_6_EXMPLR, 
      outputRegPage2_5_EXMPLR, outputRegPage2_4_EXMPLR, 
      outputRegPage2_3_EXMPLR, outputRegPage2_2_EXMPLR, 
      outputRegPage2_1_EXMPLR, outputRegPage2_0_EXMPLR, outFilter_7_EXMPLR, 
      outFilter_6_EXMPLR, outFilter_5_EXMPLR, outFilter_4_EXMPLR, 
      outFilter_3_EXMPLR, outFilter_2_EXMPLR, outFilter_1_EXMPLR, 
      outFilter_0_EXMPLR, nx133, nx143, nx153, nx163, nx173, nx183, nx193, 
      nx203, nx213, nx223, nx233, nx243, nx253, nx263, nx273, nx283, nx293, 
      nx303, nx313, nx323, nx333, nx343, nx353, nx363, nx373, nx383, nx393, 
      nx403, nx413, nx423, nx433, nx443, nx453, nx463, nx473, nx483, nx493, 
      nx503, nx513, nx523, nx535, nx539, nx544, nx546, nx551, nx553, nx558, 
      nx560, nx565, nx567, nx572, nx574, nx579, nx581, nx586, nx588, nx593, 
      nx595, nx597, nx599, nx601, nx604, nx606, nx608, nx611, nx613, nx615, 
      nx618, nx620, nx622, nx625, nx627, nx629, nx632, nx634, nx636, nx639, 
      nx641, nx643, nx646, nx648, nx650, nx653, nx655, nx657, nx660, nx662, 
      nx664, nx667, nx669, nx671, nx674, nx676, nx678, nx681, nx683, nx685, 
      nx688, nx690, nx692, nx695, nx697, nx699, nx702, nx704, nx706, nx709, 
      nx711, nx713, nx715, nx717, nx720, nx722, nx724, nx727, nx729, nx731, 
      nx734, nx736, nx738, nx741, nx743, nx745, nx748, nx750, nx752, nx755, 
      nx757, nx759, nx762, nx764, nx766, nx769, nx771, nx773, nx776, nx778, 
      nx780, nx783, nx785, nx787, nx790, nx792, nx794, nx797, nx799, nx801, 
      nx804, nx806, nx808, nx811, nx813, nx815, nx818, nx820, nx822, nx846, 
      nx848, nx850, nx852, nx854, nx856, nx858, nx860, nx862, nx868, nx870, 
      nx872, nx874, nx876, nx878, nx880, nx882, nx884, nx886, nx888, nx890: 
   std_logic ;

begin
   outputRegPage1(15) <= outputRegPage1_15_EXMPLR ;
   outputRegPage1(14) <= outputRegPage1_14_EXMPLR ;
   outputRegPage1(13) <= outputRegPage1_13_EXMPLR ;
   outputRegPage1(12) <= outputRegPage1_12_EXMPLR ;
   outputRegPage1(11) <= outputRegPage1_11_EXMPLR ;
   outputRegPage1(10) <= outputRegPage1_10_EXMPLR ;
   outputRegPage1(9) <= outputRegPage1_9_EXMPLR ;
   outputRegPage1(8) <= outputRegPage1_8_EXMPLR ;
   outputRegPage1(7) <= outputRegPage1_7_EXMPLR ;
   outputRegPage1(6) <= outputRegPage1_6_EXMPLR ;
   outputRegPage1(5) <= outputRegPage1_5_EXMPLR ;
   outputRegPage1(4) <= outputRegPage1_4_EXMPLR ;
   outputRegPage1(3) <= outputRegPage1_3_EXMPLR ;
   outputRegPage1(2) <= outputRegPage1_2_EXMPLR ;
   outputRegPage1(1) <= outputRegPage1_1_EXMPLR ;
   outputRegPage1(0) <= outputRegPage1_0_EXMPLR ;
   outputRegPage2(15) <= outputRegPage2_15_EXMPLR ;
   outputRegPage2(14) <= outputRegPage2_14_EXMPLR ;
   outputRegPage2(13) <= outputRegPage2_13_EXMPLR ;
   outputRegPage2(12) <= outputRegPage2_12_EXMPLR ;
   outputRegPage2(11) <= outputRegPage2_11_EXMPLR ;
   outputRegPage2(10) <= outputRegPage2_10_EXMPLR ;
   outputRegPage2(9) <= outputRegPage2_9_EXMPLR ;
   outputRegPage2(8) <= outputRegPage2_8_EXMPLR ;
   outputRegPage2(7) <= outputRegPage2_7_EXMPLR ;
   outputRegPage2(6) <= outputRegPage2_6_EXMPLR ;
   outputRegPage2(5) <= outputRegPage2_5_EXMPLR ;
   outputRegPage2(4) <= outputRegPage2_4_EXMPLR ;
   outputRegPage2(3) <= outputRegPage2_3_EXMPLR ;
   outputRegPage2(2) <= outputRegPage2_2_EXMPLR ;
   outputRegPage2(1) <= outputRegPage2_1_EXMPLR ;
   outputRegPage2(0) <= outputRegPage2_0_EXMPLR ;
   outFilter(7) <= outFilter_7_EXMPLR ;
   outFilter(6) <= outFilter_6_EXMPLR ;
   outFilter(5) <= outFilter_5_EXMPLR ;
   outFilter(4) <= outFilter_4_EXMPLR ;
   outFilter(3) <= outFilter_3_EXMPLR ;
   outFilter(2) <= outFilter_2_EXMPLR ;
   outFilter(1) <= outFilter_1_EXMPLR ;
   outFilter(0) <= outFilter_0_EXMPLR ;
   regFilterMap_reg_Q_0 : dffr port map ( Q=>outFilter_0_EXMPLR, QB=>OPEN, D
      =>nx453, CLK=>clk, R=>rst);
   ix454 : nand02 port map ( Y=>nx453, A0=>nx535, A1=>nx539);
   ix536 : nand02 port map ( Y=>nx535, A0=>outFilter_0_EXMPLR, A1=>nx888);
   ix540 : nand02 port map ( Y=>nx539, A0=>filterBus(0), A1=>nx884);
   regFilterMap_reg_Q_1 : dffr port map ( Q=>outFilter_1_EXMPLR, QB=>OPEN, D
      =>nx463, CLK=>clk, R=>rst);
   ix464 : nand02 port map ( Y=>nx463, A0=>nx544, A1=>nx546);
   ix545 : nand02 port map ( Y=>nx544, A0=>outFilter_1_EXMPLR, A1=>nx888);
   ix547 : nand02 port map ( Y=>nx546, A0=>filterBus(1), A1=>nx884);
   regFilterMap_reg_Q_2 : dffr port map ( Q=>outFilter_2_EXMPLR, QB=>OPEN, D
      =>nx473, CLK=>clk, R=>rst);
   ix474 : nand02 port map ( Y=>nx473, A0=>nx551, A1=>nx553);
   ix552 : nand02 port map ( Y=>nx551, A0=>outFilter_2_EXMPLR, A1=>nx888);
   ix554 : nand02 port map ( Y=>nx553, A0=>filterBus(2), A1=>nx884);
   regFilterMap_reg_Q_3 : dffr port map ( Q=>outFilter_3_EXMPLR, QB=>OPEN, D
      =>nx483, CLK=>clk, R=>rst);
   ix484 : nand02 port map ( Y=>nx483, A0=>nx558, A1=>nx560);
   ix559 : nand02 port map ( Y=>nx558, A0=>outFilter_3_EXMPLR, A1=>nx888);
   ix561 : nand02 port map ( Y=>nx560, A0=>filterBus(3), A1=>nx884);
   regFilterMap_reg_Q_4 : dffr port map ( Q=>outFilter_4_EXMPLR, QB=>OPEN, D
      =>nx493, CLK=>clk, R=>rst);
   ix494 : nand02 port map ( Y=>nx493, A0=>nx565, A1=>nx567);
   ix566 : nand02 port map ( Y=>nx565, A0=>outFilter_4_EXMPLR, A1=>nx888);
   ix568 : nand02 port map ( Y=>nx567, A0=>filterBus(4), A1=>nx884);
   regFilterMap_reg_Q_5 : dffr port map ( Q=>outFilter_5_EXMPLR, QB=>OPEN, D
      =>nx503, CLK=>clk, R=>rst);
   ix504 : nand02 port map ( Y=>nx503, A0=>nx572, A1=>nx574);
   ix573 : nand02 port map ( Y=>nx572, A0=>outFilter_5_EXMPLR, A1=>nx888);
   ix575 : nand02 port map ( Y=>nx574, A0=>filterBus(5), A1=>nx884);
   regFilterMap_reg_Q_6 : dffr port map ( Q=>outFilter_6_EXMPLR, QB=>OPEN, D
      =>nx513, CLK=>clk, R=>rst);
   ix514 : nand02 port map ( Y=>nx513, A0=>nx579, A1=>nx581);
   ix580 : nand02 port map ( Y=>nx579, A0=>outFilter_6_EXMPLR, A1=>nx888);
   ix582 : nand02 port map ( Y=>nx581, A0=>filterBus(6), A1=>nx884);
   regFilterMap_reg_Q_7 : dffr port map ( Q=>outFilter_7_EXMPLR, QB=>OPEN, D
      =>nx523, CLK=>clk, R=>rst);
   ix524 : nand02 port map ( Y=>nx523, A0=>nx586, A1=>nx588);
   ix587 : nand02 port map ( Y=>nx586, A0=>outFilter_7_EXMPLR, A1=>nx846);
   ix589 : nand02 port map ( Y=>nx588, A0=>filterBus(7), A1=>nx886);
   regPage2Map_reg_Q_0 : dffr port map ( Q=>outputRegPage2_0_EXMPLR, QB=>
      nx601, D=>nx143, CLK=>clk, R=>rst);
   ix144 : nand02 port map ( Y=>nx143, A0=>nx593, A1=>nx597);
   ix594 : nand02 port map ( Y=>nx593, A0=>outputRegPage2_0_EXMPLR, A1=>
      nx848);
   ix596 : nor02_2x port map ( Y=>nx595, A0=>nx878, A1=>page2ReadBusOrPage1
   );
   ix598 : nand03 port map ( Y=>nx597, A0=>windowBus(0), A1=>nx852, A2=>
      nx878);
   ix600 : inv01 port map ( Y=>nx599, A=>page2ReadBusOrPage1);
   regPage2Map_reg_Q_1 : dffr port map ( Q=>outputRegPage2_1_EXMPLR, QB=>
      nx608, D=>nx163, CLK=>clk, R=>rst);
   ix164 : nand02 port map ( Y=>nx163, A0=>nx604, A1=>nx606);
   ix605 : nand02 port map ( Y=>nx604, A0=>outputRegPage2_1_EXMPLR, A1=>
      nx848);
   ix607 : nand03 port map ( Y=>nx606, A0=>windowBus(1), A1=>nx852, A2=>
      nx878);
   regPage2Map_reg_Q_2 : dffr port map ( Q=>outputRegPage2_2_EXMPLR, QB=>
      nx615, D=>nx183, CLK=>clk, R=>rst);
   ix184 : nand02 port map ( Y=>nx183, A0=>nx611, A1=>nx613);
   ix612 : nand02 port map ( Y=>nx611, A0=>outputRegPage2_2_EXMPLR, A1=>
      nx848);
   ix614 : nand03 port map ( Y=>nx613, A0=>windowBus(2), A1=>nx852, A2=>
      nx878);
   regPage2Map_reg_Q_3 : dffr port map ( Q=>outputRegPage2_3_EXMPLR, QB=>
      nx622, D=>nx203, CLK=>clk, R=>rst);
   ix204 : nand02 port map ( Y=>nx203, A0=>nx618, A1=>nx620);
   ix619 : nand02 port map ( Y=>nx618, A0=>outputRegPage2_3_EXMPLR, A1=>
      nx848);
   ix621 : nand03 port map ( Y=>nx620, A0=>windowBus(3), A1=>nx852, A2=>
      nx878);
   regPage2Map_reg_Q_4 : dffr port map ( Q=>outputRegPage2_4_EXMPLR, QB=>
      nx629, D=>nx223, CLK=>clk, R=>rst);
   ix224 : nand02 port map ( Y=>nx223, A0=>nx625, A1=>nx627);
   ix626 : nand02 port map ( Y=>nx625, A0=>outputRegPage2_4_EXMPLR, A1=>
      nx848);
   ix628 : nand03 port map ( Y=>nx627, A0=>windowBus(4), A1=>nx852, A2=>
      nx878);
   regPage2Map_reg_Q_5 : dffr port map ( Q=>outputRegPage2_5_EXMPLR, QB=>
      nx636, D=>nx243, CLK=>clk, R=>rst);
   ix244 : nand02 port map ( Y=>nx243, A0=>nx632, A1=>nx634);
   ix633 : nand02 port map ( Y=>nx632, A0=>outputRegPage2_5_EXMPLR, A1=>
      nx848);
   ix635 : nand03 port map ( Y=>nx634, A0=>windowBus(5), A1=>nx852, A2=>
      nx878);
   regPage2Map_reg_Q_6 : dffr port map ( Q=>outputRegPage2_6_EXMPLR, QB=>
      nx643, D=>nx263, CLK=>clk, R=>rst);
   ix264 : nand02 port map ( Y=>nx263, A0=>nx639, A1=>nx641);
   ix640 : nand02 port map ( Y=>nx639, A0=>outputRegPage2_6_EXMPLR, A1=>
      nx848);
   ix642 : nand03 port map ( Y=>nx641, A0=>windowBus(6), A1=>nx854, A2=>
      nx880);
   regPage2Map_reg_Q_7 : dffr port map ( Q=>outputRegPage2_7_EXMPLR, QB=>
      nx650, D=>nx283, CLK=>clk, R=>rst);
   ix284 : nand02 port map ( Y=>nx283, A0=>nx646, A1=>nx648);
   ix647 : nand02 port map ( Y=>nx646, A0=>outputRegPage2_7_EXMPLR, A1=>
      nx850);
   ix649 : nand03 port map ( Y=>nx648, A0=>windowBus(7), A1=>nx854, A2=>
      nx880);
   regPage2Map_reg_Q_8 : dffr port map ( Q=>outputRegPage2_8_EXMPLR, QB=>
      nx657, D=>nx303, CLK=>clk, R=>rst);
   ix304 : nand02 port map ( Y=>nx303, A0=>nx653, A1=>nx655);
   ix654 : nand02 port map ( Y=>nx653, A0=>outputRegPage2_8_EXMPLR, A1=>
      nx850);
   ix656 : nand03 port map ( Y=>nx655, A0=>windowBus(8), A1=>nx854, A2=>
      nx880);
   regPage2Map_reg_Q_9 : dffr port map ( Q=>outputRegPage2_9_EXMPLR, QB=>
      nx664, D=>nx323, CLK=>clk, R=>rst);
   ix324 : nand02 port map ( Y=>nx323, A0=>nx660, A1=>nx662);
   ix661 : nand02 port map ( Y=>nx660, A0=>outputRegPage2_9_EXMPLR, A1=>
      nx850);
   ix663 : nand03 port map ( Y=>nx662, A0=>windowBus(9), A1=>nx854, A2=>
      nx880);
   regPage2Map_reg_Q_10 : dffr port map ( Q=>outputRegPage2_10_EXMPLR, QB=>
      nx671, D=>nx343, CLK=>clk, R=>rst);
   ix344 : nand02 port map ( Y=>nx343, A0=>nx667, A1=>nx669);
   ix668 : nand02 port map ( Y=>nx667, A0=>outputRegPage2_10_EXMPLR, A1=>
      nx850);
   ix670 : nand03 port map ( Y=>nx669, A0=>windowBus(10), A1=>nx854, A2=>
      nx880);
   regPage2Map_reg_Q_11 : dffr port map ( Q=>outputRegPage2_11_EXMPLR, QB=>
      nx678, D=>nx363, CLK=>clk, R=>rst);
   ix364 : nand02 port map ( Y=>nx363, A0=>nx674, A1=>nx676);
   ix675 : nand02 port map ( Y=>nx674, A0=>outputRegPage2_11_EXMPLR, A1=>
      nx850);
   ix677 : nand03 port map ( Y=>nx676, A0=>windowBus(11), A1=>nx854, A2=>
      nx880);
   regPage2Map_reg_Q_12 : dffr port map ( Q=>outputRegPage2_12_EXMPLR, QB=>
      nx685, D=>nx383, CLK=>clk, R=>rst);
   ix384 : nand02 port map ( Y=>nx383, A0=>nx681, A1=>nx683);
   ix682 : nand02 port map ( Y=>nx681, A0=>outputRegPage2_12_EXMPLR, A1=>
      nx850);
   ix684 : nand03 port map ( Y=>nx683, A0=>windowBus(12), A1=>nx599, A2=>
      nx880);
   regPage2Map_reg_Q_13 : dffr port map ( Q=>outputRegPage2_13_EXMPLR, QB=>
      nx692, D=>nx403, CLK=>clk, R=>rst);
   ix404 : nand02 port map ( Y=>nx403, A0=>nx688, A1=>nx690);
   ix689 : nand02 port map ( Y=>nx688, A0=>outputRegPage2_13_EXMPLR, A1=>
      nx850);
   ix691 : nand03 port map ( Y=>nx690, A0=>windowBus(13), A1=>nx599, A2=>
      nx882);
   regPage2Map_reg_Q_14 : dffr port map ( Q=>outputRegPage2_14_EXMPLR, QB=>
      nx699, D=>nx423, CLK=>clk, R=>rst);
   ix424 : nand02 port map ( Y=>nx423, A0=>nx695, A1=>nx697);
   ix696 : nand02 port map ( Y=>nx695, A0=>outputRegPage2_14_EXMPLR, A1=>
      nx595);
   ix698 : nand03 port map ( Y=>nx697, A0=>windowBus(14), A1=>nx599, A2=>
      nx882);
   regPage2Map_reg_Q_15 : dffr port map ( Q=>outputRegPage2_15_EXMPLR, QB=>
      nx706, D=>nx443, CLK=>clk, R=>rst);
   ix444 : nand02 port map ( Y=>nx443, A0=>nx702, A1=>nx704);
   ix703 : nand02 port map ( Y=>nx702, A0=>outputRegPage2_15_EXMPLR, A1=>
      nx595);
   ix705 : nand03 port map ( Y=>nx704, A0=>windowBus(15), A1=>nx599, A2=>
      nx882);
   regPage1Map_reg_Q_0 : dffr port map ( Q=>outputRegPage1_0_EXMPLR, QB=>
      nx717, D=>nx133, CLK=>clk, R=>rst);
   ix134 : nand02 port map ( Y=>nx133, A0=>nx709, A1=>nx713);
   ix710 : nand02 port map ( Y=>nx709, A0=>outputRegPage1_0_EXMPLR, A1=>
      nx856);
   ix712 : nor02_2x port map ( Y=>nx711, A0=>nx870, A1=>page1ReadBusOrPage2
   );
   ix714 : nand03 port map ( Y=>nx713, A0=>windowBus(0), A1=>nx860, A2=>
      nx870);
   ix716 : inv01 port map ( Y=>nx715, A=>page1ReadBusOrPage2);
   regPage1Map_reg_Q_1 : dffr port map ( Q=>outputRegPage1_1_EXMPLR, QB=>
      nx724, D=>nx153, CLK=>clk, R=>rst);
   ix154 : nand02 port map ( Y=>nx153, A0=>nx720, A1=>nx722);
   ix721 : nand02 port map ( Y=>nx720, A0=>outputRegPage1_1_EXMPLR, A1=>
      nx856);
   ix723 : nand03 port map ( Y=>nx722, A0=>windowBus(1), A1=>nx860, A2=>
      nx870);
   regPage1Map_reg_Q_2 : dffr port map ( Q=>outputRegPage1_2_EXMPLR, QB=>
      nx731, D=>nx173, CLK=>clk, R=>rst);
   ix174 : nand02 port map ( Y=>nx173, A0=>nx727, A1=>nx729);
   ix728 : nand02 port map ( Y=>nx727, A0=>outputRegPage1_2_EXMPLR, A1=>
      nx856);
   ix730 : nand03 port map ( Y=>nx729, A0=>windowBus(2), A1=>nx860, A2=>
      nx870);
   regPage1Map_reg_Q_3 : dffr port map ( Q=>outputRegPage1_3_EXMPLR, QB=>
      nx738, D=>nx193, CLK=>clk, R=>rst);
   ix194 : nand02 port map ( Y=>nx193, A0=>nx734, A1=>nx736);
   ix735 : nand02 port map ( Y=>nx734, A0=>outputRegPage1_3_EXMPLR, A1=>
      nx856);
   ix737 : nand03 port map ( Y=>nx736, A0=>windowBus(3), A1=>nx860, A2=>
      nx870);
   regPage1Map_reg_Q_4 : dffr port map ( Q=>outputRegPage1_4_EXMPLR, QB=>
      nx745, D=>nx213, CLK=>clk, R=>rst);
   ix214 : nand02 port map ( Y=>nx213, A0=>nx741, A1=>nx743);
   ix742 : nand02 port map ( Y=>nx741, A0=>outputRegPage1_4_EXMPLR, A1=>
      nx856);
   ix744 : nand03 port map ( Y=>nx743, A0=>windowBus(4), A1=>nx860, A2=>
      nx870);
   regPage1Map_reg_Q_5 : dffr port map ( Q=>outputRegPage1_5_EXMPLR, QB=>
      nx752, D=>nx233, CLK=>clk, R=>rst);
   ix234 : nand02 port map ( Y=>nx233, A0=>nx748, A1=>nx750);
   ix749 : nand02 port map ( Y=>nx748, A0=>outputRegPage1_5_EXMPLR, A1=>
      nx856);
   ix751 : nand03 port map ( Y=>nx750, A0=>windowBus(5), A1=>nx860, A2=>
      nx870);
   regPage1Map_reg_Q_6 : dffr port map ( Q=>outputRegPage1_6_EXMPLR, QB=>
      nx759, D=>nx253, CLK=>clk, R=>rst);
   ix254 : nand02 port map ( Y=>nx253, A0=>nx755, A1=>nx757);
   ix756 : nand02 port map ( Y=>nx755, A0=>outputRegPage1_6_EXMPLR, A1=>
      nx856);
   ix758 : nand03 port map ( Y=>nx757, A0=>windowBus(6), A1=>nx862, A2=>
      nx872);
   regPage1Map_reg_Q_7 : dffr port map ( Q=>outputRegPage1_7_EXMPLR, QB=>
      nx766, D=>nx273, CLK=>clk, R=>rst);
   ix274 : nand02 port map ( Y=>nx273, A0=>nx762, A1=>nx764);
   ix763 : nand02 port map ( Y=>nx762, A0=>outputRegPage1_7_EXMPLR, A1=>
      nx858);
   ix765 : nand03 port map ( Y=>nx764, A0=>windowBus(7), A1=>nx862, A2=>
      nx872);
   regPage1Map_reg_Q_8 : dffr port map ( Q=>outputRegPage1_8_EXMPLR, QB=>
      nx773, D=>nx293, CLK=>clk, R=>rst);
   ix294 : nand02 port map ( Y=>nx293, A0=>nx769, A1=>nx771);
   ix770 : nand02 port map ( Y=>nx769, A0=>outputRegPage1_8_EXMPLR, A1=>
      nx858);
   ix772 : nand03 port map ( Y=>nx771, A0=>windowBus(8), A1=>nx862, A2=>
      nx872);
   regPage1Map_reg_Q_9 : dffr port map ( Q=>outputRegPage1_9_EXMPLR, QB=>
      nx780, D=>nx313, CLK=>clk, R=>rst);
   ix314 : nand02 port map ( Y=>nx313, A0=>nx776, A1=>nx778);
   ix777 : nand02 port map ( Y=>nx776, A0=>outputRegPage1_9_EXMPLR, A1=>
      nx858);
   ix779 : nand03 port map ( Y=>nx778, A0=>windowBus(9), A1=>nx862, A2=>
      nx872);
   regPage1Map_reg_Q_10 : dffr port map ( Q=>outputRegPage1_10_EXMPLR, QB=>
      nx787, D=>nx333, CLK=>clk, R=>rst);
   ix334 : nand02 port map ( Y=>nx333, A0=>nx783, A1=>nx785);
   ix784 : nand02 port map ( Y=>nx783, A0=>outputRegPage1_10_EXMPLR, A1=>
      nx858);
   ix786 : nand03 port map ( Y=>nx785, A0=>windowBus(10), A1=>nx862, A2=>
      nx872);
   regPage1Map_reg_Q_11 : dffr port map ( Q=>outputRegPage1_11_EXMPLR, QB=>
      nx794, D=>nx353, CLK=>clk, R=>rst);
   ix354 : nand02 port map ( Y=>nx353, A0=>nx790, A1=>nx792);
   ix791 : nand02 port map ( Y=>nx790, A0=>outputRegPage1_11_EXMPLR, A1=>
      nx858);
   ix793 : nand03 port map ( Y=>nx792, A0=>windowBus(11), A1=>nx862, A2=>
      nx872);
   regPage1Map_reg_Q_12 : dffr port map ( Q=>outputRegPage1_12_EXMPLR, QB=>
      nx801, D=>nx373, CLK=>clk, R=>rst);
   ix374 : nand02 port map ( Y=>nx373, A0=>nx797, A1=>nx799);
   ix798 : nand02 port map ( Y=>nx797, A0=>outputRegPage1_12_EXMPLR, A1=>
      nx858);
   ix800 : nand03 port map ( Y=>nx799, A0=>windowBus(12), A1=>nx715, A2=>
      nx872);
   regPage1Map_reg_Q_13 : dffr port map ( Q=>outputRegPage1_13_EXMPLR, QB=>
      nx808, D=>nx393, CLK=>clk, R=>rst);
   ix394 : nand02 port map ( Y=>nx393, A0=>nx804, A1=>nx806);
   ix805 : nand02 port map ( Y=>nx804, A0=>outputRegPage1_13_EXMPLR, A1=>
      nx858);
   ix807 : nand03 port map ( Y=>nx806, A0=>windowBus(13), A1=>nx715, A2=>
      nx874);
   regPage1Map_reg_Q_14 : dffr port map ( Q=>outputRegPage1_14_EXMPLR, QB=>
      nx815, D=>nx413, CLK=>clk, R=>rst);
   ix414 : nand02 port map ( Y=>nx413, A0=>nx811, A1=>nx813);
   ix812 : nand02 port map ( Y=>nx811, A0=>outputRegPage1_14_EXMPLR, A1=>
      nx711);
   ix814 : nand03 port map ( Y=>nx813, A0=>windowBus(14), A1=>nx715, A2=>
      nx874);
   regPage1Map_reg_Q_15 : dffr port map ( Q=>outputRegPage1_15_EXMPLR, QB=>
      nx822, D=>nx433, CLK=>clk, R=>rst);
   ix434 : nand02 port map ( Y=>nx433, A0=>nx818, A1=>nx820);
   ix819 : nand02 port map ( Y=>nx818, A0=>outputRegPage1_15_EXMPLR, A1=>
      nx711);
   ix821 : nand03 port map ( Y=>nx820, A0=>windowBus(15), A1=>nx715, A2=>
      nx874);
   ix25 : mux21 port map ( Y=>outRegPage(0), A0=>nx717, A1=>nx601, S0=>
      pageTurn);
   ix45 : mux21 port map ( Y=>outRegPage(1), A0=>nx724, A1=>nx608, S0=>
      pageTurn);
   ix65 : mux21 port map ( Y=>outRegPage(2), A0=>nx731, A1=>nx615, S0=>
      pageTurn);
   ix85 : mux21 port map ( Y=>outRegPage(3), A0=>nx738, A1=>nx622, S0=>
      pageTurn);
   ix105 : mux21 port map ( Y=>outRegPage(4), A0=>nx745, A1=>nx629, S0=>
      pageTurn);
   ix125 : mux21 port map ( Y=>outRegPage(5), A0=>nx752, A1=>nx636, S0=>
      pageTurn);
   ix145 : mux21 port map ( Y=>outRegPage(6), A0=>nx759, A1=>nx643, S0=>
      pageTurn);
   ix165 : mux21 port map ( Y=>outRegPage(7), A0=>nx766, A1=>nx650, S0=>
      pageTurn);
   ix185 : mux21 port map ( Y=>outRegPage(8), A0=>nx773, A1=>nx657, S0=>
      pageTurn);
   ix205 : mux21 port map ( Y=>outRegPage(9), A0=>nx780, A1=>nx664, S0=>
      pageTurn);
   ix225 : mux21 port map ( Y=>outRegPage(10), A0=>nx787, A1=>nx671, S0=>
      pageTurn);
   ix245 : mux21 port map ( Y=>outRegPage(11), A0=>nx794, A1=>nx678, S0=>
      pageTurn);
   ix265 : mux21 port map ( Y=>outRegPage(12), A0=>nx801, A1=>nx685, S0=>
      pageTurn);
   ix285 : mux21 port map ( Y=>outRegPage(13), A0=>nx808, A1=>nx692, S0=>
      pageTurn);
   ix305 : mux21 port map ( Y=>outRegPage(14), A0=>nx815, A1=>nx699, S0=>
      pageTurn);
   ix325 : mux21 port map ( Y=>outRegPage(15), A0=>nx822, A1=>nx706, S0=>
      pageTurn);
   ix845 : inv01 port map ( Y=>nx846, A=>nx886);
   ix847 : nor02_2x port map ( Y=>nx848, A0=>nx882, A1=>page2ReadBusOrPage1
   );
   ix849 : nor02_2x port map ( Y=>nx850, A0=>nx882, A1=>page2ReadBusOrPage1
   );
   ix851 : inv01 port map ( Y=>nx852, A=>page2ReadBusOrPage1);
   ix853 : inv01 port map ( Y=>nx854, A=>page2ReadBusOrPage1);
   ix855 : nor02_2x port map ( Y=>nx856, A0=>nx874, A1=>page1ReadBusOrPage2
   );
   ix857 : nor02_2x port map ( Y=>nx858, A0=>nx874, A1=>page1ReadBusOrPage2
   );
   ix859 : inv01 port map ( Y=>nx860, A=>page1ReadBusOrPage2);
   ix861 : inv01 port map ( Y=>nx862, A=>page1ReadBusOrPage2);
   ix867 : inv01 port map ( Y=>nx868, A=>enableRegPage1);
   ix869 : inv02 port map ( Y=>nx870, A=>nx868);
   ix871 : inv02 port map ( Y=>nx872, A=>nx868);
   ix873 : inv02 port map ( Y=>nx874, A=>nx868);
   ix875 : inv01 port map ( Y=>nx876, A=>enableRegPage2);
   ix877 : inv02 port map ( Y=>nx878, A=>nx876);
   ix879 : inv02 port map ( Y=>nx880, A=>nx876);
   ix881 : inv02 port map ( Y=>nx882, A=>nx876);
   ix883 : inv02 port map ( Y=>nx884, A=>nx890);
   ix885 : inv02 port map ( Y=>nx886, A=>nx890);
   ix887 : inv02 port map ( Y=>nx888, A=>enableRegFilter);
   ix889 : inv02 port map ( Y=>nx890, A=>enableRegFilter);
end RegUnitArch_unfold_2792_2_xmplrcopy ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity NBitAdder_16 is
   port (
      a : IN std_logic_vector (15 DOWNTO 0) ;
      b : IN std_logic_vector (15 DOWNTO 0) ;
      carryIn : IN std_logic ;
      sum : OUT std_logic_vector (15 DOWNTO 0) ;
      carryOut : OUT std_logic) ;
end NBitAdder_16 ;

architecture NBitAdderArch_unfold_2263 of NBitAdder_16 is
   signal nx2, nx8, nx10, nx18, nx24, nx26, nx34, nx40, nx42, nx50, nx56, 
      nx58, nx66, nx72, nx74, nx82, nx88, nx90, nx98, nx104, nx106, nx114, 
      nx85, nx89, nx93, nx99, nx101, nx103, nx107, nx111, nx115, nx121, 
      nx123, nx125, nx129, nx133, nx137, nx143, nx145, nx147, nx151, nx154, 
      nx157, nx161, nx163, nx165, nx168, nx171, nx174, nx178, nx180, nx182, 
      nx185, nx188, nx191, nx195, nx197, nx199, nx202, nx205, nx208, nx212, 
      nx214, nx216, nx219, nx222, nx225: std_logic ;

begin
   ix42 : fake_gnd port map ( Y=>carryOut);
   ix151 : xnor2 port map ( Y=>sum(0), A0=>b(0), A1=>nx85);
   ix86 : inv01 port map ( Y=>nx85, A=>a(0));
   ix145 : xnor2 port map ( Y=>sum(1), A0=>nx89, A1=>nx2);
   ix90 : nand02 port map ( Y=>nx89, A0=>b(0), A1=>a(0));
   ix3 : xnor2 port map ( Y=>nx2, A0=>a(1), A1=>nx93);
   ix94 : inv01 port map ( Y=>nx93, A=>b(1));
   ix143 : xnor2 port map ( Y=>sum(2), A0=>nx8, A1=>nx103);
   ix9 : oai22 port map ( Y=>nx8, A0=>nx89, A1=>nx99, B0=>nx93, B1=>nx101);
   ix100 : xnor2 port map ( Y=>nx99, A0=>a(1), A1=>b(1));
   ix102 : inv01 port map ( Y=>nx101, A=>a(1));
   ix104 : xnor2 port map ( Y=>nx103, A0=>a(2), A1=>b(2));
   ix141 : xnor2 port map ( Y=>sum(3), A0=>nx107, A1=>nx18);
   ix108 : aoi22 port map ( Y=>nx107, A0=>b(2), A1=>a(2), B0=>nx8, B1=>nx10
   );
   ix11 : xnor2 port map ( Y=>nx10, A0=>a(2), A1=>nx111);
   ix112 : inv01 port map ( Y=>nx111, A=>b(2));
   ix19 : xnor2 port map ( Y=>nx18, A0=>a(3), A1=>nx115);
   ix116 : inv01 port map ( Y=>nx115, A=>b(3));
   ix139 : xnor2 port map ( Y=>sum(4), A0=>nx24, A1=>nx125);
   ix25 : oai21 port map ( Y=>nx24, A0=>nx107, A1=>nx121, B0=>nx123);
   ix122 : xnor2 port map ( Y=>nx121, A0=>a(3), A1=>b(3));
   ix124 : nand02 port map ( Y=>nx123, A0=>b(3), A1=>a(3));
   ix126 : xnor2 port map ( Y=>nx125, A0=>a(4), A1=>b(4));
   ix137 : xnor2 port map ( Y=>sum(5), A0=>nx129, A1=>nx34);
   ix130 : aoi22 port map ( Y=>nx129, A0=>b(4), A1=>a(4), B0=>nx24, B1=>nx26
   );
   ix27 : xnor2 port map ( Y=>nx26, A0=>a(4), A1=>nx133);
   ix134 : inv01 port map ( Y=>nx133, A=>b(4));
   ix35 : xnor2 port map ( Y=>nx34, A0=>a(5), A1=>nx137);
   ix138 : inv01 port map ( Y=>nx137, A=>b(5));
   ix135 : xnor2 port map ( Y=>sum(6), A0=>nx40, A1=>nx147);
   ix41 : oai21 port map ( Y=>nx40, A0=>nx129, A1=>nx143, B0=>nx145);
   ix144 : xnor2 port map ( Y=>nx143, A0=>a(5), A1=>b(5));
   ix146 : nand02 port map ( Y=>nx145, A0=>b(5), A1=>a(5));
   ix148 : xnor2 port map ( Y=>nx147, A0=>a(6), A1=>b(6));
   ix133 : xnor2 port map ( Y=>sum(7), A0=>nx151, A1=>nx50);
   ix152 : aoi22 port map ( Y=>nx151, A0=>b(6), A1=>a(6), B0=>nx40, B1=>nx42
   );
   ix43 : xnor2 port map ( Y=>nx42, A0=>a(6), A1=>nx154);
   ix155 : inv01 port map ( Y=>nx154, A=>b(6));
   ix51 : xnor2 port map ( Y=>nx50, A0=>a(7), A1=>nx157);
   ix158 : inv01 port map ( Y=>nx157, A=>b(7));
   ix131 : xnor2 port map ( Y=>sum(8), A0=>nx56, A1=>nx165);
   ix57 : oai21 port map ( Y=>nx56, A0=>nx151, A1=>nx161, B0=>nx163);
   ix162 : xnor2 port map ( Y=>nx161, A0=>a(7), A1=>b(7));
   ix164 : nand02 port map ( Y=>nx163, A0=>b(7), A1=>a(7));
   ix166 : xnor2 port map ( Y=>nx165, A0=>a(8), A1=>b(8));
   ix129 : xnor2 port map ( Y=>sum(9), A0=>nx168, A1=>nx66);
   ix169 : aoi22 port map ( Y=>nx168, A0=>b(8), A1=>a(8), B0=>nx56, B1=>nx58
   );
   ix59 : xnor2 port map ( Y=>nx58, A0=>a(8), A1=>nx171);
   ix172 : inv01 port map ( Y=>nx171, A=>b(8));
   ix67 : xnor2 port map ( Y=>nx66, A0=>a(9), A1=>nx174);
   ix175 : inv01 port map ( Y=>nx174, A=>b(9));
   ix127 : xnor2 port map ( Y=>sum(10), A0=>nx72, A1=>nx182);
   ix73 : oai21 port map ( Y=>nx72, A0=>nx168, A1=>nx178, B0=>nx180);
   ix179 : xnor2 port map ( Y=>nx178, A0=>a(9), A1=>b(9));
   ix181 : nand02 port map ( Y=>nx180, A0=>b(9), A1=>a(9));
   ix183 : xnor2 port map ( Y=>nx182, A0=>a(10), A1=>b(10));
   ix125 : xnor2 port map ( Y=>sum(11), A0=>nx185, A1=>nx82);
   ix186 : aoi22 port map ( Y=>nx185, A0=>b(10), A1=>a(10), B0=>nx72, B1=>
      nx74);
   ix75 : xnor2 port map ( Y=>nx74, A0=>a(10), A1=>nx188);
   ix189 : inv01 port map ( Y=>nx188, A=>b(10));
   ix83 : xnor2 port map ( Y=>nx82, A0=>a(11), A1=>nx191);
   ix192 : inv01 port map ( Y=>nx191, A=>b(11));
   ix123 : xnor2 port map ( Y=>sum(12), A0=>nx88, A1=>nx199);
   ix89 : oai21 port map ( Y=>nx88, A0=>nx185, A1=>nx195, B0=>nx197);
   ix196 : xnor2 port map ( Y=>nx195, A0=>a(11), A1=>b(11));
   ix198 : nand02 port map ( Y=>nx197, A0=>b(11), A1=>a(11));
   ix200 : xnor2 port map ( Y=>nx199, A0=>a(12), A1=>b(12));
   ix121 : xnor2 port map ( Y=>sum(13), A0=>nx202, A1=>nx98);
   ix203 : aoi22 port map ( Y=>nx202, A0=>b(12), A1=>a(12), B0=>nx88, B1=>
      nx90);
   ix91 : xnor2 port map ( Y=>nx90, A0=>a(12), A1=>nx205);
   ix206 : inv01 port map ( Y=>nx205, A=>b(12));
   ix99 : xnor2 port map ( Y=>nx98, A0=>a(13), A1=>nx208);
   ix209 : inv01 port map ( Y=>nx208, A=>b(13));
   ix119 : xnor2 port map ( Y=>sum(14), A0=>nx104, A1=>nx216);
   ix105 : oai21 port map ( Y=>nx104, A0=>nx202, A1=>nx212, B0=>nx214);
   ix213 : xnor2 port map ( Y=>nx212, A0=>a(13), A1=>b(13));
   ix215 : nand02 port map ( Y=>nx214, A0=>b(13), A1=>a(13));
   ix217 : xnor2 port map ( Y=>nx216, A0=>a(14), A1=>b(14));
   ix117 : xnor2 port map ( Y=>sum(15), A0=>nx219, A1=>nx114);
   ix220 : aoi22 port map ( Y=>nx219, A0=>b(14), A1=>a(14), B0=>nx104, B1=>
      nx106);
   ix107 : xnor2 port map ( Y=>nx106, A0=>a(14), A1=>nx222);
   ix223 : inv01 port map ( Y=>nx222, A=>b(14));
   ix115 : xnor2 port map ( Y=>nx114, A0=>a(15), A1=>nx225);
   ix226 : inv01 port map ( Y=>nx225, A=>b(15));
end NBitAdderArch_unfold_2263 ;

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity CNNCores is
   port (
      filterBus : IN std_logic_vector (39 DOWNTO 0) ;
      windowBus : IN std_logic_vector (79 DOWNTO 0) ;
      decoderRow : IN std_logic_vector (2 DOWNTO 0) ;
      clk : IN std_logic ;
      rst : IN std_logic ;
      writePage1 : IN std_logic ;
      writePage2 : IN std_logic ;
      writeFilter : IN std_logic ;
      shift2To1 : IN std_logic ;
      shift1To2 : IN std_logic ;
      pageTurn : IN std_logic ;
      start : IN std_logic ;
      layerType : IN std_logic ;
      filterType : IN std_logic ;
      done : OUT std_logic ;
      finalSum : OUT std_logic_vector (15 DOWNTO 0)) ;
end CNNCores ;

architecture CNNCoresArch of CNNCores is
   component CNNMuls_25
      port (
         filter_24_7 : IN std_logic ;
         filter_24_6 : IN std_logic ;
         filter_24_5 : IN std_logic ;
         filter_24_4 : IN std_logic ;
         filter_24_3 : IN std_logic ;
         filter_24_2 : IN std_logic ;
         filter_24_1 : IN std_logic ;
         filter_24_0 : IN std_logic ;
         filter_23_7 : IN std_logic ;
         filter_23_6 : IN std_logic ;
         filter_23_5 : IN std_logic ;
         filter_23_4 : IN std_logic ;
         filter_23_3 : IN std_logic ;
         filter_23_2 : IN std_logic ;
         filter_23_1 : IN std_logic ;
         filter_23_0 : IN std_logic ;
         filter_22_7 : IN std_logic ;
         filter_22_6 : IN std_logic ;
         filter_22_5 : IN std_logic ;
         filter_22_4 : IN std_logic ;
         filter_22_3 : IN std_logic ;
         filter_22_2 : IN std_logic ;
         filter_22_1 : IN std_logic ;
         filter_22_0 : IN std_logic ;
         filter_21_7 : IN std_logic ;
         filter_21_6 : IN std_logic ;
         filter_21_5 : IN std_logic ;
         filter_21_4 : IN std_logic ;
         filter_21_3 : IN std_logic ;
         filter_21_2 : IN std_logic ;
         filter_21_1 : IN std_logic ;
         filter_21_0 : IN std_logic ;
         filter_20_7 : IN std_logic ;
         filter_20_6 : IN std_logic ;
         filter_20_5 : IN std_logic ;
         filter_20_4 : IN std_logic ;
         filter_20_3 : IN std_logic ;
         filter_20_2 : IN std_logic ;
         filter_20_1 : IN std_logic ;
         filter_20_0 : IN std_logic ;
         filter_19_7 : IN std_logic ;
         filter_19_6 : IN std_logic ;
         filter_19_5 : IN std_logic ;
         filter_19_4 : IN std_logic ;
         filter_19_3 : IN std_logic ;
         filter_19_2 : IN std_logic ;
         filter_19_1 : IN std_logic ;
         filter_19_0 : IN std_logic ;
         filter_18_7 : IN std_logic ;
         filter_18_6 : IN std_logic ;
         filter_18_5 : IN std_logic ;
         filter_18_4 : IN std_logic ;
         filter_18_3 : IN std_logic ;
         filter_18_2 : IN std_logic ;
         filter_18_1 : IN std_logic ;
         filter_18_0 : IN std_logic ;
         filter_17_7 : IN std_logic ;
         filter_17_6 : IN std_logic ;
         filter_17_5 : IN std_logic ;
         filter_17_4 : IN std_logic ;
         filter_17_3 : IN std_logic ;
         filter_17_2 : IN std_logic ;
         filter_17_1 : IN std_logic ;
         filter_17_0 : IN std_logic ;
         filter_16_7 : IN std_logic ;
         filter_16_6 : IN std_logic ;
         filter_16_5 : IN std_logic ;
         filter_16_4 : IN std_logic ;
         filter_16_3 : IN std_logic ;
         filter_16_2 : IN std_logic ;
         filter_16_1 : IN std_logic ;
         filter_16_0 : IN std_logic ;
         filter_15_7 : IN std_logic ;
         filter_15_6 : IN std_logic ;
         filter_15_5 : IN std_logic ;
         filter_15_4 : IN std_logic ;
         filter_15_3 : IN std_logic ;
         filter_15_2 : IN std_logic ;
         filter_15_1 : IN std_logic ;
         filter_15_0 : IN std_logic ;
         filter_14_7 : IN std_logic ;
         filter_14_6 : IN std_logic ;
         filter_14_5 : IN std_logic ;
         filter_14_4 : IN std_logic ;
         filter_14_3 : IN std_logic ;
         filter_14_2 : IN std_logic ;
         filter_14_1 : IN std_logic ;
         filter_14_0 : IN std_logic ;
         filter_13_7 : IN std_logic ;
         filter_13_6 : IN std_logic ;
         filter_13_5 : IN std_logic ;
         filter_13_4 : IN std_logic ;
         filter_13_3 : IN std_logic ;
         filter_13_2 : IN std_logic ;
         filter_13_1 : IN std_logic ;
         filter_13_0 : IN std_logic ;
         filter_12_7 : IN std_logic ;
         filter_12_6 : IN std_logic ;
         filter_12_5 : IN std_logic ;
         filter_12_4 : IN std_logic ;
         filter_12_3 : IN std_logic ;
         filter_12_2 : IN std_logic ;
         filter_12_1 : IN std_logic ;
         filter_12_0 : IN std_logic ;
         filter_11_7 : IN std_logic ;
         filter_11_6 : IN std_logic ;
         filter_11_5 : IN std_logic ;
         filter_11_4 : IN std_logic ;
         filter_11_3 : IN std_logic ;
         filter_11_2 : IN std_logic ;
         filter_11_1 : IN std_logic ;
         filter_11_0 : IN std_logic ;
         filter_10_7 : IN std_logic ;
         filter_10_6 : IN std_logic ;
         filter_10_5 : IN std_logic ;
         filter_10_4 : IN std_logic ;
         filter_10_3 : IN std_logic ;
         filter_10_2 : IN std_logic ;
         filter_10_1 : IN std_logic ;
         filter_10_0 : IN std_logic ;
         filter_9_7 : IN std_logic ;
         filter_9_6 : IN std_logic ;
         filter_9_5 : IN std_logic ;
         filter_9_4 : IN std_logic ;
         filter_9_3 : IN std_logic ;
         filter_9_2 : IN std_logic ;
         filter_9_1 : IN std_logic ;
         filter_9_0 : IN std_logic ;
         filter_8_7 : IN std_logic ;
         filter_8_6 : IN std_logic ;
         filter_8_5 : IN std_logic ;
         filter_8_4 : IN std_logic ;
         filter_8_3 : IN std_logic ;
         filter_8_2 : IN std_logic ;
         filter_8_1 : IN std_logic ;
         filter_8_0 : IN std_logic ;
         filter_7_7 : IN std_logic ;
         filter_7_6 : IN std_logic ;
         filter_7_5 : IN std_logic ;
         filter_7_4 : IN std_logic ;
         filter_7_3 : IN std_logic ;
         filter_7_2 : IN std_logic ;
         filter_7_1 : IN std_logic ;
         filter_7_0 : IN std_logic ;
         filter_6_7 : IN std_logic ;
         filter_6_6 : IN std_logic ;
         filter_6_5 : IN std_logic ;
         filter_6_4 : IN std_logic ;
         filter_6_3 : IN std_logic ;
         filter_6_2 : IN std_logic ;
         filter_6_1 : IN std_logic ;
         filter_6_0 : IN std_logic ;
         filter_5_7 : IN std_logic ;
         filter_5_6 : IN std_logic ;
         filter_5_5 : IN std_logic ;
         filter_5_4 : IN std_logic ;
         filter_5_3 : IN std_logic ;
         filter_5_2 : IN std_logic ;
         filter_5_1 : IN std_logic ;
         filter_5_0 : IN std_logic ;
         filter_4_7 : IN std_logic ;
         filter_4_6 : IN std_logic ;
         filter_4_5 : IN std_logic ;
         filter_4_4 : IN std_logic ;
         filter_4_3 : IN std_logic ;
         filter_4_2 : IN std_logic ;
         filter_4_1 : IN std_logic ;
         filter_4_0 : IN std_logic ;
         filter_3_7 : IN std_logic ;
         filter_3_6 : IN std_logic ;
         filter_3_5 : IN std_logic ;
         filter_3_4 : IN std_logic ;
         filter_3_3 : IN std_logic ;
         filter_3_2 : IN std_logic ;
         filter_3_1 : IN std_logic ;
         filter_3_0 : IN std_logic ;
         filter_2_7 : IN std_logic ;
         filter_2_6 : IN std_logic ;
         filter_2_5 : IN std_logic ;
         filter_2_4 : IN std_logic ;
         filter_2_3 : IN std_logic ;
         filter_2_2 : IN std_logic ;
         filter_2_1 : IN std_logic ;
         filter_2_0 : IN std_logic ;
         filter_1_7 : IN std_logic ;
         filter_1_6 : IN std_logic ;
         filter_1_5 : IN std_logic ;
         filter_1_4 : IN std_logic ;
         filter_1_3 : IN std_logic ;
         filter_1_2 : IN std_logic ;
         filter_1_1 : IN std_logic ;
         filter_1_0 : IN std_logic ;
         filter_0_7 : IN std_logic ;
         filter_0_6 : IN std_logic ;
         filter_0_5 : IN std_logic ;
         filter_0_4 : IN std_logic ;
         filter_0_3 : IN std_logic ;
         filter_0_2 : IN std_logic ;
         filter_0_1 : IN std_logic ;
         filter_0_0 : IN std_logic ;
         window_24_15 : IN std_logic ;
         window_24_14 : IN std_logic ;
         window_24_13 : IN std_logic ;
         window_24_12 : IN std_logic ;
         window_24_11 : IN std_logic ;
         window_24_10 : IN std_logic ;
         window_24_9 : IN std_logic ;
         window_24_8 : IN std_logic ;
         window_24_7 : IN std_logic ;
         window_24_6 : IN std_logic ;
         window_24_5 : IN std_logic ;
         window_24_4 : IN std_logic ;
         window_24_3 : IN std_logic ;
         window_24_2 : IN std_logic ;
         window_24_1 : IN std_logic ;
         window_24_0 : IN std_logic ;
         window_23_15 : IN std_logic ;
         window_23_14 : IN std_logic ;
         window_23_13 : IN std_logic ;
         window_23_12 : IN std_logic ;
         window_23_11 : IN std_logic ;
         window_23_10 : IN std_logic ;
         window_23_9 : IN std_logic ;
         window_23_8 : IN std_logic ;
         window_23_7 : IN std_logic ;
         window_23_6 : IN std_logic ;
         window_23_5 : IN std_logic ;
         window_23_4 : IN std_logic ;
         window_23_3 : IN std_logic ;
         window_23_2 : IN std_logic ;
         window_23_1 : IN std_logic ;
         window_23_0 : IN std_logic ;
         window_22_15 : IN std_logic ;
         window_22_14 : IN std_logic ;
         window_22_13 : IN std_logic ;
         window_22_12 : IN std_logic ;
         window_22_11 : IN std_logic ;
         window_22_10 : IN std_logic ;
         window_22_9 : IN std_logic ;
         window_22_8 : IN std_logic ;
         window_22_7 : IN std_logic ;
         window_22_6 : IN std_logic ;
         window_22_5 : IN std_logic ;
         window_22_4 : IN std_logic ;
         window_22_3 : IN std_logic ;
         window_22_2 : IN std_logic ;
         window_22_1 : IN std_logic ;
         window_22_0 : IN std_logic ;
         window_21_15 : IN std_logic ;
         window_21_14 : IN std_logic ;
         window_21_13 : IN std_logic ;
         window_21_12 : IN std_logic ;
         window_21_11 : IN std_logic ;
         window_21_10 : IN std_logic ;
         window_21_9 : IN std_logic ;
         window_21_8 : IN std_logic ;
         window_21_7 : IN std_logic ;
         window_21_6 : IN std_logic ;
         window_21_5 : IN std_logic ;
         window_21_4 : IN std_logic ;
         window_21_3 : IN std_logic ;
         window_21_2 : IN std_logic ;
         window_21_1 : IN std_logic ;
         window_21_0 : IN std_logic ;
         window_20_15 : IN std_logic ;
         window_20_14 : IN std_logic ;
         window_20_13 : IN std_logic ;
         window_20_12 : IN std_logic ;
         window_20_11 : IN std_logic ;
         window_20_10 : IN std_logic ;
         window_20_9 : IN std_logic ;
         window_20_8 : IN std_logic ;
         window_20_7 : IN std_logic ;
         window_20_6 : IN std_logic ;
         window_20_5 : IN std_logic ;
         window_20_4 : IN std_logic ;
         window_20_3 : IN std_logic ;
         window_20_2 : IN std_logic ;
         window_20_1 : IN std_logic ;
         window_20_0 : IN std_logic ;
         window_19_15 : IN std_logic ;
         window_19_14 : IN std_logic ;
         window_19_13 : IN std_logic ;
         window_19_12 : IN std_logic ;
         window_19_11 : IN std_logic ;
         window_19_10 : IN std_logic ;
         window_19_9 : IN std_logic ;
         window_19_8 : IN std_logic ;
         window_19_7 : IN std_logic ;
         window_19_6 : IN std_logic ;
         window_19_5 : IN std_logic ;
         window_19_4 : IN std_logic ;
         window_19_3 : IN std_logic ;
         window_19_2 : IN std_logic ;
         window_19_1 : IN std_logic ;
         window_19_0 : IN std_logic ;
         window_18_15 : IN std_logic ;
         window_18_14 : IN std_logic ;
         window_18_13 : IN std_logic ;
         window_18_12 : IN std_logic ;
         window_18_11 : IN std_logic ;
         window_18_10 : IN std_logic ;
         window_18_9 : IN std_logic ;
         window_18_8 : IN std_logic ;
         window_18_7 : IN std_logic ;
         window_18_6 : IN std_logic ;
         window_18_5 : IN std_logic ;
         window_18_4 : IN std_logic ;
         window_18_3 : IN std_logic ;
         window_18_2 : IN std_logic ;
         window_18_1 : IN std_logic ;
         window_18_0 : IN std_logic ;
         window_17_15 : IN std_logic ;
         window_17_14 : IN std_logic ;
         window_17_13 : IN std_logic ;
         window_17_12 : IN std_logic ;
         window_17_11 : IN std_logic ;
         window_17_10 : IN std_logic ;
         window_17_9 : IN std_logic ;
         window_17_8 : IN std_logic ;
         window_17_7 : IN std_logic ;
         window_17_6 : IN std_logic ;
         window_17_5 : IN std_logic ;
         window_17_4 : IN std_logic ;
         window_17_3 : IN std_logic ;
         window_17_2 : IN std_logic ;
         window_17_1 : IN std_logic ;
         window_17_0 : IN std_logic ;
         window_16_15 : IN std_logic ;
         window_16_14 : IN std_logic ;
         window_16_13 : IN std_logic ;
         window_16_12 : IN std_logic ;
         window_16_11 : IN std_logic ;
         window_16_10 : IN std_logic ;
         window_16_9 : IN std_logic ;
         window_16_8 : IN std_logic ;
         window_16_7 : IN std_logic ;
         window_16_6 : IN std_logic ;
         window_16_5 : IN std_logic ;
         window_16_4 : IN std_logic ;
         window_16_3 : IN std_logic ;
         window_16_2 : IN std_logic ;
         window_16_1 : IN std_logic ;
         window_16_0 : IN std_logic ;
         window_15_15 : IN std_logic ;
         window_15_14 : IN std_logic ;
         window_15_13 : IN std_logic ;
         window_15_12 : IN std_logic ;
         window_15_11 : IN std_logic ;
         window_15_10 : IN std_logic ;
         window_15_9 : IN std_logic ;
         window_15_8 : IN std_logic ;
         window_15_7 : IN std_logic ;
         window_15_6 : IN std_logic ;
         window_15_5 : IN std_logic ;
         window_15_4 : IN std_logic ;
         window_15_3 : IN std_logic ;
         window_15_2 : IN std_logic ;
         window_15_1 : IN std_logic ;
         window_15_0 : IN std_logic ;
         window_14_15 : IN std_logic ;
         window_14_14 : IN std_logic ;
         window_14_13 : IN std_logic ;
         window_14_12 : IN std_logic ;
         window_14_11 : IN std_logic ;
         window_14_10 : IN std_logic ;
         window_14_9 : IN std_logic ;
         window_14_8 : IN std_logic ;
         window_14_7 : IN std_logic ;
         window_14_6 : IN std_logic ;
         window_14_5 : IN std_logic ;
         window_14_4 : IN std_logic ;
         window_14_3 : IN std_logic ;
         window_14_2 : IN std_logic ;
         window_14_1 : IN std_logic ;
         window_14_0 : IN std_logic ;
         window_13_15 : IN std_logic ;
         window_13_14 : IN std_logic ;
         window_13_13 : IN std_logic ;
         window_13_12 : IN std_logic ;
         window_13_11 : IN std_logic ;
         window_13_10 : IN std_logic ;
         window_13_9 : IN std_logic ;
         window_13_8 : IN std_logic ;
         window_13_7 : IN std_logic ;
         window_13_6 : IN std_logic ;
         window_13_5 : IN std_logic ;
         window_13_4 : IN std_logic ;
         window_13_3 : IN std_logic ;
         window_13_2 : IN std_logic ;
         window_13_1 : IN std_logic ;
         window_13_0 : IN std_logic ;
         window_12_15 : IN std_logic ;
         window_12_14 : IN std_logic ;
         window_12_13 : IN std_logic ;
         window_12_12 : IN std_logic ;
         window_12_11 : IN std_logic ;
         window_12_10 : IN std_logic ;
         window_12_9 : IN std_logic ;
         window_12_8 : IN std_logic ;
         window_12_7 : IN std_logic ;
         window_12_6 : IN std_logic ;
         window_12_5 : IN std_logic ;
         window_12_4 : IN std_logic ;
         window_12_3 : IN std_logic ;
         window_12_2 : IN std_logic ;
         window_12_1 : IN std_logic ;
         window_12_0 : IN std_logic ;
         window_11_15 : IN std_logic ;
         window_11_14 : IN std_logic ;
         window_11_13 : IN std_logic ;
         window_11_12 : IN std_logic ;
         window_11_11 : IN std_logic ;
         window_11_10 : IN std_logic ;
         window_11_9 : IN std_logic ;
         window_11_8 : IN std_logic ;
         window_11_7 : IN std_logic ;
         window_11_6 : IN std_logic ;
         window_11_5 : IN std_logic ;
         window_11_4 : IN std_logic ;
         window_11_3 : IN std_logic ;
         window_11_2 : IN std_logic ;
         window_11_1 : IN std_logic ;
         window_11_0 : IN std_logic ;
         window_10_15 : IN std_logic ;
         window_10_14 : IN std_logic ;
         window_10_13 : IN std_logic ;
         window_10_12 : IN std_logic ;
         window_10_11 : IN std_logic ;
         window_10_10 : IN std_logic ;
         window_10_9 : IN std_logic ;
         window_10_8 : IN std_logic ;
         window_10_7 : IN std_logic ;
         window_10_6 : IN std_logic ;
         window_10_5 : IN std_logic ;
         window_10_4 : IN std_logic ;
         window_10_3 : IN std_logic ;
         window_10_2 : IN std_logic ;
         window_10_1 : IN std_logic ;
         window_10_0 : IN std_logic ;
         window_9_15 : IN std_logic ;
         window_9_14 : IN std_logic ;
         window_9_13 : IN std_logic ;
         window_9_12 : IN std_logic ;
         window_9_11 : IN std_logic ;
         window_9_10 : IN std_logic ;
         window_9_9 : IN std_logic ;
         window_9_8 : IN std_logic ;
         window_9_7 : IN std_logic ;
         window_9_6 : IN std_logic ;
         window_9_5 : IN std_logic ;
         window_9_4 : IN std_logic ;
         window_9_3 : IN std_logic ;
         window_9_2 : IN std_logic ;
         window_9_1 : IN std_logic ;
         window_9_0 : IN std_logic ;
         window_8_15 : IN std_logic ;
         window_8_14 : IN std_logic ;
         window_8_13 : IN std_logic ;
         window_8_12 : IN std_logic ;
         window_8_11 : IN std_logic ;
         window_8_10 : IN std_logic ;
         window_8_9 : IN std_logic ;
         window_8_8 : IN std_logic ;
         window_8_7 : IN std_logic ;
         window_8_6 : IN std_logic ;
         window_8_5 : IN std_logic ;
         window_8_4 : IN std_logic ;
         window_8_3 : IN std_logic ;
         window_8_2 : IN std_logic ;
         window_8_1 : IN std_logic ;
         window_8_0 : IN std_logic ;
         window_7_15 : IN std_logic ;
         window_7_14 : IN std_logic ;
         window_7_13 : IN std_logic ;
         window_7_12 : IN std_logic ;
         window_7_11 : IN std_logic ;
         window_7_10 : IN std_logic ;
         window_7_9 : IN std_logic ;
         window_7_8 : IN std_logic ;
         window_7_7 : IN std_logic ;
         window_7_6 : IN std_logic ;
         window_7_5 : IN std_logic ;
         window_7_4 : IN std_logic ;
         window_7_3 : IN std_logic ;
         window_7_2 : IN std_logic ;
         window_7_1 : IN std_logic ;
         window_7_0 : IN std_logic ;
         window_6_15 : IN std_logic ;
         window_6_14 : IN std_logic ;
         window_6_13 : IN std_logic ;
         window_6_12 : IN std_logic ;
         window_6_11 : IN std_logic ;
         window_6_10 : IN std_logic ;
         window_6_9 : IN std_logic ;
         window_6_8 : IN std_logic ;
         window_6_7 : IN std_logic ;
         window_6_6 : IN std_logic ;
         window_6_5 : IN std_logic ;
         window_6_4 : IN std_logic ;
         window_6_3 : IN std_logic ;
         window_6_2 : IN std_logic ;
         window_6_1 : IN std_logic ;
         window_6_0 : IN std_logic ;
         window_5_15 : IN std_logic ;
         window_5_14 : IN std_logic ;
         window_5_13 : IN std_logic ;
         window_5_12 : IN std_logic ;
         window_5_11 : IN std_logic ;
         window_5_10 : IN std_logic ;
         window_5_9 : IN std_logic ;
         window_5_8 : IN std_logic ;
         window_5_7 : IN std_logic ;
         window_5_6 : IN std_logic ;
         window_5_5 : IN std_logic ;
         window_5_4 : IN std_logic ;
         window_5_3 : IN std_logic ;
         window_5_2 : IN std_logic ;
         window_5_1 : IN std_logic ;
         window_5_0 : IN std_logic ;
         window_4_15 : IN std_logic ;
         window_4_14 : IN std_logic ;
         window_4_13 : IN std_logic ;
         window_4_12 : IN std_logic ;
         window_4_11 : IN std_logic ;
         window_4_10 : IN std_logic ;
         window_4_9 : IN std_logic ;
         window_4_8 : IN std_logic ;
         window_4_7 : IN std_logic ;
         window_4_6 : IN std_logic ;
         window_4_5 : IN std_logic ;
         window_4_4 : IN std_logic ;
         window_4_3 : IN std_logic ;
         window_4_2 : IN std_logic ;
         window_4_1 : IN std_logic ;
         window_4_0 : IN std_logic ;
         window_3_15 : IN std_logic ;
         window_3_14 : IN std_logic ;
         window_3_13 : IN std_logic ;
         window_3_12 : IN std_logic ;
         window_3_11 : IN std_logic ;
         window_3_10 : IN std_logic ;
         window_3_9 : IN std_logic ;
         window_3_8 : IN std_logic ;
         window_3_7 : IN std_logic ;
         window_3_6 : IN std_logic ;
         window_3_5 : IN std_logic ;
         window_3_4 : IN std_logic ;
         window_3_3 : IN std_logic ;
         window_3_2 : IN std_logic ;
         window_3_1 : IN std_logic ;
         window_3_0 : IN std_logic ;
         window_2_15 : IN std_logic ;
         window_2_14 : IN std_logic ;
         window_2_13 : IN std_logic ;
         window_2_12 : IN std_logic ;
         window_2_11 : IN std_logic ;
         window_2_10 : IN std_logic ;
         window_2_9 : IN std_logic ;
         window_2_8 : IN std_logic ;
         window_2_7 : IN std_logic ;
         window_2_6 : IN std_logic ;
         window_2_5 : IN std_logic ;
         window_2_4 : IN std_logic ;
         window_2_3 : IN std_logic ;
         window_2_2 : IN std_logic ;
         window_2_1 : IN std_logic ;
         window_2_0 : IN std_logic ;
         window_1_15 : IN std_logic ;
         window_1_14 : IN std_logic ;
         window_1_13 : IN std_logic ;
         window_1_12 : IN std_logic ;
         window_1_11 : IN std_logic ;
         window_1_10 : IN std_logic ;
         window_1_9 : IN std_logic ;
         window_1_8 : IN std_logic ;
         window_1_7 : IN std_logic ;
         window_1_6 : IN std_logic ;
         window_1_5 : IN std_logic ;
         window_1_4 : IN std_logic ;
         window_1_3 : IN std_logic ;
         window_1_2 : IN std_logic ;
         window_1_1 : IN std_logic ;
         window_1_0 : IN std_logic ;
         window_0_15 : IN std_logic ;
         window_0_14 : IN std_logic ;
         window_0_13 : IN std_logic ;
         window_0_12 : IN std_logic ;
         window_0_11 : IN std_logic ;
         window_0_10 : IN std_logic ;
         window_0_9 : IN std_logic ;
         window_0_8 : IN std_logic ;
         window_0_7 : IN std_logic ;
         window_0_6 : IN std_logic ;
         window_0_5 : IN std_logic ;
         window_0_4 : IN std_logic ;
         window_0_3 : IN std_logic ;
         window_0_2 : IN std_logic ;
         window_0_1 : IN std_logic ;
         window_0_0 : IN std_logic ;
         outputs_24_15 : INOUT std_logic ;
         outputs_24_14 : INOUT std_logic ;
         outputs_24_13 : INOUT std_logic ;
         outputs_24_12 : INOUT std_logic ;
         outputs_24_11 : INOUT std_logic ;
         outputs_24_10 : INOUT std_logic ;
         outputs_24_9 : INOUT std_logic ;
         outputs_24_8 : INOUT std_logic ;
         outputs_24_7 : INOUT std_logic ;
         outputs_24_6 : INOUT std_logic ;
         outputs_24_5 : INOUT std_logic ;
         outputs_24_4 : INOUT std_logic ;
         outputs_24_3 : INOUT std_logic ;
         outputs_24_2 : INOUT std_logic ;
         outputs_24_1 : INOUT std_logic ;
         outputs_24_0 : INOUT std_logic ;
         outputs_23_15 : INOUT std_logic ;
         outputs_23_14 : INOUT std_logic ;
         outputs_23_13 : INOUT std_logic ;
         outputs_23_12 : INOUT std_logic ;
         outputs_23_11 : INOUT std_logic ;
         outputs_23_10 : INOUT std_logic ;
         outputs_23_9 : INOUT std_logic ;
         outputs_23_8 : INOUT std_logic ;
         outputs_23_7 : INOUT std_logic ;
         outputs_23_6 : INOUT std_logic ;
         outputs_23_5 : INOUT std_logic ;
         outputs_23_4 : INOUT std_logic ;
         outputs_23_3 : INOUT std_logic ;
         outputs_23_2 : INOUT std_logic ;
         outputs_23_1 : INOUT std_logic ;
         outputs_23_0 : INOUT std_logic ;
         outputs_22_15 : INOUT std_logic ;
         outputs_22_14 : INOUT std_logic ;
         outputs_22_13 : INOUT std_logic ;
         outputs_22_12 : INOUT std_logic ;
         outputs_22_11 : INOUT std_logic ;
         outputs_22_10 : INOUT std_logic ;
         outputs_22_9 : INOUT std_logic ;
         outputs_22_8 : INOUT std_logic ;
         outputs_22_7 : INOUT std_logic ;
         outputs_22_6 : INOUT std_logic ;
         outputs_22_5 : INOUT std_logic ;
         outputs_22_4 : INOUT std_logic ;
         outputs_22_3 : INOUT std_logic ;
         outputs_22_2 : INOUT std_logic ;
         outputs_22_1 : INOUT std_logic ;
         outputs_22_0 : INOUT std_logic ;
         outputs_21_15 : INOUT std_logic ;
         outputs_21_14 : INOUT std_logic ;
         outputs_21_13 : INOUT std_logic ;
         outputs_21_12 : INOUT std_logic ;
         outputs_21_11 : INOUT std_logic ;
         outputs_21_10 : INOUT std_logic ;
         outputs_21_9 : INOUT std_logic ;
         outputs_21_8 : INOUT std_logic ;
         outputs_21_7 : INOUT std_logic ;
         outputs_21_6 : INOUT std_logic ;
         outputs_21_5 : INOUT std_logic ;
         outputs_21_4 : INOUT std_logic ;
         outputs_21_3 : INOUT std_logic ;
         outputs_21_2 : INOUT std_logic ;
         outputs_21_1 : INOUT std_logic ;
         outputs_21_0 : INOUT std_logic ;
         outputs_20_15 : INOUT std_logic ;
         outputs_20_14 : INOUT std_logic ;
         outputs_20_13 : INOUT std_logic ;
         outputs_20_12 : INOUT std_logic ;
         outputs_20_11 : INOUT std_logic ;
         outputs_20_10 : INOUT std_logic ;
         outputs_20_9 : INOUT std_logic ;
         outputs_20_8 : INOUT std_logic ;
         outputs_20_7 : INOUT std_logic ;
         outputs_20_6 : INOUT std_logic ;
         outputs_20_5 : INOUT std_logic ;
         outputs_20_4 : INOUT std_logic ;
         outputs_20_3 : INOUT std_logic ;
         outputs_20_2 : INOUT std_logic ;
         outputs_20_1 : INOUT std_logic ;
         outputs_20_0 : INOUT std_logic ;
         outputs_19_15 : INOUT std_logic ;
         outputs_19_14 : INOUT std_logic ;
         outputs_19_13 : INOUT std_logic ;
         outputs_19_12 : INOUT std_logic ;
         outputs_19_11 : INOUT std_logic ;
         outputs_19_10 : INOUT std_logic ;
         outputs_19_9 : INOUT std_logic ;
         outputs_19_8 : INOUT std_logic ;
         outputs_19_7 : INOUT std_logic ;
         outputs_19_6 : INOUT std_logic ;
         outputs_19_5 : INOUT std_logic ;
         outputs_19_4 : INOUT std_logic ;
         outputs_19_3 : INOUT std_logic ;
         outputs_19_2 : INOUT std_logic ;
         outputs_19_1 : INOUT std_logic ;
         outputs_19_0 : INOUT std_logic ;
         outputs_18_15 : INOUT std_logic ;
         outputs_18_14 : INOUT std_logic ;
         outputs_18_13 : INOUT std_logic ;
         outputs_18_12 : INOUT std_logic ;
         outputs_18_11 : INOUT std_logic ;
         outputs_18_10 : INOUT std_logic ;
         outputs_18_9 : INOUT std_logic ;
         outputs_18_8 : INOUT std_logic ;
         outputs_18_7 : INOUT std_logic ;
         outputs_18_6 : INOUT std_logic ;
         outputs_18_5 : INOUT std_logic ;
         outputs_18_4 : INOUT std_logic ;
         outputs_18_3 : INOUT std_logic ;
         outputs_18_2 : INOUT std_logic ;
         outputs_18_1 : INOUT std_logic ;
         outputs_18_0 : INOUT std_logic ;
         outputs_17_15 : INOUT std_logic ;
         outputs_17_14 : INOUT std_logic ;
         outputs_17_13 : INOUT std_logic ;
         outputs_17_12 : INOUT std_logic ;
         outputs_17_11 : INOUT std_logic ;
         outputs_17_10 : INOUT std_logic ;
         outputs_17_9 : INOUT std_logic ;
         outputs_17_8 : INOUT std_logic ;
         outputs_17_7 : INOUT std_logic ;
         outputs_17_6 : INOUT std_logic ;
         outputs_17_5 : INOUT std_logic ;
         outputs_17_4 : INOUT std_logic ;
         outputs_17_3 : INOUT std_logic ;
         outputs_17_2 : INOUT std_logic ;
         outputs_17_1 : INOUT std_logic ;
         outputs_17_0 : INOUT std_logic ;
         outputs_16_15 : INOUT std_logic ;
         outputs_16_14 : INOUT std_logic ;
         outputs_16_13 : INOUT std_logic ;
         outputs_16_12 : INOUT std_logic ;
         outputs_16_11 : INOUT std_logic ;
         outputs_16_10 : INOUT std_logic ;
         outputs_16_9 : INOUT std_logic ;
         outputs_16_8 : INOUT std_logic ;
         outputs_16_7 : INOUT std_logic ;
         outputs_16_6 : INOUT std_logic ;
         outputs_16_5 : INOUT std_logic ;
         outputs_16_4 : INOUT std_logic ;
         outputs_16_3 : INOUT std_logic ;
         outputs_16_2 : INOUT std_logic ;
         outputs_16_1 : INOUT std_logic ;
         outputs_16_0 : INOUT std_logic ;
         outputs_15_15 : INOUT std_logic ;
         outputs_15_14 : INOUT std_logic ;
         outputs_15_13 : INOUT std_logic ;
         outputs_15_12 : INOUT std_logic ;
         outputs_15_11 : INOUT std_logic ;
         outputs_15_10 : INOUT std_logic ;
         outputs_15_9 : INOUT std_logic ;
         outputs_15_8 : INOUT std_logic ;
         outputs_15_7 : INOUT std_logic ;
         outputs_15_6 : INOUT std_logic ;
         outputs_15_5 : INOUT std_logic ;
         outputs_15_4 : INOUT std_logic ;
         outputs_15_3 : INOUT std_logic ;
         outputs_15_2 : INOUT std_logic ;
         outputs_15_1 : INOUT std_logic ;
         outputs_15_0 : INOUT std_logic ;
         outputs_14_15 : INOUT std_logic ;
         outputs_14_14 : INOUT std_logic ;
         outputs_14_13 : INOUT std_logic ;
         outputs_14_12 : INOUT std_logic ;
         outputs_14_11 : INOUT std_logic ;
         outputs_14_10 : INOUT std_logic ;
         outputs_14_9 : INOUT std_logic ;
         outputs_14_8 : INOUT std_logic ;
         outputs_14_7 : INOUT std_logic ;
         outputs_14_6 : INOUT std_logic ;
         outputs_14_5 : INOUT std_logic ;
         outputs_14_4 : INOUT std_logic ;
         outputs_14_3 : INOUT std_logic ;
         outputs_14_2 : INOUT std_logic ;
         outputs_14_1 : INOUT std_logic ;
         outputs_14_0 : INOUT std_logic ;
         outputs_13_15 : INOUT std_logic ;
         outputs_13_14 : INOUT std_logic ;
         outputs_13_13 : INOUT std_logic ;
         outputs_13_12 : INOUT std_logic ;
         outputs_13_11 : INOUT std_logic ;
         outputs_13_10 : INOUT std_logic ;
         outputs_13_9 : INOUT std_logic ;
         outputs_13_8 : INOUT std_logic ;
         outputs_13_7 : INOUT std_logic ;
         outputs_13_6 : INOUT std_logic ;
         outputs_13_5 : INOUT std_logic ;
         outputs_13_4 : INOUT std_logic ;
         outputs_13_3 : INOUT std_logic ;
         outputs_13_2 : INOUT std_logic ;
         outputs_13_1 : INOUT std_logic ;
         outputs_13_0 : INOUT std_logic ;
         outputs_12_15 : INOUT std_logic ;
         outputs_12_14 : INOUT std_logic ;
         outputs_12_13 : INOUT std_logic ;
         outputs_12_12 : INOUT std_logic ;
         outputs_12_11 : INOUT std_logic ;
         outputs_12_10 : INOUT std_logic ;
         outputs_12_9 : INOUT std_logic ;
         outputs_12_8 : INOUT std_logic ;
         outputs_12_7 : INOUT std_logic ;
         outputs_12_6 : INOUT std_logic ;
         outputs_12_5 : INOUT std_logic ;
         outputs_12_4 : INOUT std_logic ;
         outputs_12_3 : INOUT std_logic ;
         outputs_12_2 : INOUT std_logic ;
         outputs_12_1 : INOUT std_logic ;
         outputs_12_0 : INOUT std_logic ;
         outputs_11_15 : INOUT std_logic ;
         outputs_11_14 : INOUT std_logic ;
         outputs_11_13 : INOUT std_logic ;
         outputs_11_12 : INOUT std_logic ;
         outputs_11_11 : INOUT std_logic ;
         outputs_11_10 : INOUT std_logic ;
         outputs_11_9 : INOUT std_logic ;
         outputs_11_8 : INOUT std_logic ;
         outputs_11_7 : INOUT std_logic ;
         outputs_11_6 : INOUT std_logic ;
         outputs_11_5 : INOUT std_logic ;
         outputs_11_4 : INOUT std_logic ;
         outputs_11_3 : INOUT std_logic ;
         outputs_11_2 : INOUT std_logic ;
         outputs_11_1 : INOUT std_logic ;
         outputs_11_0 : INOUT std_logic ;
         outputs_10_15 : INOUT std_logic ;
         outputs_10_14 : INOUT std_logic ;
         outputs_10_13 : INOUT std_logic ;
         outputs_10_12 : INOUT std_logic ;
         outputs_10_11 : INOUT std_logic ;
         outputs_10_10 : INOUT std_logic ;
         outputs_10_9 : INOUT std_logic ;
         outputs_10_8 : INOUT std_logic ;
         outputs_10_7 : INOUT std_logic ;
         outputs_10_6 : INOUT std_logic ;
         outputs_10_5 : INOUT std_logic ;
         outputs_10_4 : INOUT std_logic ;
         outputs_10_3 : INOUT std_logic ;
         outputs_10_2 : INOUT std_logic ;
         outputs_10_1 : INOUT std_logic ;
         outputs_10_0 : INOUT std_logic ;
         outputs_9_15 : INOUT std_logic ;
         outputs_9_14 : INOUT std_logic ;
         outputs_9_13 : INOUT std_logic ;
         outputs_9_12 : INOUT std_logic ;
         outputs_9_11 : INOUT std_logic ;
         outputs_9_10 : INOUT std_logic ;
         outputs_9_9 : INOUT std_logic ;
         outputs_9_8 : INOUT std_logic ;
         outputs_9_7 : INOUT std_logic ;
         outputs_9_6 : INOUT std_logic ;
         outputs_9_5 : INOUT std_logic ;
         outputs_9_4 : INOUT std_logic ;
         outputs_9_3 : INOUT std_logic ;
         outputs_9_2 : INOUT std_logic ;
         outputs_9_1 : INOUT std_logic ;
         outputs_9_0 : INOUT std_logic ;
         outputs_8_15 : INOUT std_logic ;
         outputs_8_14 : INOUT std_logic ;
         outputs_8_13 : INOUT std_logic ;
         outputs_8_12 : INOUT std_logic ;
         outputs_8_11 : INOUT std_logic ;
         outputs_8_10 : INOUT std_logic ;
         outputs_8_9 : INOUT std_logic ;
         outputs_8_8 : INOUT std_logic ;
         outputs_8_7 : INOUT std_logic ;
         outputs_8_6 : INOUT std_logic ;
         outputs_8_5 : INOUT std_logic ;
         outputs_8_4 : INOUT std_logic ;
         outputs_8_3 : INOUT std_logic ;
         outputs_8_2 : INOUT std_logic ;
         outputs_8_1 : INOUT std_logic ;
         outputs_8_0 : INOUT std_logic ;
         outputs_7_15 : INOUT std_logic ;
         outputs_7_14 : INOUT std_logic ;
         outputs_7_13 : INOUT std_logic ;
         outputs_7_12 : INOUT std_logic ;
         outputs_7_11 : INOUT std_logic ;
         outputs_7_10 : INOUT std_logic ;
         outputs_7_9 : INOUT std_logic ;
         outputs_7_8 : INOUT std_logic ;
         outputs_7_7 : INOUT std_logic ;
         outputs_7_6 : INOUT std_logic ;
         outputs_7_5 : INOUT std_logic ;
         outputs_7_4 : INOUT std_logic ;
         outputs_7_3 : INOUT std_logic ;
         outputs_7_2 : INOUT std_logic ;
         outputs_7_1 : INOUT std_logic ;
         outputs_7_0 : INOUT std_logic ;
         outputs_6_15 : INOUT std_logic ;
         outputs_6_14 : INOUT std_logic ;
         outputs_6_13 : INOUT std_logic ;
         outputs_6_12 : INOUT std_logic ;
         outputs_6_11 : INOUT std_logic ;
         outputs_6_10 : INOUT std_logic ;
         outputs_6_9 : INOUT std_logic ;
         outputs_6_8 : INOUT std_logic ;
         outputs_6_7 : INOUT std_logic ;
         outputs_6_6 : INOUT std_logic ;
         outputs_6_5 : INOUT std_logic ;
         outputs_6_4 : INOUT std_logic ;
         outputs_6_3 : INOUT std_logic ;
         outputs_6_2 : INOUT std_logic ;
         outputs_6_1 : INOUT std_logic ;
         outputs_6_0 : INOUT std_logic ;
         outputs_5_15 : INOUT std_logic ;
         outputs_5_14 : INOUT std_logic ;
         outputs_5_13 : INOUT std_logic ;
         outputs_5_12 : INOUT std_logic ;
         outputs_5_11 : INOUT std_logic ;
         outputs_5_10 : INOUT std_logic ;
         outputs_5_9 : INOUT std_logic ;
         outputs_5_8 : INOUT std_logic ;
         outputs_5_7 : INOUT std_logic ;
         outputs_5_6 : INOUT std_logic ;
         outputs_5_5 : INOUT std_logic ;
         outputs_5_4 : INOUT std_logic ;
         outputs_5_3 : INOUT std_logic ;
         outputs_5_2 : INOUT std_logic ;
         outputs_5_1 : INOUT std_logic ;
         outputs_5_0 : INOUT std_logic ;
         outputs_4_15 : INOUT std_logic ;
         outputs_4_14 : INOUT std_logic ;
         outputs_4_13 : INOUT std_logic ;
         outputs_4_12 : INOUT std_logic ;
         outputs_4_11 : INOUT std_logic ;
         outputs_4_10 : INOUT std_logic ;
         outputs_4_9 : INOUT std_logic ;
         outputs_4_8 : INOUT std_logic ;
         outputs_4_7 : INOUT std_logic ;
         outputs_4_6 : INOUT std_logic ;
         outputs_4_5 : INOUT std_logic ;
         outputs_4_4 : INOUT std_logic ;
         outputs_4_3 : INOUT std_logic ;
         outputs_4_2 : INOUT std_logic ;
         outputs_4_1 : INOUT std_logic ;
         outputs_4_0 : INOUT std_logic ;
         outputs_3_15 : INOUT std_logic ;
         outputs_3_14 : INOUT std_logic ;
         outputs_3_13 : INOUT std_logic ;
         outputs_3_12 : INOUT std_logic ;
         outputs_3_11 : INOUT std_logic ;
         outputs_3_10 : INOUT std_logic ;
         outputs_3_9 : INOUT std_logic ;
         outputs_3_8 : INOUT std_logic ;
         outputs_3_7 : INOUT std_logic ;
         outputs_3_6 : INOUT std_logic ;
         outputs_3_5 : INOUT std_logic ;
         outputs_3_4 : INOUT std_logic ;
         outputs_3_3 : INOUT std_logic ;
         outputs_3_2 : INOUT std_logic ;
         outputs_3_1 : INOUT std_logic ;
         outputs_3_0 : INOUT std_logic ;
         outputs_2_15 : INOUT std_logic ;
         outputs_2_14 : INOUT std_logic ;
         outputs_2_13 : INOUT std_logic ;
         outputs_2_12 : INOUT std_logic ;
         outputs_2_11 : INOUT std_logic ;
         outputs_2_10 : INOUT std_logic ;
         outputs_2_9 : INOUT std_logic ;
         outputs_2_8 : INOUT std_logic ;
         outputs_2_7 : INOUT std_logic ;
         outputs_2_6 : INOUT std_logic ;
         outputs_2_5 : INOUT std_logic ;
         outputs_2_4 : INOUT std_logic ;
         outputs_2_3 : INOUT std_logic ;
         outputs_2_2 : INOUT std_logic ;
         outputs_2_1 : INOUT std_logic ;
         outputs_2_0 : INOUT std_logic ;
         outputs_1_15 : INOUT std_logic ;
         outputs_1_14 : INOUT std_logic ;
         outputs_1_13 : INOUT std_logic ;
         outputs_1_12 : INOUT std_logic ;
         outputs_1_11 : INOUT std_logic ;
         outputs_1_10 : INOUT std_logic ;
         outputs_1_9 : INOUT std_logic ;
         outputs_1_8 : INOUT std_logic ;
         outputs_1_7 : INOUT std_logic ;
         outputs_1_6 : INOUT std_logic ;
         outputs_1_5 : INOUT std_logic ;
         outputs_1_4 : INOUT std_logic ;
         outputs_1_3 : INOUT std_logic ;
         outputs_1_2 : INOUT std_logic ;
         outputs_1_1 : INOUT std_logic ;
         outputs_1_0 : INOUT std_logic ;
         outputs_0_15 : INOUT std_logic ;
         outputs_0_14 : INOUT std_logic ;
         outputs_0_13 : INOUT std_logic ;
         outputs_0_12 : INOUT std_logic ;
         outputs_0_11 : INOUT std_logic ;
         outputs_0_10 : INOUT std_logic ;
         outputs_0_9 : INOUT std_logic ;
         outputs_0_8 : INOUT std_logic ;
         outputs_0_7 : INOUT std_logic ;
         outputs_0_6 : INOUT std_logic ;
         outputs_0_5 : INOUT std_logic ;
         outputs_0_4 : INOUT std_logic ;
         outputs_0_3 : INOUT std_logic ;
         outputs_0_2 : INOUT std_logic ;
         outputs_0_1 : INOUT std_logic ;
         outputs_0_0 : INOUT std_logic ;
         clk : IN std_logic ;
         start : IN std_logic ;
         rst : IN std_logic ;
         done : INOUT std_logic ;
         working : INOUT std_logic) ;
   end component ;
   component RegUnit_8_16
      port (
         filterBus : IN std_logic_vector (7 DOWNTO 0) ;
         windowBus : IN std_logic_vector (15 DOWNTO 0) ;
         regPage1NextUnit : IN std_logic_vector (15 DOWNTO 0) ;
         regPage2NextUnit : IN std_logic_vector (15 DOWNTO 0) ;
         clk : IN std_logic ;
         rst : IN std_logic ;
         enableRegPage1 : IN std_logic ;
         enableRegPage2 : IN std_logic ;
         enableRegFilter : IN std_logic ;
         page1ReadBusOrPage2 : IN std_logic ;
         page2ReadBusOrPage1 : IN std_logic ;
         pageTurn : IN std_logic ;
         outRegPage : OUT std_logic_vector (15 DOWNTO 0) ;
         outputRegPage1 : OUT std_logic_vector (15 DOWNTO 0) ;
         outputRegPage2 : OUT std_logic_vector (15 DOWNTO 0) ;
         outFilter : OUT std_logic_vector (7 DOWNTO 0)) ;
   end component ;
   component RegUnit_8_16_unfolded2
      port (
         filterBus : IN std_logic_vector (7 DOWNTO 0) ;
         windowBus : IN std_logic_vector (15 DOWNTO 0) ;
         regPage1NextUnit : IN std_logic_vector (15 DOWNTO 0) ;
         regPage2NextUnit : IN std_logic_vector (15 DOWNTO 0) ;
         clk : IN std_logic ;
         rst : IN std_logic ;
         enableRegPage1 : IN std_logic ;
         enableRegPage2 : IN std_logic ;
         enableRegFilter : IN std_logic ;
         page1ReadBusOrPage2 : IN std_logic ;
         page2ReadBusOrPage1 : IN std_logic ;
         pageTurn : IN std_logic ;
         outRegPage : OUT std_logic_vector (15 DOWNTO 0) ;
         outputRegPage1 : OUT std_logic_vector (15 DOWNTO 0) ;
         outputRegPage2 : OUT std_logic_vector (15 DOWNTO 0) ;
         outFilter : OUT std_logic_vector (7 DOWNTO 0)) ;
   end component ;
   component RegUnit_8_16_unfolded3
      port (
         filterBus : IN std_logic_vector (7 DOWNTO 0) ;
         windowBus : IN std_logic_vector (15 DOWNTO 0) ;
         regPage1NextUnit : IN std_logic_vector (15 DOWNTO 0) ;
         regPage2NextUnit : IN std_logic_vector (15 DOWNTO 0) ;
         clk : IN std_logic ;
         rst : IN std_logic ;
         enableRegPage1 : IN std_logic ;
         enableRegPage2 : IN std_logic ;
         enableRegFilter : IN std_logic ;
         page1ReadBusOrPage2 : IN std_logic ;
         page2ReadBusOrPage1 : IN std_logic ;
         pageTurn : IN std_logic ;
         outRegPage : OUT std_logic_vector (15 DOWNTO 0) ;
         outputRegPage1 : OUT std_logic_vector (15 DOWNTO 0) ;
         outputRegPage2 : OUT std_logic_vector (15 DOWNTO 0) ;
         outFilter : OUT std_logic_vector (7 DOWNTO 0)) ;
   end component ;
   component NBitAdder_16
      port (
         a : IN std_logic_vector (15 DOWNTO 0) ;
         b : IN std_logic_vector (15 DOWNTO 0) ;
         carryIn : IN std_logic ;
         sum : OUT std_logic_vector (15 DOWNTO 0) ;
         carryOut : OUT std_logic) ;
   end component ;
   signal currentPage_0_15, currentPage_0_14, currentPage_0_13, 
      currentPage_0_12, currentPage_0_11, currentPage_0_10, currentPage_0_9, 
      currentPage_0_8, currentPage_0_7, currentPage_0_6, currentPage_0_5, 
      currentPage_0_4, currentPage_0_3, currentPage_0_2, currentPage_0_1, 
      currentPage_0_0, currentPage_1_15, currentPage_1_14, currentPage_1_13, 
      currentPage_1_12, currentPage_1_11, currentPage_1_10, currentPage_1_9, 
      currentPage_1_8, currentPage_1_7, currentPage_1_6, currentPage_1_5, 
      currentPage_1_4, currentPage_1_3, currentPage_1_2, currentPage_1_1, 
      currentPage_1_0, currentPage_2_15, currentPage_2_14, currentPage_2_13, 
      currentPage_2_12, currentPage_2_11, currentPage_2_10, currentPage_2_9, 
      currentPage_2_8, currentPage_2_7, currentPage_2_6, currentPage_2_5, 
      currentPage_2_4, currentPage_2_3, currentPage_2_2, currentPage_2_1, 
      currentPage_2_0, currentPage_3_15, currentPage_3_14, currentPage_3_13, 
      currentPage_3_12, currentPage_3_11, currentPage_3_10, currentPage_3_9, 
      currentPage_3_8, currentPage_3_7, currentPage_3_6, currentPage_3_5, 
      currentPage_3_4, currentPage_3_3, currentPage_3_2, currentPage_3_1, 
      currentPage_3_0, currentPage_4_15, currentPage_4_14, currentPage_4_13, 
      currentPage_4_12, currentPage_4_11, currentPage_4_10, currentPage_4_9, 
      currentPage_4_8, currentPage_4_7, currentPage_4_6, currentPage_4_5, 
      currentPage_4_4, currentPage_4_3, currentPage_4_2, currentPage_4_1, 
      currentPage_4_0, currentPage_5_15, currentPage_5_14, currentPage_5_13, 
      currentPage_5_12, currentPage_5_11, currentPage_5_10, currentPage_5_9, 
      currentPage_5_8, currentPage_5_7, currentPage_5_6, currentPage_5_5, 
      currentPage_5_4, currentPage_5_3, currentPage_5_2, currentPage_5_1, 
      currentPage_5_0, currentPage_6_15, currentPage_6_14, currentPage_6_13, 
      currentPage_6_12, currentPage_6_11, currentPage_6_10, currentPage_6_9, 
      currentPage_6_8, currentPage_6_7, currentPage_6_6, currentPage_6_5, 
      currentPage_6_4, currentPage_6_3, currentPage_6_2, currentPage_6_1, 
      currentPage_6_0, currentPage_7_15, currentPage_7_14, currentPage_7_13, 
      currentPage_7_12, currentPage_7_11, currentPage_7_10, currentPage_7_9, 
      currentPage_7_8, currentPage_7_7, currentPage_7_6, currentPage_7_5, 
      currentPage_7_4, currentPage_7_3, currentPage_7_2, currentPage_7_1, 
      currentPage_7_0, currentPage_8_15, currentPage_8_14, currentPage_8_13, 
      currentPage_8_12, currentPage_8_11, currentPage_8_10, currentPage_8_9, 
      currentPage_8_8, currentPage_8_7, currentPage_8_6, currentPage_8_5, 
      currentPage_8_4, currentPage_8_3, currentPage_8_2, currentPage_8_1, 
      currentPage_8_0, currentPage_9_15, currentPage_9_14, currentPage_9_13, 
      currentPage_9_12, currentPage_9_11, currentPage_9_10, currentPage_9_9, 
      currentPage_9_8, currentPage_9_7, currentPage_9_6, currentPage_9_5, 
      currentPage_9_4, currentPage_9_3, currentPage_9_2, currentPage_9_1, 
      currentPage_9_0, currentPage_10_15, currentPage_10_14, 
      currentPage_10_13, currentPage_10_12, currentPage_10_11, 
      currentPage_10_10, currentPage_10_9, currentPage_10_8, 
      currentPage_10_7, currentPage_10_6, currentPage_10_5, currentPage_10_4, 
      currentPage_10_3, currentPage_10_2, currentPage_10_1, currentPage_10_0, 
      currentPage_11_15, currentPage_11_14, currentPage_11_13, 
      currentPage_11_12, currentPage_11_11, currentPage_11_10, 
      currentPage_11_9, currentPage_11_8, currentPage_11_7, currentPage_11_6, 
      currentPage_11_5, currentPage_11_4, currentPage_11_3, currentPage_11_2, 
      currentPage_11_1, currentPage_11_0, currentPage_12_15, 
      currentPage_12_14, currentPage_12_13, currentPage_12_12, 
      currentPage_12_11, currentPage_12_10, currentPage_12_9, 
      currentPage_12_8, currentPage_12_7, currentPage_12_6, currentPage_12_5, 
      currentPage_12_4, currentPage_12_3, currentPage_12_2, currentPage_12_1, 
      currentPage_12_0, currentPage_13_15, currentPage_13_14, 
      currentPage_13_13, currentPage_13_12, currentPage_13_11, 
      currentPage_13_10, currentPage_13_9, currentPage_13_8, 
      currentPage_13_7, currentPage_13_6, currentPage_13_5, currentPage_13_4, 
      currentPage_13_3, currentPage_13_2, currentPage_13_1, currentPage_13_0, 
      currentPage_14_15, currentPage_14_14, currentPage_14_13, 
      currentPage_14_12, currentPage_14_11, currentPage_14_10, 
      currentPage_14_9, currentPage_14_8, currentPage_14_7, currentPage_14_6, 
      currentPage_14_5, currentPage_14_4, currentPage_14_3, currentPage_14_2, 
      currentPage_14_1, currentPage_14_0, currentPage_15_15, 
      currentPage_15_14, currentPage_15_13, currentPage_15_12, 
      currentPage_15_11, currentPage_15_10, currentPage_15_9, 
      currentPage_15_8, currentPage_15_7, currentPage_15_6, currentPage_15_5, 
      currentPage_15_4, currentPage_15_3, currentPage_15_2, currentPage_15_1, 
      currentPage_15_0, currentPage_16_15, currentPage_16_14, 
      currentPage_16_13, currentPage_16_12, currentPage_16_11, 
      currentPage_16_10, currentPage_16_9, currentPage_16_8, 
      currentPage_16_7, currentPage_16_6, currentPage_16_5, currentPage_16_4, 
      currentPage_16_3, currentPage_16_2, currentPage_16_1, currentPage_16_0, 
      currentPage_17_15, currentPage_17_14, currentPage_17_13, 
      currentPage_17_12, currentPage_17_11, currentPage_17_10, 
      currentPage_17_9, currentPage_17_8, currentPage_17_7, currentPage_17_6, 
      currentPage_17_5, currentPage_17_4, currentPage_17_3, currentPage_17_2, 
      currentPage_17_1, currentPage_17_0, currentPage_18_15, 
      currentPage_18_14, currentPage_18_13, currentPage_18_12, 
      currentPage_18_11, currentPage_18_10, currentPage_18_9, 
      currentPage_18_8, currentPage_18_7, currentPage_18_6, currentPage_18_5, 
      currentPage_18_4, currentPage_18_3, currentPage_18_2, currentPage_18_1, 
      currentPage_18_0, currentPage_19_15, currentPage_19_14, 
      currentPage_19_13, currentPage_19_12, currentPage_19_11, 
      currentPage_19_10, currentPage_19_9, currentPage_19_8, 
      currentPage_19_7, currentPage_19_6, currentPage_19_5, currentPage_19_4, 
      currentPage_19_3, currentPage_19_2, currentPage_19_1, currentPage_19_0, 
      currentPage_20_15, currentPage_20_14, currentPage_20_13, 
      currentPage_20_12, currentPage_20_11, currentPage_20_10, 
      currentPage_20_9, currentPage_20_8, currentPage_20_7, currentPage_20_6, 
      currentPage_20_5, currentPage_20_4, currentPage_20_3, currentPage_20_2, 
      currentPage_20_1, currentPage_20_0, currentPage_21_15, 
      currentPage_21_14, currentPage_21_13, currentPage_21_12, 
      currentPage_21_11, currentPage_21_10, currentPage_21_9, 
      currentPage_21_8, currentPage_21_7, currentPage_21_6, currentPage_21_5, 
      currentPage_21_4, currentPage_21_3, currentPage_21_2, currentPage_21_1, 
      currentPage_21_0, currentPage_22_15, currentPage_22_14, 
      currentPage_22_13, currentPage_22_12, currentPage_22_11, 
      currentPage_22_10, currentPage_22_9, currentPage_22_8, 
      currentPage_22_7, currentPage_22_6, currentPage_22_5, currentPage_22_4, 
      currentPage_22_3, currentPage_22_2, currentPage_22_1, currentPage_22_0, 
      currentPage_23_15, currentPage_23_14, currentPage_23_13, 
      currentPage_23_12, currentPage_23_11, currentPage_23_10, 
      currentPage_23_9, currentPage_23_8, currentPage_23_7, currentPage_23_6, 
      currentPage_23_5, currentPage_23_4, currentPage_23_3, currentPage_23_2, 
      currentPage_23_1, currentPage_23_0, currentPage_24_15, 
      currentPage_24_14, currentPage_24_13, currentPage_24_12, 
      currentPage_24_11, currentPage_24_10, currentPage_24_9, 
      currentPage_24_8, currentPage_24_7, currentPage_24_6, currentPage_24_5, 
      currentPage_24_4, currentPage_24_3, currentPage_24_2, currentPage_24_1, 
      currentPage_24_0, outMuls_0_15, outMuls_0_14, outMuls_0_13, 
      outMuls_0_12, outMuls_0_11, outMuls_0_10, outMuls_0_9, outMuls_0_8, 
      outMuls_0_7, outMuls_0_6, outMuls_0_5, outMuls_0_4, outMuls_0_3, 
      outMuls_0_2, outMuls_0_1, outMuls_0_0, outMuls_1_15, outMuls_1_14, 
      outMuls_1_13, outMuls_1_12, outMuls_1_11, outMuls_1_10, outMuls_1_9, 
      outMuls_1_8, outMuls_1_7, outMuls_1_6, outMuls_1_5, outMuls_1_4, 
      outMuls_1_3, outMuls_1_2, outMuls_1_1, outMuls_1_0, outMuls_2_15, 
      outMuls_2_14, outMuls_2_13, outMuls_2_12, outMuls_2_11, outMuls_2_10, 
      outMuls_2_9, outMuls_2_8, outMuls_2_7, outMuls_2_6, outMuls_2_5, 
      outMuls_2_4, outMuls_2_3, outMuls_2_2, outMuls_2_1, outMuls_2_0, 
      outMuls_3_15, outMuls_3_14, outMuls_3_13, outMuls_3_12, outMuls_3_11, 
      outMuls_3_10, outMuls_3_9, outMuls_3_8, outMuls_3_7, outMuls_3_6, 
      outMuls_3_5, outMuls_3_4, outMuls_3_3, outMuls_3_2, outMuls_3_1, 
      outMuls_3_0, outMuls_4_15, outMuls_4_14, outMuls_4_13, outMuls_4_12, 
      outMuls_4_11, outMuls_4_10, outMuls_4_9, outMuls_4_8, outMuls_4_7, 
      outMuls_4_6, outMuls_4_5, outMuls_4_4, outMuls_4_3, outMuls_4_2, 
      outMuls_4_1, outMuls_4_0, outMuls_5_15, outMuls_5_14, outMuls_5_13, 
      outMuls_5_12, outMuls_5_11, outMuls_5_10, outMuls_5_9, outMuls_5_8, 
      outMuls_5_7, outMuls_5_6, outMuls_5_5, outMuls_5_4, outMuls_5_3, 
      outMuls_5_2, outMuls_5_1, outMuls_5_0, outMuls_6_15, outMuls_6_14, 
      outMuls_6_13, outMuls_6_12, outMuls_6_11, outMuls_6_10, outMuls_6_9, 
      outMuls_6_8, outMuls_6_7, outMuls_6_6, outMuls_6_5, outMuls_6_4, 
      outMuls_6_3, outMuls_6_2, outMuls_6_1, outMuls_6_0, outMuls_7_15, 
      outMuls_7_14, outMuls_7_13, outMuls_7_12, outMuls_7_11, outMuls_7_10, 
      outMuls_7_9, outMuls_7_8, outMuls_7_7, outMuls_7_6, outMuls_7_5, 
      outMuls_7_4, outMuls_7_3, outMuls_7_2, outMuls_7_1, outMuls_7_0, 
      outMuls_8_15, outMuls_8_14, outMuls_8_13, outMuls_8_12, outMuls_8_11, 
      outMuls_8_10, outMuls_8_9, outMuls_8_8, outMuls_8_7, outMuls_8_6, 
      outMuls_8_5, outMuls_8_4, outMuls_8_3, outMuls_8_2, outMuls_8_1, 
      outMuls_8_0, outMuls_9_15, outMuls_9_14, outMuls_9_13, outMuls_9_12, 
      outMuls_9_11, outMuls_9_10, outMuls_9_9, outMuls_9_8, outMuls_9_7, 
      outMuls_9_6, outMuls_9_5, outMuls_9_4, outMuls_9_3, outMuls_9_2, 
      outMuls_9_1, outMuls_9_0, outMuls_10_15, outMuls_10_14, outMuls_10_13, 
      outMuls_10_12, outMuls_10_11, outMuls_10_10, outMuls_10_9, 
      outMuls_10_8, outMuls_10_7, outMuls_10_6, outMuls_10_5, outMuls_10_4, 
      outMuls_10_3, outMuls_10_2, outMuls_10_1, outMuls_10_0, outMuls_11_15, 
      outMuls_11_14, outMuls_11_13, outMuls_11_12, outMuls_11_11, 
      outMuls_11_10, outMuls_11_9, outMuls_11_8, outMuls_11_7, outMuls_11_6, 
      outMuls_11_5, outMuls_11_4, outMuls_11_3, outMuls_11_2, outMuls_11_1, 
      outMuls_11_0, outMuls_12_15, outMuls_12_14, outMuls_12_13, 
      outMuls_12_12, outMuls_12_11, outMuls_12_10, outMuls_12_9, 
      outMuls_12_8, outMuls_12_7, outMuls_12_6, outMuls_12_5, outMuls_12_4, 
      outMuls_12_3, outMuls_12_2, outMuls_12_1, outMuls_12_0, outMuls_13_15, 
      outMuls_13_14, outMuls_13_13, outMuls_13_12, outMuls_13_11, 
      outMuls_13_10, outMuls_13_9, outMuls_13_8, outMuls_13_7, outMuls_13_6, 
      outMuls_13_5, outMuls_13_4, outMuls_13_3, outMuls_13_2, outMuls_13_1, 
      outMuls_13_0, outMuls_14_15, outMuls_14_14, outMuls_14_13, 
      outMuls_14_12, outMuls_14_11, outMuls_14_10, outMuls_14_9, 
      outMuls_14_8, outMuls_14_7, outMuls_14_6, outMuls_14_5, outMuls_14_4, 
      outMuls_14_3, outMuls_14_2, outMuls_14_1, outMuls_14_0, outMuls_15_15, 
      outMuls_15_14, outMuls_15_13, outMuls_15_12, outMuls_15_11, 
      outMuls_15_10, outMuls_15_9, outMuls_15_8, outMuls_15_7, outMuls_15_6, 
      outMuls_15_5, outMuls_15_4, outMuls_15_3, outMuls_15_2, outMuls_15_1, 
      outMuls_15_0, outMuls_16_15, outMuls_16_14, outMuls_16_13, 
      outMuls_16_12, outMuls_16_11, outMuls_16_10, outMuls_16_9, 
      outMuls_16_8, outMuls_16_7, outMuls_16_6, outMuls_16_5, outMuls_16_4, 
      outMuls_16_3, outMuls_16_2, outMuls_16_1, outMuls_16_0, outMuls_17_15, 
      outMuls_17_14, outMuls_17_13, outMuls_17_12, outMuls_17_11, 
      outMuls_17_10, outMuls_17_9, outMuls_17_8, outMuls_17_7, outMuls_17_6, 
      outMuls_17_5, outMuls_17_4, outMuls_17_3, outMuls_17_2, outMuls_17_1, 
      outMuls_17_0, outMuls_18_15, outMuls_18_14, outMuls_18_13, 
      outMuls_18_12, outMuls_18_11, outMuls_18_10, outMuls_18_9, 
      outMuls_18_8, outMuls_18_7, outMuls_18_6, outMuls_18_5, outMuls_18_4, 
      outMuls_18_3, outMuls_18_2, outMuls_18_1, outMuls_18_0, outMuls_19_15, 
      outMuls_19_14, outMuls_19_13, outMuls_19_12, outMuls_19_11, 
      outMuls_19_10, outMuls_19_9, outMuls_19_8, outMuls_19_7, outMuls_19_6, 
      outMuls_19_5, outMuls_19_4, outMuls_19_3, outMuls_19_2, outMuls_19_1, 
      outMuls_19_0, outMuls_20_15, outMuls_20_14, outMuls_20_13, 
      outMuls_20_12, outMuls_20_11, outMuls_20_10, outMuls_20_9, 
      outMuls_20_8, outMuls_20_7, outMuls_20_6, outMuls_20_5, outMuls_20_4, 
      outMuls_20_3, outMuls_20_2, outMuls_20_1, outMuls_20_0, outMuls_21_15, 
      outMuls_21_14, outMuls_21_13, outMuls_21_12, outMuls_21_11, 
      outMuls_21_10, outMuls_21_9, outMuls_21_8, outMuls_21_7, outMuls_21_6, 
      outMuls_21_5, outMuls_21_4, outMuls_21_3, outMuls_21_2, outMuls_21_1, 
      outMuls_21_0, outMuls_22_15, outMuls_22_14, outMuls_22_13, 
      outMuls_22_12, outMuls_22_11, outMuls_22_10, outMuls_22_9, 
      outMuls_22_8, outMuls_22_7, outMuls_22_6, outMuls_22_5, outMuls_22_4, 
      outMuls_22_3, outMuls_22_2, outMuls_22_1, outMuls_22_0, outMuls_23_15, 
      outMuls_23_14, outMuls_23_13, outMuls_23_12, outMuls_23_11, 
      outMuls_23_10, outMuls_23_9, outMuls_23_8, outMuls_23_7, outMuls_23_6, 
      outMuls_23_5, outMuls_23_4, outMuls_23_3, outMuls_23_2, outMuls_23_1, 
      outMuls_23_0, outMuls_24_15, outMuls_24_14, outMuls_24_13, 
      outMuls_24_12, outMuls_24_11, outMuls_24_10, outMuls_24_9, 
      outMuls_24_8, outMuls_24_7, outMuls_24_6, outMuls_24_5, outMuls_24_4, 
      outMuls_24_3, outMuls_24_2, outMuls_24_1, outMuls_24_0, 
      addersInputs_0_15, addersInputs_0_14, addersInputs_0_13, 
      addersInputs_0_12, addersInputs_0_11, addersInputs_0_10, 
      addersInputs_0_9, addersInputs_0_8, addersInputs_0_7, addersInputs_0_6, 
      addersInputs_0_5, addersInputs_0_4, addersInputs_0_3, addersInputs_0_2, 
      addersInputs_0_1, addersInputs_0_0, addersInputs_1_15, 
      addersInputs_1_14, addersInputs_1_13, addersInputs_1_12, 
      addersInputs_1_11, addersInputs_1_10, addersInputs_1_9, 
      addersInputs_1_8, addersInputs_1_7, addersInputs_1_6, addersInputs_1_5, 
      addersInputs_1_4, addersInputs_1_3, addersInputs_1_2, addersInputs_1_1, 
      addersInputs_1_0, addersInputs_2_15, addersInputs_2_14, 
      addersInputs_2_13, addersInputs_2_12, addersInputs_2_11, 
      addersInputs_2_10, addersInputs_2_9, addersInputs_2_8, 
      addersInputs_2_7, addersInputs_2_6, addersInputs_2_5, addersInputs_2_4, 
      addersInputs_2_3, addersInputs_2_2, addersInputs_2_1, addersInputs_2_0, 
      addersInputs_3_15, addersInputs_3_14, addersInputs_3_13, 
      addersInputs_3_12, addersInputs_3_11, addersInputs_3_10, 
      addersInputs_3_9, addersInputs_3_8, addersInputs_3_7, addersInputs_3_6, 
      addersInputs_3_5, addersInputs_3_4, addersInputs_3_3, addersInputs_3_2, 
      addersInputs_3_1, addersInputs_3_0, addersInputs_4_15, 
      addersInputs_4_14, addersInputs_4_13, addersInputs_4_12, 
      addersInputs_4_11, addersInputs_4_10, addersInputs_4_9, 
      addersInputs_4_8, addersInputs_4_7, addersInputs_4_6, addersInputs_4_5, 
      addersInputs_4_4, addersInputs_4_3, addersInputs_4_2, addersInputs_4_1, 
      addersInputs_4_0, addersInputs_5_15, addersInputs_5_14, 
      addersInputs_5_13, addersInputs_5_12, addersInputs_5_11, 
      addersInputs_5_10, addersInputs_5_9, addersInputs_5_8, 
      addersInputs_5_7, addersInputs_5_6, addersInputs_5_5, addersInputs_5_4, 
      addersInputs_5_3, addersInputs_5_2, addersInputs_5_1, addersInputs_5_0, 
      addersInputs_6_15, addersInputs_6_14, addersInputs_6_13, 
      addersInputs_6_12, addersInputs_6_11, addersInputs_6_10, 
      addersInputs_6_9, addersInputs_6_8, addersInputs_6_7, addersInputs_6_6, 
      addersInputs_6_5, addersInputs_6_4, addersInputs_6_3, addersInputs_6_2, 
      addersInputs_6_1, addersInputs_6_0, addersInputs_7_15, 
      addersInputs_7_14, addersInputs_7_13, addersInputs_7_12, 
      addersInputs_7_11, addersInputs_7_10, addersInputs_7_9, 
      addersInputs_7_8, addersInputs_7_7, addersInputs_7_6, addersInputs_7_5, 
      addersInputs_7_4, addersInputs_7_3, addersInputs_7_2, addersInputs_7_1, 
      addersInputs_7_0, addersInputs_8_15, addersInputs_8_14, 
      addersInputs_8_13, addersInputs_8_12, addersInputs_8_11, 
      addersInputs_8_10, addersInputs_8_9, addersInputs_8_8, 
      addersInputs_8_7, addersInputs_8_6, addersInputs_8_5, addersInputs_8_4, 
      addersInputs_8_3, addersInputs_8_2, addersInputs_8_1, addersInputs_8_0, 
      addersInputs_9_15, addersInputs_9_14, addersInputs_9_13, 
      addersInputs_9_12, addersInputs_9_11, addersInputs_9_10, 
      addersInputs_9_9, addersInputs_9_8, addersInputs_9_7, addersInputs_9_6, 
      addersInputs_9_5, addersInputs_9_4, addersInputs_9_3, addersInputs_9_2, 
      addersInputs_9_1, addersInputs_9_0, addersInputs_10_15, 
      addersInputs_10_14, addersInputs_10_13, addersInputs_10_12, 
      addersInputs_10_11, addersInputs_10_10, addersInputs_10_9, 
      addersInputs_10_8, addersInputs_10_7, addersInputs_10_6, 
      addersInputs_10_5, addersInputs_10_4, addersInputs_10_3, 
      addersInputs_10_2, addersInputs_10_1, addersInputs_10_0, 
      addersInputs_11_15, addersInputs_11_14, addersInputs_11_13, 
      addersInputs_11_12, addersInputs_11_11, addersInputs_11_10, 
      addersInputs_11_9, addersInputs_11_8, addersInputs_11_7, 
      addersInputs_11_6, addersInputs_11_5, addersInputs_11_4, 
      addersInputs_11_3, addersInputs_11_2, addersInputs_11_1, 
      addersInputs_11_0, addersInputs_12_15, addersInputs_12_14, 
      addersInputs_12_13, addersInputs_12_12, addersInputs_12_11, 
      addersInputs_12_10, addersInputs_12_9, addersInputs_12_8, 
      addersInputs_12_7, addersInputs_12_6, addersInputs_12_5, 
      addersInputs_12_4, addersInputs_12_3, addersInputs_12_2, 
      addersInputs_12_1, addersInputs_12_0, addersInputs_13_15, 
      addersInputs_13_14, addersInputs_13_13, addersInputs_13_12, 
      addersInputs_13_11, addersInputs_13_10, addersInputs_13_9, 
      addersInputs_13_8, addersInputs_13_7, addersInputs_13_6, 
      addersInputs_13_5, addersInputs_13_4, addersInputs_13_3, 
      addersInputs_13_2, addersInputs_13_1, addersInputs_13_0, 
      addersInputs_14_15, addersInputs_14_14, addersInputs_14_13, 
      addersInputs_14_12, addersInputs_14_11, addersInputs_14_10, 
      addersInputs_14_9, addersInputs_14_8, addersInputs_14_7, 
      addersInputs_14_6, addersInputs_14_5, addersInputs_14_4, 
      addersInputs_14_3, addersInputs_14_2, addersInputs_14_1, 
      addersInputs_14_0, addersInputs_15_15, addersInputs_15_14, 
      addersInputs_15_13, addersInputs_15_12, addersInputs_15_11, 
      addersInputs_15_10, addersInputs_15_9, addersInputs_15_8, 
      addersInputs_15_7, addersInputs_15_6, addersInputs_15_5, 
      addersInputs_15_4, addersInputs_15_3, addersInputs_15_2, 
      addersInputs_15_1, addersInputs_15_0, addersInputs_16_15, 
      addersInputs_16_14, addersInputs_16_13, addersInputs_16_12, 
      addersInputs_16_11, addersInputs_16_10, addersInputs_16_9, 
      addersInputs_16_8, addersInputs_16_7, addersInputs_16_6, 
      addersInputs_16_5, addersInputs_16_4, addersInputs_16_3, 
      addersInputs_16_2, addersInputs_16_1, addersInputs_16_0, 
      addersInputs_17_15, addersInputs_17_14, addersInputs_17_13, 
      addersInputs_17_12, addersInputs_17_11, addersInputs_17_10, 
      addersInputs_17_9, addersInputs_17_8, addersInputs_17_7, 
      addersInputs_17_6, addersInputs_17_5, addersInputs_17_4, 
      addersInputs_17_3, addersInputs_17_2, addersInputs_17_1, 
      addersInputs_17_0, addersInputs_18_15, addersInputs_18_14, 
      addersInputs_18_13, addersInputs_18_12, addersInputs_18_11, 
      addersInputs_18_10, addersInputs_18_9, addersInputs_18_8, 
      addersInputs_18_7, addersInputs_18_6, addersInputs_18_5, 
      addersInputs_18_4, addersInputs_18_3, addersInputs_18_2, 
      addersInputs_18_1, addersInputs_18_0, addersInputs_19_15, 
      addersInputs_19_14, addersInputs_19_13, addersInputs_19_12, 
      addersInputs_19_11, addersInputs_19_10, addersInputs_19_9, 
      addersInputs_19_8, addersInputs_19_7, addersInputs_19_6, 
      addersInputs_19_5, addersInputs_19_4, addersInputs_19_3, 
      addersInputs_19_2, addersInputs_19_1, addersInputs_19_0, 
      addersInputs_20_15, addersInputs_20_14, addersInputs_20_13, 
      addersInputs_20_12, addersInputs_20_11, addersInputs_20_10, 
      addersInputs_20_9, addersInputs_20_8, addersInputs_20_7, 
      addersInputs_20_6, addersInputs_20_5, addersInputs_20_4, 
      addersInputs_20_3, addersInputs_20_2, addersInputs_20_1, 
      addersInputs_20_0, addersInputs_21_15, addersInputs_21_14, 
      addersInputs_21_13, addersInputs_21_12, addersInputs_21_11, 
      addersInputs_21_10, addersInputs_21_9, addersInputs_21_8, 
      addersInputs_21_7, addersInputs_21_6, addersInputs_21_5, 
      addersInputs_21_4, addersInputs_21_3, addersInputs_21_2, 
      addersInputs_21_1, addersInputs_21_0, addersInputs_22_15, 
      addersInputs_22_14, addersInputs_22_13, addersInputs_22_12, 
      addersInputs_22_11, addersInputs_22_10, addersInputs_22_9, 
      addersInputs_22_8, addersInputs_22_7, addersInputs_22_6, 
      addersInputs_22_5, addersInputs_22_4, addersInputs_22_3, 
      addersInputs_22_2, addersInputs_22_1, addersInputs_22_0, 
      addersInputs_23_15, addersInputs_23_14, addersInputs_23_13, 
      addersInputs_23_12, addersInputs_23_11, addersInputs_23_10, 
      addersInputs_23_9, addersInputs_23_8, addersInputs_23_7, 
      addersInputs_23_6, addersInputs_23_5, addersInputs_23_4, 
      addersInputs_23_3, addersInputs_23_2, addersInputs_23_1, 
      addersInputs_23_0, addersInputs_24_15, addersInputs_24_14, 
      addersInputs_24_13, addersInputs_24_12, addersInputs_24_11, 
      addersInputs_24_10, addersInputs_24_9, addersInputs_24_8, 
      addersInputs_24_7, addersInputs_24_6, addersInputs_24_5, 
      addersInputs_24_4, addersInputs_24_3, addersInputs_24_2, 
      addersInputs_24_1, addersInputs_24_0, filter_0_7, filter_0_6, 
      filter_0_5, filter_0_4, filter_0_3, filter_0_2, filter_0_1, filter_0_0, 
      filter_1_7, filter_1_6, filter_1_5, filter_1_4, filter_1_3, filter_1_2, 
      filter_1_1, filter_1_0, filter_2_7, filter_2_6, filter_2_5, filter_2_4, 
      filter_2_3, filter_2_2, filter_2_1, filter_2_0, filter_3_7, filter_3_6, 
      filter_3_5, filter_3_4, filter_3_3, filter_3_2, filter_3_1, filter_3_0, 
      filter_4_7, filter_4_6, filter_4_5, filter_4_4, filter_4_3, filter_4_2, 
      filter_4_1, filter_4_0, filter_5_7, filter_5_6, filter_5_5, filter_5_4, 
      filter_5_3, filter_5_2, filter_5_1, filter_5_0, filter_6_7, filter_6_6, 
      filter_6_5, filter_6_4, filter_6_3, filter_6_2, filter_6_1, filter_6_0, 
      filter_7_7, filter_7_6, filter_7_5, filter_7_4, filter_7_3, filter_7_2, 
      filter_7_1, filter_7_0, filter_8_7, filter_8_6, filter_8_5, filter_8_4, 
      filter_8_3, filter_8_2, filter_8_1, filter_8_0, filter_9_7, filter_9_6, 
      filter_9_5, filter_9_4, filter_9_3, filter_9_2, filter_9_1, filter_9_0, 
      filter_10_7, filter_10_6, filter_10_5, filter_10_4, filter_10_3, 
      filter_10_2, filter_10_1, filter_10_0, filter_11_7, filter_11_6, 
      filter_11_5, filter_11_4, filter_11_3, filter_11_2, filter_11_1, 
      filter_11_0, filter_12_7, filter_12_6, filter_12_5, filter_12_4, 
      filter_12_3, filter_12_2, filter_12_1, filter_12_0, filter_13_7, 
      filter_13_6, filter_13_5, filter_13_4, filter_13_3, filter_13_2, 
      filter_13_1, filter_13_0, filter_14_7, filter_14_6, filter_14_5, 
      filter_14_4, filter_14_3, filter_14_2, filter_14_1, filter_14_0, 
      filter_15_7, filter_15_6, filter_15_5, filter_15_4, filter_15_3, 
      filter_15_2, filter_15_1, filter_15_0, filter_16_7, filter_16_6, 
      filter_16_5, filter_16_4, filter_16_3, filter_16_2, filter_16_1, 
      filter_16_0, filter_17_7, filter_17_6, filter_17_5, filter_17_4, 
      filter_17_3, filter_17_2, filter_17_1, filter_17_0, filter_18_7, 
      filter_18_6, filter_18_5, filter_18_4, filter_18_3, filter_18_2, 
      filter_18_1, filter_18_0, filter_19_7, filter_19_6, filter_19_5, 
      filter_19_4, filter_19_3, filter_19_2, filter_19_1, filter_19_0, 
      filter_20_7, filter_20_6, filter_20_5, filter_20_4, filter_20_3, 
      filter_20_2, filter_20_1, filter_20_0, filter_21_7, filter_21_6, 
      filter_21_5, filter_21_4, filter_21_3, filter_21_2, filter_21_1, 
      filter_21_0, filter_22_7, filter_22_6, filter_22_5, filter_22_4, 
      filter_22_3, filter_22_2, filter_22_1, filter_22_0, filter_23_7, 
      filter_23_6, filter_23_5, filter_23_4, filter_23_3, filter_23_2, 
      filter_23_1, filter_23_0, filter_24_7, filter_24_6, filter_24_5, 
      filter_24_4, filter_24_3, filter_24_2, filter_24_1, filter_24_0, 
      doneMul, regFileMap_page1Out_5_15, regFileMap_page1Out_5_14, 
      regFileMap_page1Out_5_13, regFileMap_page1Out_5_12, 
      regFileMap_page1Out_5_11, regFileMap_page1Out_5_10, 
      regFileMap_page1Out_5_9, regFileMap_page1Out_5_8, 
      regFileMap_page1Out_5_7, regFileMap_page1Out_5_6, 
      regFileMap_page1Out_5_5, regFileMap_page1Out_5_4, 
      regFileMap_page1Out_5_3, regFileMap_page1Out_5_2, 
      regFileMap_page1Out_5_1, regFileMap_page1Out_5_0, 
      regFileMap_page1Out_6_15, regFileMap_page1Out_6_14, 
      regFileMap_page1Out_6_13, regFileMap_page1Out_6_12, 
      regFileMap_page1Out_6_11, regFileMap_page1Out_6_10, 
      regFileMap_page1Out_6_9, regFileMap_page1Out_6_8, 
      regFileMap_page1Out_6_7, regFileMap_page1Out_6_6, 
      regFileMap_page1Out_6_5, regFileMap_page1Out_6_4, 
      regFileMap_page1Out_6_3, regFileMap_page1Out_6_2, 
      regFileMap_page1Out_6_1, regFileMap_page1Out_6_0, 
      regFileMap_page1Out_7_15, regFileMap_page1Out_7_14, 
      regFileMap_page1Out_7_13, regFileMap_page1Out_7_12, 
      regFileMap_page1Out_7_11, regFileMap_page1Out_7_10, 
      regFileMap_page1Out_7_9, regFileMap_page1Out_7_8, 
      regFileMap_page1Out_7_7, regFileMap_page1Out_7_6, 
      regFileMap_page1Out_7_5, regFileMap_page1Out_7_4, 
      regFileMap_page1Out_7_3, regFileMap_page1Out_7_2, 
      regFileMap_page1Out_7_1, regFileMap_page1Out_7_0, 
      regFileMap_page1Out_8_15, regFileMap_page1Out_8_14, 
      regFileMap_page1Out_8_13, regFileMap_page1Out_8_12, 
      regFileMap_page1Out_8_11, regFileMap_page1Out_8_10, 
      regFileMap_page1Out_8_9, regFileMap_page1Out_8_8, 
      regFileMap_page1Out_8_7, regFileMap_page1Out_8_6, 
      regFileMap_page1Out_8_5, regFileMap_page1Out_8_4, 
      regFileMap_page1Out_8_3, regFileMap_page1Out_8_2, 
      regFileMap_page1Out_8_1, regFileMap_page1Out_8_0, 
      regFileMap_page1Out_9_15, regFileMap_page1Out_9_14, 
      regFileMap_page1Out_9_13, regFileMap_page1Out_9_12, 
      regFileMap_page1Out_9_11, regFileMap_page1Out_9_10, 
      regFileMap_page1Out_9_9, regFileMap_page1Out_9_8, 
      regFileMap_page1Out_9_7, regFileMap_page1Out_9_6, 
      regFileMap_page1Out_9_5, regFileMap_page1Out_9_4, 
      regFileMap_page1Out_9_3, regFileMap_page1Out_9_2, 
      regFileMap_page1Out_9_1, regFileMap_page1Out_9_0, 
      regFileMap_page1Out_10_15, regFileMap_page1Out_10_14, 
      regFileMap_page1Out_10_13, regFileMap_page1Out_10_12, 
      regFileMap_page1Out_10_11, regFileMap_page1Out_10_10, 
      regFileMap_page1Out_10_9, regFileMap_page1Out_10_8, 
      regFileMap_page1Out_10_7, regFileMap_page1Out_10_6, 
      regFileMap_page1Out_10_5, regFileMap_page1Out_10_4, 
      regFileMap_page1Out_10_3, regFileMap_page1Out_10_2, 
      regFileMap_page1Out_10_1, regFileMap_page1Out_10_0, 
      regFileMap_page1Out_11_15, regFileMap_page1Out_11_14, 
      regFileMap_page1Out_11_13, regFileMap_page1Out_11_12, 
      regFileMap_page1Out_11_11, regFileMap_page1Out_11_10, 
      regFileMap_page1Out_11_9, regFileMap_page1Out_11_8, 
      regFileMap_page1Out_11_7, regFileMap_page1Out_11_6, 
      regFileMap_page1Out_11_5, regFileMap_page1Out_11_4, 
      regFileMap_page1Out_11_3, regFileMap_page1Out_11_2, 
      regFileMap_page1Out_11_1, regFileMap_page1Out_11_0, 
      regFileMap_page1Out_12_15, regFileMap_page1Out_12_14, 
      regFileMap_page1Out_12_13, regFileMap_page1Out_12_12, 
      regFileMap_page1Out_12_11, regFileMap_page1Out_12_10, 
      regFileMap_page1Out_12_9, regFileMap_page1Out_12_8, 
      regFileMap_page1Out_12_7, regFileMap_page1Out_12_6, 
      regFileMap_page1Out_12_5, regFileMap_page1Out_12_4, 
      regFileMap_page1Out_12_3, regFileMap_page1Out_12_2, 
      regFileMap_page1Out_12_1, regFileMap_page1Out_12_0, 
      regFileMap_page1Out_13_15, regFileMap_page1Out_13_14, 
      regFileMap_page1Out_13_13, regFileMap_page1Out_13_12, 
      regFileMap_page1Out_13_11, regFileMap_page1Out_13_10, 
      regFileMap_page1Out_13_9, regFileMap_page1Out_13_8, 
      regFileMap_page1Out_13_7, regFileMap_page1Out_13_6, 
      regFileMap_page1Out_13_5, regFileMap_page1Out_13_4, 
      regFileMap_page1Out_13_3, regFileMap_page1Out_13_2, 
      regFileMap_page1Out_13_1, regFileMap_page1Out_13_0, 
      regFileMap_page1Out_14_15, regFileMap_page1Out_14_14, 
      regFileMap_page1Out_14_13, regFileMap_page1Out_14_12, 
      regFileMap_page1Out_14_11, regFileMap_page1Out_14_10, 
      regFileMap_page1Out_14_9, regFileMap_page1Out_14_8, 
      regFileMap_page1Out_14_7, regFileMap_page1Out_14_6, 
      regFileMap_page1Out_14_5, regFileMap_page1Out_14_4, 
      regFileMap_page1Out_14_3, regFileMap_page1Out_14_2, 
      regFileMap_page1Out_14_1, regFileMap_page1Out_14_0, 
      regFileMap_page1Out_15_15, regFileMap_page1Out_15_14, 
      regFileMap_page1Out_15_13, regFileMap_page1Out_15_12, 
      regFileMap_page1Out_15_11, regFileMap_page1Out_15_10, 
      regFileMap_page1Out_15_9, regFileMap_page1Out_15_8, 
      regFileMap_page1Out_15_7, regFileMap_page1Out_15_6, 
      regFileMap_page1Out_15_5, regFileMap_page1Out_15_4, 
      regFileMap_page1Out_15_3, regFileMap_page1Out_15_2, 
      regFileMap_page1Out_15_1, regFileMap_page1Out_15_0, 
      regFileMap_page1Out_16_15, regFileMap_page1Out_16_14, 
      regFileMap_page1Out_16_13, regFileMap_page1Out_16_12, 
      regFileMap_page1Out_16_11, regFileMap_page1Out_16_10, 
      regFileMap_page1Out_16_9, regFileMap_page1Out_16_8, 
      regFileMap_page1Out_16_7, regFileMap_page1Out_16_6, 
      regFileMap_page1Out_16_5, regFileMap_page1Out_16_4, 
      regFileMap_page1Out_16_3, regFileMap_page1Out_16_2, 
      regFileMap_page1Out_16_1, regFileMap_page1Out_16_0, 
      regFileMap_page1Out_17_15, regFileMap_page1Out_17_14, 
      regFileMap_page1Out_17_13, regFileMap_page1Out_17_12, 
      regFileMap_page1Out_17_11, regFileMap_page1Out_17_10, 
      regFileMap_page1Out_17_9, regFileMap_page1Out_17_8, 
      regFileMap_page1Out_17_7, regFileMap_page1Out_17_6, 
      regFileMap_page1Out_17_5, regFileMap_page1Out_17_4, 
      regFileMap_page1Out_17_3, regFileMap_page1Out_17_2, 
      regFileMap_page1Out_17_1, regFileMap_page1Out_17_0, 
      regFileMap_page1Out_18_15, regFileMap_page1Out_18_14, 
      regFileMap_page1Out_18_13, regFileMap_page1Out_18_12, 
      regFileMap_page1Out_18_11, regFileMap_page1Out_18_10, 
      regFileMap_page1Out_18_9, regFileMap_page1Out_18_8, 
      regFileMap_page1Out_18_7, regFileMap_page1Out_18_6, 
      regFileMap_page1Out_18_5, regFileMap_page1Out_18_4, 
      regFileMap_page1Out_18_3, regFileMap_page1Out_18_2, 
      regFileMap_page1Out_18_1, regFileMap_page1Out_18_0, 
      regFileMap_page1Out_19_15, regFileMap_page1Out_19_14, 
      regFileMap_page1Out_19_13, regFileMap_page1Out_19_12, 
      regFileMap_page1Out_19_11, regFileMap_page1Out_19_10, 
      regFileMap_page1Out_19_9, regFileMap_page1Out_19_8, 
      regFileMap_page1Out_19_7, regFileMap_page1Out_19_6, 
      regFileMap_page1Out_19_5, regFileMap_page1Out_19_4, 
      regFileMap_page1Out_19_3, regFileMap_page1Out_19_2, 
      regFileMap_page1Out_19_1, regFileMap_page1Out_19_0, 
      regFileMap_page1Out_20_15, regFileMap_page1Out_20_14, 
      regFileMap_page1Out_20_13, regFileMap_page1Out_20_12, 
      regFileMap_page1Out_20_11, regFileMap_page1Out_20_10, 
      regFileMap_page1Out_20_9, regFileMap_page1Out_20_8, 
      regFileMap_page1Out_20_7, regFileMap_page1Out_20_6, 
      regFileMap_page1Out_20_5, regFileMap_page1Out_20_4, 
      regFileMap_page1Out_20_3, regFileMap_page1Out_20_2, 
      regFileMap_page1Out_20_1, regFileMap_page1Out_20_0, 
      regFileMap_page1Out_21_15, regFileMap_page1Out_21_14, 
      regFileMap_page1Out_21_13, regFileMap_page1Out_21_12, 
      regFileMap_page1Out_21_11, regFileMap_page1Out_21_10, 
      regFileMap_page1Out_21_9, regFileMap_page1Out_21_8, 
      regFileMap_page1Out_21_7, regFileMap_page1Out_21_6, 
      regFileMap_page1Out_21_5, regFileMap_page1Out_21_4, 
      regFileMap_page1Out_21_3, regFileMap_page1Out_21_2, 
      regFileMap_page1Out_21_1, regFileMap_page1Out_21_0, 
      regFileMap_page1Out_22_15, regFileMap_page1Out_22_14, 
      regFileMap_page1Out_22_13, regFileMap_page1Out_22_12, 
      regFileMap_page1Out_22_11, regFileMap_page1Out_22_10, 
      regFileMap_page1Out_22_9, regFileMap_page1Out_22_8, 
      regFileMap_page1Out_22_7, regFileMap_page1Out_22_6, 
      regFileMap_page1Out_22_5, regFileMap_page1Out_22_4, 
      regFileMap_page1Out_22_3, regFileMap_page1Out_22_2, 
      regFileMap_page1Out_22_1, regFileMap_page1Out_22_0, 
      regFileMap_page1Out_23_15, regFileMap_page1Out_23_14, 
      regFileMap_page1Out_23_13, regFileMap_page1Out_23_12, 
      regFileMap_page1Out_23_11, regFileMap_page1Out_23_10, 
      regFileMap_page1Out_23_9, regFileMap_page1Out_23_8, 
      regFileMap_page1Out_23_7, regFileMap_page1Out_23_6, 
      regFileMap_page1Out_23_5, regFileMap_page1Out_23_4, 
      regFileMap_page1Out_23_3, regFileMap_page1Out_23_2, 
      regFileMap_page1Out_23_1, regFileMap_page1Out_23_0, 
      regFileMap_page1Out_24_15, regFileMap_page1Out_24_14, 
      regFileMap_page1Out_24_13, regFileMap_page1Out_24_12, 
      regFileMap_page1Out_24_11, regFileMap_page1Out_24_10, 
      regFileMap_page1Out_24_9, regFileMap_page1Out_24_8, 
      regFileMap_page1Out_24_7, regFileMap_page1Out_24_6, 
      regFileMap_page1Out_24_5, regFileMap_page1Out_24_4, 
      regFileMap_page1Out_24_3, regFileMap_page1Out_24_2, 
      regFileMap_page1Out_24_1, regFileMap_page1Out_24_0, 
      regFileMap_page2Out_5_15, regFileMap_page2Out_5_14, 
      regFileMap_page2Out_5_13, regFileMap_page2Out_5_12, 
      regFileMap_page2Out_5_11, regFileMap_page2Out_5_10, 
      regFileMap_page2Out_5_9, regFileMap_page2Out_5_8, 
      regFileMap_page2Out_5_7, regFileMap_page2Out_5_6, 
      regFileMap_page2Out_5_5, regFileMap_page2Out_5_4, 
      regFileMap_page2Out_5_3, regFileMap_page2Out_5_2, 
      regFileMap_page2Out_5_1, regFileMap_page2Out_5_0, 
      regFileMap_page2Out_6_15, regFileMap_page2Out_6_14, 
      regFileMap_page2Out_6_13, regFileMap_page2Out_6_12, 
      regFileMap_page2Out_6_11, regFileMap_page2Out_6_10, 
      regFileMap_page2Out_6_9, regFileMap_page2Out_6_8, 
      regFileMap_page2Out_6_7, regFileMap_page2Out_6_6, 
      regFileMap_page2Out_6_5, regFileMap_page2Out_6_4, 
      regFileMap_page2Out_6_3, regFileMap_page2Out_6_2, 
      regFileMap_page2Out_6_1, regFileMap_page2Out_6_0, 
      regFileMap_page2Out_7_15, regFileMap_page2Out_7_14, 
      regFileMap_page2Out_7_13, regFileMap_page2Out_7_12, 
      regFileMap_page2Out_7_11, regFileMap_page2Out_7_10, 
      regFileMap_page2Out_7_9, regFileMap_page2Out_7_8, 
      regFileMap_page2Out_7_7, regFileMap_page2Out_7_6, 
      regFileMap_page2Out_7_5, regFileMap_page2Out_7_4, 
      regFileMap_page2Out_7_3, regFileMap_page2Out_7_2, 
      regFileMap_page2Out_7_1, regFileMap_page2Out_7_0, 
      regFileMap_page2Out_8_15, regFileMap_page2Out_8_14, 
      regFileMap_page2Out_8_13, regFileMap_page2Out_8_12, 
      regFileMap_page2Out_8_11, regFileMap_page2Out_8_10, 
      regFileMap_page2Out_8_9, regFileMap_page2Out_8_8, 
      regFileMap_page2Out_8_7, regFileMap_page2Out_8_6, 
      regFileMap_page2Out_8_5, regFileMap_page2Out_8_4, 
      regFileMap_page2Out_8_3, regFileMap_page2Out_8_2, 
      regFileMap_page2Out_8_1, regFileMap_page2Out_8_0, 
      regFileMap_page2Out_9_15, regFileMap_page2Out_9_14, 
      regFileMap_page2Out_9_13, regFileMap_page2Out_9_12, 
      regFileMap_page2Out_9_11, regFileMap_page2Out_9_10, 
      regFileMap_page2Out_9_9, regFileMap_page2Out_9_8, 
      regFileMap_page2Out_9_7, regFileMap_page2Out_9_6, 
      regFileMap_page2Out_9_5, regFileMap_page2Out_9_4, 
      regFileMap_page2Out_9_3, regFileMap_page2Out_9_2, 
      regFileMap_page2Out_9_1, regFileMap_page2Out_9_0, 
      regFileMap_page2Out_10_15, regFileMap_page2Out_10_14, 
      regFileMap_page2Out_10_13, regFileMap_page2Out_10_12, 
      regFileMap_page2Out_10_11, regFileMap_page2Out_10_10, 
      regFileMap_page2Out_10_9, regFileMap_page2Out_10_8, 
      regFileMap_page2Out_10_7, regFileMap_page2Out_10_6, 
      regFileMap_page2Out_10_5, regFileMap_page2Out_10_4, 
      regFileMap_page2Out_10_3, regFileMap_page2Out_10_2, 
      regFileMap_page2Out_10_1, regFileMap_page2Out_10_0, 
      regFileMap_page2Out_11_15, regFileMap_page2Out_11_14, 
      regFileMap_page2Out_11_13, regFileMap_page2Out_11_12, 
      regFileMap_page2Out_11_11, regFileMap_page2Out_11_10, 
      regFileMap_page2Out_11_9, regFileMap_page2Out_11_8, 
      regFileMap_page2Out_11_7, regFileMap_page2Out_11_6, 
      regFileMap_page2Out_11_5, regFileMap_page2Out_11_4, 
      regFileMap_page2Out_11_3, regFileMap_page2Out_11_2, 
      regFileMap_page2Out_11_1, regFileMap_page2Out_11_0, 
      regFileMap_page2Out_12_15, regFileMap_page2Out_12_14, 
      regFileMap_page2Out_12_13, regFileMap_page2Out_12_12, 
      regFileMap_page2Out_12_11, regFileMap_page2Out_12_10, 
      regFileMap_page2Out_12_9, regFileMap_page2Out_12_8, 
      regFileMap_page2Out_12_7, regFileMap_page2Out_12_6, 
      regFileMap_page2Out_12_5, regFileMap_page2Out_12_4, 
      regFileMap_page2Out_12_3, regFileMap_page2Out_12_2, 
      regFileMap_page2Out_12_1, regFileMap_page2Out_12_0, 
      regFileMap_page2Out_13_15, regFileMap_page2Out_13_14, 
      regFileMap_page2Out_13_13, regFileMap_page2Out_13_12, 
      regFileMap_page2Out_13_11, regFileMap_page2Out_13_10, 
      regFileMap_page2Out_13_9, regFileMap_page2Out_13_8, 
      regFileMap_page2Out_13_7, regFileMap_page2Out_13_6, 
      regFileMap_page2Out_13_5, regFileMap_page2Out_13_4, 
      regFileMap_page2Out_13_3, regFileMap_page2Out_13_2, 
      regFileMap_page2Out_13_1, regFileMap_page2Out_13_0, 
      regFileMap_page2Out_14_15, regFileMap_page2Out_14_14, 
      regFileMap_page2Out_14_13, regFileMap_page2Out_14_12, 
      regFileMap_page2Out_14_11, regFileMap_page2Out_14_10, 
      regFileMap_page2Out_14_9, regFileMap_page2Out_14_8, 
      regFileMap_page2Out_14_7, regFileMap_page2Out_14_6, 
      regFileMap_page2Out_14_5, regFileMap_page2Out_14_4, 
      regFileMap_page2Out_14_3, regFileMap_page2Out_14_2, 
      regFileMap_page2Out_14_1, regFileMap_page2Out_14_0, 
      regFileMap_page2Out_15_15, regFileMap_page2Out_15_14, 
      regFileMap_page2Out_15_13, regFileMap_page2Out_15_12, 
      regFileMap_page2Out_15_11, regFileMap_page2Out_15_10, 
      regFileMap_page2Out_15_9, regFileMap_page2Out_15_8, 
      regFileMap_page2Out_15_7, regFileMap_page2Out_15_6, 
      regFileMap_page2Out_15_5, regFileMap_page2Out_15_4, 
      regFileMap_page2Out_15_3, regFileMap_page2Out_15_2, 
      regFileMap_page2Out_15_1, regFileMap_page2Out_15_0, 
      regFileMap_page2Out_16_15, regFileMap_page2Out_16_14, 
      regFileMap_page2Out_16_13, regFileMap_page2Out_16_12, 
      regFileMap_page2Out_16_11, regFileMap_page2Out_16_10, 
      regFileMap_page2Out_16_9, regFileMap_page2Out_16_8, 
      regFileMap_page2Out_16_7, regFileMap_page2Out_16_6, 
      regFileMap_page2Out_16_5, regFileMap_page2Out_16_4, 
      regFileMap_page2Out_16_3, regFileMap_page2Out_16_2, 
      regFileMap_page2Out_16_1, regFileMap_page2Out_16_0, 
      regFileMap_page2Out_17_15, regFileMap_page2Out_17_14, 
      regFileMap_page2Out_17_13, regFileMap_page2Out_17_12, 
      regFileMap_page2Out_17_11, regFileMap_page2Out_17_10, 
      regFileMap_page2Out_17_9, regFileMap_page2Out_17_8, 
      regFileMap_page2Out_17_7, regFileMap_page2Out_17_6, 
      regFileMap_page2Out_17_5, regFileMap_page2Out_17_4, 
      regFileMap_page2Out_17_3, regFileMap_page2Out_17_2, 
      regFileMap_page2Out_17_1, regFileMap_page2Out_17_0, 
      regFileMap_page2Out_18_15, regFileMap_page2Out_18_14, 
      regFileMap_page2Out_18_13, regFileMap_page2Out_18_12, 
      regFileMap_page2Out_18_11, regFileMap_page2Out_18_10, 
      regFileMap_page2Out_18_9, regFileMap_page2Out_18_8, 
      regFileMap_page2Out_18_7, regFileMap_page2Out_18_6, 
      regFileMap_page2Out_18_5, regFileMap_page2Out_18_4, 
      regFileMap_page2Out_18_3, regFileMap_page2Out_18_2, 
      regFileMap_page2Out_18_1, regFileMap_page2Out_18_0, 
      regFileMap_page2Out_19_15, regFileMap_page2Out_19_14, 
      regFileMap_page2Out_19_13, regFileMap_page2Out_19_12, 
      regFileMap_page2Out_19_11, regFileMap_page2Out_19_10, 
      regFileMap_page2Out_19_9, regFileMap_page2Out_19_8, 
      regFileMap_page2Out_19_7, regFileMap_page2Out_19_6, 
      regFileMap_page2Out_19_5, regFileMap_page2Out_19_4, 
      regFileMap_page2Out_19_3, regFileMap_page2Out_19_2, 
      regFileMap_page2Out_19_1, regFileMap_page2Out_19_0, 
      regFileMap_page2Out_20_15, regFileMap_page2Out_20_14, 
      regFileMap_page2Out_20_13, regFileMap_page2Out_20_12, 
      regFileMap_page2Out_20_11, regFileMap_page2Out_20_10, 
      regFileMap_page2Out_20_9, regFileMap_page2Out_20_8, 
      regFileMap_page2Out_20_7, regFileMap_page2Out_20_6, 
      regFileMap_page2Out_20_5, regFileMap_page2Out_20_4, 
      regFileMap_page2Out_20_3, regFileMap_page2Out_20_2, 
      regFileMap_page2Out_20_1, regFileMap_page2Out_20_0, 
      regFileMap_page2Out_21_15, regFileMap_page2Out_21_14, 
      regFileMap_page2Out_21_13, regFileMap_page2Out_21_12, 
      regFileMap_page2Out_21_11, regFileMap_page2Out_21_10, 
      regFileMap_page2Out_21_9, regFileMap_page2Out_21_8, 
      regFileMap_page2Out_21_7, regFileMap_page2Out_21_6, 
      regFileMap_page2Out_21_5, regFileMap_page2Out_21_4, 
      regFileMap_page2Out_21_3, regFileMap_page2Out_21_2, 
      regFileMap_page2Out_21_1, regFileMap_page2Out_21_0, 
      regFileMap_page2Out_22_15, regFileMap_page2Out_22_14, 
      regFileMap_page2Out_22_13, regFileMap_page2Out_22_12, 
      regFileMap_page2Out_22_11, regFileMap_page2Out_22_10, 
      regFileMap_page2Out_22_9, regFileMap_page2Out_22_8, 
      regFileMap_page2Out_22_7, regFileMap_page2Out_22_6, 
      regFileMap_page2Out_22_5, regFileMap_page2Out_22_4, 
      regFileMap_page2Out_22_3, regFileMap_page2Out_22_2, 
      regFileMap_page2Out_22_1, regFileMap_page2Out_22_0, 
      regFileMap_page2Out_23_15, regFileMap_page2Out_23_14, 
      regFileMap_page2Out_23_13, regFileMap_page2Out_23_12, 
      regFileMap_page2Out_23_11, regFileMap_page2Out_23_10, 
      regFileMap_page2Out_23_9, regFileMap_page2Out_23_8, 
      regFileMap_page2Out_23_7, regFileMap_page2Out_23_6, 
      regFileMap_page2Out_23_5, regFileMap_page2Out_23_4, 
      regFileMap_page2Out_23_3, regFileMap_page2Out_23_2, 
      regFileMap_page2Out_23_1, regFileMap_page2Out_23_0, 
      regFileMap_page2Out_24_15, regFileMap_page2Out_24_14, 
      regFileMap_page2Out_24_13, regFileMap_page2Out_24_12, 
      regFileMap_page2Out_24_11, regFileMap_page2Out_24_10, 
      regFileMap_page2Out_24_9, regFileMap_page2Out_24_8, 
      regFileMap_page2Out_24_7, regFileMap_page2Out_24_6, 
      regFileMap_page2Out_24_5, regFileMap_page2Out_24_4, 
      regFileMap_page2Out_24_3, regFileMap_page2Out_24_2, 
      regFileMap_page2Out_24_1, regFileMap_page2Out_24_0, 
      regFileMap_page1Enables_0, regFileMap_page1Enables_1, 
      regFileMap_page1Enables_2, regFileMap_page1Enables_3, 
      regFileMap_page1Enables_4, regFileMap_page2Enables_0, 
      regFileMap_page2Enables_1, regFileMap_page2Enables_2, 
      regFileMap_page2Enables_3, regFileMap_page2Enables_4, 
      regFileMap_filterEnables_0, regFileMap_filterEnables_1, 
      regFileMap_filterEnables_2, regFileMap_filterEnables_3, 
      addersMap_sum1_15, addersMap_sum1_14, addersMap_sum1_13, 
      addersMap_sum1_12, addersMap_sum1_11, addersMap_sum1_10, 
      addersMap_sum1_9, addersMap_sum1_8, addersMap_sum1_7, addersMap_sum1_6, 
      addersMap_sum1_5, addersMap_sum1_4, addersMap_sum1_3, addersMap_sum1_2, 
      addersMap_sum1_1, addersMap_sum1_0, addersMap_sum2_15, 
      addersMap_sum2_14, addersMap_sum2_13, addersMap_sum2_12, 
      addersMap_sum2_11, addersMap_sum2_10, addersMap_sum2_9, 
      addersMap_sum2_8, addersMap_sum2_7, addersMap_sum2_6, addersMap_sum2_5, 
      addersMap_sum2_4, addersMap_sum2_3, addersMap_sum2_2, addersMap_sum2_1, 
      addersMap_sum2_0, addersMap_sum3_15, addersMap_sum3_14, 
      addersMap_sum3_13, addersMap_sum3_12, addersMap_sum3_11, 
      addersMap_sum3_10, addersMap_sum3_9, addersMap_sum3_8, 
      addersMap_sum3_7, addersMap_sum3_6, addersMap_sum3_5, addersMap_sum3_4, 
      addersMap_sum3_3, addersMap_sum3_2, addersMap_sum3_1, addersMap_sum3_0, 
      addersMap_sum3Filter_15, addersMap_sum3Filter_14, 
      addersMap_sum3Filter_13, addersMap_sum3Filter_12, 
      addersMap_sum3Filter_11, addersMap_sum3Filter_10, 
      addersMap_sum3Filter_9, addersMap_sum3Filter_8, addersMap_sum3Filter_7, 
      addersMap_sum3Filter_6, addersMap_sum3Filter_5, addersMap_sum3Filter_4, 
      addersMap_sum3Filter_3, addersMap_sum3Filter_2, addersMap_sum3Filter_1, 
      addersMap_sum3Filter_0, addersMap_sum4_15, addersMap_sum4_14, 
      addersMap_sum4_13, addersMap_sum4_12, addersMap_sum4_11, 
      addersMap_sum4_10, addersMap_sum4_9, addersMap_sum4_8, 
      addersMap_sum4_7, addersMap_sum4_6, addersMap_sum4_5, addersMap_sum4_4, 
      addersMap_sum4_3, addersMap_sum4_2, addersMap_sum4_1, addersMap_sum4_0, 
      addersMap_totalSum_15, addersMap_totalSum_14, addersMap_totalSum_13, 
      addersMap_totalSum_12, addersMap_totalSum_11, addersMap_totalSum_10, 
      addersMap_totalSum_9, addersMap_totalSum_8, addersMap_totalSum_7, 
      addersMap_totalSum_6, addersMap_totalSum_5, addersMap_totalSum_4, 
      addersMap_totalSum_3, addersMap_totalSum_2, addersMap_totalSum_1, 
      addersMap_totalSum_0, addersMap_sum1Map_sum1_15_dup_0, 
      addersMap_sum1Map_sum1_14_dup_0, addersMap_sum1Map_sum1_13_dup_0, 
      addersMap_sum1Map_sum1_12_dup_0, addersMap_sum1Map_sum1_11_dup_0, 
      addersMap_sum1Map_sum1_10_dup_0, addersMap_sum1Map_sum1_9_dup_0, 
      addersMap_sum1Map_sum1_8_dup_0, addersMap_sum1Map_sum1_7_dup_0, 
      addersMap_sum1Map_sum1_6_dup_0, addersMap_sum1Map_sum1_5_dup_0, 
      addersMap_sum1Map_sum1_4_dup_0, addersMap_sum1Map_sum1_3_dup_0, 
      addersMap_sum1Map_sum1_2_dup_0, addersMap_sum1Map_sum1_1_dup_0, 
      addersMap_sum1Map_sum1_0_dup_0, addersMap_sum1Map_sum2_15_dup_0, 
      addersMap_sum1Map_sum2_14_dup_0, addersMap_sum1Map_sum2_13_dup_0, 
      addersMap_sum1Map_sum2_12_dup_0, addersMap_sum1Map_sum2_11_dup_0, 
      addersMap_sum1Map_sum2_10_dup_0, addersMap_sum1Map_sum2_9_dup_0, 
      addersMap_sum1Map_sum2_8_dup_0, addersMap_sum1Map_sum2_7_dup_0, 
      addersMap_sum1Map_sum2_6_dup_0, addersMap_sum1Map_sum2_5_dup_0, 
      addersMap_sum1Map_sum2_4_dup_0, addersMap_sum1Map_sum2_3_dup_0, 
      addersMap_sum1Map_sum2_2_dup_0, addersMap_sum1Map_sum2_1_dup_0, 
      addersMap_sum1Map_sum2_0_dup_0, addersMap_sum1Map_sum1Map_sum1_15, 
      addersMap_sum1Map_sum1Map_sum1_14, addersMap_sum1Map_sum1Map_sum1_13, 
      addersMap_sum1Map_sum1Map_sum1_12, addersMap_sum1Map_sum1Map_sum1_11, 
      addersMap_sum1Map_sum1Map_sum1_10, addersMap_sum1Map_sum1Map_sum1_9, 
      addersMap_sum1Map_sum1Map_sum1_8, addersMap_sum1Map_sum1Map_sum1_7, 
      addersMap_sum1Map_sum1Map_sum1_6, addersMap_sum1Map_sum1Map_sum1_5, 
      addersMap_sum1Map_sum1Map_sum1_4, addersMap_sum1Map_sum1Map_sum1_3, 
      addersMap_sum1Map_sum1Map_sum1_2, addersMap_sum1Map_sum1Map_sum1_1, 
      addersMap_sum1Map_sum1Map_sum1_0, addersMap_sum1Map_sum1Map_sum2_15, 
      addersMap_sum1Map_sum1Map_sum2_14, addersMap_sum1Map_sum1Map_sum2_13, 
      addersMap_sum1Map_sum1Map_sum2_12, addersMap_sum1Map_sum1Map_sum2_11, 
      addersMap_sum1Map_sum1Map_sum2_10, addersMap_sum1Map_sum1Map_sum2_9, 
      addersMap_sum1Map_sum1Map_sum2_8, addersMap_sum1Map_sum1Map_sum2_7, 
      addersMap_sum1Map_sum1Map_sum2_6, addersMap_sum1Map_sum1Map_sum2_5, 
      addersMap_sum1Map_sum1Map_sum2_4, addersMap_sum1Map_sum1Map_sum2_3, 
      addersMap_sum1Map_sum1Map_sum2_2, addersMap_sum1Map_sum1Map_sum2_1, 
      addersMap_sum1Map_sum1Map_sum2_0, addersMap_sum1Map_sum2Map_sum1_15, 
      addersMap_sum1Map_sum2Map_sum1_14, addersMap_sum1Map_sum2Map_sum1_13, 
      addersMap_sum1Map_sum2Map_sum1_12, addersMap_sum1Map_sum2Map_sum1_11, 
      addersMap_sum1Map_sum2Map_sum1_10, addersMap_sum1Map_sum2Map_sum1_9, 
      addersMap_sum1Map_sum2Map_sum1_8, addersMap_sum1Map_sum2Map_sum1_7, 
      addersMap_sum1Map_sum2Map_sum1_6, addersMap_sum1Map_sum2Map_sum1_5, 
      addersMap_sum1Map_sum2Map_sum1_4, addersMap_sum1Map_sum2Map_sum1_3, 
      addersMap_sum1Map_sum2Map_sum1_2, addersMap_sum1Map_sum2Map_sum1_1, 
      addersMap_sum1Map_sum2Map_sum1_0, addersMap_sum1Map_sum2Map_sum2_15, 
      addersMap_sum1Map_sum2Map_sum2_14, addersMap_sum1Map_sum2Map_sum2_13, 
      addersMap_sum1Map_sum2Map_sum2_12, addersMap_sum1Map_sum2Map_sum2_11, 
      addersMap_sum1Map_sum2Map_sum2_10, addersMap_sum1Map_sum2Map_sum2_9, 
      addersMap_sum1Map_sum2Map_sum2_8, addersMap_sum1Map_sum2Map_sum2_7, 
      addersMap_sum1Map_sum2Map_sum2_6, addersMap_sum1Map_sum2Map_sum2_5, 
      addersMap_sum1Map_sum2Map_sum2_4, addersMap_sum1Map_sum2Map_sum2_3, 
      addersMap_sum1Map_sum2Map_sum2_2, addersMap_sum1Map_sum2Map_sum2_1, 
      addersMap_sum1Map_sum2Map_sum2_0, addersMap_sum2Map_sum1_15_dup_0, 
      addersMap_sum2Map_sum1_14_dup_0, addersMap_sum2Map_sum1_13_dup_0, 
      addersMap_sum2Map_sum1_12_dup_0, addersMap_sum2Map_sum1_11_dup_0, 
      addersMap_sum2Map_sum1_10_dup_0, addersMap_sum2Map_sum1_9_dup_0, 
      addersMap_sum2Map_sum1_8_dup_0, addersMap_sum2Map_sum1_7_dup_0, 
      addersMap_sum2Map_sum1_6_dup_0, addersMap_sum2Map_sum1_5_dup_0, 
      addersMap_sum2Map_sum1_4_dup_0, addersMap_sum2Map_sum1_3_dup_0, 
      addersMap_sum2Map_sum1_2_dup_0, addersMap_sum2Map_sum1_1_dup_0, 
      addersMap_sum2Map_sum1_0_dup_0, addersMap_sum2Map_sum2_15_dup_0, 
      addersMap_sum2Map_sum2_14_dup_0, addersMap_sum2Map_sum2_13_dup_0, 
      addersMap_sum2Map_sum2_12_dup_0, addersMap_sum2Map_sum2_11_dup_0, 
      addersMap_sum2Map_sum2_10_dup_0, addersMap_sum2Map_sum2_9_dup_0, 
      addersMap_sum2Map_sum2_8_dup_0, addersMap_sum2Map_sum2_7_dup_0, 
      addersMap_sum2Map_sum2_6_dup_0, addersMap_sum2Map_sum2_5_dup_0, 
      addersMap_sum2Map_sum2_4_dup_0, addersMap_sum2Map_sum2_3_dup_0, 
      addersMap_sum2Map_sum2_2_dup_0, addersMap_sum2Map_sum2_1_dup_0, 
      addersMap_sum2Map_sum2_0_dup_0, addersMap_sum2Map_sum1Map_sum1_15, 
      addersMap_sum2Map_sum1Map_sum1_14, addersMap_sum2Map_sum1Map_sum1_13, 
      addersMap_sum2Map_sum1Map_sum1_12, addersMap_sum2Map_sum1Map_sum1_11, 
      addersMap_sum2Map_sum1Map_sum1_10, addersMap_sum2Map_sum1Map_sum1_9, 
      addersMap_sum2Map_sum1Map_sum1_8, addersMap_sum2Map_sum1Map_sum1_7, 
      addersMap_sum2Map_sum1Map_sum1_6, addersMap_sum2Map_sum1Map_sum1_5, 
      addersMap_sum2Map_sum1Map_sum1_4, addersMap_sum2Map_sum1Map_sum1_3, 
      addersMap_sum2Map_sum1Map_sum1_2, addersMap_sum2Map_sum1Map_sum1_1, 
      addersMap_sum2Map_sum1Map_sum1_0, addersMap_sum2Map_sum1Map_sum2_15, 
      addersMap_sum2Map_sum1Map_sum2_14, addersMap_sum2Map_sum1Map_sum2_13, 
      addersMap_sum2Map_sum1Map_sum2_12, addersMap_sum2Map_sum1Map_sum2_11, 
      addersMap_sum2Map_sum1Map_sum2_10, addersMap_sum2Map_sum1Map_sum2_9, 
      addersMap_sum2Map_sum1Map_sum2_8, addersMap_sum2Map_sum1Map_sum2_7, 
      addersMap_sum2Map_sum1Map_sum2_6, addersMap_sum2Map_sum1Map_sum2_5, 
      addersMap_sum2Map_sum1Map_sum2_4, addersMap_sum2Map_sum1Map_sum2_3, 
      addersMap_sum2Map_sum1Map_sum2_2, addersMap_sum2Map_sum1Map_sum2_1, 
      addersMap_sum2Map_sum1Map_sum2_0, addersMap_sum2Map_sum2Map_sum1_15, 
      addersMap_sum2Map_sum2Map_sum1_14, addersMap_sum2Map_sum2Map_sum1_13, 
      addersMap_sum2Map_sum2Map_sum1_12, addersMap_sum2Map_sum2Map_sum1_11, 
      addersMap_sum2Map_sum2Map_sum1_10, addersMap_sum2Map_sum2Map_sum1_9, 
      addersMap_sum2Map_sum2Map_sum1_8, addersMap_sum2Map_sum2Map_sum1_7, 
      addersMap_sum2Map_sum2Map_sum1_6, addersMap_sum2Map_sum2Map_sum1_5, 
      addersMap_sum2Map_sum2Map_sum1_4, addersMap_sum2Map_sum2Map_sum1_3, 
      addersMap_sum2Map_sum2Map_sum1_2, addersMap_sum2Map_sum2Map_sum1_1, 
      addersMap_sum2Map_sum2Map_sum1_0, addersMap_sum2Map_sum2Map_sum2_15, 
      addersMap_sum2Map_sum2Map_sum2_14, addersMap_sum2Map_sum2Map_sum2_13, 
      addersMap_sum2Map_sum2Map_sum2_12, addersMap_sum2Map_sum2Map_sum2_11, 
      addersMap_sum2Map_sum2Map_sum2_10, addersMap_sum2Map_sum2Map_sum2_9, 
      addersMap_sum2Map_sum2Map_sum2_8, addersMap_sum2Map_sum2Map_sum2_7, 
      addersMap_sum2Map_sum2Map_sum2_6, addersMap_sum2Map_sum2Map_sum2_5, 
      addersMap_sum2Map_sum2Map_sum2_4, addersMap_sum2Map_sum2Map_sum2_3, 
      addersMap_sum2Map_sum2Map_sum2_2, addersMap_sum2Map_sum2Map_sum2_1, 
      addersMap_sum2Map_sum2Map_sum2_0, addersMap_sum3Map_sum1_15, 
      addersMap_sum3Map_sum1_14, addersMap_sum3Map_sum1_13, 
      addersMap_sum3Map_sum1_12, addersMap_sum3Map_sum1_11, 
      addersMap_sum3Map_sum1_10, addersMap_sum3Map_sum1_9, 
      addersMap_sum3Map_sum1_8, addersMap_sum3Map_sum1_7, 
      addersMap_sum3Map_sum1_6, addersMap_sum3Map_sum1_5, 
      addersMap_sum3Map_sum1_4, addersMap_sum3Map_sum1_3, 
      addersMap_sum3Map_sum1_2, addersMap_sum3Map_sum1_1, 
      addersMap_sum3Map_sum1_0, addersMap_sum3Map_sum2_15, 
      addersMap_sum3Map_sum2_14, addersMap_sum3Map_sum2_13, 
      addersMap_sum3Map_sum2_12, addersMap_sum3Map_sum2_11, 
      addersMap_sum3Map_sum2_10, addersMap_sum3Map_sum2_9, 
      addersMap_sum3Map_sum2_8, addersMap_sum3Map_sum2_7, 
      addersMap_sum3Map_sum2_6, addersMap_sum3Map_sum2_5, 
      addersMap_sum3Map_sum2_4, addersMap_sum3Map_sum2_3, 
      addersMap_sum3Map_sum2_2, addersMap_sum3Map_sum2_1, 
      addersMap_sum3Map_sum2_0, addersMap_sum3Map_sum1Map_sum1_15, 
      addersMap_sum3Map_sum1Map_sum1_14, addersMap_sum3Map_sum1Map_sum1_13, 
      addersMap_sum3Map_sum1Map_sum1_12, addersMap_sum3Map_sum1Map_sum1_11, 
      addersMap_sum3Map_sum1Map_sum1_10, addersMap_sum3Map_sum1Map_sum1_9, 
      addersMap_sum3Map_sum1Map_sum1_8, addersMap_sum3Map_sum1Map_sum1_7, 
      addersMap_sum3Map_sum1Map_sum1_6, addersMap_sum3Map_sum1Map_sum1_5, 
      addersMap_sum3Map_sum1Map_sum1_4, addersMap_sum3Map_sum1Map_sum1_3, 
      addersMap_sum3Map_sum1Map_sum1_2, addersMap_sum3Map_sum1Map_sum1_1, 
      addersMap_sum3Map_sum1Map_sum1_0, addersMap_sum3Map_sum1Map_sum2_15, 
      addersMap_sum3Map_sum1Map_sum2_14, addersMap_sum3Map_sum1Map_sum2_13, 
      addersMap_sum3Map_sum1Map_sum2_12, addersMap_sum3Map_sum1Map_sum2_11, 
      addersMap_sum3Map_sum1Map_sum2_10, addersMap_sum3Map_sum1Map_sum2_9, 
      addersMap_sum3Map_sum1Map_sum2_8, addersMap_sum3Map_sum1Map_sum2_7, 
      addersMap_sum3Map_sum1Map_sum2_6, addersMap_sum3Map_sum1Map_sum2_5, 
      addersMap_sum3Map_sum1Map_sum2_4, addersMap_sum3Map_sum1Map_sum2_3, 
      addersMap_sum3Map_sum1Map_sum2_2, addersMap_sum3Map_sum1Map_sum2_1, 
      addersMap_sum3Map_sum1Map_sum2_0, addersMap_sum3Map_sum2Map_sum1_15, 
      addersMap_sum3Map_sum2Map_sum1_14, addersMap_sum3Map_sum2Map_sum1_13, 
      addersMap_sum3Map_sum2Map_sum1_12, addersMap_sum3Map_sum2Map_sum1_11, 
      addersMap_sum3Map_sum2Map_sum1_10, addersMap_sum3Map_sum2Map_sum1_9, 
      addersMap_sum3Map_sum2Map_sum1_8, addersMap_sum3Map_sum2Map_sum1_7, 
      addersMap_sum3Map_sum2Map_sum1_6, addersMap_sum3Map_sum2Map_sum1_5, 
      addersMap_sum3Map_sum2Map_sum1_4, addersMap_sum3Map_sum2Map_sum1_3, 
      addersMap_sum3Map_sum2Map_sum1_2, addersMap_sum3Map_sum2Map_sum1_1, 
      addersMap_sum3Map_sum2Map_sum1_0, addersMap_sum3Map_sum2Map_sum2_15, 
      addersMap_sum3Map_sum2Map_sum2_14, addersMap_sum3Map_sum2Map_sum2_13, 
      addersMap_sum3Map_sum2Map_sum2_12, addersMap_sum3Map_sum2Map_sum2_11, 
      addersMap_sum3Map_sum2Map_sum2_10, addersMap_sum3Map_sum2Map_sum2_9, 
      addersMap_sum3Map_sum2Map_sum2_8, addersMap_sum3Map_sum2Map_sum2_7, 
      addersMap_sum3Map_sum2Map_sum2_6, addersMap_sum3Map_sum2Map_sum2_5, 
      addersMap_sum3Map_sum2Map_sum2_4, addersMap_sum3Map_sum2Map_sum2_3, 
      addersMap_sum3Map_sum2Map_sum2_2, addersMap_sum3Map_sum2Map_sum2_1, 
      addersMap_sum3Map_sum2Map_sum2_0, outShifter_15, nx4, nx3412, nx3470, 
      nx2917, nx2923, nx2925, nx2929, nx2931, nx2935, nx2937, nx2941, nx2947, 
      nx2951, nx2959, nx2963, nx2971, nx2973, nx2979, nx2981, nx2985, nx2987, 
      nx2991, nx2993, nx2997, nx2999, nx3003, nx3005, nx3009, nx3011, nx3015, 
      nx3017, nx3021, nx3023, nx3027, nx3029, nx3033, nx3035, nx3039, nx3041, 
      nx3045, nx3047, nx3051, nx3053, nx3057, nx3059, nx3063, nx3065, nx3069, 
      nx3071, nx3075, nx3077, nx3081, nx3083, nx3087, nx3089, nx3093, nx3095, 
      nx3099, nx3101, nx3105, nx3107, nx3111, nx3113, nx3117, nx3119, nx3123, 
      nx3125, nx3129, nx3131, nx3135, nx3137, nx3141, nx3143, nx3147, nx3149, 
      nx3153, nx3155, nx3159, nx3161, nx3165, nx3167, nx3171, nx3173, nx3177, 
      nx3179, nx3183, nx3185, nx3189, nx3191, nx3195, nx3197, nx3201, nx3203, 
      nx3207, nx3209, nx3213, nx3215, nx3219, nx3221, nx3225, nx3227, nx3231, 
      nx3233, nx3237, nx3239, nx3243, nx3245, nx3249, nx3251, nx3255, nx3257, 
      nx3261, nx3263, nx3267, nx3269, nx3273, nx3275, nx3279, nx3281, nx3285, 
      nx3287, nx3291, nx3293, nx3297, nx3299, nx3303, nx3305, nx3309, nx3311, 
      nx3315, nx3317, nx3321, nx3323, nx3327, nx3329, nx3333, nx3335, nx3339, 
      nx3341, nx3345, nx3347, nx3351, nx3353, nx3357, nx3359, nx3363, nx3365, 
      nx3369, nx3371, nx3375, nx3377, nx3381, nx3383, nx3387, nx3389, nx3393, 
      nx3395, nx3399, nx3401, nx3405, nx3407, nx3411, nx3413, nx3417, nx3419, 
      nx3423, nx3425, nx3429, nx3431, nx3435, nx3437, nx3441, nx3443, nx3447, 
      nx3449, nx3453, nx3455, nx3459, nx3461, nx3465, nx3467, nx3471, nx3473, 
      nx3477, nx3479, nx3483, nx3485, nx3488, nx3490, nx3493, nx3495, nx3498, 
      nx3500, nx3503, nx3505, nx3508, nx3510, nx3513, nx3515, nx3518, nx3520, 
      nx3523, nx3525, nx3528, nx3530, nx3533, nx3535, nx3538, nx3540, nx3543, 
      nx3545, nx3548, nx3550, nx3553, nx3555, nx3558, nx3560, nx3563, nx3565, 
      nx3568, nx3570, nx3573, nx3575, nx3578, nx3580, nx3583, nx3585, nx3588, 
      nx3590, nx3593, nx3595, nx3598, nx3600, nx3603, nx3605, nx3608, nx3610, 
      nx3613, nx3615, nx3618, nx3620, nx3623, nx3625, nx3628, nx3630, nx3633, 
      nx3635, nx3638, nx3640, nx3643, nx3645, nx3648, nx3650, nx3653, nx3655, 
      nx3658, nx3660, nx3663, nx3665, nx3668, nx3670, nx3673, nx3675, nx3678, 
      nx3680, nx3683, nx3685, nx3688, nx3690, nx3693, nx3695, nx3698, nx3700, 
      nx3703, nx3705, nx3708, nx3710, nx3713, nx3715, nx3718, nx3720, nx3723, 
      nx3725, nx3728, nx3730, nx3733, nx3735, nx3738, nx3740, nx3743, nx3745, 
      nx3748, nx3750, nx3753, nx3755, nx3758, nx3760, nx3763, nx3765, nx3768, 
      nx3770, nx3773, nx3775, nx3778, nx3780, nx3783, nx3785, nx3788, nx3790, 
      nx3793, nx3795, nx3798, nx3800, nx3803, nx3805, nx3808, nx3810, nx3813, 
      nx3815, nx3818, nx3820, nx3823, nx3825, nx3828, nx3830, nx3833, nx3835, 
      nx3838, nx3840, nx3843, nx3845, nx3848, nx3850, nx3853, nx3855, nx3858, 
      nx3860, nx3863, nx3865, nx3868, nx3870, nx3873, nx3875, nx3878, nx3880, 
      nx3883, nx3885, nx3888, nx3890, nx3893, nx3895, nx3898, nx3900, nx3903, 
      nx3905, nx3908, nx3910, nx3913, nx3915, nx3918, nx3920, nx3923, nx3925, 
      nx3928, nx3930, nx3933, nx3935, nx3938, nx3940, nx3943, nx3945, nx3948, 
      nx3950, nx3953, nx3955, nx3958, nx3960, nx3963, nx3965, nx3968, nx3970, 
      nx3973, nx3975, nx3978, nx3980, nx3983, nx3985, nx3988, nx3990, nx3993, 
      nx3995, nx3998, nx4000, nx4003, nx4005, nx4008, nx4010, nx4013, nx4015, 
      nx4018, nx4020, nx4023, nx4025, nx4028, nx4030, nx4033, nx4035, nx4038, 
      nx4040, nx4043, nx4045, nx4048, nx4050, nx4053, nx4055, nx4058, nx4060, 
      nx4063, nx4065, nx4068, nx4070, nx4073, nx4075, nx4078, nx4080, nx4083, 
      nx4085, nx4088, nx4090, nx4093, nx4095, nx4098, nx4100, nx4103, nx4105, 
      nx4108, nx4110, nx4113, nx4115, nx4118, nx4120, nx4123, nx4125, nx4128, 
      nx4130, nx4133, nx4135, nx4138, nx4140, nx4143, nx4145, nx4148, nx4150, 
      nx4153, nx4155, nx4158, nx4160, nx4163, nx4165, nx4168, nx4170, nx4173, 
      nx4175, nx4178, nx4180, nx4183, nx4185, nx4188, nx4190, nx4193, nx4195, 
      nx4198, nx4200, nx4203, nx4205, nx4208, nx4210, nx4213, nx4215, nx4218, 
      nx4220, nx4223, nx4225, nx4228, nx4230, nx4233, nx4235, nx4238, nx4240, 
      nx4243, nx4245, nx4248, nx4250, nx4253, nx4255, nx4258, nx4260, nx4263, 
      nx4265, nx4268, nx4270, nx4273, nx4275, nx4278, nx4280, nx4283, nx4285, 
      nx4288, nx4290, nx4293, nx4295, nx4298, nx4300, nx4303, nx4305, nx4308, 
      nx4310, nx4313, nx4315, nx4318, nx4320, nx4323, nx4325, nx4328, nx4330, 
      nx4333, nx4335, nx4338, nx4340, nx4343, nx4345, nx4348, nx4350, nx4353, 
      nx4355, nx4358, nx4360, nx4363, nx4365, nx4368, nx4370, nx4373, nx4375, 
      nx4378, nx4380, nx4383, nx4385, nx4388, nx4390, nx4393, nx4395, nx4398, 
      nx4400, nx4403, nx4405, nx4408, nx4410, nx4413, nx4415, nx4418, nx4420, 
      nx4423, nx4425, nx4428, nx4430, nx4433, nx4435, nx4438, nx4440, nx4443, 
      nx4445, nx4448, nx4450, nx4453, nx4455, nx4458, nx4460, nx4463, nx4465, 
      nx4468, nx4470, nx4473, nx4475, nx4478, nx4480, nx4483, nx4485, nx4488, 
      nx4490, nx4493, nx4495, nx4498, nx4500, nx4503, nx4505, nx4508, nx4510, 
      nx4513, nx4515, nx4518, nx4520, nx4523, nx4525, nx4528, nx4530, nx4533, 
      nx4535, nx4538, nx4540, nx4543, nx4545, nx4548, nx4550, nx4553, nx4555, 
      nx4558, nx4560, nx4563, nx4565, nx4568, nx4570, nx4573, nx4575, nx4578, 
      nx4580, nx4583, nx4585, nx4588, nx4590, nx4593, nx4595, nx4598, nx4600, 
      nx4603, nx4605, nx4608, nx4610, nx4613, nx4615, nx4618, nx4620, nx4623, 
      nx4625, nx4628, nx4630, nx4633, nx4635, nx4638, nx4640, nx4643, nx4645, 
      nx4648, nx4650, nx4653, nx4655, nx4658, nx4660, nx4663, nx4665, nx4668, 
      nx4670, nx4673, nx4675, nx4678, nx4680, nx4683, nx4685, nx4688, nx4690, 
      nx4693, nx4695, nx4698, nx4700, nx4703, nx4705, nx4708, nx4710, nx4713, 
      nx4715, nx4718, nx4720, nx4723, nx4725, nx4728, nx4730, nx4733, nx4735, 
      nx4738, nx4740, nx4743, nx4745, nx4748, nx4750, nx4753, nx4755, nx4758, 
      nx4760, nx4763, nx4765, nx4768, nx4770, nx4773, nx4775, nx4778, nx4780, 
      nx4783, nx4785, nx4788, nx4790, nx4793, nx4795, nx4798, nx4800, nx4803, 
      nx4805, nx4808, nx4810, nx4813, nx4815, nx4818, nx4820, nx4823, nx4825, 
      nx4828, nx4830, nx4833, nx4835, nx4838, nx4840, nx4843, nx4845, nx4848, 
      nx4850, nx4853, nx4855, nx4858, nx4860, nx4863, nx4865, nx4868, nx4870, 
      nx4873, nx4875, nx4878, nx4880, nx4883, nx4885, nx4888, nx4890, nx4893, 
      nx4895, nx4898, nx4900, nx4903, nx4905, nx4908, nx4910, nx4913, nx4915, 
      nx4918, nx4920, nx4923, nx4925, nx4928, nx4930, nx4933, nx4935, nx4938, 
      nx4940, nx4943, nx4945, nx4948, nx4950, nx4953, nx4955, nx4958, nx4960, 
      nx4963, nx4965, nx4968, nx4970, nx4973, nx4975, nx4978, nx4980, nx4983, 
      nx4985, nx4988, nx4990, nx4993, nx4995, nx4998, nx5000, nx5003, nx5005, 
      nx5008, nx5010, nx5013, nx5015, nx5018, nx5020, nx5023, nx5025, nx5028, 
      nx5030, nx5033, nx5035, nx5038, nx5040, nx5043, nx5045, nx5048, nx5050, 
      nx5053, nx5055, nx5058, nx5060, nx5063, nx5067, nx5070, nx5072, nx5074, 
      nx5076, nx5079, nx5081, nx5083, nx5085, nx5088, nx5090, nx5092, nx5094, 
      nx5097, nx5099, nx5101, nx5103, nx5106, nx5108, nx5110, nx5112, nx5115, 
      nx5117, nx5119, nx5121, nx5124, nx5126, nx5128, nx5130, nx5133, nx5135, 
      nx5137, nx5139, nx5142, nx5144, nx5146, nx5148, nx5151, nx5153, nx5155, 
      nx5157, nx5160, nx5162, nx5164, nx5167, nx5169, nx5171, nx5174, nx5176, 
      nx5179, nx5181, nx5184, nx5186, nx5189, nx5196, nx5198, nx5200, nx5202, 
      nx5204, nx5206, nx5208, nx5210, nx5212, nx5214, nx5216, nx5218, nx5220, 
      nx5222, nx5224, nx5226, nx5228, nx5230, nx5232, nx5234, nx5236, nx5238, 
      nx5240, nx5242, nx5244, nx5246, nx5248, nx5250, nx5252, nx5254, nx5256, 
      nx5258, nx5260, nx5262, nx5264, nx5266, nx5268, nx5270, nx5272, nx5274, 
      nx5276, nx5278, nx5280, nx5282, nx5284, nx5286, nx5288, nx5290, nx5292, 
      nx5294, nx5296, nx5298, nx5300, nx5302, nx5304, nx5306, nx5308, nx5310, 
      nx5312, nx5314, nx5316, nx5318, nx5320, nx5322, nx5328, nx5330, nx5332, 
      nx5334, nx5336, nx5338, nx5340, nx5342, nx5344, nx5346: std_logic ;
   
   signal DANGLING : std_logic_vector (184 downto 0 );

begin
   mulsMap : CNNMuls_25 port map ( filter_24_7=>filter_0_7, filter_24_6=>
      filter_0_6, filter_24_5=>filter_0_5, filter_24_4=>filter_0_4, 
      filter_24_3=>filter_0_3, filter_24_2=>filter_0_2, filter_24_1=>
      filter_0_1, filter_24_0=>filter_0_0, filter_23_7=>filter_1_7, 
      filter_23_6=>filter_1_6, filter_23_5=>filter_1_5, filter_23_4=>
      filter_1_4, filter_23_3=>filter_1_3, filter_23_2=>filter_1_2, 
      filter_23_1=>filter_1_1, filter_23_0=>filter_1_0, filter_22_7=>
      filter_2_7, filter_22_6=>filter_2_6, filter_22_5=>filter_2_5, 
      filter_22_4=>filter_2_4, filter_22_3=>filter_2_3, filter_22_2=>
      filter_2_2, filter_22_1=>filter_2_1, filter_22_0=>filter_2_0, 
      filter_21_7=>filter_3_7, filter_21_6=>filter_3_6, filter_21_5=>
      filter_3_5, filter_21_4=>filter_3_4, filter_21_3=>filter_3_3, 
      filter_21_2=>filter_3_2, filter_21_1=>filter_3_1, filter_21_0=>
      filter_3_0, filter_20_7=>filter_4_7, filter_20_6=>filter_4_6, 
      filter_20_5=>filter_4_5, filter_20_4=>filter_4_4, filter_20_3=>
      filter_4_3, filter_20_2=>filter_4_2, filter_20_1=>filter_4_1, 
      filter_20_0=>filter_4_0, filter_19_7=>filter_5_7, filter_19_6=>
      filter_5_6, filter_19_5=>filter_5_5, filter_19_4=>filter_5_4, 
      filter_19_3=>filter_5_3, filter_19_2=>filter_5_2, filter_19_1=>
      filter_5_1, filter_19_0=>filter_5_0, filter_18_7=>filter_6_7, 
      filter_18_6=>filter_6_6, filter_18_5=>filter_6_5, filter_18_4=>
      filter_6_4, filter_18_3=>filter_6_3, filter_18_2=>filter_6_2, 
      filter_18_1=>filter_6_1, filter_18_0=>filter_6_0, filter_17_7=>
      filter_7_7, filter_17_6=>filter_7_6, filter_17_5=>filter_7_5, 
      filter_17_4=>filter_7_4, filter_17_3=>filter_7_3, filter_17_2=>
      filter_7_2, filter_17_1=>filter_7_1, filter_17_0=>filter_7_0, 
      filter_16_7=>filter_8_7, filter_16_6=>filter_8_6, filter_16_5=>
      filter_8_5, filter_16_4=>filter_8_4, filter_16_3=>filter_8_3, 
      filter_16_2=>filter_8_2, filter_16_1=>filter_8_1, filter_16_0=>
      filter_8_0, filter_15_7=>filter_9_7, filter_15_6=>filter_9_6, 
      filter_15_5=>filter_9_5, filter_15_4=>filter_9_4, filter_15_3=>
      filter_9_3, filter_15_2=>filter_9_2, filter_15_1=>filter_9_1, 
      filter_15_0=>filter_9_0, filter_14_7=>filter_10_7, filter_14_6=>
      filter_10_6, filter_14_5=>filter_10_5, filter_14_4=>filter_10_4, 
      filter_14_3=>filter_10_3, filter_14_2=>filter_10_2, filter_14_1=>
      filter_10_1, filter_14_0=>filter_10_0, filter_13_7=>filter_11_7, 
      filter_13_6=>filter_11_6, filter_13_5=>filter_11_5, filter_13_4=>
      filter_11_4, filter_13_3=>filter_11_3, filter_13_2=>filter_11_2, 
      filter_13_1=>filter_11_1, filter_13_0=>filter_11_0, filter_12_7=>
      filter_12_7, filter_12_6=>filter_12_6, filter_12_5=>filter_12_5, 
      filter_12_4=>filter_12_4, filter_12_3=>filter_12_3, filter_12_2=>
      filter_12_2, filter_12_1=>filter_12_1, filter_12_0=>filter_12_0, 
      filter_11_7=>filter_13_7, filter_11_6=>filter_13_6, filter_11_5=>
      filter_13_5, filter_11_4=>filter_13_4, filter_11_3=>filter_13_3, 
      filter_11_2=>filter_13_2, filter_11_1=>filter_13_1, filter_11_0=>
      filter_13_0, filter_10_7=>filter_14_7, filter_10_6=>filter_14_6, 
      filter_10_5=>filter_14_5, filter_10_4=>filter_14_4, filter_10_3=>
      filter_14_3, filter_10_2=>filter_14_2, filter_10_1=>filter_14_1, 
      filter_10_0=>filter_14_0, filter_9_7=>filter_15_7, filter_9_6=>
      filter_15_6, filter_9_5=>filter_15_5, filter_9_4=>filter_15_4, 
      filter_9_3=>filter_15_3, filter_9_2=>filter_15_2, filter_9_1=>
      filter_15_1, filter_9_0=>filter_15_0, filter_8_7=>filter_16_7, 
      filter_8_6=>filter_16_6, filter_8_5=>filter_16_5, filter_8_4=>
      filter_16_4, filter_8_3=>filter_16_3, filter_8_2=>filter_16_2, 
      filter_8_1=>filter_16_1, filter_8_0=>filter_16_0, filter_7_7=>
      filter_17_7, filter_7_6=>filter_17_6, filter_7_5=>filter_17_5, 
      filter_7_4=>filter_17_4, filter_7_3=>filter_17_3, filter_7_2=>
      filter_17_2, filter_7_1=>filter_17_1, filter_7_0=>filter_17_0, 
      filter_6_7=>filter_18_7, filter_6_6=>filter_18_6, filter_6_5=>
      filter_18_5, filter_6_4=>filter_18_4, filter_6_3=>filter_18_3, 
      filter_6_2=>filter_18_2, filter_6_1=>filter_18_1, filter_6_0=>
      filter_18_0, filter_5_7=>filter_19_7, filter_5_6=>filter_19_6, 
      filter_5_5=>filter_19_5, filter_5_4=>filter_19_4, filter_5_3=>
      filter_19_3, filter_5_2=>filter_19_2, filter_5_1=>filter_19_1, 
      filter_5_0=>filter_19_0, filter_4_7=>filter_20_7, filter_4_6=>
      filter_20_6, filter_4_5=>filter_20_5, filter_4_4=>filter_20_4, 
      filter_4_3=>filter_20_3, filter_4_2=>filter_20_2, filter_4_1=>
      filter_20_1, filter_4_0=>filter_20_0, filter_3_7=>filter_21_7, 
      filter_3_6=>filter_21_6, filter_3_5=>filter_21_5, filter_3_4=>
      filter_21_4, filter_3_3=>filter_21_3, filter_3_2=>filter_21_2, 
      filter_3_1=>filter_21_1, filter_3_0=>filter_21_0, filter_2_7=>
      filter_22_7, filter_2_6=>filter_22_6, filter_2_5=>filter_22_5, 
      filter_2_4=>filter_22_4, filter_2_3=>filter_22_3, filter_2_2=>
      filter_22_2, filter_2_1=>filter_22_1, filter_2_0=>filter_22_0, 
      filter_1_7=>filter_23_7, filter_1_6=>filter_23_6, filter_1_5=>
      filter_23_5, filter_1_4=>filter_23_4, filter_1_3=>filter_23_3, 
      filter_1_2=>filter_23_2, filter_1_1=>filter_23_1, filter_1_0=>
      filter_23_0, filter_0_7=>filter_24_7, filter_0_6=>filter_24_6, 
      filter_0_5=>filter_24_5, filter_0_4=>filter_24_4, filter_0_3=>
      filter_24_3, filter_0_2=>filter_24_2, filter_0_1=>filter_24_1, 
      filter_0_0=>filter_24_0, window_24_15=>currentPage_0_15, window_24_14
      =>currentPage_0_14, window_24_13=>currentPage_0_13, window_24_12=>
      currentPage_0_12, window_24_11=>currentPage_0_11, window_24_10=>
      currentPage_0_10, window_24_9=>currentPage_0_9, window_24_8=>
      currentPage_0_8, window_24_7=>currentPage_0_7, window_24_6=>
      currentPage_0_6, window_24_5=>currentPage_0_5, window_24_4=>
      currentPage_0_4, window_24_3=>currentPage_0_3, window_24_2=>
      currentPage_0_2, window_24_1=>currentPage_0_1, window_24_0=>
      currentPage_0_0, window_23_15=>currentPage_1_15, window_23_14=>
      currentPage_1_14, window_23_13=>currentPage_1_13, window_23_12=>
      currentPage_1_12, window_23_11=>currentPage_1_11, window_23_10=>
      currentPage_1_10, window_23_9=>currentPage_1_9, window_23_8=>
      currentPage_1_8, window_23_7=>currentPage_1_7, window_23_6=>
      currentPage_1_6, window_23_5=>currentPage_1_5, window_23_4=>
      currentPage_1_4, window_23_3=>currentPage_1_3, window_23_2=>
      currentPage_1_2, window_23_1=>currentPage_1_1, window_23_0=>
      currentPage_1_0, window_22_15=>currentPage_2_15, window_22_14=>
      currentPage_2_14, window_22_13=>currentPage_2_13, window_22_12=>
      currentPage_2_12, window_22_11=>currentPage_2_11, window_22_10=>
      currentPage_2_10, window_22_9=>currentPage_2_9, window_22_8=>
      currentPage_2_8, window_22_7=>currentPage_2_7, window_22_6=>
      currentPage_2_6, window_22_5=>currentPage_2_5, window_22_4=>
      currentPage_2_4, window_22_3=>currentPage_2_3, window_22_2=>
      currentPage_2_2, window_22_1=>currentPage_2_1, window_22_0=>
      currentPage_2_0, window_21_15=>currentPage_3_15, window_21_14=>
      currentPage_3_14, window_21_13=>currentPage_3_13, window_21_12=>
      currentPage_3_12, window_21_11=>currentPage_3_11, window_21_10=>
      currentPage_3_10, window_21_9=>currentPage_3_9, window_21_8=>
      currentPage_3_8, window_21_7=>currentPage_3_7, window_21_6=>
      currentPage_3_6, window_21_5=>currentPage_3_5, window_21_4=>
      currentPage_3_4, window_21_3=>currentPage_3_3, window_21_2=>
      currentPage_3_2, window_21_1=>currentPage_3_1, window_21_0=>
      currentPage_3_0, window_20_15=>currentPage_4_15, window_20_14=>
      currentPage_4_14, window_20_13=>currentPage_4_13, window_20_12=>
      currentPage_4_12, window_20_11=>currentPage_4_11, window_20_10=>
      currentPage_4_10, window_20_9=>currentPage_4_9, window_20_8=>
      currentPage_4_8, window_20_7=>currentPage_4_7, window_20_6=>
      currentPage_4_6, window_20_5=>currentPage_4_5, window_20_4=>
      currentPage_4_4, window_20_3=>currentPage_4_3, window_20_2=>
      currentPage_4_2, window_20_1=>currentPage_4_1, window_20_0=>
      currentPage_4_0, window_19_15=>currentPage_5_15, window_19_14=>
      currentPage_5_14, window_19_13=>currentPage_5_13, window_19_12=>
      currentPage_5_12, window_19_11=>currentPage_5_11, window_19_10=>
      currentPage_5_10, window_19_9=>currentPage_5_9, window_19_8=>
      currentPage_5_8, window_19_7=>currentPage_5_7, window_19_6=>
      currentPage_5_6, window_19_5=>currentPage_5_5, window_19_4=>
      currentPage_5_4, window_19_3=>currentPage_5_3, window_19_2=>
      currentPage_5_2, window_19_1=>currentPage_5_1, window_19_0=>
      currentPage_5_0, window_18_15=>currentPage_6_15, window_18_14=>
      currentPage_6_14, window_18_13=>currentPage_6_13, window_18_12=>
      currentPage_6_12, window_18_11=>currentPage_6_11, window_18_10=>
      currentPage_6_10, window_18_9=>currentPage_6_9, window_18_8=>
      currentPage_6_8, window_18_7=>currentPage_6_7, window_18_6=>
      currentPage_6_6, window_18_5=>currentPage_6_5, window_18_4=>
      currentPage_6_4, window_18_3=>currentPage_6_3, window_18_2=>
      currentPage_6_2, window_18_1=>currentPage_6_1, window_18_0=>
      currentPage_6_0, window_17_15=>currentPage_7_15, window_17_14=>
      currentPage_7_14, window_17_13=>currentPage_7_13, window_17_12=>
      currentPage_7_12, window_17_11=>currentPage_7_11, window_17_10=>
      currentPage_7_10, window_17_9=>currentPage_7_9, window_17_8=>
      currentPage_7_8, window_17_7=>currentPage_7_7, window_17_6=>
      currentPage_7_6, window_17_5=>currentPage_7_5, window_17_4=>
      currentPage_7_4, window_17_3=>currentPage_7_3, window_17_2=>
      currentPage_7_2, window_17_1=>currentPage_7_1, window_17_0=>
      currentPage_7_0, window_16_15=>currentPage_8_15, window_16_14=>
      currentPage_8_14, window_16_13=>currentPage_8_13, window_16_12=>
      currentPage_8_12, window_16_11=>currentPage_8_11, window_16_10=>
      currentPage_8_10, window_16_9=>currentPage_8_9, window_16_8=>
      currentPage_8_8, window_16_7=>currentPage_8_7, window_16_6=>
      currentPage_8_6, window_16_5=>currentPage_8_5, window_16_4=>
      currentPage_8_4, window_16_3=>currentPage_8_3, window_16_2=>
      currentPage_8_2, window_16_1=>currentPage_8_1, window_16_0=>
      currentPage_8_0, window_15_15=>currentPage_9_15, window_15_14=>
      currentPage_9_14, window_15_13=>currentPage_9_13, window_15_12=>
      currentPage_9_12, window_15_11=>currentPage_9_11, window_15_10=>
      currentPage_9_10, window_15_9=>currentPage_9_9, window_15_8=>
      currentPage_9_8, window_15_7=>currentPage_9_7, window_15_6=>
      currentPage_9_6, window_15_5=>currentPage_9_5, window_15_4=>
      currentPage_9_4, window_15_3=>currentPage_9_3, window_15_2=>
      currentPage_9_2, window_15_1=>currentPage_9_1, window_15_0=>
      currentPage_9_0, window_14_15=>currentPage_10_15, window_14_14=>
      currentPage_10_14, window_14_13=>currentPage_10_13, window_14_12=>
      currentPage_10_12, window_14_11=>currentPage_10_11, window_14_10=>
      currentPage_10_10, window_14_9=>currentPage_10_9, window_14_8=>
      currentPage_10_8, window_14_7=>currentPage_10_7, window_14_6=>
      currentPage_10_6, window_14_5=>currentPage_10_5, window_14_4=>
      currentPage_10_4, window_14_3=>currentPage_10_3, window_14_2=>
      currentPage_10_2, window_14_1=>currentPage_10_1, window_14_0=>
      currentPage_10_0, window_13_15=>currentPage_11_15, window_13_14=>
      currentPage_11_14, window_13_13=>currentPage_11_13, window_13_12=>
      currentPage_11_12, window_13_11=>currentPage_11_11, window_13_10=>
      currentPage_11_10, window_13_9=>currentPage_11_9, window_13_8=>
      currentPage_11_8, window_13_7=>currentPage_11_7, window_13_6=>
      currentPage_11_6, window_13_5=>currentPage_11_5, window_13_4=>
      currentPage_11_4, window_13_3=>currentPage_11_3, window_13_2=>
      currentPage_11_2, window_13_1=>currentPage_11_1, window_13_0=>
      currentPage_11_0, window_12_15=>currentPage_12_15, window_12_14=>
      currentPage_12_14, window_12_13=>currentPage_12_13, window_12_12=>
      currentPage_12_12, window_12_11=>currentPage_12_11, window_12_10=>
      currentPage_12_10, window_12_9=>currentPage_12_9, window_12_8=>
      currentPage_12_8, window_12_7=>currentPage_12_7, window_12_6=>
      currentPage_12_6, window_12_5=>currentPage_12_5, window_12_4=>
      currentPage_12_4, window_12_3=>currentPage_12_3, window_12_2=>
      currentPage_12_2, window_12_1=>currentPage_12_1, window_12_0=>
      currentPage_12_0, window_11_15=>currentPage_13_15, window_11_14=>
      currentPage_13_14, window_11_13=>currentPage_13_13, window_11_12=>
      currentPage_13_12, window_11_11=>currentPage_13_11, window_11_10=>
      currentPage_13_10, window_11_9=>currentPage_13_9, window_11_8=>
      currentPage_13_8, window_11_7=>currentPage_13_7, window_11_6=>
      currentPage_13_6, window_11_5=>currentPage_13_5, window_11_4=>
      currentPage_13_4, window_11_3=>currentPage_13_3, window_11_2=>
      currentPage_13_2, window_11_1=>currentPage_13_1, window_11_0=>
      currentPage_13_0, window_10_15=>currentPage_14_15, window_10_14=>
      currentPage_14_14, window_10_13=>currentPage_14_13, window_10_12=>
      currentPage_14_12, window_10_11=>currentPage_14_11, window_10_10=>
      currentPage_14_10, window_10_9=>currentPage_14_9, window_10_8=>
      currentPage_14_8, window_10_7=>currentPage_14_7, window_10_6=>
      currentPage_14_6, window_10_5=>currentPage_14_5, window_10_4=>
      currentPage_14_4, window_10_3=>currentPage_14_3, window_10_2=>
      currentPage_14_2, window_10_1=>currentPage_14_1, window_10_0=>
      currentPage_14_0, window_9_15=>currentPage_15_15, window_9_14=>
      currentPage_15_14, window_9_13=>currentPage_15_13, window_9_12=>
      currentPage_15_12, window_9_11=>currentPage_15_11, window_9_10=>
      currentPage_15_10, window_9_9=>currentPage_15_9, window_9_8=>
      currentPage_15_8, window_9_7=>currentPage_15_7, window_9_6=>
      currentPage_15_6, window_9_5=>currentPage_15_5, window_9_4=>
      currentPage_15_4, window_9_3=>currentPage_15_3, window_9_2=>
      currentPage_15_2, window_9_1=>currentPage_15_1, window_9_0=>
      currentPage_15_0, window_8_15=>currentPage_16_15, window_8_14=>
      currentPage_16_14, window_8_13=>currentPage_16_13, window_8_12=>
      currentPage_16_12, window_8_11=>currentPage_16_11, window_8_10=>
      currentPage_16_10, window_8_9=>currentPage_16_9, window_8_8=>
      currentPage_16_8, window_8_7=>currentPage_16_7, window_8_6=>
      currentPage_16_6, window_8_5=>currentPage_16_5, window_8_4=>
      currentPage_16_4, window_8_3=>currentPage_16_3, window_8_2=>
      currentPage_16_2, window_8_1=>currentPage_16_1, window_8_0=>
      currentPage_16_0, window_7_15=>currentPage_17_15, window_7_14=>
      currentPage_17_14, window_7_13=>currentPage_17_13, window_7_12=>
      currentPage_17_12, window_7_11=>currentPage_17_11, window_7_10=>
      currentPage_17_10, window_7_9=>currentPage_17_9, window_7_8=>
      currentPage_17_8, window_7_7=>currentPage_17_7, window_7_6=>
      currentPage_17_6, window_7_5=>currentPage_17_5, window_7_4=>
      currentPage_17_4, window_7_3=>currentPage_17_3, window_7_2=>
      currentPage_17_2, window_7_1=>currentPage_17_1, window_7_0=>
      currentPage_17_0, window_6_15=>currentPage_18_15, window_6_14=>
      currentPage_18_14, window_6_13=>currentPage_18_13, window_6_12=>
      currentPage_18_12, window_6_11=>currentPage_18_11, window_6_10=>
      currentPage_18_10, window_6_9=>currentPage_18_9, window_6_8=>
      currentPage_18_8, window_6_7=>currentPage_18_7, window_6_6=>
      currentPage_18_6, window_6_5=>currentPage_18_5, window_6_4=>
      currentPage_18_4, window_6_3=>currentPage_18_3, window_6_2=>
      currentPage_18_2, window_6_1=>currentPage_18_1, window_6_0=>
      currentPage_18_0, window_5_15=>currentPage_19_15, window_5_14=>
      currentPage_19_14, window_5_13=>currentPage_19_13, window_5_12=>
      currentPage_19_12, window_5_11=>currentPage_19_11, window_5_10=>
      currentPage_19_10, window_5_9=>currentPage_19_9, window_5_8=>
      currentPage_19_8, window_5_7=>currentPage_19_7, window_5_6=>
      currentPage_19_6, window_5_5=>currentPage_19_5, window_5_4=>
      currentPage_19_4, window_5_3=>currentPage_19_3, window_5_2=>
      currentPage_19_2, window_5_1=>currentPage_19_1, window_5_0=>
      currentPage_19_0, window_4_15=>currentPage_20_15, window_4_14=>
      currentPage_20_14, window_4_13=>currentPage_20_13, window_4_12=>
      currentPage_20_12, window_4_11=>currentPage_20_11, window_4_10=>
      currentPage_20_10, window_4_9=>currentPage_20_9, window_4_8=>
      currentPage_20_8, window_4_7=>currentPage_20_7, window_4_6=>
      currentPage_20_6, window_4_5=>currentPage_20_5, window_4_4=>
      currentPage_20_4, window_4_3=>currentPage_20_3, window_4_2=>
      currentPage_20_2, window_4_1=>currentPage_20_1, window_4_0=>
      currentPage_20_0, window_3_15=>currentPage_21_15, window_3_14=>
      currentPage_21_14, window_3_13=>currentPage_21_13, window_3_12=>
      currentPage_21_12, window_3_11=>currentPage_21_11, window_3_10=>
      currentPage_21_10, window_3_9=>currentPage_21_9, window_3_8=>
      currentPage_21_8, window_3_7=>currentPage_21_7, window_3_6=>
      currentPage_21_6, window_3_5=>currentPage_21_5, window_3_4=>
      currentPage_21_4, window_3_3=>currentPage_21_3, window_3_2=>
      currentPage_21_2, window_3_1=>currentPage_21_1, window_3_0=>
      currentPage_21_0, window_2_15=>currentPage_22_15, window_2_14=>
      currentPage_22_14, window_2_13=>currentPage_22_13, window_2_12=>
      currentPage_22_12, window_2_11=>currentPage_22_11, window_2_10=>
      currentPage_22_10, window_2_9=>currentPage_22_9, window_2_8=>
      currentPage_22_8, window_2_7=>currentPage_22_7, window_2_6=>
      currentPage_22_6, window_2_5=>currentPage_22_5, window_2_4=>
      currentPage_22_4, window_2_3=>currentPage_22_3, window_2_2=>
      currentPage_22_2, window_2_1=>currentPage_22_1, window_2_0=>
      currentPage_22_0, window_1_15=>currentPage_23_15, window_1_14=>
      currentPage_23_14, window_1_13=>currentPage_23_13, window_1_12=>
      currentPage_23_12, window_1_11=>currentPage_23_11, window_1_10=>
      currentPage_23_10, window_1_9=>currentPage_23_9, window_1_8=>
      currentPage_23_8, window_1_7=>currentPage_23_7, window_1_6=>
      currentPage_23_6, window_1_5=>currentPage_23_5, window_1_4=>
      currentPage_23_4, window_1_3=>currentPage_23_3, window_1_2=>
      currentPage_23_2, window_1_1=>currentPage_23_1, window_1_0=>
      currentPage_23_0, window_0_15=>currentPage_24_15, window_0_14=>
      currentPage_24_14, window_0_13=>currentPage_24_13, window_0_12=>
      currentPage_24_12, window_0_11=>currentPage_24_11, window_0_10=>
      currentPage_24_10, window_0_9=>currentPage_24_9, window_0_8=>
      currentPage_24_8, window_0_7=>currentPage_24_7, window_0_6=>
      currentPage_24_6, window_0_5=>currentPage_24_5, window_0_4=>
      currentPage_24_4, window_0_3=>currentPage_24_3, window_0_2=>
      currentPage_24_2, window_0_1=>currentPage_24_1, window_0_0=>
      currentPage_24_0, outputs_24_15=>outMuls_0_15, outputs_24_14=>
      outMuls_0_14, outputs_24_13=>outMuls_0_13, outputs_24_12=>outMuls_0_12, 
      outputs_24_11=>outMuls_0_11, outputs_24_10=>outMuls_0_10, outputs_24_9
      =>outMuls_0_9, outputs_24_8=>outMuls_0_8, outputs_24_7=>outMuls_0_7, 
      outputs_24_6=>outMuls_0_6, outputs_24_5=>outMuls_0_5, outputs_24_4=>
      outMuls_0_4, outputs_24_3=>outMuls_0_3, outputs_24_2=>outMuls_0_2, 
      outputs_24_1=>outMuls_0_1, outputs_24_0=>outMuls_0_0, outputs_23_15=>
      outMuls_1_15, outputs_23_14=>outMuls_1_14, outputs_23_13=>outMuls_1_13, 
      outputs_23_12=>outMuls_1_12, outputs_23_11=>outMuls_1_11, 
      outputs_23_10=>outMuls_1_10, outputs_23_9=>outMuls_1_9, outputs_23_8=>
      outMuls_1_8, outputs_23_7=>outMuls_1_7, outputs_23_6=>outMuls_1_6, 
      outputs_23_5=>outMuls_1_5, outputs_23_4=>outMuls_1_4, outputs_23_3=>
      outMuls_1_3, outputs_23_2=>outMuls_1_2, outputs_23_1=>outMuls_1_1, 
      outputs_23_0=>outMuls_1_0, outputs_22_15=>outMuls_2_15, outputs_22_14
      =>outMuls_2_14, outputs_22_13=>outMuls_2_13, outputs_22_12=>
      outMuls_2_12, outputs_22_11=>outMuls_2_11, outputs_22_10=>outMuls_2_10, 
      outputs_22_9=>outMuls_2_9, outputs_22_8=>outMuls_2_8, outputs_22_7=>
      outMuls_2_7, outputs_22_6=>outMuls_2_6, outputs_22_5=>outMuls_2_5, 
      outputs_22_4=>outMuls_2_4, outputs_22_3=>outMuls_2_3, outputs_22_2=>
      outMuls_2_2, outputs_22_1=>outMuls_2_1, outputs_22_0=>outMuls_2_0, 
      outputs_21_15=>outMuls_3_15, outputs_21_14=>outMuls_3_14, 
      outputs_21_13=>outMuls_3_13, outputs_21_12=>outMuls_3_12, 
      outputs_21_11=>outMuls_3_11, outputs_21_10=>outMuls_3_10, outputs_21_9
      =>outMuls_3_9, outputs_21_8=>outMuls_3_8, outputs_21_7=>outMuls_3_7, 
      outputs_21_6=>outMuls_3_6, outputs_21_5=>outMuls_3_5, outputs_21_4=>
      outMuls_3_4, outputs_21_3=>outMuls_3_3, outputs_21_2=>outMuls_3_2, 
      outputs_21_1=>outMuls_3_1, outputs_21_0=>outMuls_3_0, outputs_20_15=>
      outMuls_4_15, outputs_20_14=>outMuls_4_14, outputs_20_13=>outMuls_4_13, 
      outputs_20_12=>outMuls_4_12, outputs_20_11=>outMuls_4_11, 
      outputs_20_10=>outMuls_4_10, outputs_20_9=>outMuls_4_9, outputs_20_8=>
      outMuls_4_8, outputs_20_7=>outMuls_4_7, outputs_20_6=>outMuls_4_6, 
      outputs_20_5=>outMuls_4_5, outputs_20_4=>outMuls_4_4, outputs_20_3=>
      outMuls_4_3, outputs_20_2=>outMuls_4_2, outputs_20_1=>outMuls_4_1, 
      outputs_20_0=>outMuls_4_0, outputs_19_15=>outMuls_5_15, outputs_19_14
      =>outMuls_5_14, outputs_19_13=>outMuls_5_13, outputs_19_12=>
      outMuls_5_12, outputs_19_11=>outMuls_5_11, outputs_19_10=>outMuls_5_10, 
      outputs_19_9=>outMuls_5_9, outputs_19_8=>outMuls_5_8, outputs_19_7=>
      outMuls_5_7, outputs_19_6=>outMuls_5_6, outputs_19_5=>outMuls_5_5, 
      outputs_19_4=>outMuls_5_4, outputs_19_3=>outMuls_5_3, outputs_19_2=>
      outMuls_5_2, outputs_19_1=>outMuls_5_1, outputs_19_0=>outMuls_5_0, 
      outputs_18_15=>outMuls_6_15, outputs_18_14=>outMuls_6_14, 
      outputs_18_13=>outMuls_6_13, outputs_18_12=>outMuls_6_12, 
      outputs_18_11=>outMuls_6_11, outputs_18_10=>outMuls_6_10, outputs_18_9
      =>outMuls_6_9, outputs_18_8=>outMuls_6_8, outputs_18_7=>outMuls_6_7, 
      outputs_18_6=>outMuls_6_6, outputs_18_5=>outMuls_6_5, outputs_18_4=>
      outMuls_6_4, outputs_18_3=>outMuls_6_3, outputs_18_2=>outMuls_6_2, 
      outputs_18_1=>outMuls_6_1, outputs_18_0=>outMuls_6_0, outputs_17_15=>
      outMuls_7_15, outputs_17_14=>outMuls_7_14, outputs_17_13=>outMuls_7_13, 
      outputs_17_12=>outMuls_7_12, outputs_17_11=>outMuls_7_11, 
      outputs_17_10=>outMuls_7_10, outputs_17_9=>outMuls_7_9, outputs_17_8=>
      outMuls_7_8, outputs_17_7=>outMuls_7_7, outputs_17_6=>outMuls_7_6, 
      outputs_17_5=>outMuls_7_5, outputs_17_4=>outMuls_7_4, outputs_17_3=>
      outMuls_7_3, outputs_17_2=>outMuls_7_2, outputs_17_1=>outMuls_7_1, 
      outputs_17_0=>outMuls_7_0, outputs_16_15=>outMuls_8_15, outputs_16_14
      =>outMuls_8_14, outputs_16_13=>outMuls_8_13, outputs_16_12=>
      outMuls_8_12, outputs_16_11=>outMuls_8_11, outputs_16_10=>outMuls_8_10, 
      outputs_16_9=>outMuls_8_9, outputs_16_8=>outMuls_8_8, outputs_16_7=>
      outMuls_8_7, outputs_16_6=>outMuls_8_6, outputs_16_5=>outMuls_8_5, 
      outputs_16_4=>outMuls_8_4, outputs_16_3=>outMuls_8_3, outputs_16_2=>
      outMuls_8_2, outputs_16_1=>outMuls_8_1, outputs_16_0=>outMuls_8_0, 
      outputs_15_15=>outMuls_9_15, outputs_15_14=>outMuls_9_14, 
      outputs_15_13=>outMuls_9_13, outputs_15_12=>outMuls_9_12, 
      outputs_15_11=>outMuls_9_11, outputs_15_10=>outMuls_9_10, outputs_15_9
      =>outMuls_9_9, outputs_15_8=>outMuls_9_8, outputs_15_7=>outMuls_9_7, 
      outputs_15_6=>outMuls_9_6, outputs_15_5=>outMuls_9_5, outputs_15_4=>
      outMuls_9_4, outputs_15_3=>outMuls_9_3, outputs_15_2=>outMuls_9_2, 
      outputs_15_1=>outMuls_9_1, outputs_15_0=>outMuls_9_0, outputs_14_15=>
      outMuls_10_15, outputs_14_14=>outMuls_10_14, outputs_14_13=>
      outMuls_10_13, outputs_14_12=>outMuls_10_12, outputs_14_11=>
      outMuls_10_11, outputs_14_10=>outMuls_10_10, outputs_14_9=>
      outMuls_10_9, outputs_14_8=>outMuls_10_8, outputs_14_7=>outMuls_10_7, 
      outputs_14_6=>outMuls_10_6, outputs_14_5=>outMuls_10_5, outputs_14_4=>
      outMuls_10_4, outputs_14_3=>outMuls_10_3, outputs_14_2=>outMuls_10_2, 
      outputs_14_1=>outMuls_10_1, outputs_14_0=>outMuls_10_0, outputs_13_15
      =>outMuls_11_15, outputs_13_14=>outMuls_11_14, outputs_13_13=>
      outMuls_11_13, outputs_13_12=>outMuls_11_12, outputs_13_11=>
      outMuls_11_11, outputs_13_10=>outMuls_11_10, outputs_13_9=>
      outMuls_11_9, outputs_13_8=>outMuls_11_8, outputs_13_7=>outMuls_11_7, 
      outputs_13_6=>outMuls_11_6, outputs_13_5=>outMuls_11_5, outputs_13_4=>
      outMuls_11_4, outputs_13_3=>outMuls_11_3, outputs_13_2=>outMuls_11_2, 
      outputs_13_1=>outMuls_11_1, outputs_13_0=>outMuls_11_0, outputs_12_15
      =>outMuls_12_15, outputs_12_14=>outMuls_12_14, outputs_12_13=>
      outMuls_12_13, outputs_12_12=>outMuls_12_12, outputs_12_11=>
      outMuls_12_11, outputs_12_10=>outMuls_12_10, outputs_12_9=>
      outMuls_12_9, outputs_12_8=>outMuls_12_8, outputs_12_7=>outMuls_12_7, 
      outputs_12_6=>outMuls_12_6, outputs_12_5=>outMuls_12_5, outputs_12_4=>
      outMuls_12_4, outputs_12_3=>outMuls_12_3, outputs_12_2=>outMuls_12_2, 
      outputs_12_1=>outMuls_12_1, outputs_12_0=>outMuls_12_0, outputs_11_15
      =>outMuls_13_15, outputs_11_14=>outMuls_13_14, outputs_11_13=>
      outMuls_13_13, outputs_11_12=>outMuls_13_12, outputs_11_11=>
      outMuls_13_11, outputs_11_10=>outMuls_13_10, outputs_11_9=>
      outMuls_13_9, outputs_11_8=>outMuls_13_8, outputs_11_7=>outMuls_13_7, 
      outputs_11_6=>outMuls_13_6, outputs_11_5=>outMuls_13_5, outputs_11_4=>
      outMuls_13_4, outputs_11_3=>outMuls_13_3, outputs_11_2=>outMuls_13_2, 
      outputs_11_1=>outMuls_13_1, outputs_11_0=>outMuls_13_0, outputs_10_15
      =>outMuls_14_15, outputs_10_14=>outMuls_14_14, outputs_10_13=>
      outMuls_14_13, outputs_10_12=>outMuls_14_12, outputs_10_11=>
      outMuls_14_11, outputs_10_10=>outMuls_14_10, outputs_10_9=>
      outMuls_14_9, outputs_10_8=>outMuls_14_8, outputs_10_7=>outMuls_14_7, 
      outputs_10_6=>outMuls_14_6, outputs_10_5=>outMuls_14_5, outputs_10_4=>
      outMuls_14_4, outputs_10_3=>outMuls_14_3, outputs_10_2=>outMuls_14_2, 
      outputs_10_1=>outMuls_14_1, outputs_10_0=>outMuls_14_0, outputs_9_15=>
      outMuls_15_15, outputs_9_14=>outMuls_15_14, outputs_9_13=>
      outMuls_15_13, outputs_9_12=>outMuls_15_12, outputs_9_11=>
      outMuls_15_11, outputs_9_10=>outMuls_15_10, outputs_9_9=>outMuls_15_9, 
      outputs_9_8=>outMuls_15_8, outputs_9_7=>outMuls_15_7, outputs_9_6=>
      outMuls_15_6, outputs_9_5=>outMuls_15_5, outputs_9_4=>outMuls_15_4, 
      outputs_9_3=>outMuls_15_3, outputs_9_2=>outMuls_15_2, outputs_9_1=>
      outMuls_15_1, outputs_9_0=>outMuls_15_0, outputs_8_15=>outMuls_16_15, 
      outputs_8_14=>outMuls_16_14, outputs_8_13=>outMuls_16_13, outputs_8_12
      =>outMuls_16_12, outputs_8_11=>outMuls_16_11, outputs_8_10=>
      outMuls_16_10, outputs_8_9=>outMuls_16_9, outputs_8_8=>outMuls_16_8, 
      outputs_8_7=>outMuls_16_7, outputs_8_6=>outMuls_16_6, outputs_8_5=>
      outMuls_16_5, outputs_8_4=>outMuls_16_4, outputs_8_3=>outMuls_16_3, 
      outputs_8_2=>outMuls_16_2, outputs_8_1=>outMuls_16_1, outputs_8_0=>
      outMuls_16_0, outputs_7_15=>outMuls_17_15, outputs_7_14=>outMuls_17_14, 
      outputs_7_13=>outMuls_17_13, outputs_7_12=>outMuls_17_12, outputs_7_11
      =>outMuls_17_11, outputs_7_10=>outMuls_17_10, outputs_7_9=>
      outMuls_17_9, outputs_7_8=>outMuls_17_8, outputs_7_7=>outMuls_17_7, 
      outputs_7_6=>outMuls_17_6, outputs_7_5=>outMuls_17_5, outputs_7_4=>
      outMuls_17_4, outputs_7_3=>outMuls_17_3, outputs_7_2=>outMuls_17_2, 
      outputs_7_1=>outMuls_17_1, outputs_7_0=>outMuls_17_0, outputs_6_15=>
      outMuls_18_15, outputs_6_14=>outMuls_18_14, outputs_6_13=>
      outMuls_18_13, outputs_6_12=>outMuls_18_12, outputs_6_11=>
      outMuls_18_11, outputs_6_10=>outMuls_18_10, outputs_6_9=>outMuls_18_9, 
      outputs_6_8=>outMuls_18_8, outputs_6_7=>outMuls_18_7, outputs_6_6=>
      outMuls_18_6, outputs_6_5=>outMuls_18_5, outputs_6_4=>outMuls_18_4, 
      outputs_6_3=>outMuls_18_3, outputs_6_2=>outMuls_18_2, outputs_6_1=>
      outMuls_18_1, outputs_6_0=>outMuls_18_0, outputs_5_15=>outMuls_19_15, 
      outputs_5_14=>outMuls_19_14, outputs_5_13=>outMuls_19_13, outputs_5_12
      =>outMuls_19_12, outputs_5_11=>outMuls_19_11, outputs_5_10=>
      outMuls_19_10, outputs_5_9=>outMuls_19_9, outputs_5_8=>outMuls_19_8, 
      outputs_5_7=>outMuls_19_7, outputs_5_6=>outMuls_19_6, outputs_5_5=>
      outMuls_19_5, outputs_5_4=>outMuls_19_4, outputs_5_3=>outMuls_19_3, 
      outputs_5_2=>outMuls_19_2, outputs_5_1=>outMuls_19_1, outputs_5_0=>
      outMuls_19_0, outputs_4_15=>outMuls_20_15, outputs_4_14=>outMuls_20_14, 
      outputs_4_13=>outMuls_20_13, outputs_4_12=>outMuls_20_12, outputs_4_11
      =>outMuls_20_11, outputs_4_10=>outMuls_20_10, outputs_4_9=>
      outMuls_20_9, outputs_4_8=>outMuls_20_8, outputs_4_7=>outMuls_20_7, 
      outputs_4_6=>outMuls_20_6, outputs_4_5=>outMuls_20_5, outputs_4_4=>
      outMuls_20_4, outputs_4_3=>outMuls_20_3, outputs_4_2=>outMuls_20_2, 
      outputs_4_1=>outMuls_20_1, outputs_4_0=>outMuls_20_0, outputs_3_15=>
      outMuls_21_15, outputs_3_14=>outMuls_21_14, outputs_3_13=>
      outMuls_21_13, outputs_3_12=>outMuls_21_12, outputs_3_11=>
      outMuls_21_11, outputs_3_10=>outMuls_21_10, outputs_3_9=>outMuls_21_9, 
      outputs_3_8=>outMuls_21_8, outputs_3_7=>outMuls_21_7, outputs_3_6=>
      outMuls_21_6, outputs_3_5=>outMuls_21_5, outputs_3_4=>outMuls_21_4, 
      outputs_3_3=>outMuls_21_3, outputs_3_2=>outMuls_21_2, outputs_3_1=>
      outMuls_21_1, outputs_3_0=>outMuls_21_0, outputs_2_15=>outMuls_22_15, 
      outputs_2_14=>outMuls_22_14, outputs_2_13=>outMuls_22_13, outputs_2_12
      =>outMuls_22_12, outputs_2_11=>outMuls_22_11, outputs_2_10=>
      outMuls_22_10, outputs_2_9=>outMuls_22_9, outputs_2_8=>outMuls_22_8, 
      outputs_2_7=>outMuls_22_7, outputs_2_6=>outMuls_22_6, outputs_2_5=>
      outMuls_22_5, outputs_2_4=>outMuls_22_4, outputs_2_3=>outMuls_22_3, 
      outputs_2_2=>outMuls_22_2, outputs_2_1=>outMuls_22_1, outputs_2_0=>
      outMuls_22_0, outputs_1_15=>outMuls_23_15, outputs_1_14=>outMuls_23_14, 
      outputs_1_13=>outMuls_23_13, outputs_1_12=>outMuls_23_12, outputs_1_11
      =>outMuls_23_11, outputs_1_10=>outMuls_23_10, outputs_1_9=>
      outMuls_23_9, outputs_1_8=>outMuls_23_8, outputs_1_7=>outMuls_23_7, 
      outputs_1_6=>outMuls_23_6, outputs_1_5=>outMuls_23_5, outputs_1_4=>
      outMuls_23_4, outputs_1_3=>outMuls_23_3, outputs_1_2=>outMuls_23_2, 
      outputs_1_1=>outMuls_23_1, outputs_1_0=>outMuls_23_0, outputs_0_15=>
      outMuls_24_15, outputs_0_14=>outMuls_24_14, outputs_0_13=>
      outMuls_24_13, outputs_0_12=>outMuls_24_12, outputs_0_11=>
      outMuls_24_11, outputs_0_10=>outMuls_24_10, outputs_0_9=>outMuls_24_9, 
      outputs_0_8=>outMuls_24_8, outputs_0_7=>outMuls_24_7, outputs_0_6=>
      outMuls_24_6, outputs_0_5=>outMuls_24_5, outputs_0_4=>outMuls_24_4, 
      outputs_0_3=>outMuls_24_3, outputs_0_2=>outMuls_24_2, outputs_0_1=>
      outMuls_24_1, outputs_0_0=>outMuls_24_0, clk=>clk, start=>start, rst=>
      rst, done=>doneMul, working=>DANGLING(0));
   regFileMap_loop1_0_regRowMap_loop1_0_regUnitMap : RegUnit_8_16
       port map ( filterBus(7)=>filterBus(7), filterBus(6)=>filterBus(6), 
      filterBus(5)=>filterBus(5), filterBus(4)=>filterBus(4), filterBus(3)=>
      filterBus(3), filterBus(2)=>filterBus(2), filterBus(1)=>filterBus(1), 
      filterBus(0)=>filterBus(0), windowBus(15)=>windowBus(15), 
      windowBus(14)=>windowBus(14), windowBus(13)=>windowBus(13), 
      windowBus(12)=>windowBus(12), windowBus(11)=>windowBus(11), 
      windowBus(10)=>windowBus(10), windowBus(9)=>windowBus(9), windowBus(8)
      =>windowBus(8), windowBus(7)=>windowBus(7), windowBus(6)=>windowBus(6), 
      windowBus(5)=>windowBus(5), windowBus(4)=>windowBus(4), windowBus(3)=>
      windowBus(3), windowBus(2)=>windowBus(2), windowBus(1)=>windowBus(1), 
      windowBus(0)=>windowBus(0), regPage1NextUnit(15)=>
      regFileMap_page1Out_5_15, regPage1NextUnit(14)=>
      regFileMap_page1Out_5_14, regPage1NextUnit(13)=>
      regFileMap_page1Out_5_13, regPage1NextUnit(12)=>
      regFileMap_page1Out_5_12, regPage1NextUnit(11)=>
      regFileMap_page1Out_5_11, regPage1NextUnit(10)=>
      regFileMap_page1Out_5_10, regPage1NextUnit(9)=>regFileMap_page1Out_5_9, 
      regPage1NextUnit(8)=>regFileMap_page1Out_5_8, regPage1NextUnit(7)=>
      regFileMap_page1Out_5_7, regPage1NextUnit(6)=>regFileMap_page1Out_5_6, 
      regPage1NextUnit(5)=>regFileMap_page1Out_5_5, regPage1NextUnit(4)=>
      regFileMap_page1Out_5_4, regPage1NextUnit(3)=>regFileMap_page1Out_5_3, 
      regPage1NextUnit(2)=>regFileMap_page1Out_5_2, regPage1NextUnit(1)=>
      regFileMap_page1Out_5_1, regPage1NextUnit(0)=>regFileMap_page1Out_5_0, 
      regPage2NextUnit(15)=>regFileMap_page2Out_5_15, regPage2NextUnit(14)=>
      regFileMap_page2Out_5_14, regPage2NextUnit(13)=>
      regFileMap_page2Out_5_13, regPage2NextUnit(12)=>
      regFileMap_page2Out_5_12, regPage2NextUnit(11)=>
      regFileMap_page2Out_5_11, regPage2NextUnit(10)=>
      regFileMap_page2Out_5_10, regPage2NextUnit(9)=>regFileMap_page2Out_5_9, 
      regPage2NextUnit(8)=>regFileMap_page2Out_5_8, regPage2NextUnit(7)=>
      regFileMap_page2Out_5_7, regPage2NextUnit(6)=>regFileMap_page2Out_5_6, 
      regPage2NextUnit(5)=>regFileMap_page2Out_5_5, regPage2NextUnit(4)=>
      regFileMap_page2Out_5_4, regPage2NextUnit(3)=>regFileMap_page2Out_5_3, 
      regPage2NextUnit(2)=>regFileMap_page2Out_5_2, regPage2NextUnit(1)=>
      regFileMap_page2Out_5_1, regPage2NextUnit(0)=>regFileMap_page2Out_5_0, 
      clk=>clk, rst=>rst, enableRegPage1=>regFileMap_page1Enables_0, 
      enableRegPage2=>regFileMap_page2Enables_0, enableRegFilter=>nx5328, 
      page1ReadBusOrPage2=>shift2To1, page2ReadBusOrPage1=>shift1To2, 
      pageTurn=>pageTurn, outRegPage(15)=>currentPage_0_15, outRegPage(14)=>
      currentPage_0_14, outRegPage(13)=>currentPage_0_13, outRegPage(12)=>
      currentPage_0_12, outRegPage(11)=>currentPage_0_11, outRegPage(10)=>
      currentPage_0_10, outRegPage(9)=>currentPage_0_9, outRegPage(8)=>
      currentPage_0_8, outRegPage(7)=>currentPage_0_7, outRegPage(6)=>
      currentPage_0_6, outRegPage(5)=>currentPage_0_5, outRegPage(4)=>
      currentPage_0_4, outRegPage(3)=>currentPage_0_3, outRegPage(2)=>
      currentPage_0_2, outRegPage(1)=>currentPage_0_1, outRegPage(0)=>
      currentPage_0_0, outputRegPage1(15)=>DANGLING(1), outputRegPage1(14)=>
      DANGLING(2), outputRegPage1(13)=>DANGLING(3), outputRegPage1(12)=>
      DANGLING(4), outputRegPage1(11)=>DANGLING(5), outputRegPage1(10)=>
      DANGLING(6), outputRegPage1(9)=>DANGLING(7), outputRegPage1(8)=>
      DANGLING(8), outputRegPage1(7)=>DANGLING(9), outputRegPage1(6)=>
      DANGLING(10), outputRegPage1(5)=>DANGLING(11), outputRegPage1(4)=>
      DANGLING(12), outputRegPage1(3)=>DANGLING(13), outputRegPage1(2)=>
      DANGLING(14), outputRegPage1(1)=>DANGLING(15), outputRegPage1(0)=>
      DANGLING(16), outputRegPage2(15)=>DANGLING(17), outputRegPage2(14)=>
      DANGLING(18), outputRegPage2(13)=>DANGLING(19), outputRegPage2(12)=>
      DANGLING(20), outputRegPage2(11)=>DANGLING(21), outputRegPage2(10)=>
      DANGLING(22), outputRegPage2(9)=>DANGLING(23), outputRegPage2(8)=>
      DANGLING(24), outputRegPage2(7)=>DANGLING(25), outputRegPage2(6)=>
      DANGLING(26), outputRegPage2(5)=>DANGLING(27), outputRegPage2(4)=>
      DANGLING(28), outputRegPage2(3)=>DANGLING(29), outputRegPage2(2)=>
      DANGLING(30), outputRegPage2(1)=>DANGLING(31), outputRegPage2(0)=>
      DANGLING(32), outFilter(7)=>filter_0_7, outFilter(6)=>filter_0_6, 
      outFilter(5)=>filter_0_5, outFilter(4)=>filter_0_4, outFilter(3)=>
      filter_0_3, outFilter(2)=>filter_0_2, outFilter(1)=>filter_0_1, 
      outFilter(0)=>filter_0_0);
   regFileMap_loop1_0_regRowMap_loop1_1_regUnitMap : RegUnit_8_16
       port map ( filterBus(7)=>filterBus(15), filterBus(6)=>filterBus(14), 
      filterBus(5)=>filterBus(13), filterBus(4)=>filterBus(12), filterBus(3)
      =>filterBus(11), filterBus(2)=>filterBus(10), filterBus(1)=>
      filterBus(9), filterBus(0)=>filterBus(8), windowBus(15)=>windowBus(31), 
      windowBus(14)=>windowBus(30), windowBus(13)=>windowBus(29), 
      windowBus(12)=>windowBus(28), windowBus(11)=>windowBus(27), 
      windowBus(10)=>windowBus(26), windowBus(9)=>windowBus(25), 
      windowBus(8)=>windowBus(24), windowBus(7)=>windowBus(23), windowBus(6)
      =>windowBus(22), windowBus(5)=>windowBus(21), windowBus(4)=>
      windowBus(20), windowBus(3)=>windowBus(19), windowBus(2)=>
      windowBus(18), windowBus(1)=>windowBus(17), windowBus(0)=>
      windowBus(16), regPage1NextUnit(15)=>regFileMap_page1Out_6_15, 
      regPage1NextUnit(14)=>regFileMap_page1Out_6_14, regPage1NextUnit(13)=>
      regFileMap_page1Out_6_13, regPage1NextUnit(12)=>
      regFileMap_page1Out_6_12, regPage1NextUnit(11)=>
      regFileMap_page1Out_6_11, regPage1NextUnit(10)=>
      regFileMap_page1Out_6_10, regPage1NextUnit(9)=>regFileMap_page1Out_6_9, 
      regPage1NextUnit(8)=>regFileMap_page1Out_6_8, regPage1NextUnit(7)=>
      regFileMap_page1Out_6_7, regPage1NextUnit(6)=>regFileMap_page1Out_6_6, 
      regPage1NextUnit(5)=>regFileMap_page1Out_6_5, regPage1NextUnit(4)=>
      regFileMap_page1Out_6_4, regPage1NextUnit(3)=>regFileMap_page1Out_6_3, 
      regPage1NextUnit(2)=>regFileMap_page1Out_6_2, regPage1NextUnit(1)=>
      regFileMap_page1Out_6_1, regPage1NextUnit(0)=>regFileMap_page1Out_6_0, 
      regPage2NextUnit(15)=>regFileMap_page2Out_6_15, regPage2NextUnit(14)=>
      regFileMap_page2Out_6_14, regPage2NextUnit(13)=>
      regFileMap_page2Out_6_13, regPage2NextUnit(12)=>
      regFileMap_page2Out_6_12, regPage2NextUnit(11)=>
      regFileMap_page2Out_6_11, regPage2NextUnit(10)=>
      regFileMap_page2Out_6_10, regPage2NextUnit(9)=>regFileMap_page2Out_6_9, 
      regPage2NextUnit(8)=>regFileMap_page2Out_6_8, regPage2NextUnit(7)=>
      regFileMap_page2Out_6_7, regPage2NextUnit(6)=>regFileMap_page2Out_6_6, 
      regPage2NextUnit(5)=>regFileMap_page2Out_6_5, regPage2NextUnit(4)=>
      regFileMap_page2Out_6_4, regPage2NextUnit(3)=>regFileMap_page2Out_6_3, 
      regPage2NextUnit(2)=>regFileMap_page2Out_6_2, regPage2NextUnit(1)=>
      regFileMap_page2Out_6_1, regPage2NextUnit(0)=>regFileMap_page2Out_6_0, 
      clk=>clk, rst=>rst, enableRegPage1=>regFileMap_page1Enables_0, 
      enableRegPage2=>regFileMap_page2Enables_0, enableRegFilter=>nx5328, 
      page1ReadBusOrPage2=>shift2To1, page2ReadBusOrPage1=>shift1To2, 
      pageTurn=>pageTurn, outRegPage(15)=>currentPage_1_15, outRegPage(14)=>
      currentPage_1_14, outRegPage(13)=>currentPage_1_13, outRegPage(12)=>
      currentPage_1_12, outRegPage(11)=>currentPage_1_11, outRegPage(10)=>
      currentPage_1_10, outRegPage(9)=>currentPage_1_9, outRegPage(8)=>
      currentPage_1_8, outRegPage(7)=>currentPage_1_7, outRegPage(6)=>
      currentPage_1_6, outRegPage(5)=>currentPage_1_5, outRegPage(4)=>
      currentPage_1_4, outRegPage(3)=>currentPage_1_3, outRegPage(2)=>
      currentPage_1_2, outRegPage(1)=>currentPage_1_1, outRegPage(0)=>
      currentPage_1_0, outputRegPage1(15)=>DANGLING(33), outputRegPage1(14)
      =>DANGLING(34), outputRegPage1(13)=>DANGLING(35), outputRegPage1(12)=>
      DANGLING(36), outputRegPage1(11)=>DANGLING(37), outputRegPage1(10)=>
      DANGLING(38), outputRegPage1(9)=>DANGLING(39), outputRegPage1(8)=>
      DANGLING(40), outputRegPage1(7)=>DANGLING(41), outputRegPage1(6)=>
      DANGLING(42), outputRegPage1(5)=>DANGLING(43), outputRegPage1(4)=>
      DANGLING(44), outputRegPage1(3)=>DANGLING(45), outputRegPage1(2)=>
      DANGLING(46), outputRegPage1(1)=>DANGLING(47), outputRegPage1(0)=>
      DANGLING(48), outputRegPage2(15)=>DANGLING(49), outputRegPage2(14)=>
      DANGLING(50), outputRegPage2(13)=>DANGLING(51), outputRegPage2(12)=>
      DANGLING(52), outputRegPage2(11)=>DANGLING(53), outputRegPage2(10)=>
      DANGLING(54), outputRegPage2(9)=>DANGLING(55), outputRegPage2(8)=>
      DANGLING(56), outputRegPage2(7)=>DANGLING(57), outputRegPage2(6)=>
      DANGLING(58), outputRegPage2(5)=>DANGLING(59), outputRegPage2(4)=>
      DANGLING(60), outputRegPage2(3)=>DANGLING(61), outputRegPage2(2)=>
      DANGLING(62), outputRegPage2(1)=>DANGLING(63), outputRegPage2(0)=>
      DANGLING(64), outFilter(7)=>filter_1_7, outFilter(6)=>filter_1_6, 
      outFilter(5)=>filter_1_5, outFilter(4)=>filter_1_4, outFilter(3)=>
      filter_1_3, outFilter(2)=>filter_1_2, outFilter(1)=>filter_1_1, 
      outFilter(0)=>filter_1_0);
   regFileMap_loop1_0_regRowMap_loop1_2_regUnitMap : RegUnit_8_16
       port map ( filterBus(7)=>filterBus(23), filterBus(6)=>filterBus(22), 
      filterBus(5)=>filterBus(21), filterBus(4)=>filterBus(20), filterBus(3)
      =>filterBus(19), filterBus(2)=>filterBus(18), filterBus(1)=>
      filterBus(17), filterBus(0)=>filterBus(16), windowBus(15)=>
      windowBus(47), windowBus(14)=>windowBus(46), windowBus(13)=>
      windowBus(45), windowBus(12)=>windowBus(44), windowBus(11)=>
      windowBus(43), windowBus(10)=>windowBus(42), windowBus(9)=>
      windowBus(41), windowBus(8)=>windowBus(40), windowBus(7)=>
      windowBus(39), windowBus(6)=>windowBus(38), windowBus(5)=>
      windowBus(37), windowBus(4)=>windowBus(36), windowBus(3)=>
      windowBus(35), windowBus(2)=>windowBus(34), windowBus(1)=>
      windowBus(33), windowBus(0)=>windowBus(32), regPage1NextUnit(15)=>
      regFileMap_page1Out_7_15, regPage1NextUnit(14)=>
      regFileMap_page1Out_7_14, regPage1NextUnit(13)=>
      regFileMap_page1Out_7_13, regPage1NextUnit(12)=>
      regFileMap_page1Out_7_12, regPage1NextUnit(11)=>
      regFileMap_page1Out_7_11, regPage1NextUnit(10)=>
      regFileMap_page1Out_7_10, regPage1NextUnit(9)=>regFileMap_page1Out_7_9, 
      regPage1NextUnit(8)=>regFileMap_page1Out_7_8, regPage1NextUnit(7)=>
      regFileMap_page1Out_7_7, regPage1NextUnit(6)=>regFileMap_page1Out_7_6, 
      regPage1NextUnit(5)=>regFileMap_page1Out_7_5, regPage1NextUnit(4)=>
      regFileMap_page1Out_7_4, regPage1NextUnit(3)=>regFileMap_page1Out_7_3, 
      regPage1NextUnit(2)=>regFileMap_page1Out_7_2, regPage1NextUnit(1)=>
      regFileMap_page1Out_7_1, regPage1NextUnit(0)=>regFileMap_page1Out_7_0, 
      regPage2NextUnit(15)=>regFileMap_page2Out_7_15, regPage2NextUnit(14)=>
      regFileMap_page2Out_7_14, regPage2NextUnit(13)=>
      regFileMap_page2Out_7_13, regPage2NextUnit(12)=>
      regFileMap_page2Out_7_12, regPage2NextUnit(11)=>
      regFileMap_page2Out_7_11, regPage2NextUnit(10)=>
      regFileMap_page2Out_7_10, regPage2NextUnit(9)=>regFileMap_page2Out_7_9, 
      regPage2NextUnit(8)=>regFileMap_page2Out_7_8, regPage2NextUnit(7)=>
      regFileMap_page2Out_7_7, regPage2NextUnit(6)=>regFileMap_page2Out_7_6, 
      regPage2NextUnit(5)=>regFileMap_page2Out_7_5, regPage2NextUnit(4)=>
      regFileMap_page2Out_7_4, regPage2NextUnit(3)=>regFileMap_page2Out_7_3, 
      regPage2NextUnit(2)=>regFileMap_page2Out_7_2, regPage2NextUnit(1)=>
      regFileMap_page2Out_7_1, regPage2NextUnit(0)=>regFileMap_page2Out_7_0, 
      clk=>clk, rst=>rst, enableRegPage1=>regFileMap_page1Enables_0, 
      enableRegPage2=>regFileMap_page2Enables_0, enableRegFilter=>nx5328, 
      page1ReadBusOrPage2=>shift2To1, page2ReadBusOrPage1=>shift1To2, 
      pageTurn=>pageTurn, outRegPage(15)=>currentPage_2_15, outRegPage(14)=>
      currentPage_2_14, outRegPage(13)=>currentPage_2_13, outRegPage(12)=>
      currentPage_2_12, outRegPage(11)=>currentPage_2_11, outRegPage(10)=>
      currentPage_2_10, outRegPage(9)=>currentPage_2_9, outRegPage(8)=>
      currentPage_2_8, outRegPage(7)=>currentPage_2_7, outRegPage(6)=>
      currentPage_2_6, outRegPage(5)=>currentPage_2_5, outRegPage(4)=>
      currentPage_2_4, outRegPage(3)=>currentPage_2_3, outRegPage(2)=>
      currentPage_2_2, outRegPage(1)=>currentPage_2_1, outRegPage(0)=>
      currentPage_2_0, outputRegPage1(15)=>DANGLING(65), outputRegPage1(14)
      =>DANGLING(66), outputRegPage1(13)=>DANGLING(67), outputRegPage1(12)=>
      DANGLING(68), outputRegPage1(11)=>DANGLING(69), outputRegPage1(10)=>
      DANGLING(70), outputRegPage1(9)=>DANGLING(71), outputRegPage1(8)=>
      DANGLING(72), outputRegPage1(7)=>DANGLING(73), outputRegPage1(6)=>
      DANGLING(74), outputRegPage1(5)=>DANGLING(75), outputRegPage1(4)=>
      DANGLING(76), outputRegPage1(3)=>DANGLING(77), outputRegPage1(2)=>
      DANGLING(78), outputRegPage1(1)=>DANGLING(79), outputRegPage1(0)=>
      DANGLING(80), outputRegPage2(15)=>DANGLING(81), outputRegPage2(14)=>
      DANGLING(82), outputRegPage2(13)=>DANGLING(83), outputRegPage2(12)=>
      DANGLING(84), outputRegPage2(11)=>DANGLING(85), outputRegPage2(10)=>
      DANGLING(86), outputRegPage2(9)=>DANGLING(87), outputRegPage2(8)=>
      DANGLING(88), outputRegPage2(7)=>DANGLING(89), outputRegPage2(6)=>
      DANGLING(90), outputRegPage2(5)=>DANGLING(91), outputRegPage2(4)=>
      DANGLING(92), outputRegPage2(3)=>DANGLING(93), outputRegPage2(2)=>
      DANGLING(94), outputRegPage2(1)=>DANGLING(95), outputRegPage2(0)=>
      DANGLING(96), outFilter(7)=>filter_2_7, outFilter(6)=>filter_2_6, 
      outFilter(5)=>filter_2_5, outFilter(4)=>filter_2_4, outFilter(3)=>
      filter_2_3, outFilter(2)=>filter_2_2, outFilter(1)=>filter_2_1, 
      outFilter(0)=>filter_2_0);
   regFileMap_loop1_0_regRowMap_loop1_3_regUnitMap : RegUnit_8_16
       port map ( filterBus(7)=>filterBus(31), filterBus(6)=>filterBus(30), 
      filterBus(5)=>filterBus(29), filterBus(4)=>filterBus(28), filterBus(3)
      =>filterBus(27), filterBus(2)=>filterBus(26), filterBus(1)=>
      filterBus(25), filterBus(0)=>filterBus(24), windowBus(15)=>
      windowBus(63), windowBus(14)=>windowBus(62), windowBus(13)=>
      windowBus(61), windowBus(12)=>windowBus(60), windowBus(11)=>
      windowBus(59), windowBus(10)=>windowBus(58), windowBus(9)=>
      windowBus(57), windowBus(8)=>windowBus(56), windowBus(7)=>
      windowBus(55), windowBus(6)=>windowBus(54), windowBus(5)=>
      windowBus(53), windowBus(4)=>windowBus(52), windowBus(3)=>
      windowBus(51), windowBus(2)=>windowBus(50), windowBus(1)=>
      windowBus(49), windowBus(0)=>windowBus(48), regPage1NextUnit(15)=>
      regFileMap_page1Out_8_15, regPage1NextUnit(14)=>
      regFileMap_page1Out_8_14, regPage1NextUnit(13)=>
      regFileMap_page1Out_8_13, regPage1NextUnit(12)=>
      regFileMap_page1Out_8_12, regPage1NextUnit(11)=>
      regFileMap_page1Out_8_11, regPage1NextUnit(10)=>
      regFileMap_page1Out_8_10, regPage1NextUnit(9)=>regFileMap_page1Out_8_9, 
      regPage1NextUnit(8)=>regFileMap_page1Out_8_8, regPage1NextUnit(7)=>
      regFileMap_page1Out_8_7, regPage1NextUnit(6)=>regFileMap_page1Out_8_6, 
      regPage1NextUnit(5)=>regFileMap_page1Out_8_5, regPage1NextUnit(4)=>
      regFileMap_page1Out_8_4, regPage1NextUnit(3)=>regFileMap_page1Out_8_3, 
      regPage1NextUnit(2)=>regFileMap_page1Out_8_2, regPage1NextUnit(1)=>
      regFileMap_page1Out_8_1, regPage1NextUnit(0)=>regFileMap_page1Out_8_0, 
      regPage2NextUnit(15)=>regFileMap_page2Out_8_15, regPage2NextUnit(14)=>
      regFileMap_page2Out_8_14, regPage2NextUnit(13)=>
      regFileMap_page2Out_8_13, regPage2NextUnit(12)=>
      regFileMap_page2Out_8_12, regPage2NextUnit(11)=>
      regFileMap_page2Out_8_11, regPage2NextUnit(10)=>
      regFileMap_page2Out_8_10, regPage2NextUnit(9)=>regFileMap_page2Out_8_9, 
      regPage2NextUnit(8)=>regFileMap_page2Out_8_8, regPage2NextUnit(7)=>
      regFileMap_page2Out_8_7, regPage2NextUnit(6)=>regFileMap_page2Out_8_6, 
      regPage2NextUnit(5)=>regFileMap_page2Out_8_5, regPage2NextUnit(4)=>
      regFileMap_page2Out_8_4, regPage2NextUnit(3)=>regFileMap_page2Out_8_3, 
      regPage2NextUnit(2)=>regFileMap_page2Out_8_2, regPage2NextUnit(1)=>
      regFileMap_page2Out_8_1, regPage2NextUnit(0)=>regFileMap_page2Out_8_0, 
      clk=>clk, rst=>rst, enableRegPage1=>regFileMap_page1Enables_0, 
      enableRegPage2=>regFileMap_page2Enables_0, enableRegFilter=>nx5330, 
      page1ReadBusOrPage2=>shift2To1, page2ReadBusOrPage1=>shift1To2, 
      pageTurn=>pageTurn, outRegPage(15)=>currentPage_15_15, outRegPage(14)
      =>currentPage_15_14, outRegPage(13)=>currentPage_15_13, outRegPage(12)
      =>currentPage_15_12, outRegPage(11)=>currentPage_15_11, outRegPage(10)
      =>currentPage_15_10, outRegPage(9)=>currentPage_15_9, outRegPage(8)=>
      currentPage_15_8, outRegPage(7)=>currentPage_15_7, outRegPage(6)=>
      currentPage_15_6, outRegPage(5)=>currentPage_15_5, outRegPage(4)=>
      currentPage_15_4, outRegPage(3)=>currentPage_15_3, outRegPage(2)=>
      currentPage_15_2, outRegPage(1)=>currentPage_15_1, outRegPage(0)=>
      currentPage_15_0, outputRegPage1(15)=>DANGLING(97), outputRegPage1(14)
      =>DANGLING(98), outputRegPage1(13)=>DANGLING(99), outputRegPage1(12)=>
      DANGLING(100), outputRegPage1(11)=>DANGLING(101), outputRegPage1(10)=>
      DANGLING(102), outputRegPage1(9)=>DANGLING(103), outputRegPage1(8)=>
      DANGLING(104), outputRegPage1(7)=>DANGLING(105), outputRegPage1(6)=>
      DANGLING(106), outputRegPage1(5)=>DANGLING(107), outputRegPage1(4)=>
      DANGLING(108), outputRegPage1(3)=>DANGLING(109), outputRegPage1(2)=>
      DANGLING(110), outputRegPage1(1)=>DANGLING(111), outputRegPage1(0)=>
      DANGLING(112), outputRegPage2(15)=>DANGLING(113), outputRegPage2(14)=>
      DANGLING(114), outputRegPage2(13)=>DANGLING(115), outputRegPage2(12)=>
      DANGLING(116), outputRegPage2(11)=>DANGLING(117), outputRegPage2(10)=>
      DANGLING(118), outputRegPage2(9)=>DANGLING(119), outputRegPage2(8)=>
      DANGLING(120), outputRegPage2(7)=>DANGLING(121), outputRegPage2(6)=>
      DANGLING(122), outputRegPage2(5)=>DANGLING(123), outputRegPage2(4)=>
      DANGLING(124), outputRegPage2(3)=>DANGLING(125), outputRegPage2(2)=>
      DANGLING(126), outputRegPage2(1)=>DANGLING(127), outputRegPage2(0)=>
      DANGLING(128), outFilter(7)=>filter_15_7, outFilter(6)=>filter_15_6, 
      outFilter(5)=>filter_15_5, outFilter(4)=>filter_15_4, outFilter(3)=>
      filter_15_3, outFilter(2)=>filter_15_2, outFilter(1)=>filter_15_1, 
      outFilter(0)=>filter_15_0);
   regFileMap_loop1_0_regRowMap_loop1_4_regUnitMap : RegUnit_8_16
       port map ( filterBus(7)=>filterBus(39), filterBus(6)=>filterBus(38), 
      filterBus(5)=>filterBus(37), filterBus(4)=>filterBus(36), filterBus(3)
      =>filterBus(35), filterBus(2)=>filterBus(34), filterBus(1)=>
      filterBus(33), filterBus(0)=>filterBus(32), windowBus(15)=>
      windowBus(79), windowBus(14)=>windowBus(78), windowBus(13)=>
      windowBus(77), windowBus(12)=>windowBus(76), windowBus(11)=>
      windowBus(75), windowBus(10)=>windowBus(74), windowBus(9)=>
      windowBus(73), windowBus(8)=>windowBus(72), windowBus(7)=>
      windowBus(71), windowBus(6)=>windowBus(70), windowBus(5)=>
      windowBus(69), windowBus(4)=>windowBus(68), windowBus(3)=>
      windowBus(67), windowBus(2)=>windowBus(66), windowBus(1)=>
      windowBus(65), windowBus(0)=>windowBus(64), regPage1NextUnit(15)=>
      regFileMap_page1Out_9_15, regPage1NextUnit(14)=>
      regFileMap_page1Out_9_14, regPage1NextUnit(13)=>
      regFileMap_page1Out_9_13, regPage1NextUnit(12)=>
      regFileMap_page1Out_9_12, regPage1NextUnit(11)=>
      regFileMap_page1Out_9_11, regPage1NextUnit(10)=>
      regFileMap_page1Out_9_10, regPage1NextUnit(9)=>regFileMap_page1Out_9_9, 
      regPage1NextUnit(8)=>regFileMap_page1Out_9_8, regPage1NextUnit(7)=>
      regFileMap_page1Out_9_7, regPage1NextUnit(6)=>regFileMap_page1Out_9_6, 
      regPage1NextUnit(5)=>regFileMap_page1Out_9_5, regPage1NextUnit(4)=>
      regFileMap_page1Out_9_4, regPage1NextUnit(3)=>regFileMap_page1Out_9_3, 
      regPage1NextUnit(2)=>regFileMap_page1Out_9_2, regPage1NextUnit(1)=>
      regFileMap_page1Out_9_1, regPage1NextUnit(0)=>regFileMap_page1Out_9_0, 
      regPage2NextUnit(15)=>regFileMap_page2Out_9_15, regPage2NextUnit(14)=>
      regFileMap_page2Out_9_14, regPage2NextUnit(13)=>
      regFileMap_page2Out_9_13, regPage2NextUnit(12)=>
      regFileMap_page2Out_9_12, regPage2NextUnit(11)=>
      regFileMap_page2Out_9_11, regPage2NextUnit(10)=>
      regFileMap_page2Out_9_10, regPage2NextUnit(9)=>regFileMap_page2Out_9_9, 
      regPage2NextUnit(8)=>regFileMap_page2Out_9_8, regPage2NextUnit(7)=>
      regFileMap_page2Out_9_7, regPage2NextUnit(6)=>regFileMap_page2Out_9_6, 
      regPage2NextUnit(5)=>regFileMap_page2Out_9_5, regPage2NextUnit(4)=>
      regFileMap_page2Out_9_4, regPage2NextUnit(3)=>regFileMap_page2Out_9_3, 
      regPage2NextUnit(2)=>regFileMap_page2Out_9_2, regPage2NextUnit(1)=>
      regFileMap_page2Out_9_1, regPage2NextUnit(0)=>regFileMap_page2Out_9_0, 
      clk=>clk, rst=>rst, enableRegPage1=>regFileMap_page1Enables_0, 
      enableRegPage2=>regFileMap_page2Enables_0, enableRegFilter=>nx5330, 
      page1ReadBusOrPage2=>shift2To1, page2ReadBusOrPage1=>shift1To2, 
      pageTurn=>pageTurn, outRegPage(15)=>currentPage_16_15, outRegPage(14)
      =>currentPage_16_14, outRegPage(13)=>currentPage_16_13, outRegPage(12)
      =>currentPage_16_12, outRegPage(11)=>currentPage_16_11, outRegPage(10)
      =>currentPage_16_10, outRegPage(9)=>currentPage_16_9, outRegPage(8)=>
      currentPage_16_8, outRegPage(7)=>currentPage_16_7, outRegPage(6)=>
      currentPage_16_6, outRegPage(5)=>currentPage_16_5, outRegPage(4)=>
      currentPage_16_4, outRegPage(3)=>currentPage_16_3, outRegPage(2)=>
      currentPage_16_2, outRegPage(1)=>currentPage_16_1, outRegPage(0)=>
      currentPage_16_0, outputRegPage1(15)=>DANGLING(129), 
      outputRegPage1(14)=>DANGLING(130), outputRegPage1(13)=>DANGLING(131), 
      outputRegPage1(12)=>DANGLING(132), outputRegPage1(11)=>DANGLING(133), 
      outputRegPage1(10)=>DANGLING(134), outputRegPage1(9)=>DANGLING(135), 
      outputRegPage1(8)=>DANGLING(136), outputRegPage1(7)=>DANGLING(137), 
      outputRegPage1(6)=>DANGLING(138), outputRegPage1(5)=>DANGLING(139), 
      outputRegPage1(4)=>DANGLING(140), outputRegPage1(3)=>DANGLING(141), 
      outputRegPage1(2)=>DANGLING(142), outputRegPage1(1)=>DANGLING(143), 
      outputRegPage1(0)=>DANGLING(144), outputRegPage2(15)=>DANGLING(145), 
      outputRegPage2(14)=>DANGLING(146), outputRegPage2(13)=>DANGLING(147), 
      outputRegPage2(12)=>DANGLING(148), outputRegPage2(11)=>DANGLING(149), 
      outputRegPage2(10)=>DANGLING(150), outputRegPage2(9)=>DANGLING(151), 
      outputRegPage2(8)=>DANGLING(152), outputRegPage2(7)=>DANGLING(153), 
      outputRegPage2(6)=>DANGLING(154), outputRegPage2(5)=>DANGLING(155), 
      outputRegPage2(4)=>DANGLING(156), outputRegPage2(3)=>DANGLING(157), 
      outputRegPage2(2)=>DANGLING(158), outputRegPage2(1)=>DANGLING(159), 
      outputRegPage2(0)=>DANGLING(160), outFilter(7)=>filter_16_7, 
      outFilter(6)=>filter_16_6, outFilter(5)=>filter_16_5, outFilter(4)=>
      filter_16_4, outFilter(3)=>filter_16_3, outFilter(2)=>filter_16_2, 
      outFilter(1)=>filter_16_1, outFilter(0)=>filter_16_0);
   regFileMap_loop1_1_regRowMap_loop1_0_regUnitMap : RegUnit_8_16_unfolded2
       port map ( filterBus(7)=>filterBus(7), filterBus(6)=>filterBus(6), 
      filterBus(5)=>filterBus(5), filterBus(4)=>filterBus(4), filterBus(3)=>
      filterBus(3), filterBus(2)=>filterBus(2), filterBus(1)=>filterBus(1), 
      filterBus(0)=>filterBus(0), windowBus(15)=>windowBus(15), 
      windowBus(14)=>windowBus(14), windowBus(13)=>windowBus(13), 
      windowBus(12)=>windowBus(12), windowBus(11)=>windowBus(11), 
      windowBus(10)=>windowBus(10), windowBus(9)=>windowBus(9), windowBus(8)
      =>windowBus(8), windowBus(7)=>windowBus(7), windowBus(6)=>windowBus(6), 
      windowBus(5)=>windowBus(5), windowBus(4)=>windowBus(4), windowBus(3)=>
      windowBus(3), windowBus(2)=>windowBus(2), windowBus(1)=>windowBus(1), 
      windowBus(0)=>windowBus(0), regPage1NextUnit(15)=>
      regFileMap_page1Out_10_15, regPage1NextUnit(14)=>
      regFileMap_page1Out_10_14, regPage1NextUnit(13)=>
      regFileMap_page1Out_10_13, regPage1NextUnit(12)=>
      regFileMap_page1Out_10_12, regPage1NextUnit(11)=>
      regFileMap_page1Out_10_11, regPage1NextUnit(10)=>
      regFileMap_page1Out_10_10, regPage1NextUnit(9)=>
      regFileMap_page1Out_10_9, regPage1NextUnit(8)=>
      regFileMap_page1Out_10_8, regPage1NextUnit(7)=>
      regFileMap_page1Out_10_7, regPage1NextUnit(6)=>
      regFileMap_page1Out_10_6, regPage1NextUnit(5)=>
      regFileMap_page1Out_10_5, regPage1NextUnit(4)=>
      regFileMap_page1Out_10_4, regPage1NextUnit(3)=>
      regFileMap_page1Out_10_3, regPage1NextUnit(2)=>
      regFileMap_page1Out_10_2, regPage1NextUnit(1)=>
      regFileMap_page1Out_10_1, regPage1NextUnit(0)=>
      regFileMap_page1Out_10_0, regPage2NextUnit(15)=>
      regFileMap_page2Out_10_15, regPage2NextUnit(14)=>
      regFileMap_page2Out_10_14, regPage2NextUnit(13)=>
      regFileMap_page2Out_10_13, regPage2NextUnit(12)=>
      regFileMap_page2Out_10_12, regPage2NextUnit(11)=>
      regFileMap_page2Out_10_11, regPage2NextUnit(10)=>
      regFileMap_page2Out_10_10, regPage2NextUnit(9)=>
      regFileMap_page2Out_10_9, regPage2NextUnit(8)=>
      regFileMap_page2Out_10_8, regPage2NextUnit(7)=>
      regFileMap_page2Out_10_7, regPage2NextUnit(6)=>
      regFileMap_page2Out_10_6, regPage2NextUnit(5)=>
      regFileMap_page2Out_10_5, regPage2NextUnit(4)=>
      regFileMap_page2Out_10_4, regPage2NextUnit(3)=>
      regFileMap_page2Out_10_3, regPage2NextUnit(2)=>
      regFileMap_page2Out_10_2, regPage2NextUnit(1)=>
      regFileMap_page2Out_10_1, regPage2NextUnit(0)=>
      regFileMap_page2Out_10_0, clk=>clk, rst=>rst, enableRegPage1=>
      regFileMap_page1Enables_1, enableRegPage2=>regFileMap_page2Enables_1, 
      enableRegFilter=>nx5332, page1ReadBusOrPage2=>shift2To1, 
      page2ReadBusOrPage1=>shift1To2, pageTurn=>pageTurn, outRegPage(15)=>
      currentPage_3_15, outRegPage(14)=>currentPage_3_14, outRegPage(13)=>
      currentPage_3_13, outRegPage(12)=>currentPage_3_12, outRegPage(11)=>
      currentPage_3_11, outRegPage(10)=>currentPage_3_10, outRegPage(9)=>
      currentPage_3_9, outRegPage(8)=>currentPage_3_8, outRegPage(7)=>
      currentPage_3_7, outRegPage(6)=>currentPage_3_6, outRegPage(5)=>
      currentPage_3_5, outRegPage(4)=>currentPage_3_4, outRegPage(3)=>
      currentPage_3_3, outRegPage(2)=>currentPage_3_2, outRegPage(1)=>
      currentPage_3_1, outRegPage(0)=>currentPage_3_0, outputRegPage1(15)=>
      regFileMap_page1Out_5_15, outputRegPage1(14)=>regFileMap_page1Out_5_14, 
      outputRegPage1(13)=>regFileMap_page1Out_5_13, outputRegPage1(12)=>
      regFileMap_page1Out_5_12, outputRegPage1(11)=>regFileMap_page1Out_5_11, 
      outputRegPage1(10)=>regFileMap_page1Out_5_10, outputRegPage1(9)=>
      regFileMap_page1Out_5_9, outputRegPage1(8)=>regFileMap_page1Out_5_8, 
      outputRegPage1(7)=>regFileMap_page1Out_5_7, outputRegPage1(6)=>
      regFileMap_page1Out_5_6, outputRegPage1(5)=>regFileMap_page1Out_5_5, 
      outputRegPage1(4)=>regFileMap_page1Out_5_4, outputRegPage1(3)=>
      regFileMap_page1Out_5_3, outputRegPage1(2)=>regFileMap_page1Out_5_2, 
      outputRegPage1(1)=>regFileMap_page1Out_5_1, outputRegPage1(0)=>
      regFileMap_page1Out_5_0, outputRegPage2(15)=>regFileMap_page2Out_5_15, 
      outputRegPage2(14)=>regFileMap_page2Out_5_14, outputRegPage2(13)=>
      regFileMap_page2Out_5_13, outputRegPage2(12)=>regFileMap_page2Out_5_12, 
      outputRegPage2(11)=>regFileMap_page2Out_5_11, outputRegPage2(10)=>
      regFileMap_page2Out_5_10, outputRegPage2(9)=>regFileMap_page2Out_5_9, 
      outputRegPage2(8)=>regFileMap_page2Out_5_8, outputRegPage2(7)=>
      regFileMap_page2Out_5_7, outputRegPage2(6)=>regFileMap_page2Out_5_6, 
      outputRegPage2(5)=>regFileMap_page2Out_5_5, outputRegPage2(4)=>
      regFileMap_page2Out_5_4, outputRegPage2(3)=>regFileMap_page2Out_5_3, 
      outputRegPage2(2)=>regFileMap_page2Out_5_2, outputRegPage2(1)=>
      regFileMap_page2Out_5_1, outputRegPage2(0)=>regFileMap_page2Out_5_0, 
      outFilter(7)=>filter_3_7, outFilter(6)=>filter_3_6, outFilter(5)=>
      filter_3_5, outFilter(4)=>filter_3_4, outFilter(3)=>filter_3_3, 
      outFilter(2)=>filter_3_2, outFilter(1)=>filter_3_1, outFilter(0)=>
      filter_3_0);
   regFileMap_loop1_1_regRowMap_loop1_1_regUnitMap : RegUnit_8_16_unfolded2
       port map ( filterBus(7)=>filterBus(15), filterBus(6)=>filterBus(14), 
      filterBus(5)=>filterBus(13), filterBus(4)=>filterBus(12), filterBus(3)
      =>filterBus(11), filterBus(2)=>filterBus(10), filterBus(1)=>
      filterBus(9), filterBus(0)=>filterBus(8), windowBus(15)=>windowBus(31), 
      windowBus(14)=>windowBus(30), windowBus(13)=>windowBus(29), 
      windowBus(12)=>windowBus(28), windowBus(11)=>windowBus(27), 
      windowBus(10)=>windowBus(26), windowBus(9)=>windowBus(25), 
      windowBus(8)=>windowBus(24), windowBus(7)=>windowBus(23), windowBus(6)
      =>windowBus(22), windowBus(5)=>windowBus(21), windowBus(4)=>
      windowBus(20), windowBus(3)=>windowBus(19), windowBus(2)=>
      windowBus(18), windowBus(1)=>windowBus(17), windowBus(0)=>
      windowBus(16), regPage1NextUnit(15)=>regFileMap_page1Out_11_15, 
      regPage1NextUnit(14)=>regFileMap_page1Out_11_14, regPage1NextUnit(13)
      =>regFileMap_page1Out_11_13, regPage1NextUnit(12)=>
      regFileMap_page1Out_11_12, regPage1NextUnit(11)=>
      regFileMap_page1Out_11_11, regPage1NextUnit(10)=>
      regFileMap_page1Out_11_10, regPage1NextUnit(9)=>
      regFileMap_page1Out_11_9, regPage1NextUnit(8)=>
      regFileMap_page1Out_11_8, regPage1NextUnit(7)=>
      regFileMap_page1Out_11_7, regPage1NextUnit(6)=>
      regFileMap_page1Out_11_6, regPage1NextUnit(5)=>
      regFileMap_page1Out_11_5, regPage1NextUnit(4)=>
      regFileMap_page1Out_11_4, regPage1NextUnit(3)=>
      regFileMap_page1Out_11_3, regPage1NextUnit(2)=>
      regFileMap_page1Out_11_2, regPage1NextUnit(1)=>
      regFileMap_page1Out_11_1, regPage1NextUnit(0)=>
      regFileMap_page1Out_11_0, regPage2NextUnit(15)=>
      regFileMap_page2Out_11_15, regPage2NextUnit(14)=>
      regFileMap_page2Out_11_14, regPage2NextUnit(13)=>
      regFileMap_page2Out_11_13, regPage2NextUnit(12)=>
      regFileMap_page2Out_11_12, regPage2NextUnit(11)=>
      regFileMap_page2Out_11_11, regPage2NextUnit(10)=>
      regFileMap_page2Out_11_10, regPage2NextUnit(9)=>
      regFileMap_page2Out_11_9, regPage2NextUnit(8)=>
      regFileMap_page2Out_11_8, regPage2NextUnit(7)=>
      regFileMap_page2Out_11_7, regPage2NextUnit(6)=>
      regFileMap_page2Out_11_6, regPage2NextUnit(5)=>
      regFileMap_page2Out_11_5, regPage2NextUnit(4)=>
      regFileMap_page2Out_11_4, regPage2NextUnit(3)=>
      regFileMap_page2Out_11_3, regPage2NextUnit(2)=>
      regFileMap_page2Out_11_2, regPage2NextUnit(1)=>
      regFileMap_page2Out_11_1, regPage2NextUnit(0)=>
      regFileMap_page2Out_11_0, clk=>clk, rst=>rst, enableRegPage1=>
      regFileMap_page1Enables_1, enableRegPage2=>regFileMap_page2Enables_1, 
      enableRegFilter=>nx5332, page1ReadBusOrPage2=>shift2To1, 
      page2ReadBusOrPage1=>shift1To2, pageTurn=>pageTurn, outRegPage(15)=>
      currentPage_4_15, outRegPage(14)=>currentPage_4_14, outRegPage(13)=>
      currentPage_4_13, outRegPage(12)=>currentPage_4_12, outRegPage(11)=>
      currentPage_4_11, outRegPage(10)=>currentPage_4_10, outRegPage(9)=>
      currentPage_4_9, outRegPage(8)=>currentPage_4_8, outRegPage(7)=>
      currentPage_4_7, outRegPage(6)=>currentPage_4_6, outRegPage(5)=>
      currentPage_4_5, outRegPage(4)=>currentPage_4_4, outRegPage(3)=>
      currentPage_4_3, outRegPage(2)=>currentPage_4_2, outRegPage(1)=>
      currentPage_4_1, outRegPage(0)=>currentPage_4_0, outputRegPage1(15)=>
      regFileMap_page1Out_6_15, outputRegPage1(14)=>regFileMap_page1Out_6_14, 
      outputRegPage1(13)=>regFileMap_page1Out_6_13, outputRegPage1(12)=>
      regFileMap_page1Out_6_12, outputRegPage1(11)=>regFileMap_page1Out_6_11, 
      outputRegPage1(10)=>regFileMap_page1Out_6_10, outputRegPage1(9)=>
      regFileMap_page1Out_6_9, outputRegPage1(8)=>regFileMap_page1Out_6_8, 
      outputRegPage1(7)=>regFileMap_page1Out_6_7, outputRegPage1(6)=>
      regFileMap_page1Out_6_6, outputRegPage1(5)=>regFileMap_page1Out_6_5, 
      outputRegPage1(4)=>regFileMap_page1Out_6_4, outputRegPage1(3)=>
      regFileMap_page1Out_6_3, outputRegPage1(2)=>regFileMap_page1Out_6_2, 
      outputRegPage1(1)=>regFileMap_page1Out_6_1, outputRegPage1(0)=>
      regFileMap_page1Out_6_0, outputRegPage2(15)=>regFileMap_page2Out_6_15, 
      outputRegPage2(14)=>regFileMap_page2Out_6_14, outputRegPage2(13)=>
      regFileMap_page2Out_6_13, outputRegPage2(12)=>regFileMap_page2Out_6_12, 
      outputRegPage2(11)=>regFileMap_page2Out_6_11, outputRegPage2(10)=>
      regFileMap_page2Out_6_10, outputRegPage2(9)=>regFileMap_page2Out_6_9, 
      outputRegPage2(8)=>regFileMap_page2Out_6_8, outputRegPage2(7)=>
      regFileMap_page2Out_6_7, outputRegPage2(6)=>regFileMap_page2Out_6_6, 
      outputRegPage2(5)=>regFileMap_page2Out_6_5, outputRegPage2(4)=>
      regFileMap_page2Out_6_4, outputRegPage2(3)=>regFileMap_page2Out_6_3, 
      outputRegPage2(2)=>regFileMap_page2Out_6_2, outputRegPage2(1)=>
      regFileMap_page2Out_6_1, outputRegPage2(0)=>regFileMap_page2Out_6_0, 
      outFilter(7)=>filter_4_7, outFilter(6)=>filter_4_6, outFilter(5)=>
      filter_4_5, outFilter(4)=>filter_4_4, outFilter(3)=>filter_4_3, 
      outFilter(2)=>filter_4_2, outFilter(1)=>filter_4_1, outFilter(0)=>
      filter_4_0);
   regFileMap_loop1_1_regRowMap_loop1_2_regUnitMap : RegUnit_8_16_unfolded2
       port map ( filterBus(7)=>filterBus(23), filterBus(6)=>filterBus(22), 
      filterBus(5)=>filterBus(21), filterBus(4)=>filterBus(20), filterBus(3)
      =>filterBus(19), filterBus(2)=>filterBus(18), filterBus(1)=>
      filterBus(17), filterBus(0)=>filterBus(16), windowBus(15)=>
      windowBus(47), windowBus(14)=>windowBus(46), windowBus(13)=>
      windowBus(45), windowBus(12)=>windowBus(44), windowBus(11)=>
      windowBus(43), windowBus(10)=>windowBus(42), windowBus(9)=>
      windowBus(41), windowBus(8)=>windowBus(40), windowBus(7)=>
      windowBus(39), windowBus(6)=>windowBus(38), windowBus(5)=>
      windowBus(37), windowBus(4)=>windowBus(36), windowBus(3)=>
      windowBus(35), windowBus(2)=>windowBus(34), windowBus(1)=>
      windowBus(33), windowBus(0)=>windowBus(32), regPage1NextUnit(15)=>
      regFileMap_page1Out_12_15, regPage1NextUnit(14)=>
      regFileMap_page1Out_12_14, regPage1NextUnit(13)=>
      regFileMap_page1Out_12_13, regPage1NextUnit(12)=>
      regFileMap_page1Out_12_12, regPage1NextUnit(11)=>
      regFileMap_page1Out_12_11, regPage1NextUnit(10)=>
      regFileMap_page1Out_12_10, regPage1NextUnit(9)=>
      regFileMap_page1Out_12_9, regPage1NextUnit(8)=>
      regFileMap_page1Out_12_8, regPage1NextUnit(7)=>
      regFileMap_page1Out_12_7, regPage1NextUnit(6)=>
      regFileMap_page1Out_12_6, regPage1NextUnit(5)=>
      regFileMap_page1Out_12_5, regPage1NextUnit(4)=>
      regFileMap_page1Out_12_4, regPage1NextUnit(3)=>
      regFileMap_page1Out_12_3, regPage1NextUnit(2)=>
      regFileMap_page1Out_12_2, regPage1NextUnit(1)=>
      regFileMap_page1Out_12_1, regPage1NextUnit(0)=>
      regFileMap_page1Out_12_0, regPage2NextUnit(15)=>
      regFileMap_page2Out_12_15, regPage2NextUnit(14)=>
      regFileMap_page2Out_12_14, regPage2NextUnit(13)=>
      regFileMap_page2Out_12_13, regPage2NextUnit(12)=>
      regFileMap_page2Out_12_12, regPage2NextUnit(11)=>
      regFileMap_page2Out_12_11, regPage2NextUnit(10)=>
      regFileMap_page2Out_12_10, regPage2NextUnit(9)=>
      regFileMap_page2Out_12_9, regPage2NextUnit(8)=>
      regFileMap_page2Out_12_8, regPage2NextUnit(7)=>
      regFileMap_page2Out_12_7, regPage2NextUnit(6)=>
      regFileMap_page2Out_12_6, regPage2NextUnit(5)=>
      regFileMap_page2Out_12_5, regPage2NextUnit(4)=>
      regFileMap_page2Out_12_4, regPage2NextUnit(3)=>
      regFileMap_page2Out_12_3, regPage2NextUnit(2)=>
      regFileMap_page2Out_12_2, regPage2NextUnit(1)=>
      regFileMap_page2Out_12_1, regPage2NextUnit(0)=>
      regFileMap_page2Out_12_0, clk=>clk, rst=>rst, enableRegPage1=>
      regFileMap_page1Enables_1, enableRegPage2=>regFileMap_page2Enables_1, 
      enableRegFilter=>nx5332, page1ReadBusOrPage2=>shift2To1, 
      page2ReadBusOrPage1=>shift1To2, pageTurn=>pageTurn, outRegPage(15)=>
      currentPage_5_15, outRegPage(14)=>currentPage_5_14, outRegPage(13)=>
      currentPage_5_13, outRegPage(12)=>currentPage_5_12, outRegPage(11)=>
      currentPage_5_11, outRegPage(10)=>currentPage_5_10, outRegPage(9)=>
      currentPage_5_9, outRegPage(8)=>currentPage_5_8, outRegPage(7)=>
      currentPage_5_7, outRegPage(6)=>currentPage_5_6, outRegPage(5)=>
      currentPage_5_5, outRegPage(4)=>currentPage_5_4, outRegPage(3)=>
      currentPage_5_3, outRegPage(2)=>currentPage_5_2, outRegPage(1)=>
      currentPage_5_1, outRegPage(0)=>currentPage_5_0, outputRegPage1(15)=>
      regFileMap_page1Out_7_15, outputRegPage1(14)=>regFileMap_page1Out_7_14, 
      outputRegPage1(13)=>regFileMap_page1Out_7_13, outputRegPage1(12)=>
      regFileMap_page1Out_7_12, outputRegPage1(11)=>regFileMap_page1Out_7_11, 
      outputRegPage1(10)=>regFileMap_page1Out_7_10, outputRegPage1(9)=>
      regFileMap_page1Out_7_9, outputRegPage1(8)=>regFileMap_page1Out_7_8, 
      outputRegPage1(7)=>regFileMap_page1Out_7_7, outputRegPage1(6)=>
      regFileMap_page1Out_7_6, outputRegPage1(5)=>regFileMap_page1Out_7_5, 
      outputRegPage1(4)=>regFileMap_page1Out_7_4, outputRegPage1(3)=>
      regFileMap_page1Out_7_3, outputRegPage1(2)=>regFileMap_page1Out_7_2, 
      outputRegPage1(1)=>regFileMap_page1Out_7_1, outputRegPage1(0)=>
      regFileMap_page1Out_7_0, outputRegPage2(15)=>regFileMap_page2Out_7_15, 
      outputRegPage2(14)=>regFileMap_page2Out_7_14, outputRegPage2(13)=>
      regFileMap_page2Out_7_13, outputRegPage2(12)=>regFileMap_page2Out_7_12, 
      outputRegPage2(11)=>regFileMap_page2Out_7_11, outputRegPage2(10)=>
      regFileMap_page2Out_7_10, outputRegPage2(9)=>regFileMap_page2Out_7_9, 
      outputRegPage2(8)=>regFileMap_page2Out_7_8, outputRegPage2(7)=>
      regFileMap_page2Out_7_7, outputRegPage2(6)=>regFileMap_page2Out_7_6, 
      outputRegPage2(5)=>regFileMap_page2Out_7_5, outputRegPage2(4)=>
      regFileMap_page2Out_7_4, outputRegPage2(3)=>regFileMap_page2Out_7_3, 
      outputRegPage2(2)=>regFileMap_page2Out_7_2, outputRegPage2(1)=>
      regFileMap_page2Out_7_1, outputRegPage2(0)=>regFileMap_page2Out_7_0, 
      outFilter(7)=>filter_5_7, outFilter(6)=>filter_5_6, outFilter(5)=>
      filter_5_5, outFilter(4)=>filter_5_4, outFilter(3)=>filter_5_3, 
      outFilter(2)=>filter_5_2, outFilter(1)=>filter_5_1, outFilter(0)=>
      filter_5_0);
   regFileMap_loop1_1_regRowMap_loop1_3_regUnitMap : RegUnit_8_16_unfolded2
       port map ( filterBus(7)=>filterBus(31), filterBus(6)=>filterBus(30), 
      filterBus(5)=>filterBus(29), filterBus(4)=>filterBus(28), filterBus(3)
      =>filterBus(27), filterBus(2)=>filterBus(26), filterBus(1)=>
      filterBus(25), filterBus(0)=>filterBus(24), windowBus(15)=>
      windowBus(63), windowBus(14)=>windowBus(62), windowBus(13)=>
      windowBus(61), windowBus(12)=>windowBus(60), windowBus(11)=>
      windowBus(59), windowBus(10)=>windowBus(58), windowBus(9)=>
      windowBus(57), windowBus(8)=>windowBus(56), windowBus(7)=>
      windowBus(55), windowBus(6)=>windowBus(54), windowBus(5)=>
      windowBus(53), windowBus(4)=>windowBus(52), windowBus(3)=>
      windowBus(51), windowBus(2)=>windowBus(50), windowBus(1)=>
      windowBus(49), windowBus(0)=>windowBus(48), regPage1NextUnit(15)=>
      regFileMap_page1Out_13_15, regPage1NextUnit(14)=>
      regFileMap_page1Out_13_14, regPage1NextUnit(13)=>
      regFileMap_page1Out_13_13, regPage1NextUnit(12)=>
      regFileMap_page1Out_13_12, regPage1NextUnit(11)=>
      regFileMap_page1Out_13_11, regPage1NextUnit(10)=>
      regFileMap_page1Out_13_10, regPage1NextUnit(9)=>
      regFileMap_page1Out_13_9, regPage1NextUnit(8)=>
      regFileMap_page1Out_13_8, regPage1NextUnit(7)=>
      regFileMap_page1Out_13_7, regPage1NextUnit(6)=>
      regFileMap_page1Out_13_6, regPage1NextUnit(5)=>
      regFileMap_page1Out_13_5, regPage1NextUnit(4)=>
      regFileMap_page1Out_13_4, regPage1NextUnit(3)=>
      regFileMap_page1Out_13_3, regPage1NextUnit(2)=>
      regFileMap_page1Out_13_2, regPage1NextUnit(1)=>
      regFileMap_page1Out_13_1, regPage1NextUnit(0)=>
      regFileMap_page1Out_13_0, regPage2NextUnit(15)=>
      regFileMap_page2Out_13_15, regPage2NextUnit(14)=>
      regFileMap_page2Out_13_14, regPage2NextUnit(13)=>
      regFileMap_page2Out_13_13, regPage2NextUnit(12)=>
      regFileMap_page2Out_13_12, regPage2NextUnit(11)=>
      regFileMap_page2Out_13_11, regPage2NextUnit(10)=>
      regFileMap_page2Out_13_10, regPage2NextUnit(9)=>
      regFileMap_page2Out_13_9, regPage2NextUnit(8)=>
      regFileMap_page2Out_13_8, regPage2NextUnit(7)=>
      regFileMap_page2Out_13_7, regPage2NextUnit(6)=>
      regFileMap_page2Out_13_6, regPage2NextUnit(5)=>
      regFileMap_page2Out_13_5, regPage2NextUnit(4)=>
      regFileMap_page2Out_13_4, regPage2NextUnit(3)=>
      regFileMap_page2Out_13_3, regPage2NextUnit(2)=>
      regFileMap_page2Out_13_2, regPage2NextUnit(1)=>
      regFileMap_page2Out_13_1, regPage2NextUnit(0)=>
      regFileMap_page2Out_13_0, clk=>clk, rst=>rst, enableRegPage1=>
      regFileMap_page1Enables_1, enableRegPage2=>regFileMap_page2Enables_1, 
      enableRegFilter=>nx5334, page1ReadBusOrPage2=>shift2To1, 
      page2ReadBusOrPage1=>shift1To2, pageTurn=>pageTurn, outRegPage(15)=>
      currentPage_17_15, outRegPage(14)=>currentPage_17_14, outRegPage(13)=>
      currentPage_17_13, outRegPage(12)=>currentPage_17_12, outRegPage(11)=>
      currentPage_17_11, outRegPage(10)=>currentPage_17_10, outRegPage(9)=>
      currentPage_17_9, outRegPage(8)=>currentPage_17_8, outRegPage(7)=>
      currentPage_17_7, outRegPage(6)=>currentPage_17_6, outRegPage(5)=>
      currentPage_17_5, outRegPage(4)=>currentPage_17_4, outRegPage(3)=>
      currentPage_17_3, outRegPage(2)=>currentPage_17_2, outRegPage(1)=>
      currentPage_17_1, outRegPage(0)=>currentPage_17_0, outputRegPage1(15)
      =>regFileMap_page1Out_8_15, outputRegPage1(14)=>
      regFileMap_page1Out_8_14, outputRegPage1(13)=>regFileMap_page1Out_8_13, 
      outputRegPage1(12)=>regFileMap_page1Out_8_12, outputRegPage1(11)=>
      regFileMap_page1Out_8_11, outputRegPage1(10)=>regFileMap_page1Out_8_10, 
      outputRegPage1(9)=>regFileMap_page1Out_8_9, outputRegPage1(8)=>
      regFileMap_page1Out_8_8, outputRegPage1(7)=>regFileMap_page1Out_8_7, 
      outputRegPage1(6)=>regFileMap_page1Out_8_6, outputRegPage1(5)=>
      regFileMap_page1Out_8_5, outputRegPage1(4)=>regFileMap_page1Out_8_4, 
      outputRegPage1(3)=>regFileMap_page1Out_8_3, outputRegPage1(2)=>
      regFileMap_page1Out_8_2, outputRegPage1(1)=>regFileMap_page1Out_8_1, 
      outputRegPage1(0)=>regFileMap_page1Out_8_0, outputRegPage2(15)=>
      regFileMap_page2Out_8_15, outputRegPage2(14)=>regFileMap_page2Out_8_14, 
      outputRegPage2(13)=>regFileMap_page2Out_8_13, outputRegPage2(12)=>
      regFileMap_page2Out_8_12, outputRegPage2(11)=>regFileMap_page2Out_8_11, 
      outputRegPage2(10)=>regFileMap_page2Out_8_10, outputRegPage2(9)=>
      regFileMap_page2Out_8_9, outputRegPage2(8)=>regFileMap_page2Out_8_8, 
      outputRegPage2(7)=>regFileMap_page2Out_8_7, outputRegPage2(6)=>
      regFileMap_page2Out_8_6, outputRegPage2(5)=>regFileMap_page2Out_8_5, 
      outputRegPage2(4)=>regFileMap_page2Out_8_4, outputRegPage2(3)=>
      regFileMap_page2Out_8_3, outputRegPage2(2)=>regFileMap_page2Out_8_2, 
      outputRegPage2(1)=>regFileMap_page2Out_8_1, outputRegPage2(0)=>
      regFileMap_page2Out_8_0, outFilter(7)=>filter_17_7, outFilter(6)=>
      filter_17_6, outFilter(5)=>filter_17_5, outFilter(4)=>filter_17_4, 
      outFilter(3)=>filter_17_3, outFilter(2)=>filter_17_2, outFilter(1)=>
      filter_17_1, outFilter(0)=>filter_17_0);
   regFileMap_loop1_1_regRowMap_loop1_4_regUnitMap : RegUnit_8_16_unfolded2
       port map ( filterBus(7)=>filterBus(39), filterBus(6)=>filterBus(38), 
      filterBus(5)=>filterBus(37), filterBus(4)=>filterBus(36), filterBus(3)
      =>filterBus(35), filterBus(2)=>filterBus(34), filterBus(1)=>
      filterBus(33), filterBus(0)=>filterBus(32), windowBus(15)=>
      windowBus(79), windowBus(14)=>windowBus(78), windowBus(13)=>
      windowBus(77), windowBus(12)=>windowBus(76), windowBus(11)=>
      windowBus(75), windowBus(10)=>windowBus(74), windowBus(9)=>
      windowBus(73), windowBus(8)=>windowBus(72), windowBus(7)=>
      windowBus(71), windowBus(6)=>windowBus(70), windowBus(5)=>
      windowBus(69), windowBus(4)=>windowBus(68), windowBus(3)=>
      windowBus(67), windowBus(2)=>windowBus(66), windowBus(1)=>
      windowBus(65), windowBus(0)=>windowBus(64), regPage1NextUnit(15)=>
      regFileMap_page1Out_14_15, regPage1NextUnit(14)=>
      regFileMap_page1Out_14_14, regPage1NextUnit(13)=>
      regFileMap_page1Out_14_13, regPage1NextUnit(12)=>
      regFileMap_page1Out_14_12, regPage1NextUnit(11)=>
      regFileMap_page1Out_14_11, regPage1NextUnit(10)=>
      regFileMap_page1Out_14_10, regPage1NextUnit(9)=>
      regFileMap_page1Out_14_9, regPage1NextUnit(8)=>
      regFileMap_page1Out_14_8, regPage1NextUnit(7)=>
      regFileMap_page1Out_14_7, regPage1NextUnit(6)=>
      regFileMap_page1Out_14_6, regPage1NextUnit(5)=>
      regFileMap_page1Out_14_5, regPage1NextUnit(4)=>
      regFileMap_page1Out_14_4, regPage1NextUnit(3)=>
      regFileMap_page1Out_14_3, regPage1NextUnit(2)=>
      regFileMap_page1Out_14_2, regPage1NextUnit(1)=>
      regFileMap_page1Out_14_1, regPage1NextUnit(0)=>
      regFileMap_page1Out_14_0, regPage2NextUnit(15)=>
      regFileMap_page2Out_14_15, regPage2NextUnit(14)=>
      regFileMap_page2Out_14_14, regPage2NextUnit(13)=>
      regFileMap_page2Out_14_13, regPage2NextUnit(12)=>
      regFileMap_page2Out_14_12, regPage2NextUnit(11)=>
      regFileMap_page2Out_14_11, regPage2NextUnit(10)=>
      regFileMap_page2Out_14_10, regPage2NextUnit(9)=>
      regFileMap_page2Out_14_9, regPage2NextUnit(8)=>
      regFileMap_page2Out_14_8, regPage2NextUnit(7)=>
      regFileMap_page2Out_14_7, regPage2NextUnit(6)=>
      regFileMap_page2Out_14_6, regPage2NextUnit(5)=>
      regFileMap_page2Out_14_5, regPage2NextUnit(4)=>
      regFileMap_page2Out_14_4, regPage2NextUnit(3)=>
      regFileMap_page2Out_14_3, regPage2NextUnit(2)=>
      regFileMap_page2Out_14_2, regPage2NextUnit(1)=>
      regFileMap_page2Out_14_1, regPage2NextUnit(0)=>
      regFileMap_page2Out_14_0, clk=>clk, rst=>rst, enableRegPage1=>
      regFileMap_page1Enables_1, enableRegPage2=>regFileMap_page2Enables_1, 
      enableRegFilter=>nx5334, page1ReadBusOrPage2=>shift2To1, 
      page2ReadBusOrPage1=>shift1To2, pageTurn=>pageTurn, outRegPage(15)=>
      currentPage_18_15, outRegPage(14)=>currentPage_18_14, outRegPage(13)=>
      currentPage_18_13, outRegPage(12)=>currentPage_18_12, outRegPage(11)=>
      currentPage_18_11, outRegPage(10)=>currentPage_18_10, outRegPage(9)=>
      currentPage_18_9, outRegPage(8)=>currentPage_18_8, outRegPage(7)=>
      currentPage_18_7, outRegPage(6)=>currentPage_18_6, outRegPage(5)=>
      currentPage_18_5, outRegPage(4)=>currentPage_18_4, outRegPage(3)=>
      currentPage_18_3, outRegPage(2)=>currentPage_18_2, outRegPage(1)=>
      currentPage_18_1, outRegPage(0)=>currentPage_18_0, outputRegPage1(15)
      =>regFileMap_page1Out_9_15, outputRegPage1(14)=>
      regFileMap_page1Out_9_14, outputRegPage1(13)=>regFileMap_page1Out_9_13, 
      outputRegPage1(12)=>regFileMap_page1Out_9_12, outputRegPage1(11)=>
      regFileMap_page1Out_9_11, outputRegPage1(10)=>regFileMap_page1Out_9_10, 
      outputRegPage1(9)=>regFileMap_page1Out_9_9, outputRegPage1(8)=>
      regFileMap_page1Out_9_8, outputRegPage1(7)=>regFileMap_page1Out_9_7, 
      outputRegPage1(6)=>regFileMap_page1Out_9_6, outputRegPage1(5)=>
      regFileMap_page1Out_9_5, outputRegPage1(4)=>regFileMap_page1Out_9_4, 
      outputRegPage1(3)=>regFileMap_page1Out_9_3, outputRegPage1(2)=>
      regFileMap_page1Out_9_2, outputRegPage1(1)=>regFileMap_page1Out_9_1, 
      outputRegPage1(0)=>regFileMap_page1Out_9_0, outputRegPage2(15)=>
      regFileMap_page2Out_9_15, outputRegPage2(14)=>regFileMap_page2Out_9_14, 
      outputRegPage2(13)=>regFileMap_page2Out_9_13, outputRegPage2(12)=>
      regFileMap_page2Out_9_12, outputRegPage2(11)=>regFileMap_page2Out_9_11, 
      outputRegPage2(10)=>regFileMap_page2Out_9_10, outputRegPage2(9)=>
      regFileMap_page2Out_9_9, outputRegPage2(8)=>regFileMap_page2Out_9_8, 
      outputRegPage2(7)=>regFileMap_page2Out_9_7, outputRegPage2(6)=>
      regFileMap_page2Out_9_6, outputRegPage2(5)=>regFileMap_page2Out_9_5, 
      outputRegPage2(4)=>regFileMap_page2Out_9_4, outputRegPage2(3)=>
      regFileMap_page2Out_9_3, outputRegPage2(2)=>regFileMap_page2Out_9_2, 
      outputRegPage2(1)=>regFileMap_page2Out_9_1, outputRegPage2(0)=>
      regFileMap_page2Out_9_0, outFilter(7)=>filter_18_7, outFilter(6)=>
      filter_18_6, outFilter(5)=>filter_18_5, outFilter(4)=>filter_18_4, 
      outFilter(3)=>filter_18_3, outFilter(2)=>filter_18_2, outFilter(1)=>
      filter_18_1, outFilter(0)=>filter_18_0);
   regFileMap_loop1_2_regRowMap_loop1_0_regUnitMap : RegUnit_8_16_unfolded2
       port map ( filterBus(7)=>filterBus(7), filterBus(6)=>filterBus(6), 
      filterBus(5)=>filterBus(5), filterBus(4)=>filterBus(4), filterBus(3)=>
      filterBus(3), filterBus(2)=>filterBus(2), filterBus(1)=>filterBus(1), 
      filterBus(0)=>filterBus(0), windowBus(15)=>windowBus(15), 
      windowBus(14)=>windowBus(14), windowBus(13)=>windowBus(13), 
      windowBus(12)=>windowBus(12), windowBus(11)=>windowBus(11), 
      windowBus(10)=>windowBus(10), windowBus(9)=>windowBus(9), windowBus(8)
      =>windowBus(8), windowBus(7)=>windowBus(7), windowBus(6)=>windowBus(6), 
      windowBus(5)=>windowBus(5), windowBus(4)=>windowBus(4), windowBus(3)=>
      windowBus(3), windowBus(2)=>windowBus(2), windowBus(1)=>windowBus(1), 
      windowBus(0)=>windowBus(0), regPage1NextUnit(15)=>
      regFileMap_page1Out_15_15, regPage1NextUnit(14)=>
      regFileMap_page1Out_15_14, regPage1NextUnit(13)=>
      regFileMap_page1Out_15_13, regPage1NextUnit(12)=>
      regFileMap_page1Out_15_12, regPage1NextUnit(11)=>
      regFileMap_page1Out_15_11, regPage1NextUnit(10)=>
      regFileMap_page1Out_15_10, regPage1NextUnit(9)=>
      regFileMap_page1Out_15_9, regPage1NextUnit(8)=>
      regFileMap_page1Out_15_8, regPage1NextUnit(7)=>
      regFileMap_page1Out_15_7, regPage1NextUnit(6)=>
      regFileMap_page1Out_15_6, regPage1NextUnit(5)=>
      regFileMap_page1Out_15_5, regPage1NextUnit(4)=>
      regFileMap_page1Out_15_4, regPage1NextUnit(3)=>
      regFileMap_page1Out_15_3, regPage1NextUnit(2)=>
      regFileMap_page1Out_15_2, regPage1NextUnit(1)=>
      regFileMap_page1Out_15_1, regPage1NextUnit(0)=>
      regFileMap_page1Out_15_0, regPage2NextUnit(15)=>
      regFileMap_page2Out_15_15, regPage2NextUnit(14)=>
      regFileMap_page2Out_15_14, regPage2NextUnit(13)=>
      regFileMap_page2Out_15_13, regPage2NextUnit(12)=>
      regFileMap_page2Out_15_12, regPage2NextUnit(11)=>
      regFileMap_page2Out_15_11, regPage2NextUnit(10)=>
      regFileMap_page2Out_15_10, regPage2NextUnit(9)=>
      regFileMap_page2Out_15_9, regPage2NextUnit(8)=>
      regFileMap_page2Out_15_8, regPage2NextUnit(7)=>
      regFileMap_page2Out_15_7, regPage2NextUnit(6)=>
      regFileMap_page2Out_15_6, regPage2NextUnit(5)=>
      regFileMap_page2Out_15_5, regPage2NextUnit(4)=>
      regFileMap_page2Out_15_4, regPage2NextUnit(3)=>
      regFileMap_page2Out_15_3, regPage2NextUnit(2)=>
      regFileMap_page2Out_15_2, regPage2NextUnit(1)=>
      regFileMap_page2Out_15_1, regPage2NextUnit(0)=>
      regFileMap_page2Out_15_0, clk=>clk, rst=>rst, enableRegPage1=>
      regFileMap_page1Enables_2, enableRegPage2=>regFileMap_page2Enables_2, 
      enableRegFilter=>nx5336, page1ReadBusOrPage2=>shift2To1, 
      page2ReadBusOrPage1=>shift1To2, pageTurn=>pageTurn, outRegPage(15)=>
      currentPage_6_15, outRegPage(14)=>currentPage_6_14, outRegPage(13)=>
      currentPage_6_13, outRegPage(12)=>currentPage_6_12, outRegPage(11)=>
      currentPage_6_11, outRegPage(10)=>currentPage_6_10, outRegPage(9)=>
      currentPage_6_9, outRegPage(8)=>currentPage_6_8, outRegPage(7)=>
      currentPage_6_7, outRegPage(6)=>currentPage_6_6, outRegPage(5)=>
      currentPage_6_5, outRegPage(4)=>currentPage_6_4, outRegPage(3)=>
      currentPage_6_3, outRegPage(2)=>currentPage_6_2, outRegPage(1)=>
      currentPage_6_1, outRegPage(0)=>currentPage_6_0, outputRegPage1(15)=>
      regFileMap_page1Out_10_15, outputRegPage1(14)=>
      regFileMap_page1Out_10_14, outputRegPage1(13)=>
      regFileMap_page1Out_10_13, outputRegPage1(12)=>
      regFileMap_page1Out_10_12, outputRegPage1(11)=>
      regFileMap_page1Out_10_11, outputRegPage1(10)=>
      regFileMap_page1Out_10_10, outputRegPage1(9)=>regFileMap_page1Out_10_9, 
      outputRegPage1(8)=>regFileMap_page1Out_10_8, outputRegPage1(7)=>
      regFileMap_page1Out_10_7, outputRegPage1(6)=>regFileMap_page1Out_10_6, 
      outputRegPage1(5)=>regFileMap_page1Out_10_5, outputRegPage1(4)=>
      regFileMap_page1Out_10_4, outputRegPage1(3)=>regFileMap_page1Out_10_3, 
      outputRegPage1(2)=>regFileMap_page1Out_10_2, outputRegPage1(1)=>
      regFileMap_page1Out_10_1, outputRegPage1(0)=>regFileMap_page1Out_10_0, 
      outputRegPage2(15)=>regFileMap_page2Out_10_15, outputRegPage2(14)=>
      regFileMap_page2Out_10_14, outputRegPage2(13)=>
      regFileMap_page2Out_10_13, outputRegPage2(12)=>
      regFileMap_page2Out_10_12, outputRegPage2(11)=>
      regFileMap_page2Out_10_11, outputRegPage2(10)=>
      regFileMap_page2Out_10_10, outputRegPage2(9)=>regFileMap_page2Out_10_9, 
      outputRegPage2(8)=>regFileMap_page2Out_10_8, outputRegPage2(7)=>
      regFileMap_page2Out_10_7, outputRegPage2(6)=>regFileMap_page2Out_10_6, 
      outputRegPage2(5)=>regFileMap_page2Out_10_5, outputRegPage2(4)=>
      regFileMap_page2Out_10_4, outputRegPage2(3)=>regFileMap_page2Out_10_3, 
      outputRegPage2(2)=>regFileMap_page2Out_10_2, outputRegPage2(1)=>
      regFileMap_page2Out_10_1, outputRegPage2(0)=>regFileMap_page2Out_10_0, 
      outFilter(7)=>filter_6_7, outFilter(6)=>filter_6_6, outFilter(5)=>
      filter_6_5, outFilter(4)=>filter_6_4, outFilter(3)=>filter_6_3, 
      outFilter(2)=>filter_6_2, outFilter(1)=>filter_6_1, outFilter(0)=>
      filter_6_0);
   regFileMap_loop1_2_regRowMap_loop1_1_regUnitMap : RegUnit_8_16_unfolded2
       port map ( filterBus(7)=>filterBus(15), filterBus(6)=>filterBus(14), 
      filterBus(5)=>filterBus(13), filterBus(4)=>filterBus(12), filterBus(3)
      =>filterBus(11), filterBus(2)=>filterBus(10), filterBus(1)=>
      filterBus(9), filterBus(0)=>filterBus(8), windowBus(15)=>windowBus(31), 
      windowBus(14)=>windowBus(30), windowBus(13)=>windowBus(29), 
      windowBus(12)=>windowBus(28), windowBus(11)=>windowBus(27), 
      windowBus(10)=>windowBus(26), windowBus(9)=>windowBus(25), 
      windowBus(8)=>windowBus(24), windowBus(7)=>windowBus(23), windowBus(6)
      =>windowBus(22), windowBus(5)=>windowBus(21), windowBus(4)=>
      windowBus(20), windowBus(3)=>windowBus(19), windowBus(2)=>
      windowBus(18), windowBus(1)=>windowBus(17), windowBus(0)=>
      windowBus(16), regPage1NextUnit(15)=>regFileMap_page1Out_16_15, 
      regPage1NextUnit(14)=>regFileMap_page1Out_16_14, regPage1NextUnit(13)
      =>regFileMap_page1Out_16_13, regPage1NextUnit(12)=>
      regFileMap_page1Out_16_12, regPage1NextUnit(11)=>
      regFileMap_page1Out_16_11, regPage1NextUnit(10)=>
      regFileMap_page1Out_16_10, regPage1NextUnit(9)=>
      regFileMap_page1Out_16_9, regPage1NextUnit(8)=>
      regFileMap_page1Out_16_8, regPage1NextUnit(7)=>
      regFileMap_page1Out_16_7, regPage1NextUnit(6)=>
      regFileMap_page1Out_16_6, regPage1NextUnit(5)=>
      regFileMap_page1Out_16_5, regPage1NextUnit(4)=>
      regFileMap_page1Out_16_4, regPage1NextUnit(3)=>
      regFileMap_page1Out_16_3, regPage1NextUnit(2)=>
      regFileMap_page1Out_16_2, regPage1NextUnit(1)=>
      regFileMap_page1Out_16_1, regPage1NextUnit(0)=>
      regFileMap_page1Out_16_0, regPage2NextUnit(15)=>
      regFileMap_page2Out_16_15, regPage2NextUnit(14)=>
      regFileMap_page2Out_16_14, regPage2NextUnit(13)=>
      regFileMap_page2Out_16_13, regPage2NextUnit(12)=>
      regFileMap_page2Out_16_12, regPage2NextUnit(11)=>
      regFileMap_page2Out_16_11, regPage2NextUnit(10)=>
      regFileMap_page2Out_16_10, regPage2NextUnit(9)=>
      regFileMap_page2Out_16_9, regPage2NextUnit(8)=>
      regFileMap_page2Out_16_8, regPage2NextUnit(7)=>
      regFileMap_page2Out_16_7, regPage2NextUnit(6)=>
      regFileMap_page2Out_16_6, regPage2NextUnit(5)=>
      regFileMap_page2Out_16_5, regPage2NextUnit(4)=>
      regFileMap_page2Out_16_4, regPage2NextUnit(3)=>
      regFileMap_page2Out_16_3, regPage2NextUnit(2)=>
      regFileMap_page2Out_16_2, regPage2NextUnit(1)=>
      regFileMap_page2Out_16_1, regPage2NextUnit(0)=>
      regFileMap_page2Out_16_0, clk=>clk, rst=>rst, enableRegPage1=>
      regFileMap_page1Enables_2, enableRegPage2=>regFileMap_page2Enables_2, 
      enableRegFilter=>nx5336, page1ReadBusOrPage2=>shift2To1, 
      page2ReadBusOrPage1=>shift1To2, pageTurn=>pageTurn, outRegPage(15)=>
      currentPage_7_15, outRegPage(14)=>currentPage_7_14, outRegPage(13)=>
      currentPage_7_13, outRegPage(12)=>currentPage_7_12, outRegPage(11)=>
      currentPage_7_11, outRegPage(10)=>currentPage_7_10, outRegPage(9)=>
      currentPage_7_9, outRegPage(8)=>currentPage_7_8, outRegPage(7)=>
      currentPage_7_7, outRegPage(6)=>currentPage_7_6, outRegPage(5)=>
      currentPage_7_5, outRegPage(4)=>currentPage_7_4, outRegPage(3)=>
      currentPage_7_3, outRegPage(2)=>currentPage_7_2, outRegPage(1)=>
      currentPage_7_1, outRegPage(0)=>currentPage_7_0, outputRegPage1(15)=>
      regFileMap_page1Out_11_15, outputRegPage1(14)=>
      regFileMap_page1Out_11_14, outputRegPage1(13)=>
      regFileMap_page1Out_11_13, outputRegPage1(12)=>
      regFileMap_page1Out_11_12, outputRegPage1(11)=>
      regFileMap_page1Out_11_11, outputRegPage1(10)=>
      regFileMap_page1Out_11_10, outputRegPage1(9)=>regFileMap_page1Out_11_9, 
      outputRegPage1(8)=>regFileMap_page1Out_11_8, outputRegPage1(7)=>
      regFileMap_page1Out_11_7, outputRegPage1(6)=>regFileMap_page1Out_11_6, 
      outputRegPage1(5)=>regFileMap_page1Out_11_5, outputRegPage1(4)=>
      regFileMap_page1Out_11_4, outputRegPage1(3)=>regFileMap_page1Out_11_3, 
      outputRegPage1(2)=>regFileMap_page1Out_11_2, outputRegPage1(1)=>
      regFileMap_page1Out_11_1, outputRegPage1(0)=>regFileMap_page1Out_11_0, 
      outputRegPage2(15)=>regFileMap_page2Out_11_15, outputRegPage2(14)=>
      regFileMap_page2Out_11_14, outputRegPage2(13)=>
      regFileMap_page2Out_11_13, outputRegPage2(12)=>
      regFileMap_page2Out_11_12, outputRegPage2(11)=>
      regFileMap_page2Out_11_11, outputRegPage2(10)=>
      regFileMap_page2Out_11_10, outputRegPage2(9)=>regFileMap_page2Out_11_9, 
      outputRegPage2(8)=>regFileMap_page2Out_11_8, outputRegPage2(7)=>
      regFileMap_page2Out_11_7, outputRegPage2(6)=>regFileMap_page2Out_11_6, 
      outputRegPage2(5)=>regFileMap_page2Out_11_5, outputRegPage2(4)=>
      regFileMap_page2Out_11_4, outputRegPage2(3)=>regFileMap_page2Out_11_3, 
      outputRegPage2(2)=>regFileMap_page2Out_11_2, outputRegPage2(1)=>
      regFileMap_page2Out_11_1, outputRegPage2(0)=>regFileMap_page2Out_11_0, 
      outFilter(7)=>filter_7_7, outFilter(6)=>filter_7_6, outFilter(5)=>
      filter_7_5, outFilter(4)=>filter_7_4, outFilter(3)=>filter_7_3, 
      outFilter(2)=>filter_7_2, outFilter(1)=>filter_7_1, outFilter(0)=>
      filter_7_0);
   regFileMap_loop1_2_regRowMap_loop1_2_regUnitMap : RegUnit_8_16_unfolded2
       port map ( filterBus(7)=>filterBus(23), filterBus(6)=>filterBus(22), 
      filterBus(5)=>filterBus(21), filterBus(4)=>filterBus(20), filterBus(3)
      =>filterBus(19), filterBus(2)=>filterBus(18), filterBus(1)=>
      filterBus(17), filterBus(0)=>filterBus(16), windowBus(15)=>
      windowBus(47), windowBus(14)=>windowBus(46), windowBus(13)=>
      windowBus(45), windowBus(12)=>windowBus(44), windowBus(11)=>
      windowBus(43), windowBus(10)=>windowBus(42), windowBus(9)=>
      windowBus(41), windowBus(8)=>windowBus(40), windowBus(7)=>
      windowBus(39), windowBus(6)=>windowBus(38), windowBus(5)=>
      windowBus(37), windowBus(4)=>windowBus(36), windowBus(3)=>
      windowBus(35), windowBus(2)=>windowBus(34), windowBus(1)=>
      windowBus(33), windowBus(0)=>windowBus(32), regPage1NextUnit(15)=>
      regFileMap_page1Out_17_15, regPage1NextUnit(14)=>
      regFileMap_page1Out_17_14, regPage1NextUnit(13)=>
      regFileMap_page1Out_17_13, regPage1NextUnit(12)=>
      regFileMap_page1Out_17_12, regPage1NextUnit(11)=>
      regFileMap_page1Out_17_11, regPage1NextUnit(10)=>
      regFileMap_page1Out_17_10, regPage1NextUnit(9)=>
      regFileMap_page1Out_17_9, regPage1NextUnit(8)=>
      regFileMap_page1Out_17_8, regPage1NextUnit(7)=>
      regFileMap_page1Out_17_7, regPage1NextUnit(6)=>
      regFileMap_page1Out_17_6, regPage1NextUnit(5)=>
      regFileMap_page1Out_17_5, regPage1NextUnit(4)=>
      regFileMap_page1Out_17_4, regPage1NextUnit(3)=>
      regFileMap_page1Out_17_3, regPage1NextUnit(2)=>
      regFileMap_page1Out_17_2, regPage1NextUnit(1)=>
      regFileMap_page1Out_17_1, regPage1NextUnit(0)=>
      regFileMap_page1Out_17_0, regPage2NextUnit(15)=>
      regFileMap_page2Out_17_15, regPage2NextUnit(14)=>
      regFileMap_page2Out_17_14, regPage2NextUnit(13)=>
      regFileMap_page2Out_17_13, regPage2NextUnit(12)=>
      regFileMap_page2Out_17_12, regPage2NextUnit(11)=>
      regFileMap_page2Out_17_11, regPage2NextUnit(10)=>
      regFileMap_page2Out_17_10, regPage2NextUnit(9)=>
      regFileMap_page2Out_17_9, regPage2NextUnit(8)=>
      regFileMap_page2Out_17_8, regPage2NextUnit(7)=>
      regFileMap_page2Out_17_7, regPage2NextUnit(6)=>
      regFileMap_page2Out_17_6, regPage2NextUnit(5)=>
      regFileMap_page2Out_17_5, regPage2NextUnit(4)=>
      regFileMap_page2Out_17_4, regPage2NextUnit(3)=>
      regFileMap_page2Out_17_3, regPage2NextUnit(2)=>
      regFileMap_page2Out_17_2, regPage2NextUnit(1)=>
      regFileMap_page2Out_17_1, regPage2NextUnit(0)=>
      regFileMap_page2Out_17_0, clk=>clk, rst=>rst, enableRegPage1=>
      regFileMap_page1Enables_2, enableRegPage2=>regFileMap_page2Enables_2, 
      enableRegFilter=>nx5336, page1ReadBusOrPage2=>shift2To1, 
      page2ReadBusOrPage1=>shift1To2, pageTurn=>pageTurn, outRegPage(15)=>
      currentPage_8_15, outRegPage(14)=>currentPage_8_14, outRegPage(13)=>
      currentPage_8_13, outRegPage(12)=>currentPage_8_12, outRegPage(11)=>
      currentPage_8_11, outRegPage(10)=>currentPage_8_10, outRegPage(9)=>
      currentPage_8_9, outRegPage(8)=>currentPage_8_8, outRegPage(7)=>
      currentPage_8_7, outRegPage(6)=>currentPage_8_6, outRegPage(5)=>
      currentPage_8_5, outRegPage(4)=>currentPage_8_4, outRegPage(3)=>
      currentPage_8_3, outRegPage(2)=>currentPage_8_2, outRegPage(1)=>
      currentPage_8_1, outRegPage(0)=>currentPage_8_0, outputRegPage1(15)=>
      regFileMap_page1Out_12_15, outputRegPage1(14)=>
      regFileMap_page1Out_12_14, outputRegPage1(13)=>
      regFileMap_page1Out_12_13, outputRegPage1(12)=>
      regFileMap_page1Out_12_12, outputRegPage1(11)=>
      regFileMap_page1Out_12_11, outputRegPage1(10)=>
      regFileMap_page1Out_12_10, outputRegPage1(9)=>regFileMap_page1Out_12_9, 
      outputRegPage1(8)=>regFileMap_page1Out_12_8, outputRegPage1(7)=>
      regFileMap_page1Out_12_7, outputRegPage1(6)=>regFileMap_page1Out_12_6, 
      outputRegPage1(5)=>regFileMap_page1Out_12_5, outputRegPage1(4)=>
      regFileMap_page1Out_12_4, outputRegPage1(3)=>regFileMap_page1Out_12_3, 
      outputRegPage1(2)=>regFileMap_page1Out_12_2, outputRegPage1(1)=>
      regFileMap_page1Out_12_1, outputRegPage1(0)=>regFileMap_page1Out_12_0, 
      outputRegPage2(15)=>regFileMap_page2Out_12_15, outputRegPage2(14)=>
      regFileMap_page2Out_12_14, outputRegPage2(13)=>
      regFileMap_page2Out_12_13, outputRegPage2(12)=>
      regFileMap_page2Out_12_12, outputRegPage2(11)=>
      regFileMap_page2Out_12_11, outputRegPage2(10)=>
      regFileMap_page2Out_12_10, outputRegPage2(9)=>regFileMap_page2Out_12_9, 
      outputRegPage2(8)=>regFileMap_page2Out_12_8, outputRegPage2(7)=>
      regFileMap_page2Out_12_7, outputRegPage2(6)=>regFileMap_page2Out_12_6, 
      outputRegPage2(5)=>regFileMap_page2Out_12_5, outputRegPage2(4)=>
      regFileMap_page2Out_12_4, outputRegPage2(3)=>regFileMap_page2Out_12_3, 
      outputRegPage2(2)=>regFileMap_page2Out_12_2, outputRegPage2(1)=>
      regFileMap_page2Out_12_1, outputRegPage2(0)=>regFileMap_page2Out_12_0, 
      outFilter(7)=>filter_8_7, outFilter(6)=>filter_8_6, outFilter(5)=>
      filter_8_5, outFilter(4)=>filter_8_4, outFilter(3)=>filter_8_3, 
      outFilter(2)=>filter_8_2, outFilter(1)=>filter_8_1, outFilter(0)=>
      filter_8_0);
   regFileMap_loop1_2_regRowMap_loop1_3_regUnitMap : RegUnit_8_16_unfolded2
       port map ( filterBus(7)=>filterBus(31), filterBus(6)=>filterBus(30), 
      filterBus(5)=>filterBus(29), filterBus(4)=>filterBus(28), filterBus(3)
      =>filterBus(27), filterBus(2)=>filterBus(26), filterBus(1)=>
      filterBus(25), filterBus(0)=>filterBus(24), windowBus(15)=>
      windowBus(63), windowBus(14)=>windowBus(62), windowBus(13)=>
      windowBus(61), windowBus(12)=>windowBus(60), windowBus(11)=>
      windowBus(59), windowBus(10)=>windowBus(58), windowBus(9)=>
      windowBus(57), windowBus(8)=>windowBus(56), windowBus(7)=>
      windowBus(55), windowBus(6)=>windowBus(54), windowBus(5)=>
      windowBus(53), windowBus(4)=>windowBus(52), windowBus(3)=>
      windowBus(51), windowBus(2)=>windowBus(50), windowBus(1)=>
      windowBus(49), windowBus(0)=>windowBus(48), regPage1NextUnit(15)=>
      regFileMap_page1Out_18_15, regPage1NextUnit(14)=>
      regFileMap_page1Out_18_14, regPage1NextUnit(13)=>
      regFileMap_page1Out_18_13, regPage1NextUnit(12)=>
      regFileMap_page1Out_18_12, regPage1NextUnit(11)=>
      regFileMap_page1Out_18_11, regPage1NextUnit(10)=>
      regFileMap_page1Out_18_10, regPage1NextUnit(9)=>
      regFileMap_page1Out_18_9, regPage1NextUnit(8)=>
      regFileMap_page1Out_18_8, regPage1NextUnit(7)=>
      regFileMap_page1Out_18_7, regPage1NextUnit(6)=>
      regFileMap_page1Out_18_6, regPage1NextUnit(5)=>
      regFileMap_page1Out_18_5, regPage1NextUnit(4)=>
      regFileMap_page1Out_18_4, regPage1NextUnit(3)=>
      regFileMap_page1Out_18_3, regPage1NextUnit(2)=>
      regFileMap_page1Out_18_2, regPage1NextUnit(1)=>
      regFileMap_page1Out_18_1, regPage1NextUnit(0)=>
      regFileMap_page1Out_18_0, regPage2NextUnit(15)=>
      regFileMap_page2Out_18_15, regPage2NextUnit(14)=>
      regFileMap_page2Out_18_14, regPage2NextUnit(13)=>
      regFileMap_page2Out_18_13, regPage2NextUnit(12)=>
      regFileMap_page2Out_18_12, regPage2NextUnit(11)=>
      regFileMap_page2Out_18_11, regPage2NextUnit(10)=>
      regFileMap_page2Out_18_10, regPage2NextUnit(9)=>
      regFileMap_page2Out_18_9, regPage2NextUnit(8)=>
      regFileMap_page2Out_18_8, regPage2NextUnit(7)=>
      regFileMap_page2Out_18_7, regPage2NextUnit(6)=>
      regFileMap_page2Out_18_6, regPage2NextUnit(5)=>
      regFileMap_page2Out_18_5, regPage2NextUnit(4)=>
      regFileMap_page2Out_18_4, regPage2NextUnit(3)=>
      regFileMap_page2Out_18_3, regPage2NextUnit(2)=>
      regFileMap_page2Out_18_2, regPage2NextUnit(1)=>
      regFileMap_page2Out_18_1, regPage2NextUnit(0)=>
      regFileMap_page2Out_18_0, clk=>clk, rst=>rst, enableRegPage1=>
      regFileMap_page1Enables_2, enableRegPage2=>regFileMap_page2Enables_2, 
      enableRegFilter=>nx5338, page1ReadBusOrPage2=>shift2To1, 
      page2ReadBusOrPage1=>shift1To2, pageTurn=>pageTurn, outRegPage(15)=>
      currentPage_19_15, outRegPage(14)=>currentPage_19_14, outRegPage(13)=>
      currentPage_19_13, outRegPage(12)=>currentPage_19_12, outRegPage(11)=>
      currentPage_19_11, outRegPage(10)=>currentPage_19_10, outRegPage(9)=>
      currentPage_19_9, outRegPage(8)=>currentPage_19_8, outRegPage(7)=>
      currentPage_19_7, outRegPage(6)=>currentPage_19_6, outRegPage(5)=>
      currentPage_19_5, outRegPage(4)=>currentPage_19_4, outRegPage(3)=>
      currentPage_19_3, outRegPage(2)=>currentPage_19_2, outRegPage(1)=>
      currentPage_19_1, outRegPage(0)=>currentPage_19_0, outputRegPage1(15)
      =>regFileMap_page1Out_13_15, outputRegPage1(14)=>
      regFileMap_page1Out_13_14, outputRegPage1(13)=>
      regFileMap_page1Out_13_13, outputRegPage1(12)=>
      regFileMap_page1Out_13_12, outputRegPage1(11)=>
      regFileMap_page1Out_13_11, outputRegPage1(10)=>
      regFileMap_page1Out_13_10, outputRegPage1(9)=>regFileMap_page1Out_13_9, 
      outputRegPage1(8)=>regFileMap_page1Out_13_8, outputRegPage1(7)=>
      regFileMap_page1Out_13_7, outputRegPage1(6)=>regFileMap_page1Out_13_6, 
      outputRegPage1(5)=>regFileMap_page1Out_13_5, outputRegPage1(4)=>
      regFileMap_page1Out_13_4, outputRegPage1(3)=>regFileMap_page1Out_13_3, 
      outputRegPage1(2)=>regFileMap_page1Out_13_2, outputRegPage1(1)=>
      regFileMap_page1Out_13_1, outputRegPage1(0)=>regFileMap_page1Out_13_0, 
      outputRegPage2(15)=>regFileMap_page2Out_13_15, outputRegPage2(14)=>
      regFileMap_page2Out_13_14, outputRegPage2(13)=>
      regFileMap_page2Out_13_13, outputRegPage2(12)=>
      regFileMap_page2Out_13_12, outputRegPage2(11)=>
      regFileMap_page2Out_13_11, outputRegPage2(10)=>
      regFileMap_page2Out_13_10, outputRegPage2(9)=>regFileMap_page2Out_13_9, 
      outputRegPage2(8)=>regFileMap_page2Out_13_8, outputRegPage2(7)=>
      regFileMap_page2Out_13_7, outputRegPage2(6)=>regFileMap_page2Out_13_6, 
      outputRegPage2(5)=>regFileMap_page2Out_13_5, outputRegPage2(4)=>
      regFileMap_page2Out_13_4, outputRegPage2(3)=>regFileMap_page2Out_13_3, 
      outputRegPage2(2)=>regFileMap_page2Out_13_2, outputRegPage2(1)=>
      regFileMap_page2Out_13_1, outputRegPage2(0)=>regFileMap_page2Out_13_0, 
      outFilter(7)=>filter_19_7, outFilter(6)=>filter_19_6, outFilter(5)=>
      filter_19_5, outFilter(4)=>filter_19_4, outFilter(3)=>filter_19_3, 
      outFilter(2)=>filter_19_2, outFilter(1)=>filter_19_1, outFilter(0)=>
      filter_19_0);
   regFileMap_loop1_2_regRowMap_loop1_4_regUnitMap : RegUnit_8_16_unfolded2
       port map ( filterBus(7)=>filterBus(39), filterBus(6)=>filterBus(38), 
      filterBus(5)=>filterBus(37), filterBus(4)=>filterBus(36), filterBus(3)
      =>filterBus(35), filterBus(2)=>filterBus(34), filterBus(1)=>
      filterBus(33), filterBus(0)=>filterBus(32), windowBus(15)=>
      windowBus(79), windowBus(14)=>windowBus(78), windowBus(13)=>
      windowBus(77), windowBus(12)=>windowBus(76), windowBus(11)=>
      windowBus(75), windowBus(10)=>windowBus(74), windowBus(9)=>
      windowBus(73), windowBus(8)=>windowBus(72), windowBus(7)=>
      windowBus(71), windowBus(6)=>windowBus(70), windowBus(5)=>
      windowBus(69), windowBus(4)=>windowBus(68), windowBus(3)=>
      windowBus(67), windowBus(2)=>windowBus(66), windowBus(1)=>
      windowBus(65), windowBus(0)=>windowBus(64), regPage1NextUnit(15)=>
      regFileMap_page1Out_19_15, regPage1NextUnit(14)=>
      regFileMap_page1Out_19_14, regPage1NextUnit(13)=>
      regFileMap_page1Out_19_13, regPage1NextUnit(12)=>
      regFileMap_page1Out_19_12, regPage1NextUnit(11)=>
      regFileMap_page1Out_19_11, regPage1NextUnit(10)=>
      regFileMap_page1Out_19_10, regPage1NextUnit(9)=>
      regFileMap_page1Out_19_9, regPage1NextUnit(8)=>
      regFileMap_page1Out_19_8, regPage1NextUnit(7)=>
      regFileMap_page1Out_19_7, regPage1NextUnit(6)=>
      regFileMap_page1Out_19_6, regPage1NextUnit(5)=>
      regFileMap_page1Out_19_5, regPage1NextUnit(4)=>
      regFileMap_page1Out_19_4, regPage1NextUnit(3)=>
      regFileMap_page1Out_19_3, regPage1NextUnit(2)=>
      regFileMap_page1Out_19_2, regPage1NextUnit(1)=>
      regFileMap_page1Out_19_1, regPage1NextUnit(0)=>
      regFileMap_page1Out_19_0, regPage2NextUnit(15)=>
      regFileMap_page2Out_19_15, regPage2NextUnit(14)=>
      regFileMap_page2Out_19_14, regPage2NextUnit(13)=>
      regFileMap_page2Out_19_13, regPage2NextUnit(12)=>
      regFileMap_page2Out_19_12, regPage2NextUnit(11)=>
      regFileMap_page2Out_19_11, regPage2NextUnit(10)=>
      regFileMap_page2Out_19_10, regPage2NextUnit(9)=>
      regFileMap_page2Out_19_9, regPage2NextUnit(8)=>
      regFileMap_page2Out_19_8, regPage2NextUnit(7)=>
      regFileMap_page2Out_19_7, regPage2NextUnit(6)=>
      regFileMap_page2Out_19_6, regPage2NextUnit(5)=>
      regFileMap_page2Out_19_5, regPage2NextUnit(4)=>
      regFileMap_page2Out_19_4, regPage2NextUnit(3)=>
      regFileMap_page2Out_19_3, regPage2NextUnit(2)=>
      regFileMap_page2Out_19_2, regPage2NextUnit(1)=>
      regFileMap_page2Out_19_1, regPage2NextUnit(0)=>
      regFileMap_page2Out_19_0, clk=>clk, rst=>rst, enableRegPage1=>
      regFileMap_page1Enables_2, enableRegPage2=>regFileMap_page2Enables_2, 
      enableRegFilter=>nx5338, page1ReadBusOrPage2=>shift2To1, 
      page2ReadBusOrPage1=>shift1To2, pageTurn=>pageTurn, outRegPage(15)=>
      currentPage_20_15, outRegPage(14)=>currentPage_20_14, outRegPage(13)=>
      currentPage_20_13, outRegPage(12)=>currentPage_20_12, outRegPage(11)=>
      currentPage_20_11, outRegPage(10)=>currentPage_20_10, outRegPage(9)=>
      currentPage_20_9, outRegPage(8)=>currentPage_20_8, outRegPage(7)=>
      currentPage_20_7, outRegPage(6)=>currentPage_20_6, outRegPage(5)=>
      currentPage_20_5, outRegPage(4)=>currentPage_20_4, outRegPage(3)=>
      currentPage_20_3, outRegPage(2)=>currentPage_20_2, outRegPage(1)=>
      currentPage_20_1, outRegPage(0)=>currentPage_20_0, outputRegPage1(15)
      =>regFileMap_page1Out_14_15, outputRegPage1(14)=>
      regFileMap_page1Out_14_14, outputRegPage1(13)=>
      regFileMap_page1Out_14_13, outputRegPage1(12)=>
      regFileMap_page1Out_14_12, outputRegPage1(11)=>
      regFileMap_page1Out_14_11, outputRegPage1(10)=>
      regFileMap_page1Out_14_10, outputRegPage1(9)=>regFileMap_page1Out_14_9, 
      outputRegPage1(8)=>regFileMap_page1Out_14_8, outputRegPage1(7)=>
      regFileMap_page1Out_14_7, outputRegPage1(6)=>regFileMap_page1Out_14_6, 
      outputRegPage1(5)=>regFileMap_page1Out_14_5, outputRegPage1(4)=>
      regFileMap_page1Out_14_4, outputRegPage1(3)=>regFileMap_page1Out_14_3, 
      outputRegPage1(2)=>regFileMap_page1Out_14_2, outputRegPage1(1)=>
      regFileMap_page1Out_14_1, outputRegPage1(0)=>regFileMap_page1Out_14_0, 
      outputRegPage2(15)=>regFileMap_page2Out_14_15, outputRegPage2(14)=>
      regFileMap_page2Out_14_14, outputRegPage2(13)=>
      regFileMap_page2Out_14_13, outputRegPage2(12)=>
      regFileMap_page2Out_14_12, outputRegPage2(11)=>
      regFileMap_page2Out_14_11, outputRegPage2(10)=>
      regFileMap_page2Out_14_10, outputRegPage2(9)=>regFileMap_page2Out_14_9, 
      outputRegPage2(8)=>regFileMap_page2Out_14_8, outputRegPage2(7)=>
      regFileMap_page2Out_14_7, outputRegPage2(6)=>regFileMap_page2Out_14_6, 
      outputRegPage2(5)=>regFileMap_page2Out_14_5, outputRegPage2(4)=>
      regFileMap_page2Out_14_4, outputRegPage2(3)=>regFileMap_page2Out_14_3, 
      outputRegPage2(2)=>regFileMap_page2Out_14_2, outputRegPage2(1)=>
      regFileMap_page2Out_14_1, outputRegPage2(0)=>regFileMap_page2Out_14_0, 
      outFilter(7)=>filter_20_7, outFilter(6)=>filter_20_6, outFilter(5)=>
      filter_20_5, outFilter(4)=>filter_20_4, outFilter(3)=>filter_20_3, 
      outFilter(2)=>filter_20_2, outFilter(1)=>filter_20_1, outFilter(0)=>
      filter_20_0);
   regFileMap_loop1_3_regRowMap_loop1_0_regUnitMap : RegUnit_8_16_unfolded2
       port map ( filterBus(7)=>filterBus(7), filterBus(6)=>filterBus(6), 
      filterBus(5)=>filterBus(5), filterBus(4)=>filterBus(4), filterBus(3)=>
      filterBus(3), filterBus(2)=>filterBus(2), filterBus(1)=>filterBus(1), 
      filterBus(0)=>filterBus(0), windowBus(15)=>windowBus(15), 
      windowBus(14)=>windowBus(14), windowBus(13)=>windowBus(13), 
      windowBus(12)=>windowBus(12), windowBus(11)=>windowBus(11), 
      windowBus(10)=>windowBus(10), windowBus(9)=>windowBus(9), windowBus(8)
      =>windowBus(8), windowBus(7)=>windowBus(7), windowBus(6)=>windowBus(6), 
      windowBus(5)=>windowBus(5), windowBus(4)=>windowBus(4), windowBus(3)=>
      windowBus(3), windowBus(2)=>windowBus(2), windowBus(1)=>windowBus(1), 
      windowBus(0)=>windowBus(0), regPage1NextUnit(15)=>
      regFileMap_page1Out_20_15, regPage1NextUnit(14)=>
      regFileMap_page1Out_20_14, regPage1NextUnit(13)=>
      regFileMap_page1Out_20_13, regPage1NextUnit(12)=>
      regFileMap_page1Out_20_12, regPage1NextUnit(11)=>
      regFileMap_page1Out_20_11, regPage1NextUnit(10)=>
      regFileMap_page1Out_20_10, regPage1NextUnit(9)=>
      regFileMap_page1Out_20_9, regPage1NextUnit(8)=>
      regFileMap_page1Out_20_8, regPage1NextUnit(7)=>
      regFileMap_page1Out_20_7, regPage1NextUnit(6)=>
      regFileMap_page1Out_20_6, regPage1NextUnit(5)=>
      regFileMap_page1Out_20_5, regPage1NextUnit(4)=>
      regFileMap_page1Out_20_4, regPage1NextUnit(3)=>
      regFileMap_page1Out_20_3, regPage1NextUnit(2)=>
      regFileMap_page1Out_20_2, regPage1NextUnit(1)=>
      regFileMap_page1Out_20_1, regPage1NextUnit(0)=>
      regFileMap_page1Out_20_0, regPage2NextUnit(15)=>
      regFileMap_page2Out_20_15, regPage2NextUnit(14)=>
      regFileMap_page2Out_20_14, regPage2NextUnit(13)=>
      regFileMap_page2Out_20_13, regPage2NextUnit(12)=>
      regFileMap_page2Out_20_12, regPage2NextUnit(11)=>
      regFileMap_page2Out_20_11, regPage2NextUnit(10)=>
      regFileMap_page2Out_20_10, regPage2NextUnit(9)=>
      regFileMap_page2Out_20_9, regPage2NextUnit(8)=>
      regFileMap_page2Out_20_8, regPage2NextUnit(7)=>
      regFileMap_page2Out_20_7, regPage2NextUnit(6)=>
      regFileMap_page2Out_20_6, regPage2NextUnit(5)=>
      regFileMap_page2Out_20_5, regPage2NextUnit(4)=>
      regFileMap_page2Out_20_4, regPage2NextUnit(3)=>
      regFileMap_page2Out_20_3, regPage2NextUnit(2)=>
      regFileMap_page2Out_20_2, regPage2NextUnit(1)=>
      regFileMap_page2Out_20_1, regPage2NextUnit(0)=>
      regFileMap_page2Out_20_0, clk=>clk, rst=>rst, enableRegPage1=>
      regFileMap_page1Enables_3, enableRegPage2=>regFileMap_page2Enables_3, 
      enableRegFilter=>nx5340, page1ReadBusOrPage2=>shift2To1, 
      page2ReadBusOrPage1=>shift1To2, pageTurn=>pageTurn, outRegPage(15)=>
      currentPage_9_15, outRegPage(14)=>currentPage_9_14, outRegPage(13)=>
      currentPage_9_13, outRegPage(12)=>currentPage_9_12, outRegPage(11)=>
      currentPage_9_11, outRegPage(10)=>currentPage_9_10, outRegPage(9)=>
      currentPage_9_9, outRegPage(8)=>currentPage_9_8, outRegPage(7)=>
      currentPage_9_7, outRegPage(6)=>currentPage_9_6, outRegPage(5)=>
      currentPage_9_5, outRegPage(4)=>currentPage_9_4, outRegPage(3)=>
      currentPage_9_3, outRegPage(2)=>currentPage_9_2, outRegPage(1)=>
      currentPage_9_1, outRegPage(0)=>currentPage_9_0, outputRegPage1(15)=>
      regFileMap_page1Out_15_15, outputRegPage1(14)=>
      regFileMap_page1Out_15_14, outputRegPage1(13)=>
      regFileMap_page1Out_15_13, outputRegPage1(12)=>
      regFileMap_page1Out_15_12, outputRegPage1(11)=>
      regFileMap_page1Out_15_11, outputRegPage1(10)=>
      regFileMap_page1Out_15_10, outputRegPage1(9)=>regFileMap_page1Out_15_9, 
      outputRegPage1(8)=>regFileMap_page1Out_15_8, outputRegPage1(7)=>
      regFileMap_page1Out_15_7, outputRegPage1(6)=>regFileMap_page1Out_15_6, 
      outputRegPage1(5)=>regFileMap_page1Out_15_5, outputRegPage1(4)=>
      regFileMap_page1Out_15_4, outputRegPage1(3)=>regFileMap_page1Out_15_3, 
      outputRegPage1(2)=>regFileMap_page1Out_15_2, outputRegPage1(1)=>
      regFileMap_page1Out_15_1, outputRegPage1(0)=>regFileMap_page1Out_15_0, 
      outputRegPage2(15)=>regFileMap_page2Out_15_15, outputRegPage2(14)=>
      regFileMap_page2Out_15_14, outputRegPage2(13)=>
      regFileMap_page2Out_15_13, outputRegPage2(12)=>
      regFileMap_page2Out_15_12, outputRegPage2(11)=>
      regFileMap_page2Out_15_11, outputRegPage2(10)=>
      regFileMap_page2Out_15_10, outputRegPage2(9)=>regFileMap_page2Out_15_9, 
      outputRegPage2(8)=>regFileMap_page2Out_15_8, outputRegPage2(7)=>
      regFileMap_page2Out_15_7, outputRegPage2(6)=>regFileMap_page2Out_15_6, 
      outputRegPage2(5)=>regFileMap_page2Out_15_5, outputRegPage2(4)=>
      regFileMap_page2Out_15_4, outputRegPage2(3)=>regFileMap_page2Out_15_3, 
      outputRegPage2(2)=>regFileMap_page2Out_15_2, outputRegPage2(1)=>
      regFileMap_page2Out_15_1, outputRegPage2(0)=>regFileMap_page2Out_15_0, 
      outFilter(7)=>filter_9_7, outFilter(6)=>filter_9_6, outFilter(5)=>
      filter_9_5, outFilter(4)=>filter_9_4, outFilter(3)=>filter_9_3, 
      outFilter(2)=>filter_9_2, outFilter(1)=>filter_9_1, outFilter(0)=>
      filter_9_0);
   regFileMap_loop1_3_regRowMap_loop1_1_regUnitMap : RegUnit_8_16_unfolded2
       port map ( filterBus(7)=>filterBus(15), filterBus(6)=>filterBus(14), 
      filterBus(5)=>filterBus(13), filterBus(4)=>filterBus(12), filterBus(3)
      =>filterBus(11), filterBus(2)=>filterBus(10), filterBus(1)=>
      filterBus(9), filterBus(0)=>filterBus(8), windowBus(15)=>windowBus(31), 
      windowBus(14)=>windowBus(30), windowBus(13)=>windowBus(29), 
      windowBus(12)=>windowBus(28), windowBus(11)=>windowBus(27), 
      windowBus(10)=>windowBus(26), windowBus(9)=>windowBus(25), 
      windowBus(8)=>windowBus(24), windowBus(7)=>windowBus(23), windowBus(6)
      =>windowBus(22), windowBus(5)=>windowBus(21), windowBus(4)=>
      windowBus(20), windowBus(3)=>windowBus(19), windowBus(2)=>
      windowBus(18), windowBus(1)=>windowBus(17), windowBus(0)=>
      windowBus(16), regPage1NextUnit(15)=>regFileMap_page1Out_21_15, 
      regPage1NextUnit(14)=>regFileMap_page1Out_21_14, regPage1NextUnit(13)
      =>regFileMap_page1Out_21_13, regPage1NextUnit(12)=>
      regFileMap_page1Out_21_12, regPage1NextUnit(11)=>
      regFileMap_page1Out_21_11, regPage1NextUnit(10)=>
      regFileMap_page1Out_21_10, regPage1NextUnit(9)=>
      regFileMap_page1Out_21_9, regPage1NextUnit(8)=>
      regFileMap_page1Out_21_8, regPage1NextUnit(7)=>
      regFileMap_page1Out_21_7, regPage1NextUnit(6)=>
      regFileMap_page1Out_21_6, regPage1NextUnit(5)=>
      regFileMap_page1Out_21_5, regPage1NextUnit(4)=>
      regFileMap_page1Out_21_4, regPage1NextUnit(3)=>
      regFileMap_page1Out_21_3, regPage1NextUnit(2)=>
      regFileMap_page1Out_21_2, regPage1NextUnit(1)=>
      regFileMap_page1Out_21_1, regPage1NextUnit(0)=>
      regFileMap_page1Out_21_0, regPage2NextUnit(15)=>
      regFileMap_page2Out_21_15, regPage2NextUnit(14)=>
      regFileMap_page2Out_21_14, regPage2NextUnit(13)=>
      regFileMap_page2Out_21_13, regPage2NextUnit(12)=>
      regFileMap_page2Out_21_12, regPage2NextUnit(11)=>
      regFileMap_page2Out_21_11, regPage2NextUnit(10)=>
      regFileMap_page2Out_21_10, regPage2NextUnit(9)=>
      regFileMap_page2Out_21_9, regPage2NextUnit(8)=>
      regFileMap_page2Out_21_8, regPage2NextUnit(7)=>
      regFileMap_page2Out_21_7, regPage2NextUnit(6)=>
      regFileMap_page2Out_21_6, regPage2NextUnit(5)=>
      regFileMap_page2Out_21_5, regPage2NextUnit(4)=>
      regFileMap_page2Out_21_4, regPage2NextUnit(3)=>
      regFileMap_page2Out_21_3, regPage2NextUnit(2)=>
      regFileMap_page2Out_21_2, regPage2NextUnit(1)=>
      regFileMap_page2Out_21_1, regPage2NextUnit(0)=>
      regFileMap_page2Out_21_0, clk=>clk, rst=>rst, enableRegPage1=>
      regFileMap_page1Enables_3, enableRegPage2=>regFileMap_page2Enables_3, 
      enableRegFilter=>nx5340, page1ReadBusOrPage2=>shift2To1, 
      page2ReadBusOrPage1=>shift1To2, pageTurn=>pageTurn, outRegPage(15)=>
      currentPage_10_15, outRegPage(14)=>currentPage_10_14, outRegPage(13)=>
      currentPage_10_13, outRegPage(12)=>currentPage_10_12, outRegPage(11)=>
      currentPage_10_11, outRegPage(10)=>currentPage_10_10, outRegPage(9)=>
      currentPage_10_9, outRegPage(8)=>currentPage_10_8, outRegPage(7)=>
      currentPage_10_7, outRegPage(6)=>currentPage_10_6, outRegPage(5)=>
      currentPage_10_5, outRegPage(4)=>currentPage_10_4, outRegPage(3)=>
      currentPage_10_3, outRegPage(2)=>currentPage_10_2, outRegPage(1)=>
      currentPage_10_1, outRegPage(0)=>currentPage_10_0, outputRegPage1(15)
      =>regFileMap_page1Out_16_15, outputRegPage1(14)=>
      regFileMap_page1Out_16_14, outputRegPage1(13)=>
      regFileMap_page1Out_16_13, outputRegPage1(12)=>
      regFileMap_page1Out_16_12, outputRegPage1(11)=>
      regFileMap_page1Out_16_11, outputRegPage1(10)=>
      regFileMap_page1Out_16_10, outputRegPage1(9)=>regFileMap_page1Out_16_9, 
      outputRegPage1(8)=>regFileMap_page1Out_16_8, outputRegPage1(7)=>
      regFileMap_page1Out_16_7, outputRegPage1(6)=>regFileMap_page1Out_16_6, 
      outputRegPage1(5)=>regFileMap_page1Out_16_5, outputRegPage1(4)=>
      regFileMap_page1Out_16_4, outputRegPage1(3)=>regFileMap_page1Out_16_3, 
      outputRegPage1(2)=>regFileMap_page1Out_16_2, outputRegPage1(1)=>
      regFileMap_page1Out_16_1, outputRegPage1(0)=>regFileMap_page1Out_16_0, 
      outputRegPage2(15)=>regFileMap_page2Out_16_15, outputRegPage2(14)=>
      regFileMap_page2Out_16_14, outputRegPage2(13)=>
      regFileMap_page2Out_16_13, outputRegPage2(12)=>
      regFileMap_page2Out_16_12, outputRegPage2(11)=>
      regFileMap_page2Out_16_11, outputRegPage2(10)=>
      regFileMap_page2Out_16_10, outputRegPage2(9)=>regFileMap_page2Out_16_9, 
      outputRegPage2(8)=>regFileMap_page2Out_16_8, outputRegPage2(7)=>
      regFileMap_page2Out_16_7, outputRegPage2(6)=>regFileMap_page2Out_16_6, 
      outputRegPage2(5)=>regFileMap_page2Out_16_5, outputRegPage2(4)=>
      regFileMap_page2Out_16_4, outputRegPage2(3)=>regFileMap_page2Out_16_3, 
      outputRegPage2(2)=>regFileMap_page2Out_16_2, outputRegPage2(1)=>
      regFileMap_page2Out_16_1, outputRegPage2(0)=>regFileMap_page2Out_16_0, 
      outFilter(7)=>filter_10_7, outFilter(6)=>filter_10_6, outFilter(5)=>
      filter_10_5, outFilter(4)=>filter_10_4, outFilter(3)=>filter_10_3, 
      outFilter(2)=>filter_10_2, outFilter(1)=>filter_10_1, outFilter(0)=>
      filter_10_0);
   regFileMap_loop1_3_regRowMap_loop1_2_regUnitMap : RegUnit_8_16_unfolded2
       port map ( filterBus(7)=>filterBus(23), filterBus(6)=>filterBus(22), 
      filterBus(5)=>filterBus(21), filterBus(4)=>filterBus(20), filterBus(3)
      =>filterBus(19), filterBus(2)=>filterBus(18), filterBus(1)=>
      filterBus(17), filterBus(0)=>filterBus(16), windowBus(15)=>
      windowBus(47), windowBus(14)=>windowBus(46), windowBus(13)=>
      windowBus(45), windowBus(12)=>windowBus(44), windowBus(11)=>
      windowBus(43), windowBus(10)=>windowBus(42), windowBus(9)=>
      windowBus(41), windowBus(8)=>windowBus(40), windowBus(7)=>
      windowBus(39), windowBus(6)=>windowBus(38), windowBus(5)=>
      windowBus(37), windowBus(4)=>windowBus(36), windowBus(3)=>
      windowBus(35), windowBus(2)=>windowBus(34), windowBus(1)=>
      windowBus(33), windowBus(0)=>windowBus(32), regPage1NextUnit(15)=>
      regFileMap_page1Out_22_15, regPage1NextUnit(14)=>
      regFileMap_page1Out_22_14, regPage1NextUnit(13)=>
      regFileMap_page1Out_22_13, regPage1NextUnit(12)=>
      regFileMap_page1Out_22_12, regPage1NextUnit(11)=>
      regFileMap_page1Out_22_11, regPage1NextUnit(10)=>
      regFileMap_page1Out_22_10, regPage1NextUnit(9)=>
      regFileMap_page1Out_22_9, regPage1NextUnit(8)=>
      regFileMap_page1Out_22_8, regPage1NextUnit(7)=>
      regFileMap_page1Out_22_7, regPage1NextUnit(6)=>
      regFileMap_page1Out_22_6, regPage1NextUnit(5)=>
      regFileMap_page1Out_22_5, regPage1NextUnit(4)=>
      regFileMap_page1Out_22_4, regPage1NextUnit(3)=>
      regFileMap_page1Out_22_3, regPage1NextUnit(2)=>
      regFileMap_page1Out_22_2, regPage1NextUnit(1)=>
      regFileMap_page1Out_22_1, regPage1NextUnit(0)=>
      regFileMap_page1Out_22_0, regPage2NextUnit(15)=>
      regFileMap_page2Out_22_15, regPage2NextUnit(14)=>
      regFileMap_page2Out_22_14, regPage2NextUnit(13)=>
      regFileMap_page2Out_22_13, regPage2NextUnit(12)=>
      regFileMap_page2Out_22_12, regPage2NextUnit(11)=>
      regFileMap_page2Out_22_11, regPage2NextUnit(10)=>
      regFileMap_page2Out_22_10, regPage2NextUnit(9)=>
      regFileMap_page2Out_22_9, regPage2NextUnit(8)=>
      regFileMap_page2Out_22_8, regPage2NextUnit(7)=>
      regFileMap_page2Out_22_7, regPage2NextUnit(6)=>
      regFileMap_page2Out_22_6, regPage2NextUnit(5)=>
      regFileMap_page2Out_22_5, regPage2NextUnit(4)=>
      regFileMap_page2Out_22_4, regPage2NextUnit(3)=>
      regFileMap_page2Out_22_3, regPage2NextUnit(2)=>
      regFileMap_page2Out_22_2, regPage2NextUnit(1)=>
      regFileMap_page2Out_22_1, regPage2NextUnit(0)=>
      regFileMap_page2Out_22_0, clk=>clk, rst=>rst, enableRegPage1=>
      regFileMap_page1Enables_3, enableRegPage2=>regFileMap_page2Enables_3, 
      enableRegFilter=>nx5340, page1ReadBusOrPage2=>shift2To1, 
      page2ReadBusOrPage1=>shift1To2, pageTurn=>pageTurn, outRegPage(15)=>
      currentPage_11_15, outRegPage(14)=>currentPage_11_14, outRegPage(13)=>
      currentPage_11_13, outRegPage(12)=>currentPage_11_12, outRegPage(11)=>
      currentPage_11_11, outRegPage(10)=>currentPage_11_10, outRegPage(9)=>
      currentPage_11_9, outRegPage(8)=>currentPage_11_8, outRegPage(7)=>
      currentPage_11_7, outRegPage(6)=>currentPage_11_6, outRegPage(5)=>
      currentPage_11_5, outRegPage(4)=>currentPage_11_4, outRegPage(3)=>
      currentPage_11_3, outRegPage(2)=>currentPage_11_2, outRegPage(1)=>
      currentPage_11_1, outRegPage(0)=>currentPage_11_0, outputRegPage1(15)
      =>regFileMap_page1Out_17_15, outputRegPage1(14)=>
      regFileMap_page1Out_17_14, outputRegPage1(13)=>
      regFileMap_page1Out_17_13, outputRegPage1(12)=>
      regFileMap_page1Out_17_12, outputRegPage1(11)=>
      regFileMap_page1Out_17_11, outputRegPage1(10)=>
      regFileMap_page1Out_17_10, outputRegPage1(9)=>regFileMap_page1Out_17_9, 
      outputRegPage1(8)=>regFileMap_page1Out_17_8, outputRegPage1(7)=>
      regFileMap_page1Out_17_7, outputRegPage1(6)=>regFileMap_page1Out_17_6, 
      outputRegPage1(5)=>regFileMap_page1Out_17_5, outputRegPage1(4)=>
      regFileMap_page1Out_17_4, outputRegPage1(3)=>regFileMap_page1Out_17_3, 
      outputRegPage1(2)=>regFileMap_page1Out_17_2, outputRegPage1(1)=>
      regFileMap_page1Out_17_1, outputRegPage1(0)=>regFileMap_page1Out_17_0, 
      outputRegPage2(15)=>regFileMap_page2Out_17_15, outputRegPage2(14)=>
      regFileMap_page2Out_17_14, outputRegPage2(13)=>
      regFileMap_page2Out_17_13, outputRegPage2(12)=>
      regFileMap_page2Out_17_12, outputRegPage2(11)=>
      regFileMap_page2Out_17_11, outputRegPage2(10)=>
      regFileMap_page2Out_17_10, outputRegPage2(9)=>regFileMap_page2Out_17_9, 
      outputRegPage2(8)=>regFileMap_page2Out_17_8, outputRegPage2(7)=>
      regFileMap_page2Out_17_7, outputRegPage2(6)=>regFileMap_page2Out_17_6, 
      outputRegPage2(5)=>regFileMap_page2Out_17_5, outputRegPage2(4)=>
      regFileMap_page2Out_17_4, outputRegPage2(3)=>regFileMap_page2Out_17_3, 
      outputRegPage2(2)=>regFileMap_page2Out_17_2, outputRegPage2(1)=>
      regFileMap_page2Out_17_1, outputRegPage2(0)=>regFileMap_page2Out_17_0, 
      outFilter(7)=>filter_11_7, outFilter(6)=>filter_11_6, outFilter(5)=>
      filter_11_5, outFilter(4)=>filter_11_4, outFilter(3)=>filter_11_3, 
      outFilter(2)=>filter_11_2, outFilter(1)=>filter_11_1, outFilter(0)=>
      filter_11_0);
   regFileMap_loop1_3_regRowMap_loop1_3_regUnitMap : RegUnit_8_16_unfolded2
       port map ( filterBus(7)=>filterBus(31), filterBus(6)=>filterBus(30), 
      filterBus(5)=>filterBus(29), filterBus(4)=>filterBus(28), filterBus(3)
      =>filterBus(27), filterBus(2)=>filterBus(26), filterBus(1)=>
      filterBus(25), filterBus(0)=>filterBus(24), windowBus(15)=>
      windowBus(63), windowBus(14)=>windowBus(62), windowBus(13)=>
      windowBus(61), windowBus(12)=>windowBus(60), windowBus(11)=>
      windowBus(59), windowBus(10)=>windowBus(58), windowBus(9)=>
      windowBus(57), windowBus(8)=>windowBus(56), windowBus(7)=>
      windowBus(55), windowBus(6)=>windowBus(54), windowBus(5)=>
      windowBus(53), windowBus(4)=>windowBus(52), windowBus(3)=>
      windowBus(51), windowBus(2)=>windowBus(50), windowBus(1)=>
      windowBus(49), windowBus(0)=>windowBus(48), regPage1NextUnit(15)=>
      regFileMap_page1Out_23_15, regPage1NextUnit(14)=>
      regFileMap_page1Out_23_14, regPage1NextUnit(13)=>
      regFileMap_page1Out_23_13, regPage1NextUnit(12)=>
      regFileMap_page1Out_23_12, regPage1NextUnit(11)=>
      regFileMap_page1Out_23_11, regPage1NextUnit(10)=>
      regFileMap_page1Out_23_10, regPage1NextUnit(9)=>
      regFileMap_page1Out_23_9, regPage1NextUnit(8)=>
      regFileMap_page1Out_23_8, regPage1NextUnit(7)=>
      regFileMap_page1Out_23_7, regPage1NextUnit(6)=>
      regFileMap_page1Out_23_6, regPage1NextUnit(5)=>
      regFileMap_page1Out_23_5, regPage1NextUnit(4)=>
      regFileMap_page1Out_23_4, regPage1NextUnit(3)=>
      regFileMap_page1Out_23_3, regPage1NextUnit(2)=>
      regFileMap_page1Out_23_2, regPage1NextUnit(1)=>
      regFileMap_page1Out_23_1, regPage1NextUnit(0)=>
      regFileMap_page1Out_23_0, regPage2NextUnit(15)=>
      regFileMap_page2Out_23_15, regPage2NextUnit(14)=>
      regFileMap_page2Out_23_14, regPage2NextUnit(13)=>
      regFileMap_page2Out_23_13, regPage2NextUnit(12)=>
      regFileMap_page2Out_23_12, regPage2NextUnit(11)=>
      regFileMap_page2Out_23_11, regPage2NextUnit(10)=>
      regFileMap_page2Out_23_10, regPage2NextUnit(9)=>
      regFileMap_page2Out_23_9, regPage2NextUnit(8)=>
      regFileMap_page2Out_23_8, regPage2NextUnit(7)=>
      regFileMap_page2Out_23_7, regPage2NextUnit(6)=>
      regFileMap_page2Out_23_6, regPage2NextUnit(5)=>
      regFileMap_page2Out_23_5, regPage2NextUnit(4)=>
      regFileMap_page2Out_23_4, regPage2NextUnit(3)=>
      regFileMap_page2Out_23_3, regPage2NextUnit(2)=>
      regFileMap_page2Out_23_2, regPage2NextUnit(1)=>
      regFileMap_page2Out_23_1, regPage2NextUnit(0)=>
      regFileMap_page2Out_23_0, clk=>clk, rst=>rst, enableRegPage1=>
      regFileMap_page1Enables_3, enableRegPage2=>regFileMap_page2Enables_3, 
      enableRegFilter=>nx5342, page1ReadBusOrPage2=>shift2To1, 
      page2ReadBusOrPage1=>shift1To2, pageTurn=>pageTurn, outRegPage(15)=>
      currentPage_21_15, outRegPage(14)=>currentPage_21_14, outRegPage(13)=>
      currentPage_21_13, outRegPage(12)=>currentPage_21_12, outRegPage(11)=>
      currentPage_21_11, outRegPage(10)=>currentPage_21_10, outRegPage(9)=>
      currentPage_21_9, outRegPage(8)=>currentPage_21_8, outRegPage(7)=>
      currentPage_21_7, outRegPage(6)=>currentPage_21_6, outRegPage(5)=>
      currentPage_21_5, outRegPage(4)=>currentPage_21_4, outRegPage(3)=>
      currentPage_21_3, outRegPage(2)=>currentPage_21_2, outRegPage(1)=>
      currentPage_21_1, outRegPage(0)=>currentPage_21_0, outputRegPage1(15)
      =>regFileMap_page1Out_18_15, outputRegPage1(14)=>
      regFileMap_page1Out_18_14, outputRegPage1(13)=>
      regFileMap_page1Out_18_13, outputRegPage1(12)=>
      regFileMap_page1Out_18_12, outputRegPage1(11)=>
      regFileMap_page1Out_18_11, outputRegPage1(10)=>
      regFileMap_page1Out_18_10, outputRegPage1(9)=>regFileMap_page1Out_18_9, 
      outputRegPage1(8)=>regFileMap_page1Out_18_8, outputRegPage1(7)=>
      regFileMap_page1Out_18_7, outputRegPage1(6)=>regFileMap_page1Out_18_6, 
      outputRegPage1(5)=>regFileMap_page1Out_18_5, outputRegPage1(4)=>
      regFileMap_page1Out_18_4, outputRegPage1(3)=>regFileMap_page1Out_18_3, 
      outputRegPage1(2)=>regFileMap_page1Out_18_2, outputRegPage1(1)=>
      regFileMap_page1Out_18_1, outputRegPage1(0)=>regFileMap_page1Out_18_0, 
      outputRegPage2(15)=>regFileMap_page2Out_18_15, outputRegPage2(14)=>
      regFileMap_page2Out_18_14, outputRegPage2(13)=>
      regFileMap_page2Out_18_13, outputRegPage2(12)=>
      regFileMap_page2Out_18_12, outputRegPage2(11)=>
      regFileMap_page2Out_18_11, outputRegPage2(10)=>
      regFileMap_page2Out_18_10, outputRegPage2(9)=>regFileMap_page2Out_18_9, 
      outputRegPage2(8)=>regFileMap_page2Out_18_8, outputRegPage2(7)=>
      regFileMap_page2Out_18_7, outputRegPage2(6)=>regFileMap_page2Out_18_6, 
      outputRegPage2(5)=>regFileMap_page2Out_18_5, outputRegPage2(4)=>
      regFileMap_page2Out_18_4, outputRegPage2(3)=>regFileMap_page2Out_18_3, 
      outputRegPage2(2)=>regFileMap_page2Out_18_2, outputRegPage2(1)=>
      regFileMap_page2Out_18_1, outputRegPage2(0)=>regFileMap_page2Out_18_0, 
      outFilter(7)=>filter_21_7, outFilter(6)=>filter_21_6, outFilter(5)=>
      filter_21_5, outFilter(4)=>filter_21_4, outFilter(3)=>filter_21_3, 
      outFilter(2)=>filter_21_2, outFilter(1)=>filter_21_1, outFilter(0)=>
      filter_21_0);
   regFileMap_loop1_3_regRowMap_loop1_4_regUnitMap : RegUnit_8_16_unfolded2
       port map ( filterBus(7)=>filterBus(39), filterBus(6)=>filterBus(38), 
      filterBus(5)=>filterBus(37), filterBus(4)=>filterBus(36), filterBus(3)
      =>filterBus(35), filterBus(2)=>filterBus(34), filterBus(1)=>
      filterBus(33), filterBus(0)=>filterBus(32), windowBus(15)=>
      windowBus(79), windowBus(14)=>windowBus(78), windowBus(13)=>
      windowBus(77), windowBus(12)=>windowBus(76), windowBus(11)=>
      windowBus(75), windowBus(10)=>windowBus(74), windowBus(9)=>
      windowBus(73), windowBus(8)=>windowBus(72), windowBus(7)=>
      windowBus(71), windowBus(6)=>windowBus(70), windowBus(5)=>
      windowBus(69), windowBus(4)=>windowBus(68), windowBus(3)=>
      windowBus(67), windowBus(2)=>windowBus(66), windowBus(1)=>
      windowBus(65), windowBus(0)=>windowBus(64), regPage1NextUnit(15)=>
      regFileMap_page1Out_24_15, regPage1NextUnit(14)=>
      regFileMap_page1Out_24_14, regPage1NextUnit(13)=>
      regFileMap_page1Out_24_13, regPage1NextUnit(12)=>
      regFileMap_page1Out_24_12, regPage1NextUnit(11)=>
      regFileMap_page1Out_24_11, regPage1NextUnit(10)=>
      regFileMap_page1Out_24_10, regPage1NextUnit(9)=>
      regFileMap_page1Out_24_9, regPage1NextUnit(8)=>
      regFileMap_page1Out_24_8, regPage1NextUnit(7)=>
      regFileMap_page1Out_24_7, regPage1NextUnit(6)=>
      regFileMap_page1Out_24_6, regPage1NextUnit(5)=>
      regFileMap_page1Out_24_5, regPage1NextUnit(4)=>
      regFileMap_page1Out_24_4, regPage1NextUnit(3)=>
      regFileMap_page1Out_24_3, regPage1NextUnit(2)=>
      regFileMap_page1Out_24_2, regPage1NextUnit(1)=>
      regFileMap_page1Out_24_1, regPage1NextUnit(0)=>
      regFileMap_page1Out_24_0, regPage2NextUnit(15)=>
      regFileMap_page2Out_24_15, regPage2NextUnit(14)=>
      regFileMap_page2Out_24_14, regPage2NextUnit(13)=>
      regFileMap_page2Out_24_13, regPage2NextUnit(12)=>
      regFileMap_page2Out_24_12, regPage2NextUnit(11)=>
      regFileMap_page2Out_24_11, regPage2NextUnit(10)=>
      regFileMap_page2Out_24_10, regPage2NextUnit(9)=>
      regFileMap_page2Out_24_9, regPage2NextUnit(8)=>
      regFileMap_page2Out_24_8, regPage2NextUnit(7)=>
      regFileMap_page2Out_24_7, regPage2NextUnit(6)=>
      regFileMap_page2Out_24_6, regPage2NextUnit(5)=>
      regFileMap_page2Out_24_5, regPage2NextUnit(4)=>
      regFileMap_page2Out_24_4, regPage2NextUnit(3)=>
      regFileMap_page2Out_24_3, regPage2NextUnit(2)=>
      regFileMap_page2Out_24_2, regPage2NextUnit(1)=>
      regFileMap_page2Out_24_1, regPage2NextUnit(0)=>
      regFileMap_page2Out_24_0, clk=>clk, rst=>rst, enableRegPage1=>
      regFileMap_page1Enables_3, enableRegPage2=>regFileMap_page2Enables_3, 
      enableRegFilter=>nx5342, page1ReadBusOrPage2=>shift2To1, 
      page2ReadBusOrPage1=>shift1To2, pageTurn=>pageTurn, outRegPage(15)=>
      currentPage_22_15, outRegPage(14)=>currentPage_22_14, outRegPage(13)=>
      currentPage_22_13, outRegPage(12)=>currentPage_22_12, outRegPage(11)=>
      currentPage_22_11, outRegPage(10)=>currentPage_22_10, outRegPage(9)=>
      currentPage_22_9, outRegPage(8)=>currentPage_22_8, outRegPage(7)=>
      currentPage_22_7, outRegPage(6)=>currentPage_22_6, outRegPage(5)=>
      currentPage_22_5, outRegPage(4)=>currentPage_22_4, outRegPage(3)=>
      currentPage_22_3, outRegPage(2)=>currentPage_22_2, outRegPage(1)=>
      currentPage_22_1, outRegPage(0)=>currentPage_22_0, outputRegPage1(15)
      =>regFileMap_page1Out_19_15, outputRegPage1(14)=>
      regFileMap_page1Out_19_14, outputRegPage1(13)=>
      regFileMap_page1Out_19_13, outputRegPage1(12)=>
      regFileMap_page1Out_19_12, outputRegPage1(11)=>
      regFileMap_page1Out_19_11, outputRegPage1(10)=>
      regFileMap_page1Out_19_10, outputRegPage1(9)=>regFileMap_page1Out_19_9, 
      outputRegPage1(8)=>regFileMap_page1Out_19_8, outputRegPage1(7)=>
      regFileMap_page1Out_19_7, outputRegPage1(6)=>regFileMap_page1Out_19_6, 
      outputRegPage1(5)=>regFileMap_page1Out_19_5, outputRegPage1(4)=>
      regFileMap_page1Out_19_4, outputRegPage1(3)=>regFileMap_page1Out_19_3, 
      outputRegPage1(2)=>regFileMap_page1Out_19_2, outputRegPage1(1)=>
      regFileMap_page1Out_19_1, outputRegPage1(0)=>regFileMap_page1Out_19_0, 
      outputRegPage2(15)=>regFileMap_page2Out_19_15, outputRegPage2(14)=>
      regFileMap_page2Out_19_14, outputRegPage2(13)=>
      regFileMap_page2Out_19_13, outputRegPage2(12)=>
      regFileMap_page2Out_19_12, outputRegPage2(11)=>
      regFileMap_page2Out_19_11, outputRegPage2(10)=>
      regFileMap_page2Out_19_10, outputRegPage2(9)=>regFileMap_page2Out_19_9, 
      outputRegPage2(8)=>regFileMap_page2Out_19_8, outputRegPage2(7)=>
      regFileMap_page2Out_19_7, outputRegPage2(6)=>regFileMap_page2Out_19_6, 
      outputRegPage2(5)=>regFileMap_page2Out_19_5, outputRegPage2(4)=>
      regFileMap_page2Out_19_4, outputRegPage2(3)=>regFileMap_page2Out_19_3, 
      outputRegPage2(2)=>regFileMap_page2Out_19_2, outputRegPage2(1)=>
      regFileMap_page2Out_19_1, outputRegPage2(0)=>regFileMap_page2Out_19_0, 
      outFilter(7)=>filter_22_7, outFilter(6)=>filter_22_6, outFilter(5)=>
      filter_22_5, outFilter(4)=>filter_22_4, outFilter(3)=>filter_22_3, 
      outFilter(2)=>filter_22_2, outFilter(1)=>filter_22_1, outFilter(0)=>
      filter_22_0);
   regFileMap_loop1_4_regRowMap_loop1_0_regUnitMap : RegUnit_8_16_unfolded3
       port map ( filterBus(7)=>filterBus(7), filterBus(6)=>filterBus(6), 
      filterBus(5)=>filterBus(5), filterBus(4)=>filterBus(4), filterBus(3)=>
      filterBus(3), filterBus(2)=>filterBus(2), filterBus(1)=>filterBus(1), 
      filterBus(0)=>filterBus(0), windowBus(15)=>windowBus(15), 
      windowBus(14)=>windowBus(14), windowBus(13)=>windowBus(13), 
      windowBus(12)=>windowBus(12), windowBus(11)=>windowBus(11), 
      windowBus(10)=>windowBus(10), windowBus(9)=>windowBus(9), windowBus(8)
      =>windowBus(8), windowBus(7)=>windowBus(7), windowBus(6)=>windowBus(6), 
      windowBus(5)=>windowBus(5), windowBus(4)=>windowBus(4), windowBus(3)=>
      windowBus(3), windowBus(2)=>windowBus(2), windowBus(1)=>windowBus(1), 
      windowBus(0)=>windowBus(0), regPage1NextUnit(15)=>outShifter_15, 
      regPage1NextUnit(14)=>outShifter_15, regPage1NextUnit(13)=>
      outShifter_15, regPage1NextUnit(12)=>outShifter_15, 
      regPage1NextUnit(11)=>outShifter_15, regPage1NextUnit(10)=>
      outShifter_15, regPage1NextUnit(9)=>outShifter_15, regPage1NextUnit(8)
      =>outShifter_15, regPage1NextUnit(7)=>outShifter_15, 
      regPage1NextUnit(6)=>outShifter_15, regPage1NextUnit(5)=>outShifter_15, 
      regPage1NextUnit(4)=>outShifter_15, regPage1NextUnit(3)=>outShifter_15, 
      regPage1NextUnit(2)=>outShifter_15, regPage1NextUnit(1)=>outShifter_15, 
      regPage1NextUnit(0)=>outShifter_15, regPage2NextUnit(15)=>
      outShifter_15, regPage2NextUnit(14)=>outShifter_15, 
      regPage2NextUnit(13)=>outShifter_15, regPage2NextUnit(12)=>
      outShifter_15, regPage2NextUnit(11)=>outShifter_15, 
      regPage2NextUnit(10)=>outShifter_15, regPage2NextUnit(9)=>
      outShifter_15, regPage2NextUnit(8)=>outShifter_15, regPage2NextUnit(7)
      =>outShifter_15, regPage2NextUnit(6)=>outShifter_15, 
      regPage2NextUnit(5)=>outShifter_15, regPage2NextUnit(4)=>outShifter_15, 
      regPage2NextUnit(3)=>outShifter_15, regPage2NextUnit(2)=>outShifter_15, 
      regPage2NextUnit(1)=>outShifter_15, regPage2NextUnit(0)=>outShifter_15, 
      clk=>clk, rst=>rst, enableRegPage1=>regFileMap_page1Enables_4, 
      enableRegPage2=>regFileMap_page2Enables_4, enableRegFilter=>nx5344, 
      page1ReadBusOrPage2=>shift2To1, page2ReadBusOrPage1=>shift1To2, 
      pageTurn=>pageTurn, outRegPage(15)=>currentPage_12_15, outRegPage(14)
      =>currentPage_12_14, outRegPage(13)=>currentPage_12_13, outRegPage(12)
      =>currentPage_12_12, outRegPage(11)=>currentPage_12_11, outRegPage(10)
      =>currentPage_12_10, outRegPage(9)=>currentPage_12_9, outRegPage(8)=>
      currentPage_12_8, outRegPage(7)=>currentPage_12_7, outRegPage(6)=>
      currentPage_12_6, outRegPage(5)=>currentPage_12_5, outRegPage(4)=>
      currentPage_12_4, outRegPage(3)=>currentPage_12_3, outRegPage(2)=>
      currentPage_12_2, outRegPage(1)=>currentPage_12_1, outRegPage(0)=>
      currentPage_12_0, outputRegPage1(15)=>regFileMap_page1Out_20_15, 
      outputRegPage1(14)=>regFileMap_page1Out_20_14, outputRegPage1(13)=>
      regFileMap_page1Out_20_13, outputRegPage1(12)=>
      regFileMap_page1Out_20_12, outputRegPage1(11)=>
      regFileMap_page1Out_20_11, outputRegPage1(10)=>
      regFileMap_page1Out_20_10, outputRegPage1(9)=>regFileMap_page1Out_20_9, 
      outputRegPage1(8)=>regFileMap_page1Out_20_8, outputRegPage1(7)=>
      regFileMap_page1Out_20_7, outputRegPage1(6)=>regFileMap_page1Out_20_6, 
      outputRegPage1(5)=>regFileMap_page1Out_20_5, outputRegPage1(4)=>
      regFileMap_page1Out_20_4, outputRegPage1(3)=>regFileMap_page1Out_20_3, 
      outputRegPage1(2)=>regFileMap_page1Out_20_2, outputRegPage1(1)=>
      regFileMap_page1Out_20_1, outputRegPage1(0)=>regFileMap_page1Out_20_0, 
      outputRegPage2(15)=>regFileMap_page2Out_20_15, outputRegPage2(14)=>
      regFileMap_page2Out_20_14, outputRegPage2(13)=>
      regFileMap_page2Out_20_13, outputRegPage2(12)=>
      regFileMap_page2Out_20_12, outputRegPage2(11)=>
      regFileMap_page2Out_20_11, outputRegPage2(10)=>
      regFileMap_page2Out_20_10, outputRegPage2(9)=>regFileMap_page2Out_20_9, 
      outputRegPage2(8)=>regFileMap_page2Out_20_8, outputRegPage2(7)=>
      regFileMap_page2Out_20_7, outputRegPage2(6)=>regFileMap_page2Out_20_6, 
      outputRegPage2(5)=>regFileMap_page2Out_20_5, outputRegPage2(4)=>
      regFileMap_page2Out_20_4, outputRegPage2(3)=>regFileMap_page2Out_20_3, 
      outputRegPage2(2)=>regFileMap_page2Out_20_2, outputRegPage2(1)=>
      regFileMap_page2Out_20_1, outputRegPage2(0)=>regFileMap_page2Out_20_0, 
      outFilter(7)=>filter_12_7, outFilter(6)=>filter_12_6, outFilter(5)=>
      filter_12_5, outFilter(4)=>filter_12_4, outFilter(3)=>filter_12_3, 
      outFilter(2)=>filter_12_2, outFilter(1)=>filter_12_1, outFilter(0)=>
      filter_12_0);
   regFileMap_loop1_4_regRowMap_loop1_1_regUnitMap : RegUnit_8_16_unfolded3
       port map ( filterBus(7)=>filterBus(15), filterBus(6)=>filterBus(14), 
      filterBus(5)=>filterBus(13), filterBus(4)=>filterBus(12), filterBus(3)
      =>filterBus(11), filterBus(2)=>filterBus(10), filterBus(1)=>
      filterBus(9), filterBus(0)=>filterBus(8), windowBus(15)=>windowBus(31), 
      windowBus(14)=>windowBus(30), windowBus(13)=>windowBus(29), 
      windowBus(12)=>windowBus(28), windowBus(11)=>windowBus(27), 
      windowBus(10)=>windowBus(26), windowBus(9)=>windowBus(25), 
      windowBus(8)=>windowBus(24), windowBus(7)=>windowBus(23), windowBus(6)
      =>windowBus(22), windowBus(5)=>windowBus(21), windowBus(4)=>
      windowBus(20), windowBus(3)=>windowBus(19), windowBus(2)=>
      windowBus(18), windowBus(1)=>windowBus(17), windowBus(0)=>
      windowBus(16), regPage1NextUnit(15)=>outShifter_15, 
      regPage1NextUnit(14)=>outShifter_15, regPage1NextUnit(13)=>
      outShifter_15, regPage1NextUnit(12)=>outShifter_15, 
      regPage1NextUnit(11)=>outShifter_15, regPage1NextUnit(10)=>
      outShifter_15, regPage1NextUnit(9)=>outShifter_15, regPage1NextUnit(8)
      =>outShifter_15, regPage1NextUnit(7)=>outShifter_15, 
      regPage1NextUnit(6)=>outShifter_15, regPage1NextUnit(5)=>outShifter_15, 
      regPage1NextUnit(4)=>outShifter_15, regPage1NextUnit(3)=>outShifter_15, 
      regPage1NextUnit(2)=>outShifter_15, regPage1NextUnit(1)=>outShifter_15, 
      regPage1NextUnit(0)=>outShifter_15, regPage2NextUnit(15)=>
      outShifter_15, regPage2NextUnit(14)=>outShifter_15, 
      regPage2NextUnit(13)=>outShifter_15, regPage2NextUnit(12)=>
      outShifter_15, regPage2NextUnit(11)=>outShifter_15, 
      regPage2NextUnit(10)=>outShifter_15, regPage2NextUnit(9)=>
      outShifter_15, regPage2NextUnit(8)=>outShifter_15, regPage2NextUnit(7)
      =>outShifter_15, regPage2NextUnit(6)=>outShifter_15, 
      regPage2NextUnit(5)=>outShifter_15, regPage2NextUnit(4)=>outShifter_15, 
      regPage2NextUnit(3)=>outShifter_15, regPage2NextUnit(2)=>outShifter_15, 
      regPage2NextUnit(1)=>outShifter_15, regPage2NextUnit(0)=>outShifter_15, 
      clk=>clk, rst=>rst, enableRegPage1=>regFileMap_page1Enables_4, 
      enableRegPage2=>regFileMap_page2Enables_4, enableRegFilter=>nx5344, 
      page1ReadBusOrPage2=>shift2To1, page2ReadBusOrPage1=>shift1To2, 
      pageTurn=>pageTurn, outRegPage(15)=>currentPage_13_15, outRegPage(14)
      =>currentPage_13_14, outRegPage(13)=>currentPage_13_13, outRegPage(12)
      =>currentPage_13_12, outRegPage(11)=>currentPage_13_11, outRegPage(10)
      =>currentPage_13_10, outRegPage(9)=>currentPage_13_9, outRegPage(8)=>
      currentPage_13_8, outRegPage(7)=>currentPage_13_7, outRegPage(6)=>
      currentPage_13_6, outRegPage(5)=>currentPage_13_5, outRegPage(4)=>
      currentPage_13_4, outRegPage(3)=>currentPage_13_3, outRegPage(2)=>
      currentPage_13_2, outRegPage(1)=>currentPage_13_1, outRegPage(0)=>
      currentPage_13_0, outputRegPage1(15)=>regFileMap_page1Out_21_15, 
      outputRegPage1(14)=>regFileMap_page1Out_21_14, outputRegPage1(13)=>
      regFileMap_page1Out_21_13, outputRegPage1(12)=>
      regFileMap_page1Out_21_12, outputRegPage1(11)=>
      regFileMap_page1Out_21_11, outputRegPage1(10)=>
      regFileMap_page1Out_21_10, outputRegPage1(9)=>regFileMap_page1Out_21_9, 
      outputRegPage1(8)=>regFileMap_page1Out_21_8, outputRegPage1(7)=>
      regFileMap_page1Out_21_7, outputRegPage1(6)=>regFileMap_page1Out_21_6, 
      outputRegPage1(5)=>regFileMap_page1Out_21_5, outputRegPage1(4)=>
      regFileMap_page1Out_21_4, outputRegPage1(3)=>regFileMap_page1Out_21_3, 
      outputRegPage1(2)=>regFileMap_page1Out_21_2, outputRegPage1(1)=>
      regFileMap_page1Out_21_1, outputRegPage1(0)=>regFileMap_page1Out_21_0, 
      outputRegPage2(15)=>regFileMap_page2Out_21_15, outputRegPage2(14)=>
      regFileMap_page2Out_21_14, outputRegPage2(13)=>
      regFileMap_page2Out_21_13, outputRegPage2(12)=>
      regFileMap_page2Out_21_12, outputRegPage2(11)=>
      regFileMap_page2Out_21_11, outputRegPage2(10)=>
      regFileMap_page2Out_21_10, outputRegPage2(9)=>regFileMap_page2Out_21_9, 
      outputRegPage2(8)=>regFileMap_page2Out_21_8, outputRegPage2(7)=>
      regFileMap_page2Out_21_7, outputRegPage2(6)=>regFileMap_page2Out_21_6, 
      outputRegPage2(5)=>regFileMap_page2Out_21_5, outputRegPage2(4)=>
      regFileMap_page2Out_21_4, outputRegPage2(3)=>regFileMap_page2Out_21_3, 
      outputRegPage2(2)=>regFileMap_page2Out_21_2, outputRegPage2(1)=>
      regFileMap_page2Out_21_1, outputRegPage2(0)=>regFileMap_page2Out_21_0, 
      outFilter(7)=>filter_13_7, outFilter(6)=>filter_13_6, outFilter(5)=>
      filter_13_5, outFilter(4)=>filter_13_4, outFilter(3)=>filter_13_3, 
      outFilter(2)=>filter_13_2, outFilter(1)=>filter_13_1, outFilter(0)=>
      filter_13_0);
   regFileMap_loop1_4_regRowMap_loop1_2_regUnitMap : RegUnit_8_16_unfolded3
       port map ( filterBus(7)=>filterBus(23), filterBus(6)=>filterBus(22), 
      filterBus(5)=>filterBus(21), filterBus(4)=>filterBus(20), filterBus(3)
      =>filterBus(19), filterBus(2)=>filterBus(18), filterBus(1)=>
      filterBus(17), filterBus(0)=>filterBus(16), windowBus(15)=>
      windowBus(47), windowBus(14)=>windowBus(46), windowBus(13)=>
      windowBus(45), windowBus(12)=>windowBus(44), windowBus(11)=>
      windowBus(43), windowBus(10)=>windowBus(42), windowBus(9)=>
      windowBus(41), windowBus(8)=>windowBus(40), windowBus(7)=>
      windowBus(39), windowBus(6)=>windowBus(38), windowBus(5)=>
      windowBus(37), windowBus(4)=>windowBus(36), windowBus(3)=>
      windowBus(35), windowBus(2)=>windowBus(34), windowBus(1)=>
      windowBus(33), windowBus(0)=>windowBus(32), regPage1NextUnit(15)=>
      outShifter_15, regPage1NextUnit(14)=>outShifter_15, 
      regPage1NextUnit(13)=>outShifter_15, regPage1NextUnit(12)=>
      outShifter_15, regPage1NextUnit(11)=>outShifter_15, 
      regPage1NextUnit(10)=>outShifter_15, regPage1NextUnit(9)=>
      outShifter_15, regPage1NextUnit(8)=>outShifter_15, regPage1NextUnit(7)
      =>outShifter_15, regPage1NextUnit(6)=>outShifter_15, 
      regPage1NextUnit(5)=>outShifter_15, regPage1NextUnit(4)=>outShifter_15, 
      regPage1NextUnit(3)=>outShifter_15, regPage1NextUnit(2)=>outShifter_15, 
      regPage1NextUnit(1)=>outShifter_15, regPage1NextUnit(0)=>outShifter_15, 
      regPage2NextUnit(15)=>outShifter_15, regPage2NextUnit(14)=>
      outShifter_15, regPage2NextUnit(13)=>outShifter_15, 
      regPage2NextUnit(12)=>outShifter_15, regPage2NextUnit(11)=>
      outShifter_15, regPage2NextUnit(10)=>outShifter_15, 
      regPage2NextUnit(9)=>outShifter_15, regPage2NextUnit(8)=>outShifter_15, 
      regPage2NextUnit(7)=>outShifter_15, regPage2NextUnit(6)=>outShifter_15, 
      regPage2NextUnit(5)=>outShifter_15, regPage2NextUnit(4)=>outShifter_15, 
      regPage2NextUnit(3)=>outShifter_15, regPage2NextUnit(2)=>outShifter_15, 
      regPage2NextUnit(1)=>outShifter_15, regPage2NextUnit(0)=>outShifter_15, 
      clk=>clk, rst=>rst, enableRegPage1=>regFileMap_page1Enables_4, 
      enableRegPage2=>regFileMap_page2Enables_4, enableRegFilter=>nx5344, 
      page1ReadBusOrPage2=>shift2To1, page2ReadBusOrPage1=>shift1To2, 
      pageTurn=>pageTurn, outRegPage(15)=>currentPage_14_15, outRegPage(14)
      =>currentPage_14_14, outRegPage(13)=>currentPage_14_13, outRegPage(12)
      =>currentPage_14_12, outRegPage(11)=>currentPage_14_11, outRegPage(10)
      =>currentPage_14_10, outRegPage(9)=>currentPage_14_9, outRegPage(8)=>
      currentPage_14_8, outRegPage(7)=>currentPage_14_7, outRegPage(6)=>
      currentPage_14_6, outRegPage(5)=>currentPage_14_5, outRegPage(4)=>
      currentPage_14_4, outRegPage(3)=>currentPage_14_3, outRegPage(2)=>
      currentPage_14_2, outRegPage(1)=>currentPage_14_1, outRegPage(0)=>
      currentPage_14_0, outputRegPage1(15)=>regFileMap_page1Out_22_15, 
      outputRegPage1(14)=>regFileMap_page1Out_22_14, outputRegPage1(13)=>
      regFileMap_page1Out_22_13, outputRegPage1(12)=>
      regFileMap_page1Out_22_12, outputRegPage1(11)=>
      regFileMap_page1Out_22_11, outputRegPage1(10)=>
      regFileMap_page1Out_22_10, outputRegPage1(9)=>regFileMap_page1Out_22_9, 
      outputRegPage1(8)=>regFileMap_page1Out_22_8, outputRegPage1(7)=>
      regFileMap_page1Out_22_7, outputRegPage1(6)=>regFileMap_page1Out_22_6, 
      outputRegPage1(5)=>regFileMap_page1Out_22_5, outputRegPage1(4)=>
      regFileMap_page1Out_22_4, outputRegPage1(3)=>regFileMap_page1Out_22_3, 
      outputRegPage1(2)=>regFileMap_page1Out_22_2, outputRegPage1(1)=>
      regFileMap_page1Out_22_1, outputRegPage1(0)=>regFileMap_page1Out_22_0, 
      outputRegPage2(15)=>regFileMap_page2Out_22_15, outputRegPage2(14)=>
      regFileMap_page2Out_22_14, outputRegPage2(13)=>
      regFileMap_page2Out_22_13, outputRegPage2(12)=>
      regFileMap_page2Out_22_12, outputRegPage2(11)=>
      regFileMap_page2Out_22_11, outputRegPage2(10)=>
      regFileMap_page2Out_22_10, outputRegPage2(9)=>regFileMap_page2Out_22_9, 
      outputRegPage2(8)=>regFileMap_page2Out_22_8, outputRegPage2(7)=>
      regFileMap_page2Out_22_7, outputRegPage2(6)=>regFileMap_page2Out_22_6, 
      outputRegPage2(5)=>regFileMap_page2Out_22_5, outputRegPage2(4)=>
      regFileMap_page2Out_22_4, outputRegPage2(3)=>regFileMap_page2Out_22_3, 
      outputRegPage2(2)=>regFileMap_page2Out_22_2, outputRegPage2(1)=>
      regFileMap_page2Out_22_1, outputRegPage2(0)=>regFileMap_page2Out_22_0, 
      outFilter(7)=>filter_14_7, outFilter(6)=>filter_14_6, outFilter(5)=>
      filter_14_5, outFilter(4)=>filter_14_4, outFilter(3)=>filter_14_3, 
      outFilter(2)=>filter_14_2, outFilter(1)=>filter_14_1, outFilter(0)=>
      filter_14_0);
   regFileMap_loop1_4_regRowMap_loop1_3_regUnitMap : RegUnit_8_16_unfolded3
       port map ( filterBus(7)=>filterBus(31), filterBus(6)=>filterBus(30), 
      filterBus(5)=>filterBus(29), filterBus(4)=>filterBus(28), filterBus(3)
      =>filterBus(27), filterBus(2)=>filterBus(26), filterBus(1)=>
      filterBus(25), filterBus(0)=>filterBus(24), windowBus(15)=>
      windowBus(63), windowBus(14)=>windowBus(62), windowBus(13)=>
      windowBus(61), windowBus(12)=>windowBus(60), windowBus(11)=>
      windowBus(59), windowBus(10)=>windowBus(58), windowBus(9)=>
      windowBus(57), windowBus(8)=>windowBus(56), windowBus(7)=>
      windowBus(55), windowBus(6)=>windowBus(54), windowBus(5)=>
      windowBus(53), windowBus(4)=>windowBus(52), windowBus(3)=>
      windowBus(51), windowBus(2)=>windowBus(50), windowBus(1)=>
      windowBus(49), windowBus(0)=>windowBus(48), regPage1NextUnit(15)=>
      outShifter_15, regPage1NextUnit(14)=>outShifter_15, 
      regPage1NextUnit(13)=>outShifter_15, regPage1NextUnit(12)=>
      outShifter_15, regPage1NextUnit(11)=>outShifter_15, 
      regPage1NextUnit(10)=>outShifter_15, regPage1NextUnit(9)=>
      outShifter_15, regPage1NextUnit(8)=>outShifter_15, regPage1NextUnit(7)
      =>outShifter_15, regPage1NextUnit(6)=>outShifter_15, 
      regPage1NextUnit(5)=>outShifter_15, regPage1NextUnit(4)=>outShifter_15, 
      regPage1NextUnit(3)=>outShifter_15, regPage1NextUnit(2)=>outShifter_15, 
      regPage1NextUnit(1)=>outShifter_15, regPage1NextUnit(0)=>outShifter_15, 
      regPage2NextUnit(15)=>outShifter_15, regPage2NextUnit(14)=>
      outShifter_15, regPage2NextUnit(13)=>outShifter_15, 
      regPage2NextUnit(12)=>outShifter_15, regPage2NextUnit(11)=>
      outShifter_15, regPage2NextUnit(10)=>outShifter_15, 
      regPage2NextUnit(9)=>outShifter_15, regPage2NextUnit(8)=>outShifter_15, 
      regPage2NextUnit(7)=>outShifter_15, regPage2NextUnit(6)=>outShifter_15, 
      regPage2NextUnit(5)=>outShifter_15, regPage2NextUnit(4)=>outShifter_15, 
      regPage2NextUnit(3)=>outShifter_15, regPage2NextUnit(2)=>outShifter_15, 
      regPage2NextUnit(1)=>outShifter_15, regPage2NextUnit(0)=>outShifter_15, 
      clk=>clk, rst=>rst, enableRegPage1=>regFileMap_page1Enables_4, 
      enableRegPage2=>regFileMap_page2Enables_4, enableRegFilter=>nx5346, 
      page1ReadBusOrPage2=>shift2To1, page2ReadBusOrPage1=>shift1To2, 
      pageTurn=>pageTurn, outRegPage(15)=>currentPage_23_15, outRegPage(14)
      =>currentPage_23_14, outRegPage(13)=>currentPage_23_13, outRegPage(12)
      =>currentPage_23_12, outRegPage(11)=>currentPage_23_11, outRegPage(10)
      =>currentPage_23_10, outRegPage(9)=>currentPage_23_9, outRegPage(8)=>
      currentPage_23_8, outRegPage(7)=>currentPage_23_7, outRegPage(6)=>
      currentPage_23_6, outRegPage(5)=>currentPage_23_5, outRegPage(4)=>
      currentPage_23_4, outRegPage(3)=>currentPage_23_3, outRegPage(2)=>
      currentPage_23_2, outRegPage(1)=>currentPage_23_1, outRegPage(0)=>
      currentPage_23_0, outputRegPage1(15)=>regFileMap_page1Out_23_15, 
      outputRegPage1(14)=>regFileMap_page1Out_23_14, outputRegPage1(13)=>
      regFileMap_page1Out_23_13, outputRegPage1(12)=>
      regFileMap_page1Out_23_12, outputRegPage1(11)=>
      regFileMap_page1Out_23_11, outputRegPage1(10)=>
      regFileMap_page1Out_23_10, outputRegPage1(9)=>regFileMap_page1Out_23_9, 
      outputRegPage1(8)=>regFileMap_page1Out_23_8, outputRegPage1(7)=>
      regFileMap_page1Out_23_7, outputRegPage1(6)=>regFileMap_page1Out_23_6, 
      outputRegPage1(5)=>regFileMap_page1Out_23_5, outputRegPage1(4)=>
      regFileMap_page1Out_23_4, outputRegPage1(3)=>regFileMap_page1Out_23_3, 
      outputRegPage1(2)=>regFileMap_page1Out_23_2, outputRegPage1(1)=>
      regFileMap_page1Out_23_1, outputRegPage1(0)=>regFileMap_page1Out_23_0, 
      outputRegPage2(15)=>regFileMap_page2Out_23_15, outputRegPage2(14)=>
      regFileMap_page2Out_23_14, outputRegPage2(13)=>
      regFileMap_page2Out_23_13, outputRegPage2(12)=>
      regFileMap_page2Out_23_12, outputRegPage2(11)=>
      regFileMap_page2Out_23_11, outputRegPage2(10)=>
      regFileMap_page2Out_23_10, outputRegPage2(9)=>regFileMap_page2Out_23_9, 
      outputRegPage2(8)=>regFileMap_page2Out_23_8, outputRegPage2(7)=>
      regFileMap_page2Out_23_7, outputRegPage2(6)=>regFileMap_page2Out_23_6, 
      outputRegPage2(5)=>regFileMap_page2Out_23_5, outputRegPage2(4)=>
      regFileMap_page2Out_23_4, outputRegPage2(3)=>regFileMap_page2Out_23_3, 
      outputRegPage2(2)=>regFileMap_page2Out_23_2, outputRegPage2(1)=>
      regFileMap_page2Out_23_1, outputRegPage2(0)=>regFileMap_page2Out_23_0, 
      outFilter(7)=>filter_23_7, outFilter(6)=>filter_23_6, outFilter(5)=>
      filter_23_5, outFilter(4)=>filter_23_4, outFilter(3)=>filter_23_3, 
      outFilter(2)=>filter_23_2, outFilter(1)=>filter_23_1, outFilter(0)=>
      filter_23_0);
   regFileMap_loop1_4_regRowMap_loop1_4_regUnitMap : RegUnit_8_16_unfolded3
       port map ( filterBus(7)=>filterBus(39), filterBus(6)=>filterBus(38), 
      filterBus(5)=>filterBus(37), filterBus(4)=>filterBus(36), filterBus(3)
      =>filterBus(35), filterBus(2)=>filterBus(34), filterBus(1)=>
      filterBus(33), filterBus(0)=>filterBus(32), windowBus(15)=>
      windowBus(79), windowBus(14)=>windowBus(78), windowBus(13)=>
      windowBus(77), windowBus(12)=>windowBus(76), windowBus(11)=>
      windowBus(75), windowBus(10)=>windowBus(74), windowBus(9)=>
      windowBus(73), windowBus(8)=>windowBus(72), windowBus(7)=>
      windowBus(71), windowBus(6)=>windowBus(70), windowBus(5)=>
      windowBus(69), windowBus(4)=>windowBus(68), windowBus(3)=>
      windowBus(67), windowBus(2)=>windowBus(66), windowBus(1)=>
      windowBus(65), windowBus(0)=>windowBus(64), regPage1NextUnit(15)=>
      outShifter_15, regPage1NextUnit(14)=>outShifter_15, 
      regPage1NextUnit(13)=>outShifter_15, regPage1NextUnit(12)=>
      outShifter_15, regPage1NextUnit(11)=>outShifter_15, 
      regPage1NextUnit(10)=>outShifter_15, regPage1NextUnit(9)=>
      outShifter_15, regPage1NextUnit(8)=>outShifter_15, regPage1NextUnit(7)
      =>outShifter_15, regPage1NextUnit(6)=>outShifter_15, 
      regPage1NextUnit(5)=>outShifter_15, regPage1NextUnit(4)=>outShifter_15, 
      regPage1NextUnit(3)=>outShifter_15, regPage1NextUnit(2)=>outShifter_15, 
      regPage1NextUnit(1)=>outShifter_15, regPage1NextUnit(0)=>outShifter_15, 
      regPage2NextUnit(15)=>outShifter_15, regPage2NextUnit(14)=>
      outShifter_15, regPage2NextUnit(13)=>outShifter_15, 
      regPage2NextUnit(12)=>outShifter_15, regPage2NextUnit(11)=>
      outShifter_15, regPage2NextUnit(10)=>outShifter_15, 
      regPage2NextUnit(9)=>outShifter_15, regPage2NextUnit(8)=>outShifter_15, 
      regPage2NextUnit(7)=>outShifter_15, regPage2NextUnit(6)=>outShifter_15, 
      regPage2NextUnit(5)=>outShifter_15, regPage2NextUnit(4)=>outShifter_15, 
      regPage2NextUnit(3)=>outShifter_15, regPage2NextUnit(2)=>outShifter_15, 
      regPage2NextUnit(1)=>outShifter_15, regPage2NextUnit(0)=>outShifter_15, 
      clk=>clk, rst=>rst, enableRegPage1=>regFileMap_page1Enables_4, 
      enableRegPage2=>regFileMap_page2Enables_4, enableRegFilter=>nx5346, 
      page1ReadBusOrPage2=>shift2To1, page2ReadBusOrPage1=>shift1To2, 
      pageTurn=>pageTurn, outRegPage(15)=>currentPage_24_15, outRegPage(14)
      =>currentPage_24_14, outRegPage(13)=>currentPage_24_13, outRegPage(12)
      =>currentPage_24_12, outRegPage(11)=>currentPage_24_11, outRegPage(10)
      =>currentPage_24_10, outRegPage(9)=>currentPage_24_9, outRegPage(8)=>
      currentPage_24_8, outRegPage(7)=>currentPage_24_7, outRegPage(6)=>
      currentPage_24_6, outRegPage(5)=>currentPage_24_5, outRegPage(4)=>
      currentPage_24_4, outRegPage(3)=>currentPage_24_3, outRegPage(2)=>
      currentPage_24_2, outRegPage(1)=>currentPage_24_1, outRegPage(0)=>
      currentPage_24_0, outputRegPage1(15)=>regFileMap_page1Out_24_15, 
      outputRegPage1(14)=>regFileMap_page1Out_24_14, outputRegPage1(13)=>
      regFileMap_page1Out_24_13, outputRegPage1(12)=>
      regFileMap_page1Out_24_12, outputRegPage1(11)=>
      regFileMap_page1Out_24_11, outputRegPage1(10)=>
      regFileMap_page1Out_24_10, outputRegPage1(9)=>regFileMap_page1Out_24_9, 
      outputRegPage1(8)=>regFileMap_page1Out_24_8, outputRegPage1(7)=>
      regFileMap_page1Out_24_7, outputRegPage1(6)=>regFileMap_page1Out_24_6, 
      outputRegPage1(5)=>regFileMap_page1Out_24_5, outputRegPage1(4)=>
      regFileMap_page1Out_24_4, outputRegPage1(3)=>regFileMap_page1Out_24_3, 
      outputRegPage1(2)=>regFileMap_page1Out_24_2, outputRegPage1(1)=>
      regFileMap_page1Out_24_1, outputRegPage1(0)=>regFileMap_page1Out_24_0, 
      outputRegPage2(15)=>regFileMap_page2Out_24_15, outputRegPage2(14)=>
      regFileMap_page2Out_24_14, outputRegPage2(13)=>
      regFileMap_page2Out_24_13, outputRegPage2(12)=>
      regFileMap_page2Out_24_12, outputRegPage2(11)=>
      regFileMap_page2Out_24_11, outputRegPage2(10)=>
      regFileMap_page2Out_24_10, outputRegPage2(9)=>regFileMap_page2Out_24_9, 
      outputRegPage2(8)=>regFileMap_page2Out_24_8, outputRegPage2(7)=>
      regFileMap_page2Out_24_7, outputRegPage2(6)=>regFileMap_page2Out_24_6, 
      outputRegPage2(5)=>regFileMap_page2Out_24_5, outputRegPage2(4)=>
      regFileMap_page2Out_24_4, outputRegPage2(3)=>regFileMap_page2Out_24_3, 
      outputRegPage2(2)=>regFileMap_page2Out_24_2, outputRegPage2(1)=>
      regFileMap_page2Out_24_1, outputRegPage2(0)=>regFileMap_page2Out_24_0, 
      outFilter(7)=>filter_24_7, outFilter(6)=>filter_24_6, outFilter(5)=>
      filter_24_5, outFilter(4)=>filter_24_4, outFilter(3)=>filter_24_3, 
      outFilter(2)=>filter_24_2, outFilter(1)=>filter_24_1, outFilter(0)=>
      filter_24_0);
   addersMap_sum3FilterMap : NBitAdder_16 port map ( a(15)=>
      addersMap_sum1_15, a(14)=>addersMap_sum1_14, a(13)=>addersMap_sum1_13, 
      a(12)=>addersMap_sum1_12, a(11)=>addersMap_sum1_11, a(10)=>
      addersMap_sum1_10, a(9)=>addersMap_sum1_9, a(8)=>addersMap_sum1_8, 
      a(7)=>addersMap_sum1_7, a(6)=>addersMap_sum1_6, a(5)=>addersMap_sum1_5, 
      a(4)=>addersMap_sum1_4, a(3)=>addersMap_sum1_3, a(2)=>addersMap_sum1_2, 
      a(1)=>addersMap_sum1_1, a(0)=>addersMap_sum1_0, b(15)=>
      addersInputs_8_15, b(14)=>addersInputs_8_14, b(13)=>addersInputs_8_13, 
      b(12)=>addersInputs_8_12, b(11)=>addersInputs_8_11, b(10)=>
      addersInputs_8_10, b(9)=>addersInputs_8_9, b(8)=>addersInputs_8_8, 
      b(7)=>addersInputs_8_7, b(6)=>addersInputs_8_6, b(5)=>addersInputs_8_5, 
      b(4)=>addersInputs_8_4, b(3)=>addersInputs_8_3, b(2)=>addersInputs_8_2, 
      b(1)=>addersInputs_8_1, b(0)=>addersInputs_8_0, carryIn=>outShifter_15, 
      sum(15)=>addersMap_sum3Filter_15, sum(14)=>addersMap_sum3Filter_14, 
      sum(13)=>addersMap_sum3Filter_13, sum(12)=>addersMap_sum3Filter_12, 
      sum(11)=>addersMap_sum3Filter_11, sum(10)=>addersMap_sum3Filter_10, 
      sum(9)=>addersMap_sum3Filter_9, sum(8)=>addersMap_sum3Filter_8, sum(7)
      =>addersMap_sum3Filter_7, sum(6)=>addersMap_sum3Filter_6, sum(5)=>
      addersMap_sum3Filter_5, sum(4)=>addersMap_sum3Filter_4, sum(3)=>
      addersMap_sum3Filter_3, sum(2)=>addersMap_sum3Filter_2, sum(1)=>
      addersMap_sum3Filter_1, sum(0)=>addersMap_sum3Filter_0, carryOut=>
      DANGLING(161));
   addersMap_sumRestMap : NBitAdder_16 port map ( a(15)=>addersMap_sum2_15, 
      a(14)=>addersMap_sum2_14, a(13)=>addersMap_sum2_13, a(12)=>
      addersMap_sum2_12, a(11)=>addersMap_sum2_11, a(10)=>addersMap_sum2_10, 
      a(9)=>addersMap_sum2_9, a(8)=>addersMap_sum2_8, a(7)=>addersMap_sum2_7, 
      a(6)=>addersMap_sum2_6, a(5)=>addersMap_sum2_5, a(4)=>addersMap_sum2_4, 
      a(3)=>addersMap_sum2_3, a(2)=>addersMap_sum2_2, a(1)=>addersMap_sum2_1, 
      a(0)=>addersMap_sum2_0, b(15)=>addersMap_sum3_15, b(14)=>
      addersMap_sum3_14, b(13)=>addersMap_sum3_13, b(12)=>addersMap_sum3_12, 
      b(11)=>addersMap_sum3_11, b(10)=>addersMap_sum3_10, b(9)=>
      addersMap_sum3_9, b(8)=>addersMap_sum3_8, b(7)=>addersMap_sum3_7, b(6)
      =>addersMap_sum3_6, b(5)=>addersMap_sum3_5, b(4)=>addersMap_sum3_4, 
      b(3)=>addersMap_sum3_3, b(2)=>addersMap_sum3_2, b(1)=>addersMap_sum3_1, 
      b(0)=>addersMap_sum3_0, carryIn=>outShifter_15, sum(15)=>
      addersMap_sum4_15, sum(14)=>addersMap_sum4_14, sum(13)=>
      addersMap_sum4_13, sum(12)=>addersMap_sum4_12, sum(11)=>
      addersMap_sum4_11, sum(10)=>addersMap_sum4_10, sum(9)=>
      addersMap_sum4_9, sum(8)=>addersMap_sum4_8, sum(7)=>addersMap_sum4_7, 
      sum(6)=>addersMap_sum4_6, sum(5)=>addersMap_sum4_5, sum(4)=>
      addersMap_sum4_4, sum(3)=>addersMap_sum4_3, sum(2)=>addersMap_sum4_2, 
      sum(1)=>addersMap_sum4_1, sum(0)=>addersMap_sum4_0, carryOut=>DANGLING
      (162));
   addersMap_sumFinalMap : NBitAdder_16 port map ( a(15)=>
      addersMap_sum3Filter_15, a(14)=>addersMap_sum3Filter_14, a(13)=>
      addersMap_sum3Filter_13, a(12)=>addersMap_sum3Filter_12, a(11)=>
      addersMap_sum3Filter_11, a(10)=>addersMap_sum3Filter_10, a(9)=>
      addersMap_sum3Filter_9, a(8)=>addersMap_sum3Filter_8, a(7)=>
      addersMap_sum3Filter_7, a(6)=>addersMap_sum3Filter_6, a(5)=>
      addersMap_sum3Filter_5, a(4)=>addersMap_sum3Filter_4, a(3)=>
      addersMap_sum3Filter_3, a(2)=>addersMap_sum3Filter_2, a(1)=>
      addersMap_sum3Filter_1, a(0)=>addersMap_sum3Filter_0, b(15)=>
      addersMap_sum4_15, b(14)=>addersMap_sum4_14, b(13)=>addersMap_sum4_13, 
      b(12)=>addersMap_sum4_12, b(11)=>addersMap_sum4_11, b(10)=>
      addersMap_sum4_10, b(9)=>addersMap_sum4_9, b(8)=>addersMap_sum4_8, 
      b(7)=>addersMap_sum4_7, b(6)=>addersMap_sum4_6, b(5)=>addersMap_sum4_5, 
      b(4)=>addersMap_sum4_4, b(3)=>addersMap_sum4_3, b(2)=>addersMap_sum4_2, 
      b(1)=>addersMap_sum4_1, b(0)=>addersMap_sum4_0, carryIn=>outShifter_15, 
      sum(15)=>addersMap_totalSum_15, sum(14)=>addersMap_totalSum_14, 
      sum(13)=>addersMap_totalSum_13, sum(12)=>addersMap_totalSum_12, 
      sum(11)=>addersMap_totalSum_11, sum(10)=>addersMap_totalSum_10, sum(9)
      =>addersMap_totalSum_9, sum(8)=>addersMap_totalSum_8, sum(7)=>
      addersMap_totalSum_7, sum(6)=>addersMap_totalSum_6, sum(5)=>
      addersMap_totalSum_5, sum(4)=>addersMap_totalSum_4, sum(3)=>
      addersMap_totalSum_3, sum(2)=>addersMap_totalSum_2, sum(1)=>
      addersMap_totalSum_1, sum(0)=>addersMap_totalSum_0, carryOut=>DANGLING
      (163));
   addersMap_sum1Map_sumFinalMap_dup_0 : NBitAdder_16 port map ( a(15)=>
      addersMap_sum1Map_sum1_15_dup_0, a(14)=>
      addersMap_sum1Map_sum1_14_dup_0, a(13)=>
      addersMap_sum1Map_sum1_13_dup_0, a(12)=>
      addersMap_sum1Map_sum1_12_dup_0, a(11)=>
      addersMap_sum1Map_sum1_11_dup_0, a(10)=>
      addersMap_sum1Map_sum1_10_dup_0, a(9)=>addersMap_sum1Map_sum1_9_dup_0, 
      a(8)=>addersMap_sum1Map_sum1_8_dup_0, a(7)=>
      addersMap_sum1Map_sum1_7_dup_0, a(6)=>addersMap_sum1Map_sum1_6_dup_0, 
      a(5)=>addersMap_sum1Map_sum1_5_dup_0, a(4)=>
      addersMap_sum1Map_sum1_4_dup_0, a(3)=>addersMap_sum1Map_sum1_3_dup_0, 
      a(2)=>addersMap_sum1Map_sum1_2_dup_0, a(1)=>
      addersMap_sum1Map_sum1_1_dup_0, a(0)=>addersMap_sum1Map_sum1_0_dup_0, 
      b(15)=>addersMap_sum1Map_sum2_15_dup_0, b(14)=>
      addersMap_sum1Map_sum2_14_dup_0, b(13)=>
      addersMap_sum1Map_sum2_13_dup_0, b(12)=>
      addersMap_sum1Map_sum2_12_dup_0, b(11)=>
      addersMap_sum1Map_sum2_11_dup_0, b(10)=>
      addersMap_sum1Map_sum2_10_dup_0, b(9)=>addersMap_sum1Map_sum2_9_dup_0, 
      b(8)=>addersMap_sum1Map_sum2_8_dup_0, b(7)=>
      addersMap_sum1Map_sum2_7_dup_0, b(6)=>addersMap_sum1Map_sum2_6_dup_0, 
      b(5)=>addersMap_sum1Map_sum2_5_dup_0, b(4)=>
      addersMap_sum1Map_sum2_4_dup_0, b(3)=>addersMap_sum1Map_sum2_3_dup_0, 
      b(2)=>addersMap_sum1Map_sum2_2_dup_0, b(1)=>
      addersMap_sum1Map_sum2_1_dup_0, b(0)=>addersMap_sum1Map_sum2_0_dup_0, 
      carryIn=>outShifter_15, sum(15)=>addersMap_sum1_15, sum(14)=>
      addersMap_sum1_14, sum(13)=>addersMap_sum1_13, sum(12)=>
      addersMap_sum1_12, sum(11)=>addersMap_sum1_11, sum(10)=>
      addersMap_sum1_10, sum(9)=>addersMap_sum1_9, sum(8)=>addersMap_sum1_8, 
      sum(7)=>addersMap_sum1_7, sum(6)=>addersMap_sum1_6, sum(5)=>
      addersMap_sum1_5, sum(4)=>addersMap_sum1_4, sum(3)=>addersMap_sum1_3, 
      sum(2)=>addersMap_sum1_2, sum(1)=>addersMap_sum1_1, sum(0)=>
      addersMap_sum1_0, carryOut=>DANGLING(164));
   addersMap_sum1Map_sum1Map_sum1Map : NBitAdder_16 port map ( a(15)=>
      addersInputs_0_15, a(14)=>addersInputs_0_14, a(13)=>addersInputs_0_13, 
      a(12)=>addersInputs_0_12, a(11)=>addersInputs_0_11, a(10)=>
      addersInputs_0_10, a(9)=>addersInputs_0_9, a(8)=>addersInputs_0_8, 
      a(7)=>addersInputs_0_7, a(6)=>addersInputs_0_6, a(5)=>addersInputs_0_5, 
      a(4)=>addersInputs_0_4, a(3)=>addersInputs_0_3, a(2)=>addersInputs_0_2, 
      a(1)=>addersInputs_0_1, a(0)=>addersInputs_0_0, b(15)=>
      addersInputs_1_15, b(14)=>addersInputs_1_14, b(13)=>addersInputs_1_13, 
      b(12)=>addersInputs_1_12, b(11)=>addersInputs_1_11, b(10)=>
      addersInputs_1_10, b(9)=>addersInputs_1_9, b(8)=>addersInputs_1_8, 
      b(7)=>addersInputs_1_7, b(6)=>addersInputs_1_6, b(5)=>addersInputs_1_5, 
      b(4)=>addersInputs_1_4, b(3)=>addersInputs_1_3, b(2)=>addersInputs_1_2, 
      b(1)=>addersInputs_1_1, b(0)=>addersInputs_1_0, carryIn=>outShifter_15, 
      sum(15)=>addersMap_sum1Map_sum1Map_sum1_15, sum(14)=>
      addersMap_sum1Map_sum1Map_sum1_14, sum(13)=>
      addersMap_sum1Map_sum1Map_sum1_13, sum(12)=>
      addersMap_sum1Map_sum1Map_sum1_12, sum(11)=>
      addersMap_sum1Map_sum1Map_sum1_11, sum(10)=>
      addersMap_sum1Map_sum1Map_sum1_10, sum(9)=>
      addersMap_sum1Map_sum1Map_sum1_9, sum(8)=>
      addersMap_sum1Map_sum1Map_sum1_8, sum(7)=>
      addersMap_sum1Map_sum1Map_sum1_7, sum(6)=>
      addersMap_sum1Map_sum1Map_sum1_6, sum(5)=>
      addersMap_sum1Map_sum1Map_sum1_5, sum(4)=>
      addersMap_sum1Map_sum1Map_sum1_4, sum(3)=>
      addersMap_sum1Map_sum1Map_sum1_3, sum(2)=>
      addersMap_sum1Map_sum1Map_sum1_2, sum(1)=>
      addersMap_sum1Map_sum1Map_sum1_1, sum(0)=>
      addersMap_sum1Map_sum1Map_sum1_0, carryOut=>DANGLING(165));
   addersMap_sum1Map_sum1Map_sum2Map : NBitAdder_16 port map ( a(15)=>
      addersInputs_2_15, a(14)=>addersInputs_2_14, a(13)=>addersInputs_2_13, 
      a(12)=>addersInputs_2_12, a(11)=>addersInputs_2_11, a(10)=>
      addersInputs_2_10, a(9)=>addersInputs_2_9, a(8)=>addersInputs_2_8, 
      a(7)=>addersInputs_2_7, a(6)=>addersInputs_2_6, a(5)=>addersInputs_2_5, 
      a(4)=>addersInputs_2_4, a(3)=>addersInputs_2_3, a(2)=>addersInputs_2_2, 
      a(1)=>addersInputs_2_1, a(0)=>addersInputs_2_0, b(15)=>
      addersInputs_3_15, b(14)=>addersInputs_3_14, b(13)=>addersInputs_3_13, 
      b(12)=>addersInputs_3_12, b(11)=>addersInputs_3_11, b(10)=>
      addersInputs_3_10, b(9)=>addersInputs_3_9, b(8)=>addersInputs_3_8, 
      b(7)=>addersInputs_3_7, b(6)=>addersInputs_3_6, b(5)=>addersInputs_3_5, 
      b(4)=>addersInputs_3_4, b(3)=>addersInputs_3_3, b(2)=>addersInputs_3_2, 
      b(1)=>addersInputs_3_1, b(0)=>addersInputs_3_0, carryIn=>outShifter_15, 
      sum(15)=>addersMap_sum1Map_sum1Map_sum2_15, sum(14)=>
      addersMap_sum1Map_sum1Map_sum2_14, sum(13)=>
      addersMap_sum1Map_sum1Map_sum2_13, sum(12)=>
      addersMap_sum1Map_sum1Map_sum2_12, sum(11)=>
      addersMap_sum1Map_sum1Map_sum2_11, sum(10)=>
      addersMap_sum1Map_sum1Map_sum2_10, sum(9)=>
      addersMap_sum1Map_sum1Map_sum2_9, sum(8)=>
      addersMap_sum1Map_sum1Map_sum2_8, sum(7)=>
      addersMap_sum1Map_sum1Map_sum2_7, sum(6)=>
      addersMap_sum1Map_sum1Map_sum2_6, sum(5)=>
      addersMap_sum1Map_sum1Map_sum2_5, sum(4)=>
      addersMap_sum1Map_sum1Map_sum2_4, sum(3)=>
      addersMap_sum1Map_sum1Map_sum2_3, sum(2)=>
      addersMap_sum1Map_sum1Map_sum2_2, sum(1)=>
      addersMap_sum1Map_sum1Map_sum2_1, sum(0)=>
      addersMap_sum1Map_sum1Map_sum2_0, carryOut=>DANGLING(166));
   addersMap_sum1Map_sum1Map_sumFinalMap : NBitAdder_16 port map ( a(15)=>
      addersMap_sum1Map_sum1Map_sum1_15, a(14)=>
      addersMap_sum1Map_sum1Map_sum1_14, a(13)=>
      addersMap_sum1Map_sum1Map_sum1_13, a(12)=>
      addersMap_sum1Map_sum1Map_sum1_12, a(11)=>
      addersMap_sum1Map_sum1Map_sum1_11, a(10)=>
      addersMap_sum1Map_sum1Map_sum1_10, a(9)=>
      addersMap_sum1Map_sum1Map_sum1_9, a(8)=>
      addersMap_sum1Map_sum1Map_sum1_8, a(7)=>
      addersMap_sum1Map_sum1Map_sum1_7, a(6)=>
      addersMap_sum1Map_sum1Map_sum1_6, a(5)=>
      addersMap_sum1Map_sum1Map_sum1_5, a(4)=>
      addersMap_sum1Map_sum1Map_sum1_4, a(3)=>
      addersMap_sum1Map_sum1Map_sum1_3, a(2)=>
      addersMap_sum1Map_sum1Map_sum1_2, a(1)=>
      addersMap_sum1Map_sum1Map_sum1_1, a(0)=>
      addersMap_sum1Map_sum1Map_sum1_0, b(15)=>
      addersMap_sum1Map_sum1Map_sum2_15, b(14)=>
      addersMap_sum1Map_sum1Map_sum2_14, b(13)=>
      addersMap_sum1Map_sum1Map_sum2_13, b(12)=>
      addersMap_sum1Map_sum1Map_sum2_12, b(11)=>
      addersMap_sum1Map_sum1Map_sum2_11, b(10)=>
      addersMap_sum1Map_sum1Map_sum2_10, b(9)=>
      addersMap_sum1Map_sum1Map_sum2_9, b(8)=>
      addersMap_sum1Map_sum1Map_sum2_8, b(7)=>
      addersMap_sum1Map_sum1Map_sum2_7, b(6)=>
      addersMap_sum1Map_sum1Map_sum2_6, b(5)=>
      addersMap_sum1Map_sum1Map_sum2_5, b(4)=>
      addersMap_sum1Map_sum1Map_sum2_4, b(3)=>
      addersMap_sum1Map_sum1Map_sum2_3, b(2)=>
      addersMap_sum1Map_sum1Map_sum2_2, b(1)=>
      addersMap_sum1Map_sum1Map_sum2_1, b(0)=>
      addersMap_sum1Map_sum1Map_sum2_0, carryIn=>outShifter_15, sum(15)=>
      addersMap_sum1Map_sum1_15_dup_0, sum(14)=>
      addersMap_sum1Map_sum1_14_dup_0, sum(13)=>
      addersMap_sum1Map_sum1_13_dup_0, sum(12)=>
      addersMap_sum1Map_sum1_12_dup_0, sum(11)=>
      addersMap_sum1Map_sum1_11_dup_0, sum(10)=>
      addersMap_sum1Map_sum1_10_dup_0, sum(9)=>
      addersMap_sum1Map_sum1_9_dup_0, sum(8)=>addersMap_sum1Map_sum1_8_dup_0, 
      sum(7)=>addersMap_sum1Map_sum1_7_dup_0, sum(6)=>
      addersMap_sum1Map_sum1_6_dup_0, sum(5)=>addersMap_sum1Map_sum1_5_dup_0, 
      sum(4)=>addersMap_sum1Map_sum1_4_dup_0, sum(3)=>
      addersMap_sum1Map_sum1_3_dup_0, sum(2)=>addersMap_sum1Map_sum1_2_dup_0, 
      sum(1)=>addersMap_sum1Map_sum1_1_dup_0, sum(0)=>
      addersMap_sum1Map_sum1_0_dup_0, carryOut=>DANGLING(167));
   addersMap_sum1Map_sum2Map_sum1Map : NBitAdder_16 port map ( a(15)=>
      addersInputs_4_15, a(14)=>addersInputs_4_14, a(13)=>addersInputs_4_13, 
      a(12)=>addersInputs_4_12, a(11)=>addersInputs_4_11, a(10)=>
      addersInputs_4_10, a(9)=>addersInputs_4_9, a(8)=>addersInputs_4_8, 
      a(7)=>addersInputs_4_7, a(6)=>addersInputs_4_6, a(5)=>addersInputs_4_5, 
      a(4)=>addersInputs_4_4, a(3)=>addersInputs_4_3, a(2)=>addersInputs_4_2, 
      a(1)=>addersInputs_4_1, a(0)=>addersInputs_4_0, b(15)=>
      addersInputs_5_15, b(14)=>addersInputs_5_14, b(13)=>addersInputs_5_13, 
      b(12)=>addersInputs_5_12, b(11)=>addersInputs_5_11, b(10)=>
      addersInputs_5_10, b(9)=>addersInputs_5_9, b(8)=>addersInputs_5_8, 
      b(7)=>addersInputs_5_7, b(6)=>addersInputs_5_6, b(5)=>addersInputs_5_5, 
      b(4)=>addersInputs_5_4, b(3)=>addersInputs_5_3, b(2)=>addersInputs_5_2, 
      b(1)=>addersInputs_5_1, b(0)=>addersInputs_5_0, carryIn=>outShifter_15, 
      sum(15)=>addersMap_sum1Map_sum2Map_sum1_15, sum(14)=>
      addersMap_sum1Map_sum2Map_sum1_14, sum(13)=>
      addersMap_sum1Map_sum2Map_sum1_13, sum(12)=>
      addersMap_sum1Map_sum2Map_sum1_12, sum(11)=>
      addersMap_sum1Map_sum2Map_sum1_11, sum(10)=>
      addersMap_sum1Map_sum2Map_sum1_10, sum(9)=>
      addersMap_sum1Map_sum2Map_sum1_9, sum(8)=>
      addersMap_sum1Map_sum2Map_sum1_8, sum(7)=>
      addersMap_sum1Map_sum2Map_sum1_7, sum(6)=>
      addersMap_sum1Map_sum2Map_sum1_6, sum(5)=>
      addersMap_sum1Map_sum2Map_sum1_5, sum(4)=>
      addersMap_sum1Map_sum2Map_sum1_4, sum(3)=>
      addersMap_sum1Map_sum2Map_sum1_3, sum(2)=>
      addersMap_sum1Map_sum2Map_sum1_2, sum(1)=>
      addersMap_sum1Map_sum2Map_sum1_1, sum(0)=>
      addersMap_sum1Map_sum2Map_sum1_0, carryOut=>DANGLING(168));
   addersMap_sum1Map_sum2Map_sum2Map : NBitAdder_16 port map ( a(15)=>
      addersInputs_6_15, a(14)=>addersInputs_6_14, a(13)=>addersInputs_6_13, 
      a(12)=>addersInputs_6_12, a(11)=>addersInputs_6_11, a(10)=>
      addersInputs_6_10, a(9)=>addersInputs_6_9, a(8)=>addersInputs_6_8, 
      a(7)=>addersInputs_6_7, a(6)=>addersInputs_6_6, a(5)=>addersInputs_6_5, 
      a(4)=>addersInputs_6_4, a(3)=>addersInputs_6_3, a(2)=>addersInputs_6_2, 
      a(1)=>addersInputs_6_1, a(0)=>addersInputs_6_0, b(15)=>
      addersInputs_7_15, b(14)=>addersInputs_7_14, b(13)=>addersInputs_7_13, 
      b(12)=>addersInputs_7_12, b(11)=>addersInputs_7_11, b(10)=>
      addersInputs_7_10, b(9)=>addersInputs_7_9, b(8)=>addersInputs_7_8, 
      b(7)=>addersInputs_7_7, b(6)=>addersInputs_7_6, b(5)=>addersInputs_7_5, 
      b(4)=>addersInputs_7_4, b(3)=>addersInputs_7_3, b(2)=>addersInputs_7_2, 
      b(1)=>addersInputs_7_1, b(0)=>addersInputs_7_0, carryIn=>outShifter_15, 
      sum(15)=>addersMap_sum1Map_sum2Map_sum2_15, sum(14)=>
      addersMap_sum1Map_sum2Map_sum2_14, sum(13)=>
      addersMap_sum1Map_sum2Map_sum2_13, sum(12)=>
      addersMap_sum1Map_sum2Map_sum2_12, sum(11)=>
      addersMap_sum1Map_sum2Map_sum2_11, sum(10)=>
      addersMap_sum1Map_sum2Map_sum2_10, sum(9)=>
      addersMap_sum1Map_sum2Map_sum2_9, sum(8)=>
      addersMap_sum1Map_sum2Map_sum2_8, sum(7)=>
      addersMap_sum1Map_sum2Map_sum2_7, sum(6)=>
      addersMap_sum1Map_sum2Map_sum2_6, sum(5)=>
      addersMap_sum1Map_sum2Map_sum2_5, sum(4)=>
      addersMap_sum1Map_sum2Map_sum2_4, sum(3)=>
      addersMap_sum1Map_sum2Map_sum2_3, sum(2)=>
      addersMap_sum1Map_sum2Map_sum2_2, sum(1)=>
      addersMap_sum1Map_sum2Map_sum2_1, sum(0)=>
      addersMap_sum1Map_sum2Map_sum2_0, carryOut=>DANGLING(169));
   addersMap_sum1Map_sum2Map_sumFinalMap : NBitAdder_16 port map ( a(15)=>
      addersMap_sum1Map_sum2Map_sum1_15, a(14)=>
      addersMap_sum1Map_sum2Map_sum1_14, a(13)=>
      addersMap_sum1Map_sum2Map_sum1_13, a(12)=>
      addersMap_sum1Map_sum2Map_sum1_12, a(11)=>
      addersMap_sum1Map_sum2Map_sum1_11, a(10)=>
      addersMap_sum1Map_sum2Map_sum1_10, a(9)=>
      addersMap_sum1Map_sum2Map_sum1_9, a(8)=>
      addersMap_sum1Map_sum2Map_sum1_8, a(7)=>
      addersMap_sum1Map_sum2Map_sum1_7, a(6)=>
      addersMap_sum1Map_sum2Map_sum1_6, a(5)=>
      addersMap_sum1Map_sum2Map_sum1_5, a(4)=>
      addersMap_sum1Map_sum2Map_sum1_4, a(3)=>
      addersMap_sum1Map_sum2Map_sum1_3, a(2)=>
      addersMap_sum1Map_sum2Map_sum1_2, a(1)=>
      addersMap_sum1Map_sum2Map_sum1_1, a(0)=>
      addersMap_sum1Map_sum2Map_sum1_0, b(15)=>
      addersMap_sum1Map_sum2Map_sum2_15, b(14)=>
      addersMap_sum1Map_sum2Map_sum2_14, b(13)=>
      addersMap_sum1Map_sum2Map_sum2_13, b(12)=>
      addersMap_sum1Map_sum2Map_sum2_12, b(11)=>
      addersMap_sum1Map_sum2Map_sum2_11, b(10)=>
      addersMap_sum1Map_sum2Map_sum2_10, b(9)=>
      addersMap_sum1Map_sum2Map_sum2_9, b(8)=>
      addersMap_sum1Map_sum2Map_sum2_8, b(7)=>
      addersMap_sum1Map_sum2Map_sum2_7, b(6)=>
      addersMap_sum1Map_sum2Map_sum2_6, b(5)=>
      addersMap_sum1Map_sum2Map_sum2_5, b(4)=>
      addersMap_sum1Map_sum2Map_sum2_4, b(3)=>
      addersMap_sum1Map_sum2Map_sum2_3, b(2)=>
      addersMap_sum1Map_sum2Map_sum2_2, b(1)=>
      addersMap_sum1Map_sum2Map_sum2_1, b(0)=>
      addersMap_sum1Map_sum2Map_sum2_0, carryIn=>outShifter_15, sum(15)=>
      addersMap_sum1Map_sum2_15_dup_0, sum(14)=>
      addersMap_sum1Map_sum2_14_dup_0, sum(13)=>
      addersMap_sum1Map_sum2_13_dup_0, sum(12)=>
      addersMap_sum1Map_sum2_12_dup_0, sum(11)=>
      addersMap_sum1Map_sum2_11_dup_0, sum(10)=>
      addersMap_sum1Map_sum2_10_dup_0, sum(9)=>
      addersMap_sum1Map_sum2_9_dup_0, sum(8)=>addersMap_sum1Map_sum2_8_dup_0, 
      sum(7)=>addersMap_sum1Map_sum2_7_dup_0, sum(6)=>
      addersMap_sum1Map_sum2_6_dup_0, sum(5)=>addersMap_sum1Map_sum2_5_dup_0, 
      sum(4)=>addersMap_sum1Map_sum2_4_dup_0, sum(3)=>
      addersMap_sum1Map_sum2_3_dup_0, sum(2)=>addersMap_sum1Map_sum2_2_dup_0, 
      sum(1)=>addersMap_sum1Map_sum2_1_dup_0, sum(0)=>
      addersMap_sum1Map_sum2_0_dup_0, carryOut=>DANGLING(170));
   addersMap_sum2Map_sumFinalMap_dup_0 : NBitAdder_16 port map ( a(15)=>
      addersMap_sum2Map_sum1_15_dup_0, a(14)=>
      addersMap_sum2Map_sum1_14_dup_0, a(13)=>
      addersMap_sum2Map_sum1_13_dup_0, a(12)=>
      addersMap_sum2Map_sum1_12_dup_0, a(11)=>
      addersMap_sum2Map_sum1_11_dup_0, a(10)=>
      addersMap_sum2Map_sum1_10_dup_0, a(9)=>addersMap_sum2Map_sum1_9_dup_0, 
      a(8)=>addersMap_sum2Map_sum1_8_dup_0, a(7)=>
      addersMap_sum2Map_sum1_7_dup_0, a(6)=>addersMap_sum2Map_sum1_6_dup_0, 
      a(5)=>addersMap_sum2Map_sum1_5_dup_0, a(4)=>
      addersMap_sum2Map_sum1_4_dup_0, a(3)=>addersMap_sum2Map_sum1_3_dup_0, 
      a(2)=>addersMap_sum2Map_sum1_2_dup_0, a(1)=>
      addersMap_sum2Map_sum1_1_dup_0, a(0)=>addersMap_sum2Map_sum1_0_dup_0, 
      b(15)=>addersMap_sum2Map_sum2_15_dup_0, b(14)=>
      addersMap_sum2Map_sum2_14_dup_0, b(13)=>
      addersMap_sum2Map_sum2_13_dup_0, b(12)=>
      addersMap_sum2Map_sum2_12_dup_0, b(11)=>
      addersMap_sum2Map_sum2_11_dup_0, b(10)=>
      addersMap_sum2Map_sum2_10_dup_0, b(9)=>addersMap_sum2Map_sum2_9_dup_0, 
      b(8)=>addersMap_sum2Map_sum2_8_dup_0, b(7)=>
      addersMap_sum2Map_sum2_7_dup_0, b(6)=>addersMap_sum2Map_sum2_6_dup_0, 
      b(5)=>addersMap_sum2Map_sum2_5_dup_0, b(4)=>
      addersMap_sum2Map_sum2_4_dup_0, b(3)=>addersMap_sum2Map_sum2_3_dup_0, 
      b(2)=>addersMap_sum2Map_sum2_2_dup_0, b(1)=>
      addersMap_sum2Map_sum2_1_dup_0, b(0)=>addersMap_sum2Map_sum2_0_dup_0, 
      carryIn=>outShifter_15, sum(15)=>addersMap_sum2_15, sum(14)=>
      addersMap_sum2_14, sum(13)=>addersMap_sum2_13, sum(12)=>
      addersMap_sum2_12, sum(11)=>addersMap_sum2_11, sum(10)=>
      addersMap_sum2_10, sum(9)=>addersMap_sum2_9, sum(8)=>addersMap_sum2_8, 
      sum(7)=>addersMap_sum2_7, sum(6)=>addersMap_sum2_6, sum(5)=>
      addersMap_sum2_5, sum(4)=>addersMap_sum2_4, sum(3)=>addersMap_sum2_3, 
      sum(2)=>addersMap_sum2_2, sum(1)=>addersMap_sum2_1, sum(0)=>
      addersMap_sum2_0, carryOut=>DANGLING(171));
   addersMap_sum2Map_sum1Map_sum1Map : NBitAdder_16 port map ( a(15)=>
      addersInputs_9_15, a(14)=>addersInputs_9_14, a(13)=>addersInputs_9_13, 
      a(12)=>addersInputs_9_12, a(11)=>addersInputs_9_11, a(10)=>
      addersInputs_9_10, a(9)=>addersInputs_9_9, a(8)=>addersInputs_9_8, 
      a(7)=>addersInputs_9_7, a(6)=>addersInputs_9_6, a(5)=>addersInputs_9_5, 
      a(4)=>addersInputs_9_4, a(3)=>addersInputs_9_3, a(2)=>addersInputs_9_2, 
      a(1)=>addersInputs_9_1, a(0)=>addersInputs_9_0, b(15)=>
      addersInputs_10_15, b(14)=>addersInputs_10_14, b(13)=>
      addersInputs_10_13, b(12)=>addersInputs_10_12, b(11)=>
      addersInputs_10_11, b(10)=>addersInputs_10_10, b(9)=>addersInputs_10_9, 
      b(8)=>addersInputs_10_8, b(7)=>addersInputs_10_7, b(6)=>
      addersInputs_10_6, b(5)=>addersInputs_10_5, b(4)=>addersInputs_10_4, 
      b(3)=>addersInputs_10_3, b(2)=>addersInputs_10_2, b(1)=>
      addersInputs_10_1, b(0)=>addersInputs_10_0, carryIn=>outShifter_15, 
      sum(15)=>addersMap_sum2Map_sum1Map_sum1_15, sum(14)=>
      addersMap_sum2Map_sum1Map_sum1_14, sum(13)=>
      addersMap_sum2Map_sum1Map_sum1_13, sum(12)=>
      addersMap_sum2Map_sum1Map_sum1_12, sum(11)=>
      addersMap_sum2Map_sum1Map_sum1_11, sum(10)=>
      addersMap_sum2Map_sum1Map_sum1_10, sum(9)=>
      addersMap_sum2Map_sum1Map_sum1_9, sum(8)=>
      addersMap_sum2Map_sum1Map_sum1_8, sum(7)=>
      addersMap_sum2Map_sum1Map_sum1_7, sum(6)=>
      addersMap_sum2Map_sum1Map_sum1_6, sum(5)=>
      addersMap_sum2Map_sum1Map_sum1_5, sum(4)=>
      addersMap_sum2Map_sum1Map_sum1_4, sum(3)=>
      addersMap_sum2Map_sum1Map_sum1_3, sum(2)=>
      addersMap_sum2Map_sum1Map_sum1_2, sum(1)=>
      addersMap_sum2Map_sum1Map_sum1_1, sum(0)=>
      addersMap_sum2Map_sum1Map_sum1_0, carryOut=>DANGLING(172));
   addersMap_sum2Map_sum1Map_sum2Map : NBitAdder_16 port map ( a(15)=>
      addersInputs_11_15, a(14)=>addersInputs_11_14, a(13)=>
      addersInputs_11_13, a(12)=>addersInputs_11_12, a(11)=>
      addersInputs_11_11, a(10)=>addersInputs_11_10, a(9)=>addersInputs_11_9, 
      a(8)=>addersInputs_11_8, a(7)=>addersInputs_11_7, a(6)=>
      addersInputs_11_6, a(5)=>addersInputs_11_5, a(4)=>addersInputs_11_4, 
      a(3)=>addersInputs_11_3, a(2)=>addersInputs_11_2, a(1)=>
      addersInputs_11_1, a(0)=>addersInputs_11_0, b(15)=>addersInputs_12_15, 
      b(14)=>addersInputs_12_14, b(13)=>addersInputs_12_13, b(12)=>
      addersInputs_12_12, b(11)=>addersInputs_12_11, b(10)=>
      addersInputs_12_10, b(9)=>addersInputs_12_9, b(8)=>addersInputs_12_8, 
      b(7)=>addersInputs_12_7, b(6)=>addersInputs_12_6, b(5)=>
      addersInputs_12_5, b(4)=>addersInputs_12_4, b(3)=>addersInputs_12_3, 
      b(2)=>addersInputs_12_2, b(1)=>addersInputs_12_1, b(0)=>
      addersInputs_12_0, carryIn=>outShifter_15, sum(15)=>
      addersMap_sum2Map_sum1Map_sum2_15, sum(14)=>
      addersMap_sum2Map_sum1Map_sum2_14, sum(13)=>
      addersMap_sum2Map_sum1Map_sum2_13, sum(12)=>
      addersMap_sum2Map_sum1Map_sum2_12, sum(11)=>
      addersMap_sum2Map_sum1Map_sum2_11, sum(10)=>
      addersMap_sum2Map_sum1Map_sum2_10, sum(9)=>
      addersMap_sum2Map_sum1Map_sum2_9, sum(8)=>
      addersMap_sum2Map_sum1Map_sum2_8, sum(7)=>
      addersMap_sum2Map_sum1Map_sum2_7, sum(6)=>
      addersMap_sum2Map_sum1Map_sum2_6, sum(5)=>
      addersMap_sum2Map_sum1Map_sum2_5, sum(4)=>
      addersMap_sum2Map_sum1Map_sum2_4, sum(3)=>
      addersMap_sum2Map_sum1Map_sum2_3, sum(2)=>
      addersMap_sum2Map_sum1Map_sum2_2, sum(1)=>
      addersMap_sum2Map_sum1Map_sum2_1, sum(0)=>
      addersMap_sum2Map_sum1Map_sum2_0, carryOut=>DANGLING(173));
   addersMap_sum2Map_sum1Map_sumFinalMap : NBitAdder_16 port map ( a(15)=>
      addersMap_sum2Map_sum1Map_sum1_15, a(14)=>
      addersMap_sum2Map_sum1Map_sum1_14, a(13)=>
      addersMap_sum2Map_sum1Map_sum1_13, a(12)=>
      addersMap_sum2Map_sum1Map_sum1_12, a(11)=>
      addersMap_sum2Map_sum1Map_sum1_11, a(10)=>
      addersMap_sum2Map_sum1Map_sum1_10, a(9)=>
      addersMap_sum2Map_sum1Map_sum1_9, a(8)=>
      addersMap_sum2Map_sum1Map_sum1_8, a(7)=>
      addersMap_sum2Map_sum1Map_sum1_7, a(6)=>
      addersMap_sum2Map_sum1Map_sum1_6, a(5)=>
      addersMap_sum2Map_sum1Map_sum1_5, a(4)=>
      addersMap_sum2Map_sum1Map_sum1_4, a(3)=>
      addersMap_sum2Map_sum1Map_sum1_3, a(2)=>
      addersMap_sum2Map_sum1Map_sum1_2, a(1)=>
      addersMap_sum2Map_sum1Map_sum1_1, a(0)=>
      addersMap_sum2Map_sum1Map_sum1_0, b(15)=>
      addersMap_sum2Map_sum1Map_sum2_15, b(14)=>
      addersMap_sum2Map_sum1Map_sum2_14, b(13)=>
      addersMap_sum2Map_sum1Map_sum2_13, b(12)=>
      addersMap_sum2Map_sum1Map_sum2_12, b(11)=>
      addersMap_sum2Map_sum1Map_sum2_11, b(10)=>
      addersMap_sum2Map_sum1Map_sum2_10, b(9)=>
      addersMap_sum2Map_sum1Map_sum2_9, b(8)=>
      addersMap_sum2Map_sum1Map_sum2_8, b(7)=>
      addersMap_sum2Map_sum1Map_sum2_7, b(6)=>
      addersMap_sum2Map_sum1Map_sum2_6, b(5)=>
      addersMap_sum2Map_sum1Map_sum2_5, b(4)=>
      addersMap_sum2Map_sum1Map_sum2_4, b(3)=>
      addersMap_sum2Map_sum1Map_sum2_3, b(2)=>
      addersMap_sum2Map_sum1Map_sum2_2, b(1)=>
      addersMap_sum2Map_sum1Map_sum2_1, b(0)=>
      addersMap_sum2Map_sum1Map_sum2_0, carryIn=>outShifter_15, sum(15)=>
      addersMap_sum2Map_sum1_15_dup_0, sum(14)=>
      addersMap_sum2Map_sum1_14_dup_0, sum(13)=>
      addersMap_sum2Map_sum1_13_dup_0, sum(12)=>
      addersMap_sum2Map_sum1_12_dup_0, sum(11)=>
      addersMap_sum2Map_sum1_11_dup_0, sum(10)=>
      addersMap_sum2Map_sum1_10_dup_0, sum(9)=>
      addersMap_sum2Map_sum1_9_dup_0, sum(8)=>addersMap_sum2Map_sum1_8_dup_0, 
      sum(7)=>addersMap_sum2Map_sum1_7_dup_0, sum(6)=>
      addersMap_sum2Map_sum1_6_dup_0, sum(5)=>addersMap_sum2Map_sum1_5_dup_0, 
      sum(4)=>addersMap_sum2Map_sum1_4_dup_0, sum(3)=>
      addersMap_sum2Map_sum1_3_dup_0, sum(2)=>addersMap_sum2Map_sum1_2_dup_0, 
      sum(1)=>addersMap_sum2Map_sum1_1_dup_0, sum(0)=>
      addersMap_sum2Map_sum1_0_dup_0, carryOut=>DANGLING(174));
   addersMap_sum2Map_sum2Map_sum1Map : NBitAdder_16 port map ( a(15)=>
      addersInputs_13_15, a(14)=>addersInputs_13_14, a(13)=>
      addersInputs_13_13, a(12)=>addersInputs_13_12, a(11)=>
      addersInputs_13_11, a(10)=>addersInputs_13_10, a(9)=>addersInputs_13_9, 
      a(8)=>addersInputs_13_8, a(7)=>addersInputs_13_7, a(6)=>
      addersInputs_13_6, a(5)=>addersInputs_13_5, a(4)=>addersInputs_13_4, 
      a(3)=>addersInputs_13_3, a(2)=>addersInputs_13_2, a(1)=>
      addersInputs_13_1, a(0)=>addersInputs_13_0, b(15)=>addersInputs_14_15, 
      b(14)=>addersInputs_14_14, b(13)=>addersInputs_14_13, b(12)=>
      addersInputs_14_12, b(11)=>addersInputs_14_11, b(10)=>
      addersInputs_14_10, b(9)=>addersInputs_14_9, b(8)=>addersInputs_14_8, 
      b(7)=>addersInputs_14_7, b(6)=>addersInputs_14_6, b(5)=>
      addersInputs_14_5, b(4)=>addersInputs_14_4, b(3)=>addersInputs_14_3, 
      b(2)=>addersInputs_14_2, b(1)=>addersInputs_14_1, b(0)=>
      addersInputs_14_0, carryIn=>outShifter_15, sum(15)=>
      addersMap_sum2Map_sum2Map_sum1_15, sum(14)=>
      addersMap_sum2Map_sum2Map_sum1_14, sum(13)=>
      addersMap_sum2Map_sum2Map_sum1_13, sum(12)=>
      addersMap_sum2Map_sum2Map_sum1_12, sum(11)=>
      addersMap_sum2Map_sum2Map_sum1_11, sum(10)=>
      addersMap_sum2Map_sum2Map_sum1_10, sum(9)=>
      addersMap_sum2Map_sum2Map_sum1_9, sum(8)=>
      addersMap_sum2Map_sum2Map_sum1_8, sum(7)=>
      addersMap_sum2Map_sum2Map_sum1_7, sum(6)=>
      addersMap_sum2Map_sum2Map_sum1_6, sum(5)=>
      addersMap_sum2Map_sum2Map_sum1_5, sum(4)=>
      addersMap_sum2Map_sum2Map_sum1_4, sum(3)=>
      addersMap_sum2Map_sum2Map_sum1_3, sum(2)=>
      addersMap_sum2Map_sum2Map_sum1_2, sum(1)=>
      addersMap_sum2Map_sum2Map_sum1_1, sum(0)=>
      addersMap_sum2Map_sum2Map_sum1_0, carryOut=>DANGLING(175));
   addersMap_sum2Map_sum2Map_sum2Map : NBitAdder_16 port map ( a(15)=>
      addersInputs_15_15, a(14)=>addersInputs_15_14, a(13)=>
      addersInputs_15_13, a(12)=>addersInputs_15_12, a(11)=>
      addersInputs_15_11, a(10)=>addersInputs_15_10, a(9)=>addersInputs_15_9, 
      a(8)=>addersInputs_15_8, a(7)=>addersInputs_15_7, a(6)=>
      addersInputs_15_6, a(5)=>addersInputs_15_5, a(4)=>addersInputs_15_4, 
      a(3)=>addersInputs_15_3, a(2)=>addersInputs_15_2, a(1)=>
      addersInputs_15_1, a(0)=>addersInputs_15_0, b(15)=>addersInputs_16_15, 
      b(14)=>addersInputs_16_14, b(13)=>addersInputs_16_13, b(12)=>
      addersInputs_16_12, b(11)=>addersInputs_16_11, b(10)=>
      addersInputs_16_10, b(9)=>addersInputs_16_9, b(8)=>addersInputs_16_8, 
      b(7)=>addersInputs_16_7, b(6)=>addersInputs_16_6, b(5)=>
      addersInputs_16_5, b(4)=>addersInputs_16_4, b(3)=>addersInputs_16_3, 
      b(2)=>addersInputs_16_2, b(1)=>addersInputs_16_1, b(0)=>
      addersInputs_16_0, carryIn=>outShifter_15, sum(15)=>
      addersMap_sum2Map_sum2Map_sum2_15, sum(14)=>
      addersMap_sum2Map_sum2Map_sum2_14, sum(13)=>
      addersMap_sum2Map_sum2Map_sum2_13, sum(12)=>
      addersMap_sum2Map_sum2Map_sum2_12, sum(11)=>
      addersMap_sum2Map_sum2Map_sum2_11, sum(10)=>
      addersMap_sum2Map_sum2Map_sum2_10, sum(9)=>
      addersMap_sum2Map_sum2Map_sum2_9, sum(8)=>
      addersMap_sum2Map_sum2Map_sum2_8, sum(7)=>
      addersMap_sum2Map_sum2Map_sum2_7, sum(6)=>
      addersMap_sum2Map_sum2Map_sum2_6, sum(5)=>
      addersMap_sum2Map_sum2Map_sum2_5, sum(4)=>
      addersMap_sum2Map_sum2Map_sum2_4, sum(3)=>
      addersMap_sum2Map_sum2Map_sum2_3, sum(2)=>
      addersMap_sum2Map_sum2Map_sum2_2, sum(1)=>
      addersMap_sum2Map_sum2Map_sum2_1, sum(0)=>
      addersMap_sum2Map_sum2Map_sum2_0, carryOut=>DANGLING(176));
   addersMap_sum2Map_sum2Map_sumFinalMap : NBitAdder_16 port map ( a(15)=>
      addersMap_sum2Map_sum2Map_sum1_15, a(14)=>
      addersMap_sum2Map_sum2Map_sum1_14, a(13)=>
      addersMap_sum2Map_sum2Map_sum1_13, a(12)=>
      addersMap_sum2Map_sum2Map_sum1_12, a(11)=>
      addersMap_sum2Map_sum2Map_sum1_11, a(10)=>
      addersMap_sum2Map_sum2Map_sum1_10, a(9)=>
      addersMap_sum2Map_sum2Map_sum1_9, a(8)=>
      addersMap_sum2Map_sum2Map_sum1_8, a(7)=>
      addersMap_sum2Map_sum2Map_sum1_7, a(6)=>
      addersMap_sum2Map_sum2Map_sum1_6, a(5)=>
      addersMap_sum2Map_sum2Map_sum1_5, a(4)=>
      addersMap_sum2Map_sum2Map_sum1_4, a(3)=>
      addersMap_sum2Map_sum2Map_sum1_3, a(2)=>
      addersMap_sum2Map_sum2Map_sum1_2, a(1)=>
      addersMap_sum2Map_sum2Map_sum1_1, a(0)=>
      addersMap_sum2Map_sum2Map_sum1_0, b(15)=>
      addersMap_sum2Map_sum2Map_sum2_15, b(14)=>
      addersMap_sum2Map_sum2Map_sum2_14, b(13)=>
      addersMap_sum2Map_sum2Map_sum2_13, b(12)=>
      addersMap_sum2Map_sum2Map_sum2_12, b(11)=>
      addersMap_sum2Map_sum2Map_sum2_11, b(10)=>
      addersMap_sum2Map_sum2Map_sum2_10, b(9)=>
      addersMap_sum2Map_sum2Map_sum2_9, b(8)=>
      addersMap_sum2Map_sum2Map_sum2_8, b(7)=>
      addersMap_sum2Map_sum2Map_sum2_7, b(6)=>
      addersMap_sum2Map_sum2Map_sum2_6, b(5)=>
      addersMap_sum2Map_sum2Map_sum2_5, b(4)=>
      addersMap_sum2Map_sum2Map_sum2_4, b(3)=>
      addersMap_sum2Map_sum2Map_sum2_3, b(2)=>
      addersMap_sum2Map_sum2Map_sum2_2, b(1)=>
      addersMap_sum2Map_sum2Map_sum2_1, b(0)=>
      addersMap_sum2Map_sum2Map_sum2_0, carryIn=>outShifter_15, sum(15)=>
      addersMap_sum2Map_sum2_15_dup_0, sum(14)=>
      addersMap_sum2Map_sum2_14_dup_0, sum(13)=>
      addersMap_sum2Map_sum2_13_dup_0, sum(12)=>
      addersMap_sum2Map_sum2_12_dup_0, sum(11)=>
      addersMap_sum2Map_sum2_11_dup_0, sum(10)=>
      addersMap_sum2Map_sum2_10_dup_0, sum(9)=>
      addersMap_sum2Map_sum2_9_dup_0, sum(8)=>addersMap_sum2Map_sum2_8_dup_0, 
      sum(7)=>addersMap_sum2Map_sum2_7_dup_0, sum(6)=>
      addersMap_sum2Map_sum2_6_dup_0, sum(5)=>addersMap_sum2Map_sum2_5_dup_0, 
      sum(4)=>addersMap_sum2Map_sum2_4_dup_0, sum(3)=>
      addersMap_sum2Map_sum2_3_dup_0, sum(2)=>addersMap_sum2Map_sum2_2_dup_0, 
      sum(1)=>addersMap_sum2Map_sum2_1_dup_0, sum(0)=>
      addersMap_sum2Map_sum2_0_dup_0, carryOut=>DANGLING(177));
   addersMap_sum3Map_sumFinalMap : NBitAdder_16 port map ( a(15)=>
      addersMap_sum3Map_sum1_15, a(14)=>addersMap_sum3Map_sum1_14, a(13)=>
      addersMap_sum3Map_sum1_13, a(12)=>addersMap_sum3Map_sum1_12, a(11)=>
      addersMap_sum3Map_sum1_11, a(10)=>addersMap_sum3Map_sum1_10, a(9)=>
      addersMap_sum3Map_sum1_9, a(8)=>addersMap_sum3Map_sum1_8, a(7)=>
      addersMap_sum3Map_sum1_7, a(6)=>addersMap_sum3Map_sum1_6, a(5)=>
      addersMap_sum3Map_sum1_5, a(4)=>addersMap_sum3Map_sum1_4, a(3)=>
      addersMap_sum3Map_sum1_3, a(2)=>addersMap_sum3Map_sum1_2, a(1)=>
      addersMap_sum3Map_sum1_1, a(0)=>addersMap_sum3Map_sum1_0, b(15)=>
      addersMap_sum3Map_sum2_15, b(14)=>addersMap_sum3Map_sum2_14, b(13)=>
      addersMap_sum3Map_sum2_13, b(12)=>addersMap_sum3Map_sum2_12, b(11)=>
      addersMap_sum3Map_sum2_11, b(10)=>addersMap_sum3Map_sum2_10, b(9)=>
      addersMap_sum3Map_sum2_9, b(8)=>addersMap_sum3Map_sum2_8, b(7)=>
      addersMap_sum3Map_sum2_7, b(6)=>addersMap_sum3Map_sum2_6, b(5)=>
      addersMap_sum3Map_sum2_5, b(4)=>addersMap_sum3Map_sum2_4, b(3)=>
      addersMap_sum3Map_sum2_3, b(2)=>addersMap_sum3Map_sum2_2, b(1)=>
      addersMap_sum3Map_sum2_1, b(0)=>addersMap_sum3Map_sum2_0, carryIn=>
      outShifter_15, sum(15)=>addersMap_sum3_15, sum(14)=>addersMap_sum3_14, 
      sum(13)=>addersMap_sum3_13, sum(12)=>addersMap_sum3_12, sum(11)=>
      addersMap_sum3_11, sum(10)=>addersMap_sum3_10, sum(9)=>
      addersMap_sum3_9, sum(8)=>addersMap_sum3_8, sum(7)=>addersMap_sum3_7, 
      sum(6)=>addersMap_sum3_6, sum(5)=>addersMap_sum3_5, sum(4)=>
      addersMap_sum3_4, sum(3)=>addersMap_sum3_3, sum(2)=>addersMap_sum3_2, 
      sum(1)=>addersMap_sum3_1, sum(0)=>addersMap_sum3_0, carryOut=>DANGLING
      (178));
   addersMap_sum3Map_sum1Map_sum1Map : NBitAdder_16 port map ( a(15)=>
      addersInputs_17_15, a(14)=>addersInputs_17_14, a(13)=>
      addersInputs_17_13, a(12)=>addersInputs_17_12, a(11)=>
      addersInputs_17_11, a(10)=>addersInputs_17_10, a(9)=>addersInputs_17_9, 
      a(8)=>addersInputs_17_8, a(7)=>addersInputs_17_7, a(6)=>
      addersInputs_17_6, a(5)=>addersInputs_17_5, a(4)=>addersInputs_17_4, 
      a(3)=>addersInputs_17_3, a(2)=>addersInputs_17_2, a(1)=>
      addersInputs_17_1, a(0)=>addersInputs_17_0, b(15)=>addersInputs_18_15, 
      b(14)=>addersInputs_18_14, b(13)=>addersInputs_18_13, b(12)=>
      addersInputs_18_12, b(11)=>addersInputs_18_11, b(10)=>
      addersInputs_18_10, b(9)=>addersInputs_18_9, b(8)=>addersInputs_18_8, 
      b(7)=>addersInputs_18_7, b(6)=>addersInputs_18_6, b(5)=>
      addersInputs_18_5, b(4)=>addersInputs_18_4, b(3)=>addersInputs_18_3, 
      b(2)=>addersInputs_18_2, b(1)=>addersInputs_18_1, b(0)=>
      addersInputs_18_0, carryIn=>outShifter_15, sum(15)=>
      addersMap_sum3Map_sum1Map_sum1_15, sum(14)=>
      addersMap_sum3Map_sum1Map_sum1_14, sum(13)=>
      addersMap_sum3Map_sum1Map_sum1_13, sum(12)=>
      addersMap_sum3Map_sum1Map_sum1_12, sum(11)=>
      addersMap_sum3Map_sum1Map_sum1_11, sum(10)=>
      addersMap_sum3Map_sum1Map_sum1_10, sum(9)=>
      addersMap_sum3Map_sum1Map_sum1_9, sum(8)=>
      addersMap_sum3Map_sum1Map_sum1_8, sum(7)=>
      addersMap_sum3Map_sum1Map_sum1_7, sum(6)=>
      addersMap_sum3Map_sum1Map_sum1_6, sum(5)=>
      addersMap_sum3Map_sum1Map_sum1_5, sum(4)=>
      addersMap_sum3Map_sum1Map_sum1_4, sum(3)=>
      addersMap_sum3Map_sum1Map_sum1_3, sum(2)=>
      addersMap_sum3Map_sum1Map_sum1_2, sum(1)=>
      addersMap_sum3Map_sum1Map_sum1_1, sum(0)=>
      addersMap_sum3Map_sum1Map_sum1_0, carryOut=>DANGLING(179));
   addersMap_sum3Map_sum1Map_sum2Map : NBitAdder_16 port map ( a(15)=>
      addersInputs_19_15, a(14)=>addersInputs_19_14, a(13)=>
      addersInputs_19_13, a(12)=>addersInputs_19_12, a(11)=>
      addersInputs_19_11, a(10)=>addersInputs_19_10, a(9)=>addersInputs_19_9, 
      a(8)=>addersInputs_19_8, a(7)=>addersInputs_19_7, a(6)=>
      addersInputs_19_6, a(5)=>addersInputs_19_5, a(4)=>addersInputs_19_4, 
      a(3)=>addersInputs_19_3, a(2)=>addersInputs_19_2, a(1)=>
      addersInputs_19_1, a(0)=>addersInputs_19_0, b(15)=>addersInputs_20_15, 
      b(14)=>addersInputs_20_14, b(13)=>addersInputs_20_13, b(12)=>
      addersInputs_20_12, b(11)=>addersInputs_20_11, b(10)=>
      addersInputs_20_10, b(9)=>addersInputs_20_9, b(8)=>addersInputs_20_8, 
      b(7)=>addersInputs_20_7, b(6)=>addersInputs_20_6, b(5)=>
      addersInputs_20_5, b(4)=>addersInputs_20_4, b(3)=>addersInputs_20_3, 
      b(2)=>addersInputs_20_2, b(1)=>addersInputs_20_1, b(0)=>
      addersInputs_20_0, carryIn=>outShifter_15, sum(15)=>
      addersMap_sum3Map_sum1Map_sum2_15, sum(14)=>
      addersMap_sum3Map_sum1Map_sum2_14, sum(13)=>
      addersMap_sum3Map_sum1Map_sum2_13, sum(12)=>
      addersMap_sum3Map_sum1Map_sum2_12, sum(11)=>
      addersMap_sum3Map_sum1Map_sum2_11, sum(10)=>
      addersMap_sum3Map_sum1Map_sum2_10, sum(9)=>
      addersMap_sum3Map_sum1Map_sum2_9, sum(8)=>
      addersMap_sum3Map_sum1Map_sum2_8, sum(7)=>
      addersMap_sum3Map_sum1Map_sum2_7, sum(6)=>
      addersMap_sum3Map_sum1Map_sum2_6, sum(5)=>
      addersMap_sum3Map_sum1Map_sum2_5, sum(4)=>
      addersMap_sum3Map_sum1Map_sum2_4, sum(3)=>
      addersMap_sum3Map_sum1Map_sum2_3, sum(2)=>
      addersMap_sum3Map_sum1Map_sum2_2, sum(1)=>
      addersMap_sum3Map_sum1Map_sum2_1, sum(0)=>
      addersMap_sum3Map_sum1Map_sum2_0, carryOut=>DANGLING(180));
   addersMap_sum3Map_sum1Map_sumFinalMap : NBitAdder_16 port map ( a(15)=>
      addersMap_sum3Map_sum1Map_sum1_15, a(14)=>
      addersMap_sum3Map_sum1Map_sum1_14, a(13)=>
      addersMap_sum3Map_sum1Map_sum1_13, a(12)=>
      addersMap_sum3Map_sum1Map_sum1_12, a(11)=>
      addersMap_sum3Map_sum1Map_sum1_11, a(10)=>
      addersMap_sum3Map_sum1Map_sum1_10, a(9)=>
      addersMap_sum3Map_sum1Map_sum1_9, a(8)=>
      addersMap_sum3Map_sum1Map_sum1_8, a(7)=>
      addersMap_sum3Map_sum1Map_sum1_7, a(6)=>
      addersMap_sum3Map_sum1Map_sum1_6, a(5)=>
      addersMap_sum3Map_sum1Map_sum1_5, a(4)=>
      addersMap_sum3Map_sum1Map_sum1_4, a(3)=>
      addersMap_sum3Map_sum1Map_sum1_3, a(2)=>
      addersMap_sum3Map_sum1Map_sum1_2, a(1)=>
      addersMap_sum3Map_sum1Map_sum1_1, a(0)=>
      addersMap_sum3Map_sum1Map_sum1_0, b(15)=>
      addersMap_sum3Map_sum1Map_sum2_15, b(14)=>
      addersMap_sum3Map_sum1Map_sum2_14, b(13)=>
      addersMap_sum3Map_sum1Map_sum2_13, b(12)=>
      addersMap_sum3Map_sum1Map_sum2_12, b(11)=>
      addersMap_sum3Map_sum1Map_sum2_11, b(10)=>
      addersMap_sum3Map_sum1Map_sum2_10, b(9)=>
      addersMap_sum3Map_sum1Map_sum2_9, b(8)=>
      addersMap_sum3Map_sum1Map_sum2_8, b(7)=>
      addersMap_sum3Map_sum1Map_sum2_7, b(6)=>
      addersMap_sum3Map_sum1Map_sum2_6, b(5)=>
      addersMap_sum3Map_sum1Map_sum2_5, b(4)=>
      addersMap_sum3Map_sum1Map_sum2_4, b(3)=>
      addersMap_sum3Map_sum1Map_sum2_3, b(2)=>
      addersMap_sum3Map_sum1Map_sum2_2, b(1)=>
      addersMap_sum3Map_sum1Map_sum2_1, b(0)=>
      addersMap_sum3Map_sum1Map_sum2_0, carryIn=>outShifter_15, sum(15)=>
      addersMap_sum3Map_sum1_15, sum(14)=>addersMap_sum3Map_sum1_14, sum(13)
      =>addersMap_sum3Map_sum1_13, sum(12)=>addersMap_sum3Map_sum1_12, 
      sum(11)=>addersMap_sum3Map_sum1_11, sum(10)=>addersMap_sum3Map_sum1_10, 
      sum(9)=>addersMap_sum3Map_sum1_9, sum(8)=>addersMap_sum3Map_sum1_8, 
      sum(7)=>addersMap_sum3Map_sum1_7, sum(6)=>addersMap_sum3Map_sum1_6, 
      sum(5)=>addersMap_sum3Map_sum1_5, sum(4)=>addersMap_sum3Map_sum1_4, 
      sum(3)=>addersMap_sum3Map_sum1_3, sum(2)=>addersMap_sum3Map_sum1_2, 
      sum(1)=>addersMap_sum3Map_sum1_1, sum(0)=>addersMap_sum3Map_sum1_0, 
      carryOut=>DANGLING(181));
   addersMap_sum3Map_sum2Map_sum1Map : NBitAdder_16 port map ( a(15)=>
      addersInputs_21_15, a(14)=>addersInputs_21_14, a(13)=>
      addersInputs_21_13, a(12)=>addersInputs_21_12, a(11)=>
      addersInputs_21_11, a(10)=>addersInputs_21_10, a(9)=>addersInputs_21_9, 
      a(8)=>addersInputs_21_8, a(7)=>addersInputs_21_7, a(6)=>
      addersInputs_21_6, a(5)=>addersInputs_21_5, a(4)=>addersInputs_21_4, 
      a(3)=>addersInputs_21_3, a(2)=>addersInputs_21_2, a(1)=>
      addersInputs_21_1, a(0)=>addersInputs_21_0, b(15)=>addersInputs_22_15, 
      b(14)=>addersInputs_22_14, b(13)=>addersInputs_22_13, b(12)=>
      addersInputs_22_12, b(11)=>addersInputs_22_11, b(10)=>
      addersInputs_22_10, b(9)=>addersInputs_22_9, b(8)=>addersInputs_22_8, 
      b(7)=>addersInputs_22_7, b(6)=>addersInputs_22_6, b(5)=>
      addersInputs_22_5, b(4)=>addersInputs_22_4, b(3)=>addersInputs_22_3, 
      b(2)=>addersInputs_22_2, b(1)=>addersInputs_22_1, b(0)=>
      addersInputs_22_0, carryIn=>outShifter_15, sum(15)=>
      addersMap_sum3Map_sum2Map_sum1_15, sum(14)=>
      addersMap_sum3Map_sum2Map_sum1_14, sum(13)=>
      addersMap_sum3Map_sum2Map_sum1_13, sum(12)=>
      addersMap_sum3Map_sum2Map_sum1_12, sum(11)=>
      addersMap_sum3Map_sum2Map_sum1_11, sum(10)=>
      addersMap_sum3Map_sum2Map_sum1_10, sum(9)=>
      addersMap_sum3Map_sum2Map_sum1_9, sum(8)=>
      addersMap_sum3Map_sum2Map_sum1_8, sum(7)=>
      addersMap_sum3Map_sum2Map_sum1_7, sum(6)=>
      addersMap_sum3Map_sum2Map_sum1_6, sum(5)=>
      addersMap_sum3Map_sum2Map_sum1_5, sum(4)=>
      addersMap_sum3Map_sum2Map_sum1_4, sum(3)=>
      addersMap_sum3Map_sum2Map_sum1_3, sum(2)=>
      addersMap_sum3Map_sum2Map_sum1_2, sum(1)=>
      addersMap_sum3Map_sum2Map_sum1_1, sum(0)=>
      addersMap_sum3Map_sum2Map_sum1_0, carryOut=>DANGLING(182));
   addersMap_sum3Map_sum2Map_sum2Map : NBitAdder_16 port map ( a(15)=>
      addersInputs_23_15, a(14)=>addersInputs_23_14, a(13)=>
      addersInputs_23_13, a(12)=>addersInputs_23_12, a(11)=>
      addersInputs_23_11, a(10)=>addersInputs_23_10, a(9)=>addersInputs_23_9, 
      a(8)=>addersInputs_23_8, a(7)=>addersInputs_23_7, a(6)=>
      addersInputs_23_6, a(5)=>addersInputs_23_5, a(4)=>addersInputs_23_4, 
      a(3)=>addersInputs_23_3, a(2)=>addersInputs_23_2, a(1)=>
      addersInputs_23_1, a(0)=>addersInputs_23_0, b(15)=>addersInputs_24_15, 
      b(14)=>addersInputs_24_14, b(13)=>addersInputs_24_13, b(12)=>
      addersInputs_24_12, b(11)=>addersInputs_24_11, b(10)=>
      addersInputs_24_10, b(9)=>addersInputs_24_9, b(8)=>addersInputs_24_8, 
      b(7)=>addersInputs_24_7, b(6)=>addersInputs_24_6, b(5)=>
      addersInputs_24_5, b(4)=>addersInputs_24_4, b(3)=>addersInputs_24_3, 
      b(2)=>addersInputs_24_2, b(1)=>addersInputs_24_1, b(0)=>
      addersInputs_24_0, carryIn=>outShifter_15, sum(15)=>
      addersMap_sum3Map_sum2Map_sum2_15, sum(14)=>
      addersMap_sum3Map_sum2Map_sum2_14, sum(13)=>
      addersMap_sum3Map_sum2Map_sum2_13, sum(12)=>
      addersMap_sum3Map_sum2Map_sum2_12, sum(11)=>
      addersMap_sum3Map_sum2Map_sum2_11, sum(10)=>
      addersMap_sum3Map_sum2Map_sum2_10, sum(9)=>
      addersMap_sum3Map_sum2Map_sum2_9, sum(8)=>
      addersMap_sum3Map_sum2Map_sum2_8, sum(7)=>
      addersMap_sum3Map_sum2Map_sum2_7, sum(6)=>
      addersMap_sum3Map_sum2Map_sum2_6, sum(5)=>
      addersMap_sum3Map_sum2Map_sum2_5, sum(4)=>
      addersMap_sum3Map_sum2Map_sum2_4, sum(3)=>
      addersMap_sum3Map_sum2Map_sum2_3, sum(2)=>
      addersMap_sum3Map_sum2Map_sum2_2, sum(1)=>
      addersMap_sum3Map_sum2Map_sum2_1, sum(0)=>
      addersMap_sum3Map_sum2Map_sum2_0, carryOut=>DANGLING(183));
   addersMap_sum3Map_sum2Map_sumFinalMap : NBitAdder_16 port map ( a(15)=>
      addersMap_sum3Map_sum2Map_sum1_15, a(14)=>
      addersMap_sum3Map_sum2Map_sum1_14, a(13)=>
      addersMap_sum3Map_sum2Map_sum1_13, a(12)=>
      addersMap_sum3Map_sum2Map_sum1_12, a(11)=>
      addersMap_sum3Map_sum2Map_sum1_11, a(10)=>
      addersMap_sum3Map_sum2Map_sum1_10, a(9)=>
      addersMap_sum3Map_sum2Map_sum1_9, a(8)=>
      addersMap_sum3Map_sum2Map_sum1_8, a(7)=>
      addersMap_sum3Map_sum2Map_sum1_7, a(6)=>
      addersMap_sum3Map_sum2Map_sum1_6, a(5)=>
      addersMap_sum3Map_sum2Map_sum1_5, a(4)=>
      addersMap_sum3Map_sum2Map_sum1_4, a(3)=>
      addersMap_sum3Map_sum2Map_sum1_3, a(2)=>
      addersMap_sum3Map_sum2Map_sum1_2, a(1)=>
      addersMap_sum3Map_sum2Map_sum1_1, a(0)=>
      addersMap_sum3Map_sum2Map_sum1_0, b(15)=>
      addersMap_sum3Map_sum2Map_sum2_15, b(14)=>
      addersMap_sum3Map_sum2Map_sum2_14, b(13)=>
      addersMap_sum3Map_sum2Map_sum2_13, b(12)=>
      addersMap_sum3Map_sum2Map_sum2_12, b(11)=>
      addersMap_sum3Map_sum2Map_sum2_11, b(10)=>
      addersMap_sum3Map_sum2Map_sum2_10, b(9)=>
      addersMap_sum3Map_sum2Map_sum2_9, b(8)=>
      addersMap_sum3Map_sum2Map_sum2_8, b(7)=>
      addersMap_sum3Map_sum2Map_sum2_7, b(6)=>
      addersMap_sum3Map_sum2Map_sum2_6, b(5)=>
      addersMap_sum3Map_sum2Map_sum2_5, b(4)=>
      addersMap_sum3Map_sum2Map_sum2_4, b(3)=>
      addersMap_sum3Map_sum2Map_sum2_3, b(2)=>
      addersMap_sum3Map_sum2Map_sum2_2, b(1)=>
      addersMap_sum3Map_sum2Map_sum2_1, b(0)=>
      addersMap_sum3Map_sum2Map_sum2_0, carryIn=>outShifter_15, sum(15)=>
      addersMap_sum3Map_sum2_15, sum(14)=>addersMap_sum3Map_sum2_14, sum(13)
      =>addersMap_sum3Map_sum2_13, sum(12)=>addersMap_sum3Map_sum2_12, 
      sum(11)=>addersMap_sum3Map_sum2_11, sum(10)=>addersMap_sum3Map_sum2_10, 
      sum(9)=>addersMap_sum3Map_sum2_9, sum(8)=>addersMap_sum3Map_sum2_8, 
      sum(7)=>addersMap_sum3Map_sum2_7, sum(6)=>addersMap_sum3Map_sum2_6, 
      sum(5)=>addersMap_sum3Map_sum2_5, sum(4)=>addersMap_sum3Map_sum2_4, 
      sum(3)=>addersMap_sum3Map_sum2_3, sum(2)=>addersMap_sum3Map_sum2_2, 
      sum(1)=>addersMap_sum3Map_sum2_1, sum(0)=>addersMap_sum3Map_sum2_0, 
      carryOut=>DANGLING(184));
   ix2066 : fake_gnd port map ( Y=>outShifter_15);
   ix2918 : nand03 port map ( Y=>nx2917, A0=>writeFilter, A1=>nx3412, A2=>
      decoderRow(2));
   ix3413 : nor02_2x port map ( Y=>nx3412, A0=>decoderRow(1), A1=>
      decoderRow(0));
   ix3437 : nor03_2x port map ( Y=>regFileMap_filterEnables_3, A0=>nx2923, 
      A1=>decoderRow(2), A2=>nx2925);
   ix2924 : inv02 port map ( Y=>nx2923, A=>writeFilter);
   ix2926 : nand02 port map ( Y=>nx2925, A0=>decoderRow(1), A1=>
      decoderRow(0));
   ix3449 : nor03_2x port map ( Y=>regFileMap_filterEnables_2, A0=>nx2923, 
      A1=>decoderRow(2), A2=>nx2929);
   ix2930 : nand02 port map ( Y=>nx2929, A0=>decoderRow(1), A1=>nx2931);
   ix2932 : inv01 port map ( Y=>nx2931, A=>decoderRow(0));
   ix3461 : nor03_2x port map ( Y=>regFileMap_filterEnables_1, A0=>nx2923, 
      A1=>decoderRow(2), A2=>nx2935);
   ix2936 : nand02 port map ( Y=>nx2935, A0=>nx2937, A1=>decoderRow(0));
   ix2938 : inv01 port map ( Y=>nx2937, A=>decoderRow(1));
   ix3475 : nor03_2x port map ( Y=>regFileMap_filterEnables_0, A0=>nx2923, 
      A1=>decoderRow(2), A2=>nx2941);
   ix2942 : inv01 port map ( Y=>nx2941, A=>nx3470);
   ix3471 : nor02_2x port map ( Y=>nx3470, A0=>decoderRow(1), A1=>
      decoderRow(0));
   ix3425 : inv01 port map ( Y=>regFileMap_page2Enables_4, A=>nx2947);
   ix2948 : nand03 port map ( Y=>nx2947, A0=>writePage2, A1=>nx3412, A2=>
      decoderRow(2));
   ix3439 : nor03_2x port map ( Y=>regFileMap_page2Enables_3, A0=>nx2951, A1
      =>decoderRow(2), A2=>nx2925);
   ix2952 : inv02 port map ( Y=>nx2951, A=>writePage2);
   ix3451 : nor03_2x port map ( Y=>regFileMap_page2Enables_2, A0=>nx2951, A1
      =>decoderRow(2), A2=>nx2929);
   ix3463 : nor03_2x port map ( Y=>regFileMap_page2Enables_1, A0=>nx2951, A1
      =>decoderRow(2), A2=>nx2935);
   ix3477 : nor03_2x port map ( Y=>regFileMap_page2Enables_0, A0=>nx2951, A1
      =>decoderRow(2), A2=>nx2941);
   ix3427 : inv01 port map ( Y=>regFileMap_page1Enables_4, A=>nx2959);
   ix2960 : nand03 port map ( Y=>nx2959, A0=>writePage1, A1=>nx3412, A2=>
      decoderRow(2));
   ix3441 : nor03_2x port map ( Y=>regFileMap_page1Enables_3, A0=>nx2963, A1
      =>decoderRow(2), A2=>nx2925);
   ix2964 : inv02 port map ( Y=>nx2963, A=>writePage1);
   ix3453 : nor03_2x port map ( Y=>regFileMap_page1Enables_2, A0=>nx2963, A1
      =>decoderRow(2), A2=>nx2929);
   ix3465 : nor03_2x port map ( Y=>regFileMap_page1Enables_1, A0=>nx2963, A1
      =>decoderRow(2), A2=>nx2935);
   ix3479 : nor03_2x port map ( Y=>regFileMap_page1Enables_0, A0=>nx2963, A1
      =>decoderRow(2), A2=>nx2941);
   ix215 : nand02 port map ( Y=>addersInputs_24_0, A0=>nx2971, A1=>nx2973);
   ix2972 : nand02 port map ( Y=>nx2971, A0=>currentPage_24_0, A1=>layerType
   );
   ix2974 : nand02 port map ( Y=>nx2973, A0=>outMuls_24_0, A1=>nx5200);
   ix223 : nand02 port map ( Y=>addersInputs_24_1, A0=>nx2979, A1=>nx2981);
   ix2980 : nand02 port map ( Y=>nx2979, A0=>currentPage_24_1, A1=>layerType
   );
   ix2982 : nand02 port map ( Y=>nx2981, A0=>outMuls_24_1, A1=>nx5200);
   ix231 : nand02 port map ( Y=>addersInputs_24_2, A0=>nx2985, A1=>nx2987);
   ix2986 : nand02 port map ( Y=>nx2985, A0=>currentPage_24_2, A1=>layerType
   );
   ix2988 : nand02 port map ( Y=>nx2987, A0=>outMuls_24_2, A1=>nx5200);
   ix239 : nand02 port map ( Y=>addersInputs_24_3, A0=>nx2991, A1=>nx2993);
   ix2992 : nand02 port map ( Y=>nx2991, A0=>currentPage_24_3, A1=>layerType
   );
   ix2994 : nand02 port map ( Y=>nx2993, A0=>outMuls_24_3, A1=>nx5200);
   ix247 : nand02 port map ( Y=>addersInputs_24_4, A0=>nx2997, A1=>nx2999);
   ix2998 : nand02 port map ( Y=>nx2997, A0=>currentPage_24_4, A1=>layerType
   );
   ix3000 : nand02 port map ( Y=>nx2999, A0=>outMuls_24_4, A1=>nx5200);
   ix255 : nand02 port map ( Y=>addersInputs_24_5, A0=>nx3003, A1=>nx3005);
   ix3004 : nand02 port map ( Y=>nx3003, A0=>currentPage_24_5, A1=>layerType
   );
   ix3006 : nand02 port map ( Y=>nx3005, A0=>outMuls_24_5, A1=>nx5200);
   ix263 : nand02 port map ( Y=>addersInputs_24_6, A0=>nx3009, A1=>nx3011);
   ix3010 : nand02 port map ( Y=>nx3009, A0=>currentPage_24_6, A1=>layerType
   );
   ix3012 : nand02 port map ( Y=>nx3011, A0=>outMuls_24_6, A1=>nx5200);
   ix271 : nand02 port map ( Y=>addersInputs_24_7, A0=>nx3015, A1=>nx3017);
   ix3016 : nand02 port map ( Y=>nx3015, A0=>currentPage_24_7, A1=>layerType
   );
   ix3018 : nand02 port map ( Y=>nx3017, A0=>outMuls_24_7, A1=>nx5202);
   ix279 : nand02 port map ( Y=>addersInputs_24_8, A0=>nx3021, A1=>nx3023);
   ix3022 : nand02 port map ( Y=>nx3021, A0=>currentPage_24_8, A1=>layerType
   );
   ix3024 : nand02 port map ( Y=>nx3023, A0=>outMuls_24_8, A1=>nx5202);
   ix287 : nand02 port map ( Y=>addersInputs_24_9, A0=>nx3027, A1=>nx3029);
   ix3028 : nand02 port map ( Y=>nx3027, A0=>currentPage_24_9, A1=>layerType
   );
   ix3030 : nand02 port map ( Y=>nx3029, A0=>outMuls_24_9, A1=>nx5202);
   ix295 : nand02 port map ( Y=>addersInputs_24_10, A0=>nx3033, A1=>nx3035);
   ix3034 : nand02 port map ( Y=>nx3033, A0=>currentPage_24_10, A1=>
      layerType);
   ix3036 : nand02 port map ( Y=>nx3035, A0=>outMuls_24_10, A1=>nx5202);
   ix303 : nand02 port map ( Y=>addersInputs_24_11, A0=>nx3039, A1=>nx3041);
   ix3040 : nand02 port map ( Y=>nx3039, A0=>currentPage_24_11, A1=>
      layerType);
   ix3042 : nand02 port map ( Y=>nx3041, A0=>outMuls_24_11, A1=>nx5202);
   ix311 : nand02 port map ( Y=>addersInputs_24_12, A0=>nx3045, A1=>nx3047);
   ix3046 : nand02 port map ( Y=>nx3045, A0=>currentPage_24_12, A1=>
      layerType);
   ix3048 : nand02 port map ( Y=>nx3047, A0=>outMuls_24_12, A1=>nx5202);
   ix319 : nand02 port map ( Y=>addersInputs_24_13, A0=>nx3051, A1=>nx3053);
   ix3052 : nand02 port map ( Y=>nx3051, A0=>currentPage_24_13, A1=>
      layerType);
   ix3054 : nand02 port map ( Y=>nx3053, A0=>outMuls_24_13, A1=>nx5202);
   ix327 : nand02 port map ( Y=>addersInputs_24_14, A0=>nx3057, A1=>nx3059);
   ix3058 : nand02 port map ( Y=>nx3057, A0=>currentPage_24_14, A1=>
      layerType);
   ix3060 : nand02 port map ( Y=>nx3059, A0=>outMuls_24_14, A1=>nx5204);
   ix335 : nand02 port map ( Y=>addersInputs_24_15, A0=>nx3063, A1=>nx3065);
   ix3064 : nand02 port map ( Y=>nx3063, A0=>currentPage_24_15, A1=>
      layerType);
   ix3066 : nand02 port map ( Y=>nx3065, A0=>outMuls_24_15, A1=>nx5204);
   ix343 : nand02 port map ( Y=>addersInputs_23_0, A0=>nx3069, A1=>nx3071);
   ix3070 : nand02 port map ( Y=>nx3069, A0=>currentPage_23_0, A1=>layerType
   );
   ix3072 : nand02 port map ( Y=>nx3071, A0=>outMuls_23_0, A1=>nx5204);
   ix351 : nand02 port map ( Y=>addersInputs_23_1, A0=>nx3075, A1=>nx3077);
   ix3076 : nand02 port map ( Y=>nx3075, A0=>currentPage_23_1, A1=>layerType
   );
   ix3078 : nand02 port map ( Y=>nx3077, A0=>outMuls_23_1, A1=>nx5204);
   ix359 : nand02 port map ( Y=>addersInputs_23_2, A0=>nx3081, A1=>nx3083);
   ix3082 : nand02 port map ( Y=>nx3081, A0=>currentPage_23_2, A1=>layerType
   );
   ix3084 : nand02 port map ( Y=>nx3083, A0=>outMuls_23_2, A1=>nx5204);
   ix367 : nand02 port map ( Y=>addersInputs_23_3, A0=>nx3087, A1=>nx3089);
   ix3088 : nand02 port map ( Y=>nx3087, A0=>currentPage_23_3, A1=>layerType
   );
   ix3090 : nand02 port map ( Y=>nx3089, A0=>outMuls_23_3, A1=>nx5204);
   ix375 : nand02 port map ( Y=>addersInputs_23_4, A0=>nx3093, A1=>nx3095);
   ix3094 : nand02 port map ( Y=>nx3093, A0=>currentPage_23_4, A1=>layerType
   );
   ix3096 : nand02 port map ( Y=>nx3095, A0=>outMuls_23_4, A1=>nx5204);
   ix383 : nand02 port map ( Y=>addersInputs_23_5, A0=>nx3099, A1=>nx3101);
   ix3100 : nand02 port map ( Y=>nx3099, A0=>currentPage_23_5, A1=>layerType
   );
   ix3102 : nand02 port map ( Y=>nx3101, A0=>outMuls_23_5, A1=>nx5206);
   ix391 : nand02 port map ( Y=>addersInputs_23_6, A0=>nx3105, A1=>nx3107);
   ix3106 : nand02 port map ( Y=>nx3105, A0=>currentPage_23_6, A1=>layerType
   );
   ix3108 : nand02 port map ( Y=>nx3107, A0=>outMuls_23_6, A1=>nx5206);
   ix399 : nand02 port map ( Y=>addersInputs_23_7, A0=>nx3111, A1=>nx3113);
   ix3112 : nand02 port map ( Y=>nx3111, A0=>currentPage_23_7, A1=>layerType
   );
   ix3114 : nand02 port map ( Y=>nx3113, A0=>outMuls_23_7, A1=>nx5206);
   ix407 : nand02 port map ( Y=>addersInputs_23_8, A0=>nx3117, A1=>nx3119);
   ix3118 : nand02 port map ( Y=>nx3117, A0=>currentPage_23_8, A1=>layerType
   );
   ix3120 : nand02 port map ( Y=>nx3119, A0=>outMuls_23_8, A1=>nx5206);
   ix415 : nand02 port map ( Y=>addersInputs_23_9, A0=>nx3123, A1=>nx3125);
   ix3124 : nand02 port map ( Y=>nx3123, A0=>currentPage_23_9, A1=>layerType
   );
   ix3126 : nand02 port map ( Y=>nx3125, A0=>outMuls_23_9, A1=>nx5206);
   ix423 : nand02 port map ( Y=>addersInputs_23_10, A0=>nx3129, A1=>nx3131);
   ix3130 : nand02 port map ( Y=>nx3129, A0=>currentPage_23_10, A1=>
      layerType);
   ix3132 : nand02 port map ( Y=>nx3131, A0=>outMuls_23_10, A1=>nx5206);
   ix431 : nand02 port map ( Y=>addersInputs_23_11, A0=>nx3135, A1=>nx3137);
   ix3136 : nand02 port map ( Y=>nx3135, A0=>currentPage_23_11, A1=>
      layerType);
   ix3138 : nand02 port map ( Y=>nx3137, A0=>outMuls_23_11, A1=>nx5206);
   ix439 : nand02 port map ( Y=>addersInputs_23_12, A0=>nx3141, A1=>nx3143);
   ix3142 : nand02 port map ( Y=>nx3141, A0=>currentPage_23_12, A1=>
      layerType);
   ix3144 : nand02 port map ( Y=>nx3143, A0=>outMuls_23_12, A1=>nx5208);
   ix447 : nand02 port map ( Y=>addersInputs_23_13, A0=>nx3147, A1=>nx3149);
   ix3148 : nand02 port map ( Y=>nx3147, A0=>currentPage_23_13, A1=>
      layerType);
   ix3150 : nand02 port map ( Y=>nx3149, A0=>outMuls_23_13, A1=>nx5208);
   ix455 : nand02 port map ( Y=>addersInputs_23_14, A0=>nx3153, A1=>nx3155);
   ix3154 : nand02 port map ( Y=>nx3153, A0=>currentPage_23_14, A1=>
      layerType);
   ix3156 : nand02 port map ( Y=>nx3155, A0=>outMuls_23_14, A1=>nx5208);
   ix463 : nand02 port map ( Y=>addersInputs_23_15, A0=>nx3159, A1=>nx3161);
   ix3160 : nand02 port map ( Y=>nx3159, A0=>currentPage_23_15, A1=>
      layerType);
   ix3162 : nand02 port map ( Y=>nx3161, A0=>outMuls_23_15, A1=>nx5208);
   ix471 : nand02 port map ( Y=>addersInputs_22_0, A0=>nx3165, A1=>nx3167);
   ix3166 : nand02 port map ( Y=>nx3165, A0=>currentPage_22_0, A1=>layerType
   );
   ix3168 : nand02 port map ( Y=>nx3167, A0=>outMuls_22_0, A1=>nx5208);
   ix479 : nand02 port map ( Y=>addersInputs_22_1, A0=>nx3171, A1=>nx3173);
   ix3172 : nand02 port map ( Y=>nx3171, A0=>currentPage_22_1, A1=>layerType
   );
   ix3174 : nand02 port map ( Y=>nx3173, A0=>outMuls_22_1, A1=>nx5208);
   ix487 : nand02 port map ( Y=>addersInputs_22_2, A0=>nx3177, A1=>nx3179);
   ix3178 : nand02 port map ( Y=>nx3177, A0=>currentPage_22_2, A1=>layerType
   );
   ix3180 : nand02 port map ( Y=>nx3179, A0=>outMuls_22_2, A1=>nx5208);
   ix495 : nand02 port map ( Y=>addersInputs_22_3, A0=>nx3183, A1=>nx3185);
   ix3184 : nand02 port map ( Y=>nx3183, A0=>currentPage_22_3, A1=>layerType
   );
   ix3186 : nand02 port map ( Y=>nx3185, A0=>outMuls_22_3, A1=>nx5210);
   ix503 : nand02 port map ( Y=>addersInputs_22_4, A0=>nx3189, A1=>nx3191);
   ix3190 : nand02 port map ( Y=>nx3189, A0=>currentPage_22_4, A1=>layerType
   );
   ix3192 : nand02 port map ( Y=>nx3191, A0=>outMuls_22_4, A1=>nx5210);
   ix511 : nand02 port map ( Y=>addersInputs_22_5, A0=>nx3195, A1=>nx3197);
   ix3196 : nand02 port map ( Y=>nx3195, A0=>currentPage_22_5, A1=>layerType
   );
   ix3198 : nand02 port map ( Y=>nx3197, A0=>outMuls_22_5, A1=>nx5210);
   ix519 : nand02 port map ( Y=>addersInputs_22_6, A0=>nx3201, A1=>nx3203);
   ix3202 : nand02 port map ( Y=>nx3201, A0=>currentPage_22_6, A1=>layerType
   );
   ix3204 : nand02 port map ( Y=>nx3203, A0=>outMuls_22_6, A1=>nx5210);
   ix527 : nand02 port map ( Y=>addersInputs_22_7, A0=>nx3207, A1=>nx3209);
   ix3208 : nand02 port map ( Y=>nx3207, A0=>currentPage_22_7, A1=>layerType
   );
   ix3210 : nand02 port map ( Y=>nx3209, A0=>outMuls_22_7, A1=>nx5210);
   ix535 : nand02 port map ( Y=>addersInputs_22_8, A0=>nx3213, A1=>nx3215);
   ix3214 : nand02 port map ( Y=>nx3213, A0=>currentPage_22_8, A1=>layerType
   );
   ix3216 : nand02 port map ( Y=>nx3215, A0=>outMuls_22_8, A1=>nx5210);
   ix543 : nand02 port map ( Y=>addersInputs_22_9, A0=>nx3219, A1=>nx3221);
   ix3220 : nand02 port map ( Y=>nx3219, A0=>currentPage_22_9, A1=>layerType
   );
   ix3222 : nand02 port map ( Y=>nx3221, A0=>outMuls_22_9, A1=>nx5210);
   ix551 : nand02 port map ( Y=>addersInputs_22_10, A0=>nx3225, A1=>nx3227);
   ix3226 : nand02 port map ( Y=>nx3225, A0=>currentPage_22_10, A1=>
      layerType);
   ix3228 : nand02 port map ( Y=>nx3227, A0=>outMuls_22_10, A1=>nx5212);
   ix559 : nand02 port map ( Y=>addersInputs_22_11, A0=>nx3231, A1=>nx3233);
   ix3232 : nand02 port map ( Y=>nx3231, A0=>currentPage_22_11, A1=>
      layerType);
   ix3234 : nand02 port map ( Y=>nx3233, A0=>outMuls_22_11, A1=>nx5212);
   ix567 : nand02 port map ( Y=>addersInputs_22_12, A0=>nx3237, A1=>nx3239);
   ix3238 : nand02 port map ( Y=>nx3237, A0=>currentPage_22_12, A1=>
      layerType);
   ix3240 : nand02 port map ( Y=>nx3239, A0=>outMuls_22_12, A1=>nx5212);
   ix575 : nand02 port map ( Y=>addersInputs_22_13, A0=>nx3243, A1=>nx3245);
   ix3244 : nand02 port map ( Y=>nx3243, A0=>currentPage_22_13, A1=>
      layerType);
   ix3246 : nand02 port map ( Y=>nx3245, A0=>outMuls_22_13, A1=>nx5212);
   ix583 : nand02 port map ( Y=>addersInputs_22_14, A0=>nx3249, A1=>nx3251);
   ix3250 : nand02 port map ( Y=>nx3249, A0=>currentPage_22_14, A1=>
      layerType);
   ix3252 : nand02 port map ( Y=>nx3251, A0=>outMuls_22_14, A1=>nx5212);
   ix591 : nand02 port map ( Y=>addersInputs_22_15, A0=>nx3255, A1=>nx3257);
   ix3256 : nand02 port map ( Y=>nx3255, A0=>currentPage_22_15, A1=>
      layerType);
   ix3258 : nand02 port map ( Y=>nx3257, A0=>outMuls_22_15, A1=>nx5212);
   ix599 : nand02 port map ( Y=>addersInputs_21_0, A0=>nx3261, A1=>nx3263);
   ix3262 : nand02 port map ( Y=>nx3261, A0=>currentPage_21_0, A1=>layerType
   );
   ix3264 : nand02 port map ( Y=>nx3263, A0=>outMuls_21_0, A1=>nx5212);
   ix607 : nand02 port map ( Y=>addersInputs_21_1, A0=>nx3267, A1=>nx3269);
   ix3268 : nand02 port map ( Y=>nx3267, A0=>currentPage_21_1, A1=>layerType
   );
   ix3270 : nand02 port map ( Y=>nx3269, A0=>outMuls_21_1, A1=>nx5214);
   ix615 : nand02 port map ( Y=>addersInputs_21_2, A0=>nx3273, A1=>nx3275);
   ix3274 : nand02 port map ( Y=>nx3273, A0=>currentPage_21_2, A1=>layerType
   );
   ix3276 : nand02 port map ( Y=>nx3275, A0=>outMuls_21_2, A1=>nx5214);
   ix623 : nand02 port map ( Y=>addersInputs_21_3, A0=>nx3279, A1=>nx3281);
   ix3280 : nand02 port map ( Y=>nx3279, A0=>currentPage_21_3, A1=>layerType
   );
   ix3282 : nand02 port map ( Y=>nx3281, A0=>outMuls_21_3, A1=>nx5214);
   ix631 : nand02 port map ( Y=>addersInputs_21_4, A0=>nx3285, A1=>nx3287);
   ix3286 : nand02 port map ( Y=>nx3285, A0=>currentPage_21_4, A1=>layerType
   );
   ix3288 : nand02 port map ( Y=>nx3287, A0=>outMuls_21_4, A1=>nx5214);
   ix639 : nand02 port map ( Y=>addersInputs_21_5, A0=>nx3291, A1=>nx3293);
   ix3292 : nand02 port map ( Y=>nx3291, A0=>currentPage_21_5, A1=>layerType
   );
   ix3294 : nand02 port map ( Y=>nx3293, A0=>outMuls_21_5, A1=>nx5214);
   ix647 : nand02 port map ( Y=>addersInputs_21_6, A0=>nx3297, A1=>nx3299);
   ix3298 : nand02 port map ( Y=>nx3297, A0=>currentPage_21_6, A1=>layerType
   );
   ix3300 : nand02 port map ( Y=>nx3299, A0=>outMuls_21_6, A1=>nx5214);
   ix655 : nand02 port map ( Y=>addersInputs_21_7, A0=>nx3303, A1=>nx3305);
   ix3304 : nand02 port map ( Y=>nx3303, A0=>currentPage_21_7, A1=>layerType
   );
   ix3306 : nand02 port map ( Y=>nx3305, A0=>outMuls_21_7, A1=>nx5214);
   ix663 : nand02 port map ( Y=>addersInputs_21_8, A0=>nx3309, A1=>nx3311);
   ix3310 : nand02 port map ( Y=>nx3309, A0=>currentPage_21_8, A1=>layerType
   );
   ix3312 : nand02 port map ( Y=>nx3311, A0=>outMuls_21_8, A1=>nx5216);
   ix671 : nand02 port map ( Y=>addersInputs_21_9, A0=>nx3315, A1=>nx3317);
   ix3316 : nand02 port map ( Y=>nx3315, A0=>currentPage_21_9, A1=>layerType
   );
   ix3318 : nand02 port map ( Y=>nx3317, A0=>outMuls_21_9, A1=>nx5216);
   ix679 : nand02 port map ( Y=>addersInputs_21_10, A0=>nx3321, A1=>nx3323);
   ix3322 : nand02 port map ( Y=>nx3321, A0=>currentPage_21_10, A1=>
      layerType);
   ix3324 : nand02 port map ( Y=>nx3323, A0=>outMuls_21_10, A1=>nx5216);
   ix687 : nand02 port map ( Y=>addersInputs_21_11, A0=>nx3327, A1=>nx3329);
   ix3328 : nand02 port map ( Y=>nx3327, A0=>currentPage_21_11, A1=>
      layerType);
   ix3330 : nand02 port map ( Y=>nx3329, A0=>outMuls_21_11, A1=>nx5216);
   ix695 : nand02 port map ( Y=>addersInputs_21_12, A0=>nx3333, A1=>nx3335);
   ix3334 : nand02 port map ( Y=>nx3333, A0=>currentPage_21_12, A1=>
      layerType);
   ix3336 : nand02 port map ( Y=>nx3335, A0=>outMuls_21_12, A1=>nx5216);
   ix703 : nand02 port map ( Y=>addersInputs_21_13, A0=>nx3339, A1=>nx3341);
   ix3340 : nand02 port map ( Y=>nx3339, A0=>currentPage_21_13, A1=>
      layerType);
   ix3342 : nand02 port map ( Y=>nx3341, A0=>outMuls_21_13, A1=>nx5216);
   ix711 : nand02 port map ( Y=>addersInputs_21_14, A0=>nx3345, A1=>nx3347);
   ix3346 : nand02 port map ( Y=>nx3345, A0=>currentPage_21_14, A1=>
      layerType);
   ix3348 : nand02 port map ( Y=>nx3347, A0=>outMuls_21_14, A1=>nx5216);
   ix719 : nand02 port map ( Y=>addersInputs_21_15, A0=>nx3351, A1=>nx3353);
   ix3352 : nand02 port map ( Y=>nx3351, A0=>currentPage_21_15, A1=>
      layerType);
   ix3354 : nand02 port map ( Y=>nx3353, A0=>outMuls_21_15, A1=>nx5218);
   ix727 : nand02 port map ( Y=>addersInputs_20_0, A0=>nx3357, A1=>nx3359);
   ix3358 : nand02 port map ( Y=>nx3357, A0=>currentPage_20_0, A1=>layerType
   );
   ix3360 : nand02 port map ( Y=>nx3359, A0=>outMuls_20_0, A1=>nx5218);
   ix735 : nand02 port map ( Y=>addersInputs_20_1, A0=>nx3363, A1=>nx3365);
   ix3364 : nand02 port map ( Y=>nx3363, A0=>currentPage_20_1, A1=>layerType
   );
   ix3366 : nand02 port map ( Y=>nx3365, A0=>outMuls_20_1, A1=>nx5218);
   ix743 : nand02 port map ( Y=>addersInputs_20_2, A0=>nx3369, A1=>nx3371);
   ix3370 : nand02 port map ( Y=>nx3369, A0=>currentPage_20_2, A1=>layerType
   );
   ix3372 : nand02 port map ( Y=>nx3371, A0=>outMuls_20_2, A1=>nx5218);
   ix751 : nand02 port map ( Y=>addersInputs_20_3, A0=>nx3375, A1=>nx3377);
   ix3376 : nand02 port map ( Y=>nx3375, A0=>currentPage_20_3, A1=>layerType
   );
   ix3378 : nand02 port map ( Y=>nx3377, A0=>outMuls_20_3, A1=>nx5218);
   ix759 : nand02 port map ( Y=>addersInputs_20_4, A0=>nx3381, A1=>nx3383);
   ix3382 : nand02 port map ( Y=>nx3381, A0=>currentPage_20_4, A1=>layerType
   );
   ix3384 : nand02 port map ( Y=>nx3383, A0=>outMuls_20_4, A1=>nx5218);
   ix767 : nand02 port map ( Y=>addersInputs_20_5, A0=>nx3387, A1=>nx3389);
   ix3388 : nand02 port map ( Y=>nx3387, A0=>currentPage_20_5, A1=>layerType
   );
   ix3390 : nand02 port map ( Y=>nx3389, A0=>outMuls_20_5, A1=>nx5218);
   ix775 : nand02 port map ( Y=>addersInputs_20_6, A0=>nx3393, A1=>nx3395);
   ix3394 : nand02 port map ( Y=>nx3393, A0=>currentPage_20_6, A1=>layerType
   );
   ix3396 : nand02 port map ( Y=>nx3395, A0=>outMuls_20_6, A1=>nx5220);
   ix783 : nand02 port map ( Y=>addersInputs_20_7, A0=>nx3399, A1=>nx3401);
   ix3400 : nand02 port map ( Y=>nx3399, A0=>currentPage_20_7, A1=>layerType
   );
   ix3402 : nand02 port map ( Y=>nx3401, A0=>outMuls_20_7, A1=>nx5220);
   ix791 : nand02 port map ( Y=>addersInputs_20_8, A0=>nx3405, A1=>nx3407);
   ix3406 : nand02 port map ( Y=>nx3405, A0=>currentPage_20_8, A1=>layerType
   );
   ix3408 : nand02 port map ( Y=>nx3407, A0=>outMuls_20_8, A1=>nx5220);
   ix799 : nand02 port map ( Y=>addersInputs_20_9, A0=>nx3411, A1=>nx3413);
   ix3412 : nand02 port map ( Y=>nx3411, A0=>currentPage_20_9, A1=>layerType
   );
   ix3414 : nand02 port map ( Y=>nx3413, A0=>outMuls_20_9, A1=>nx5220);
   ix807 : nand02 port map ( Y=>addersInputs_20_10, A0=>nx3417, A1=>nx3419);
   ix3418 : nand02 port map ( Y=>nx3417, A0=>currentPage_20_10, A1=>
      layerType);
   ix3420 : nand02 port map ( Y=>nx3419, A0=>outMuls_20_10, A1=>nx5220);
   ix815 : nand02 port map ( Y=>addersInputs_20_11, A0=>nx3423, A1=>nx3425);
   ix3424 : nand02 port map ( Y=>nx3423, A0=>currentPage_20_11, A1=>
      layerType);
   ix3426 : nand02 port map ( Y=>nx3425, A0=>outMuls_20_11, A1=>nx5220);
   ix823 : nand02 port map ( Y=>addersInputs_20_12, A0=>nx3429, A1=>nx3431);
   ix3430 : nand02 port map ( Y=>nx3429, A0=>currentPage_20_12, A1=>
      layerType);
   ix3432 : nand02 port map ( Y=>nx3431, A0=>outMuls_20_12, A1=>nx5220);
   ix831 : nand02 port map ( Y=>addersInputs_20_13, A0=>nx3435, A1=>nx3437);
   ix3436 : nand02 port map ( Y=>nx3435, A0=>currentPage_20_13, A1=>
      layerType);
   ix3438 : nand02 port map ( Y=>nx3437, A0=>outMuls_20_13, A1=>nx5222);
   ix839 : nand02 port map ( Y=>addersInputs_20_14, A0=>nx3441, A1=>nx3443);
   ix3442 : nand02 port map ( Y=>nx3441, A0=>currentPage_20_14, A1=>
      layerType);
   ix3444 : nand02 port map ( Y=>nx3443, A0=>outMuls_20_14, A1=>nx5222);
   ix847 : nand02 port map ( Y=>addersInputs_20_15, A0=>nx3447, A1=>nx3449);
   ix3448 : nand02 port map ( Y=>nx3447, A0=>currentPage_20_15, A1=>
      layerType);
   ix3450 : nand02 port map ( Y=>nx3449, A0=>outMuls_20_15, A1=>nx5222);
   ix855 : nand02 port map ( Y=>addersInputs_19_0, A0=>nx3453, A1=>nx3455);
   ix3454 : nand02 port map ( Y=>nx3453, A0=>currentPage_19_0, A1=>layerType
   );
   ix3456 : nand02 port map ( Y=>nx3455, A0=>outMuls_19_0, A1=>nx5222);
   ix863 : nand02 port map ( Y=>addersInputs_19_1, A0=>nx3459, A1=>nx3461);
   ix3460 : nand02 port map ( Y=>nx3459, A0=>currentPage_19_1, A1=>layerType
   );
   ix3462 : nand02 port map ( Y=>nx3461, A0=>outMuls_19_1, A1=>nx5222);
   ix871 : nand02 port map ( Y=>addersInputs_19_2, A0=>nx3465, A1=>nx3467);
   ix3466 : nand02 port map ( Y=>nx3465, A0=>currentPage_19_2, A1=>layerType
   );
   ix3468 : nand02 port map ( Y=>nx3467, A0=>outMuls_19_2, A1=>nx5222);
   ix879 : nand02 port map ( Y=>addersInputs_19_3, A0=>nx3471, A1=>nx3473);
   ix3472 : nand02 port map ( Y=>nx3471, A0=>currentPage_19_3, A1=>layerType
   );
   ix3474 : nand02 port map ( Y=>nx3473, A0=>outMuls_19_3, A1=>nx5222);
   ix887 : nand02 port map ( Y=>addersInputs_19_4, A0=>nx3477, A1=>nx3479);
   ix3478 : nand02 port map ( Y=>nx3477, A0=>currentPage_19_4, A1=>layerType
   );
   ix3480 : nand02 port map ( Y=>nx3479, A0=>outMuls_19_4, A1=>nx5224);
   ix895 : nand02 port map ( Y=>addersInputs_19_5, A0=>nx3483, A1=>nx3485);
   ix3484 : nand02 port map ( Y=>nx3483, A0=>currentPage_19_5, A1=>layerType
   );
   ix3486 : nand02 port map ( Y=>nx3485, A0=>outMuls_19_5, A1=>nx5224);
   ix903 : nand02 port map ( Y=>addersInputs_19_6, A0=>nx3488, A1=>nx3490);
   ix3489 : nand02 port map ( Y=>nx3488, A0=>currentPage_19_6, A1=>layerType
   );
   ix3491 : nand02 port map ( Y=>nx3490, A0=>outMuls_19_6, A1=>nx5224);
   ix911 : nand02 port map ( Y=>addersInputs_19_7, A0=>nx3493, A1=>nx3495);
   ix3494 : nand02 port map ( Y=>nx3493, A0=>currentPage_19_7, A1=>layerType
   );
   ix3496 : nand02 port map ( Y=>nx3495, A0=>outMuls_19_7, A1=>nx5224);
   ix919 : nand02 port map ( Y=>addersInputs_19_8, A0=>nx3498, A1=>nx3500);
   ix3499 : nand02 port map ( Y=>nx3498, A0=>currentPage_19_8, A1=>layerType
   );
   ix3501 : nand02 port map ( Y=>nx3500, A0=>outMuls_19_8, A1=>nx5224);
   ix927 : nand02 port map ( Y=>addersInputs_19_9, A0=>nx3503, A1=>nx3505);
   ix3504 : nand02 port map ( Y=>nx3503, A0=>currentPage_19_9, A1=>layerType
   );
   ix3506 : nand02 port map ( Y=>nx3505, A0=>outMuls_19_9, A1=>nx5224);
   ix935 : nand02 port map ( Y=>addersInputs_19_10, A0=>nx3508, A1=>nx3510);
   ix3509 : nand02 port map ( Y=>nx3508, A0=>currentPage_19_10, A1=>
      layerType);
   ix3511 : nand02 port map ( Y=>nx3510, A0=>outMuls_19_10, A1=>nx5224);
   ix943 : nand02 port map ( Y=>addersInputs_19_11, A0=>nx3513, A1=>nx3515);
   ix3514 : nand02 port map ( Y=>nx3513, A0=>currentPage_19_11, A1=>
      layerType);
   ix3516 : nand02 port map ( Y=>nx3515, A0=>outMuls_19_11, A1=>nx5226);
   ix951 : nand02 port map ( Y=>addersInputs_19_12, A0=>nx3518, A1=>nx3520);
   ix3519 : nand02 port map ( Y=>nx3518, A0=>currentPage_19_12, A1=>
      layerType);
   ix3521 : nand02 port map ( Y=>nx3520, A0=>outMuls_19_12, A1=>nx5226);
   ix959 : nand02 port map ( Y=>addersInputs_19_13, A0=>nx3523, A1=>nx3525);
   ix3524 : nand02 port map ( Y=>nx3523, A0=>currentPage_19_13, A1=>
      layerType);
   ix3526 : nand02 port map ( Y=>nx3525, A0=>outMuls_19_13, A1=>nx5226);
   ix967 : nand02 port map ( Y=>addersInputs_19_14, A0=>nx3528, A1=>nx3530);
   ix3529 : nand02 port map ( Y=>nx3528, A0=>currentPage_19_14, A1=>
      layerType);
   ix3531 : nand02 port map ( Y=>nx3530, A0=>outMuls_19_14, A1=>nx5226);
   ix975 : nand02 port map ( Y=>addersInputs_19_15, A0=>nx3533, A1=>nx3535);
   ix3534 : nand02 port map ( Y=>nx3533, A0=>currentPage_19_15, A1=>
      layerType);
   ix3536 : nand02 port map ( Y=>nx3535, A0=>outMuls_19_15, A1=>nx5226);
   ix983 : nand02 port map ( Y=>addersInputs_18_0, A0=>nx3538, A1=>nx3540);
   ix3539 : nand02 port map ( Y=>nx3538, A0=>currentPage_18_0, A1=>layerType
   );
   ix3541 : nand02 port map ( Y=>nx3540, A0=>outMuls_18_0, A1=>nx5226);
   ix991 : nand02 port map ( Y=>addersInputs_18_1, A0=>nx3543, A1=>nx3545);
   ix3544 : nand02 port map ( Y=>nx3543, A0=>currentPage_18_1, A1=>layerType
   );
   ix3546 : nand02 port map ( Y=>nx3545, A0=>outMuls_18_1, A1=>nx5226);
   ix999 : nand02 port map ( Y=>addersInputs_18_2, A0=>nx3548, A1=>nx3550);
   ix3549 : nand02 port map ( Y=>nx3548, A0=>currentPage_18_2, A1=>layerType
   );
   ix3551 : nand02 port map ( Y=>nx3550, A0=>outMuls_18_2, A1=>nx5228);
   ix1007 : nand02 port map ( Y=>addersInputs_18_3, A0=>nx3553, A1=>nx3555);
   ix3554 : nand02 port map ( Y=>nx3553, A0=>currentPage_18_3, A1=>layerType
   );
   ix3556 : nand02 port map ( Y=>nx3555, A0=>outMuls_18_3, A1=>nx5228);
   ix1015 : nand02 port map ( Y=>addersInputs_18_4, A0=>nx3558, A1=>nx3560);
   ix3559 : nand02 port map ( Y=>nx3558, A0=>currentPage_18_4, A1=>layerType
   );
   ix3561 : nand02 port map ( Y=>nx3560, A0=>outMuls_18_4, A1=>nx5228);
   ix1023 : nand02 port map ( Y=>addersInputs_18_5, A0=>nx3563, A1=>nx3565);
   ix3564 : nand02 port map ( Y=>nx3563, A0=>currentPage_18_5, A1=>layerType
   );
   ix3566 : nand02 port map ( Y=>nx3565, A0=>outMuls_18_5, A1=>nx5228);
   ix1031 : nand02 port map ( Y=>addersInputs_18_6, A0=>nx3568, A1=>nx3570);
   ix3569 : nand02 port map ( Y=>nx3568, A0=>currentPage_18_6, A1=>layerType
   );
   ix3571 : nand02 port map ( Y=>nx3570, A0=>outMuls_18_6, A1=>nx5228);
   ix1039 : nand02 port map ( Y=>addersInputs_18_7, A0=>nx3573, A1=>nx3575);
   ix3574 : nand02 port map ( Y=>nx3573, A0=>currentPage_18_7, A1=>layerType
   );
   ix3576 : nand02 port map ( Y=>nx3575, A0=>outMuls_18_7, A1=>nx5228);
   ix1047 : nand02 port map ( Y=>addersInputs_18_8, A0=>nx3578, A1=>nx3580);
   ix3579 : nand02 port map ( Y=>nx3578, A0=>currentPage_18_8, A1=>layerType
   );
   ix3581 : nand02 port map ( Y=>nx3580, A0=>outMuls_18_8, A1=>nx5228);
   ix1055 : nand02 port map ( Y=>addersInputs_18_9, A0=>nx3583, A1=>nx3585);
   ix3584 : nand02 port map ( Y=>nx3583, A0=>currentPage_18_9, A1=>layerType
   );
   ix3586 : nand02 port map ( Y=>nx3585, A0=>outMuls_18_9, A1=>nx5230);
   ix1063 : nand02 port map ( Y=>addersInputs_18_10, A0=>nx3588, A1=>nx3590
   );
   ix3589 : nand02 port map ( Y=>nx3588, A0=>currentPage_18_10, A1=>
      layerType);
   ix3591 : nand02 port map ( Y=>nx3590, A0=>outMuls_18_10, A1=>nx5230);
   ix1071 : nand02 port map ( Y=>addersInputs_18_11, A0=>nx3593, A1=>nx3595
   );
   ix3594 : nand02 port map ( Y=>nx3593, A0=>currentPage_18_11, A1=>
      layerType);
   ix3596 : nand02 port map ( Y=>nx3595, A0=>outMuls_18_11, A1=>nx5230);
   ix1079 : nand02 port map ( Y=>addersInputs_18_12, A0=>nx3598, A1=>nx3600
   );
   ix3599 : nand02 port map ( Y=>nx3598, A0=>currentPage_18_12, A1=>
      layerType);
   ix3601 : nand02 port map ( Y=>nx3600, A0=>outMuls_18_12, A1=>nx5230);
   ix1087 : nand02 port map ( Y=>addersInputs_18_13, A0=>nx3603, A1=>nx3605
   );
   ix3604 : nand02 port map ( Y=>nx3603, A0=>currentPage_18_13, A1=>
      layerType);
   ix3606 : nand02 port map ( Y=>nx3605, A0=>outMuls_18_13, A1=>nx5230);
   ix1095 : nand02 port map ( Y=>addersInputs_18_14, A0=>nx3608, A1=>nx3610
   );
   ix3609 : nand02 port map ( Y=>nx3608, A0=>currentPage_18_14, A1=>
      layerType);
   ix3611 : nand02 port map ( Y=>nx3610, A0=>outMuls_18_14, A1=>nx5230);
   ix1103 : nand02 port map ( Y=>addersInputs_18_15, A0=>nx3613, A1=>nx3615
   );
   ix3614 : nand02 port map ( Y=>nx3613, A0=>currentPage_18_15, A1=>
      layerType);
   ix3616 : nand02 port map ( Y=>nx3615, A0=>outMuls_18_15, A1=>nx5230);
   ix1111 : nand02 port map ( Y=>addersInputs_17_0, A0=>nx3618, A1=>nx3620);
   ix3619 : nand02 port map ( Y=>nx3618, A0=>currentPage_17_0, A1=>layerType
   );
   ix3621 : nand02 port map ( Y=>nx3620, A0=>outMuls_17_0, A1=>nx5232);
   ix1119 : nand02 port map ( Y=>addersInputs_17_1, A0=>nx3623, A1=>nx3625);
   ix3624 : nand02 port map ( Y=>nx3623, A0=>currentPage_17_1, A1=>layerType
   );
   ix3626 : nand02 port map ( Y=>nx3625, A0=>outMuls_17_1, A1=>nx5232);
   ix1127 : nand02 port map ( Y=>addersInputs_17_2, A0=>nx3628, A1=>nx3630);
   ix3629 : nand02 port map ( Y=>nx3628, A0=>currentPage_17_2, A1=>layerType
   );
   ix3631 : nand02 port map ( Y=>nx3630, A0=>outMuls_17_2, A1=>nx5232);
   ix1135 : nand02 port map ( Y=>addersInputs_17_3, A0=>nx3633, A1=>nx3635);
   ix3634 : nand02 port map ( Y=>nx3633, A0=>currentPage_17_3, A1=>layerType
   );
   ix3636 : nand02 port map ( Y=>nx3635, A0=>outMuls_17_3, A1=>nx5232);
   ix1143 : nand02 port map ( Y=>addersInputs_17_4, A0=>nx3638, A1=>nx3640);
   ix3639 : nand02 port map ( Y=>nx3638, A0=>currentPage_17_4, A1=>layerType
   );
   ix3641 : nand02 port map ( Y=>nx3640, A0=>outMuls_17_4, A1=>nx5232);
   ix1151 : nand02 port map ( Y=>addersInputs_17_5, A0=>nx3643, A1=>nx3645);
   ix3644 : nand02 port map ( Y=>nx3643, A0=>currentPage_17_5, A1=>layerType
   );
   ix3646 : nand02 port map ( Y=>nx3645, A0=>outMuls_17_5, A1=>nx5232);
   ix1159 : nand02 port map ( Y=>addersInputs_17_6, A0=>nx3648, A1=>nx3650);
   ix3649 : nand02 port map ( Y=>nx3648, A0=>currentPage_17_6, A1=>layerType
   );
   ix3651 : nand02 port map ( Y=>nx3650, A0=>outMuls_17_6, A1=>nx5232);
   ix1167 : nand02 port map ( Y=>addersInputs_17_7, A0=>nx3653, A1=>nx3655);
   ix3654 : nand02 port map ( Y=>nx3653, A0=>currentPage_17_7, A1=>layerType
   );
   ix3656 : nand02 port map ( Y=>nx3655, A0=>outMuls_17_7, A1=>nx5234);
   ix1175 : nand02 port map ( Y=>addersInputs_17_8, A0=>nx3658, A1=>nx3660);
   ix3659 : nand02 port map ( Y=>nx3658, A0=>currentPage_17_8, A1=>layerType
   );
   ix3661 : nand02 port map ( Y=>nx3660, A0=>outMuls_17_8, A1=>nx5234);
   ix1183 : nand02 port map ( Y=>addersInputs_17_9, A0=>nx3663, A1=>nx3665);
   ix3664 : nand02 port map ( Y=>nx3663, A0=>currentPage_17_9, A1=>layerType
   );
   ix3666 : nand02 port map ( Y=>nx3665, A0=>outMuls_17_9, A1=>nx5234);
   ix1191 : nand02 port map ( Y=>addersInputs_17_10, A0=>nx3668, A1=>nx3670
   );
   ix3669 : nand02 port map ( Y=>nx3668, A0=>currentPage_17_10, A1=>
      layerType);
   ix3671 : nand02 port map ( Y=>nx3670, A0=>outMuls_17_10, A1=>nx5234);
   ix1199 : nand02 port map ( Y=>addersInputs_17_11, A0=>nx3673, A1=>nx3675
   );
   ix3674 : nand02 port map ( Y=>nx3673, A0=>currentPage_17_11, A1=>
      layerType);
   ix3676 : nand02 port map ( Y=>nx3675, A0=>outMuls_17_11, A1=>nx5234);
   ix1207 : nand02 port map ( Y=>addersInputs_17_12, A0=>nx3678, A1=>nx3680
   );
   ix3679 : nand02 port map ( Y=>nx3678, A0=>currentPage_17_12, A1=>
      layerType);
   ix3681 : nand02 port map ( Y=>nx3680, A0=>outMuls_17_12, A1=>nx5234);
   ix1215 : nand02 port map ( Y=>addersInputs_17_13, A0=>nx3683, A1=>nx3685
   );
   ix3684 : nand02 port map ( Y=>nx3683, A0=>currentPage_17_13, A1=>
      layerType);
   ix3686 : nand02 port map ( Y=>nx3685, A0=>outMuls_17_13, A1=>nx5234);
   ix1223 : nand02 port map ( Y=>addersInputs_17_14, A0=>nx3688, A1=>nx3690
   );
   ix3689 : nand02 port map ( Y=>nx3688, A0=>currentPage_17_14, A1=>
      layerType);
   ix3691 : nand02 port map ( Y=>nx3690, A0=>outMuls_17_14, A1=>nx5236);
   ix1231 : nand02 port map ( Y=>addersInputs_17_15, A0=>nx3693, A1=>nx3695
   );
   ix3694 : nand02 port map ( Y=>nx3693, A0=>currentPage_17_15, A1=>
      layerType);
   ix3696 : nand02 port map ( Y=>nx3695, A0=>outMuls_17_15, A1=>nx5236);
   ix1239 : nand02 port map ( Y=>addersInputs_16_0, A0=>nx3698, A1=>nx3700);
   ix3699 : nand02 port map ( Y=>nx3698, A0=>currentPage_16_0, A1=>layerType
   );
   ix3701 : nand02 port map ( Y=>nx3700, A0=>outMuls_16_0, A1=>nx5236);
   ix1247 : nand02 port map ( Y=>addersInputs_16_1, A0=>nx3703, A1=>nx3705);
   ix3704 : nand02 port map ( Y=>nx3703, A0=>currentPage_16_1, A1=>layerType
   );
   ix3706 : nand02 port map ( Y=>nx3705, A0=>outMuls_16_1, A1=>nx5236);
   ix1255 : nand02 port map ( Y=>addersInputs_16_2, A0=>nx3708, A1=>nx3710);
   ix3709 : nand02 port map ( Y=>nx3708, A0=>currentPage_16_2, A1=>layerType
   );
   ix3711 : nand02 port map ( Y=>nx3710, A0=>outMuls_16_2, A1=>nx5236);
   ix1263 : nand02 port map ( Y=>addersInputs_16_3, A0=>nx3713, A1=>nx3715);
   ix3714 : nand02 port map ( Y=>nx3713, A0=>currentPage_16_3, A1=>layerType
   );
   ix3716 : nand02 port map ( Y=>nx3715, A0=>outMuls_16_3, A1=>nx5236);
   ix1271 : nand02 port map ( Y=>addersInputs_16_4, A0=>nx3718, A1=>nx3720);
   ix3719 : nand02 port map ( Y=>nx3718, A0=>currentPage_16_4, A1=>layerType
   );
   ix3721 : nand02 port map ( Y=>nx3720, A0=>outMuls_16_4, A1=>nx5236);
   ix1279 : nand02 port map ( Y=>addersInputs_16_5, A0=>nx3723, A1=>nx3725);
   ix3724 : nand02 port map ( Y=>nx3723, A0=>currentPage_16_5, A1=>layerType
   );
   ix3726 : nand02 port map ( Y=>nx3725, A0=>outMuls_16_5, A1=>nx5238);
   ix1287 : nand02 port map ( Y=>addersInputs_16_6, A0=>nx3728, A1=>nx3730);
   ix3729 : nand02 port map ( Y=>nx3728, A0=>currentPage_16_6, A1=>layerType
   );
   ix3731 : nand02 port map ( Y=>nx3730, A0=>outMuls_16_6, A1=>nx5238);
   ix1295 : nand02 port map ( Y=>addersInputs_16_7, A0=>nx3733, A1=>nx3735);
   ix3734 : nand02 port map ( Y=>nx3733, A0=>currentPage_16_7, A1=>layerType
   );
   ix3736 : nand02 port map ( Y=>nx3735, A0=>outMuls_16_7, A1=>nx5238);
   ix1303 : nand02 port map ( Y=>addersInputs_16_8, A0=>nx3738, A1=>nx3740);
   ix3739 : nand02 port map ( Y=>nx3738, A0=>currentPage_16_8, A1=>layerType
   );
   ix3741 : nand02 port map ( Y=>nx3740, A0=>outMuls_16_8, A1=>nx5238);
   ix1311 : nand02 port map ( Y=>addersInputs_16_9, A0=>nx3743, A1=>nx3745);
   ix3744 : nand02 port map ( Y=>nx3743, A0=>currentPage_16_9, A1=>layerType
   );
   ix3746 : nand02 port map ( Y=>nx3745, A0=>outMuls_16_9, A1=>nx5238);
   ix1319 : nand02 port map ( Y=>addersInputs_16_10, A0=>nx3748, A1=>nx3750
   );
   ix3749 : nand02 port map ( Y=>nx3748, A0=>currentPage_16_10, A1=>
      layerType);
   ix3751 : nand02 port map ( Y=>nx3750, A0=>outMuls_16_10, A1=>nx5238);
   ix1327 : nand02 port map ( Y=>addersInputs_16_11, A0=>nx3753, A1=>nx3755
   );
   ix3754 : nand02 port map ( Y=>nx3753, A0=>currentPage_16_11, A1=>
      layerType);
   ix3756 : nand02 port map ( Y=>nx3755, A0=>outMuls_16_11, A1=>nx5238);
   ix1335 : nand02 port map ( Y=>addersInputs_16_12, A0=>nx3758, A1=>nx3760
   );
   ix3759 : nand02 port map ( Y=>nx3758, A0=>currentPage_16_12, A1=>
      layerType);
   ix3761 : nand02 port map ( Y=>nx3760, A0=>outMuls_16_12, A1=>nx5240);
   ix1343 : nand02 port map ( Y=>addersInputs_16_13, A0=>nx3763, A1=>nx3765
   );
   ix3764 : nand02 port map ( Y=>nx3763, A0=>currentPage_16_13, A1=>
      layerType);
   ix3766 : nand02 port map ( Y=>nx3765, A0=>outMuls_16_13, A1=>nx5240);
   ix1351 : nand02 port map ( Y=>addersInputs_16_14, A0=>nx3768, A1=>nx3770
   );
   ix3769 : nand02 port map ( Y=>nx3768, A0=>currentPage_16_14, A1=>
      layerType);
   ix3771 : nand02 port map ( Y=>nx3770, A0=>outMuls_16_14, A1=>nx5240);
   ix1359 : nand02 port map ( Y=>addersInputs_16_15, A0=>nx3773, A1=>nx3775
   );
   ix3774 : nand02 port map ( Y=>nx3773, A0=>currentPage_16_15, A1=>
      layerType);
   ix3776 : nand02 port map ( Y=>nx3775, A0=>outMuls_16_15, A1=>nx5240);
   ix1367 : nand02 port map ( Y=>addersInputs_15_0, A0=>nx3778, A1=>nx3780);
   ix3779 : nand02 port map ( Y=>nx3778, A0=>currentPage_15_0, A1=>layerType
   );
   ix3781 : nand02 port map ( Y=>nx3780, A0=>outMuls_15_0, A1=>nx5240);
   ix1375 : nand02 port map ( Y=>addersInputs_15_1, A0=>nx3783, A1=>nx3785);
   ix3784 : nand02 port map ( Y=>nx3783, A0=>currentPage_15_1, A1=>layerType
   );
   ix3786 : nand02 port map ( Y=>nx3785, A0=>outMuls_15_1, A1=>nx5240);
   ix1383 : nand02 port map ( Y=>addersInputs_15_2, A0=>nx3788, A1=>nx3790);
   ix3789 : nand02 port map ( Y=>nx3788, A0=>currentPage_15_2, A1=>layerType
   );
   ix3791 : nand02 port map ( Y=>nx3790, A0=>outMuls_15_2, A1=>nx5240);
   ix1391 : nand02 port map ( Y=>addersInputs_15_3, A0=>nx3793, A1=>nx3795);
   ix3794 : nand02 port map ( Y=>nx3793, A0=>currentPage_15_3, A1=>layerType
   );
   ix3796 : nand02 port map ( Y=>nx3795, A0=>outMuls_15_3, A1=>nx5242);
   ix1399 : nand02 port map ( Y=>addersInputs_15_4, A0=>nx3798, A1=>nx3800);
   ix3799 : nand02 port map ( Y=>nx3798, A0=>currentPage_15_4, A1=>layerType
   );
   ix3801 : nand02 port map ( Y=>nx3800, A0=>outMuls_15_4, A1=>nx5242);
   ix1407 : nand02 port map ( Y=>addersInputs_15_5, A0=>nx3803, A1=>nx3805);
   ix3804 : nand02 port map ( Y=>nx3803, A0=>currentPage_15_5, A1=>layerType
   );
   ix3806 : nand02 port map ( Y=>nx3805, A0=>outMuls_15_5, A1=>nx5242);
   ix1415 : nand02 port map ( Y=>addersInputs_15_6, A0=>nx3808, A1=>nx3810);
   ix3809 : nand02 port map ( Y=>nx3808, A0=>currentPage_15_6, A1=>layerType
   );
   ix3811 : nand02 port map ( Y=>nx3810, A0=>outMuls_15_6, A1=>nx5242);
   ix1423 : nand02 port map ( Y=>addersInputs_15_7, A0=>nx3813, A1=>nx3815);
   ix3814 : nand02 port map ( Y=>nx3813, A0=>currentPage_15_7, A1=>layerType
   );
   ix3816 : nand02 port map ( Y=>nx3815, A0=>outMuls_15_7, A1=>nx5242);
   ix1431 : nand02 port map ( Y=>addersInputs_15_8, A0=>nx3818, A1=>nx3820);
   ix3819 : nand02 port map ( Y=>nx3818, A0=>currentPage_15_8, A1=>layerType
   );
   ix3821 : nand02 port map ( Y=>nx3820, A0=>outMuls_15_8, A1=>nx5242);
   ix1439 : nand02 port map ( Y=>addersInputs_15_9, A0=>nx3823, A1=>nx3825);
   ix3824 : nand02 port map ( Y=>nx3823, A0=>currentPage_15_9, A1=>layerType
   );
   ix3826 : nand02 port map ( Y=>nx3825, A0=>outMuls_15_9, A1=>nx5242);
   ix1447 : nand02 port map ( Y=>addersInputs_15_10, A0=>nx3828, A1=>nx3830
   );
   ix3829 : nand02 port map ( Y=>nx3828, A0=>currentPage_15_10, A1=>
      layerType);
   ix3831 : nand02 port map ( Y=>nx3830, A0=>outMuls_15_10, A1=>nx5244);
   ix1455 : nand02 port map ( Y=>addersInputs_15_11, A0=>nx3833, A1=>nx3835
   );
   ix3834 : nand02 port map ( Y=>nx3833, A0=>currentPage_15_11, A1=>
      layerType);
   ix3836 : nand02 port map ( Y=>nx3835, A0=>outMuls_15_11, A1=>nx5244);
   ix1463 : nand02 port map ( Y=>addersInputs_15_12, A0=>nx3838, A1=>nx3840
   );
   ix3839 : nand02 port map ( Y=>nx3838, A0=>currentPage_15_12, A1=>
      layerType);
   ix3841 : nand02 port map ( Y=>nx3840, A0=>outMuls_15_12, A1=>nx5244);
   ix1471 : nand02 port map ( Y=>addersInputs_15_13, A0=>nx3843, A1=>nx3845
   );
   ix3844 : nand02 port map ( Y=>nx3843, A0=>currentPage_15_13, A1=>
      layerType);
   ix3846 : nand02 port map ( Y=>nx3845, A0=>outMuls_15_13, A1=>nx5244);
   ix1479 : nand02 port map ( Y=>addersInputs_15_14, A0=>nx3848, A1=>nx3850
   );
   ix3849 : nand02 port map ( Y=>nx3848, A0=>currentPage_15_14, A1=>
      layerType);
   ix3851 : nand02 port map ( Y=>nx3850, A0=>outMuls_15_14, A1=>nx5244);
   ix1487 : nand02 port map ( Y=>addersInputs_15_15, A0=>nx3853, A1=>nx3855
   );
   ix3854 : nand02 port map ( Y=>nx3853, A0=>currentPage_15_15, A1=>
      layerType);
   ix3856 : nand02 port map ( Y=>nx3855, A0=>outMuls_15_15, A1=>nx5244);
   ix1495 : nand02 port map ( Y=>addersInputs_14_0, A0=>nx3858, A1=>nx3860);
   ix3859 : nand02 port map ( Y=>nx3858, A0=>currentPage_14_0, A1=>layerType
   );
   ix3861 : nand02 port map ( Y=>nx3860, A0=>outMuls_14_0, A1=>nx5244);
   ix1503 : nand02 port map ( Y=>addersInputs_14_1, A0=>nx3863, A1=>nx3865);
   ix3864 : nand02 port map ( Y=>nx3863, A0=>currentPage_14_1, A1=>layerType
   );
   ix3866 : nand02 port map ( Y=>nx3865, A0=>outMuls_14_1, A1=>nx5246);
   ix1511 : nand02 port map ( Y=>addersInputs_14_2, A0=>nx3868, A1=>nx3870);
   ix3869 : nand02 port map ( Y=>nx3868, A0=>currentPage_14_2, A1=>layerType
   );
   ix3871 : nand02 port map ( Y=>nx3870, A0=>outMuls_14_2, A1=>nx5246);
   ix1519 : nand02 port map ( Y=>addersInputs_14_3, A0=>nx3873, A1=>nx3875);
   ix3874 : nand02 port map ( Y=>nx3873, A0=>currentPage_14_3, A1=>layerType
   );
   ix3876 : nand02 port map ( Y=>nx3875, A0=>outMuls_14_3, A1=>nx5246);
   ix1527 : nand02 port map ( Y=>addersInputs_14_4, A0=>nx3878, A1=>nx3880);
   ix3879 : nand02 port map ( Y=>nx3878, A0=>currentPage_14_4, A1=>layerType
   );
   ix3881 : nand02 port map ( Y=>nx3880, A0=>outMuls_14_4, A1=>nx5246);
   ix1535 : nand02 port map ( Y=>addersInputs_14_5, A0=>nx3883, A1=>nx3885);
   ix3884 : nand02 port map ( Y=>nx3883, A0=>currentPage_14_5, A1=>layerType
   );
   ix3886 : nand02 port map ( Y=>nx3885, A0=>outMuls_14_5, A1=>nx5246);
   ix1543 : nand02 port map ( Y=>addersInputs_14_6, A0=>nx3888, A1=>nx3890);
   ix3889 : nand02 port map ( Y=>nx3888, A0=>currentPage_14_6, A1=>layerType
   );
   ix3891 : nand02 port map ( Y=>nx3890, A0=>outMuls_14_6, A1=>nx5246);
   ix1551 : nand02 port map ( Y=>addersInputs_14_7, A0=>nx3893, A1=>nx3895);
   ix3894 : nand02 port map ( Y=>nx3893, A0=>currentPage_14_7, A1=>layerType
   );
   ix3896 : nand02 port map ( Y=>nx3895, A0=>outMuls_14_7, A1=>nx5246);
   ix1559 : nand02 port map ( Y=>addersInputs_14_8, A0=>nx3898, A1=>nx3900);
   ix3899 : nand02 port map ( Y=>nx3898, A0=>currentPage_14_8, A1=>layerType
   );
   ix3901 : nand02 port map ( Y=>nx3900, A0=>outMuls_14_8, A1=>nx5248);
   ix1567 : nand02 port map ( Y=>addersInputs_14_9, A0=>nx3903, A1=>nx3905);
   ix3904 : nand02 port map ( Y=>nx3903, A0=>currentPage_14_9, A1=>layerType
   );
   ix3906 : nand02 port map ( Y=>nx3905, A0=>outMuls_14_9, A1=>nx5248);
   ix1575 : nand02 port map ( Y=>addersInputs_14_10, A0=>nx3908, A1=>nx3910
   );
   ix3909 : nand02 port map ( Y=>nx3908, A0=>currentPage_14_10, A1=>
      layerType);
   ix3911 : nand02 port map ( Y=>nx3910, A0=>outMuls_14_10, A1=>nx5248);
   ix1583 : nand02 port map ( Y=>addersInputs_14_11, A0=>nx3913, A1=>nx3915
   );
   ix3914 : nand02 port map ( Y=>nx3913, A0=>currentPage_14_11, A1=>
      layerType);
   ix3916 : nand02 port map ( Y=>nx3915, A0=>outMuls_14_11, A1=>nx5248);
   ix1591 : nand02 port map ( Y=>addersInputs_14_12, A0=>nx3918, A1=>nx3920
   );
   ix3919 : nand02 port map ( Y=>nx3918, A0=>currentPage_14_12, A1=>
      layerType);
   ix3921 : nand02 port map ( Y=>nx3920, A0=>outMuls_14_12, A1=>nx5248);
   ix1599 : nand02 port map ( Y=>addersInputs_14_13, A0=>nx3923, A1=>nx3925
   );
   ix3924 : nand02 port map ( Y=>nx3923, A0=>currentPage_14_13, A1=>
      layerType);
   ix3926 : nand02 port map ( Y=>nx3925, A0=>outMuls_14_13, A1=>nx5248);
   ix1607 : nand02 port map ( Y=>addersInputs_14_14, A0=>nx3928, A1=>nx3930
   );
   ix3929 : nand02 port map ( Y=>nx3928, A0=>currentPage_14_14, A1=>
      layerType);
   ix3931 : nand02 port map ( Y=>nx3930, A0=>outMuls_14_14, A1=>nx5248);
   ix1615 : nand02 port map ( Y=>addersInputs_14_15, A0=>nx3933, A1=>nx3935
   );
   ix3934 : nand02 port map ( Y=>nx3933, A0=>currentPage_14_15, A1=>
      layerType);
   ix3936 : nand02 port map ( Y=>nx3935, A0=>outMuls_14_15, A1=>nx5250);
   ix1623 : nand02 port map ( Y=>addersInputs_13_0, A0=>nx3938, A1=>nx3940);
   ix3939 : nand02 port map ( Y=>nx3938, A0=>currentPage_13_0, A1=>layerType
   );
   ix3941 : nand02 port map ( Y=>nx3940, A0=>outMuls_13_0, A1=>nx5250);
   ix1631 : nand02 port map ( Y=>addersInputs_13_1, A0=>nx3943, A1=>nx3945);
   ix3944 : nand02 port map ( Y=>nx3943, A0=>currentPage_13_1, A1=>layerType
   );
   ix3946 : nand02 port map ( Y=>nx3945, A0=>outMuls_13_1, A1=>nx5250);
   ix1639 : nand02 port map ( Y=>addersInputs_13_2, A0=>nx3948, A1=>nx3950);
   ix3949 : nand02 port map ( Y=>nx3948, A0=>currentPage_13_2, A1=>layerType
   );
   ix3951 : nand02 port map ( Y=>nx3950, A0=>outMuls_13_2, A1=>nx5250);
   ix1647 : nand02 port map ( Y=>addersInputs_13_3, A0=>nx3953, A1=>nx3955);
   ix3954 : nand02 port map ( Y=>nx3953, A0=>currentPage_13_3, A1=>layerType
   );
   ix3956 : nand02 port map ( Y=>nx3955, A0=>outMuls_13_3, A1=>nx5250);
   ix1655 : nand02 port map ( Y=>addersInputs_13_4, A0=>nx3958, A1=>nx3960);
   ix3959 : nand02 port map ( Y=>nx3958, A0=>currentPage_13_4, A1=>layerType
   );
   ix3961 : nand02 port map ( Y=>nx3960, A0=>outMuls_13_4, A1=>nx5250);
   ix1663 : nand02 port map ( Y=>addersInputs_13_5, A0=>nx3963, A1=>nx3965);
   ix3964 : nand02 port map ( Y=>nx3963, A0=>currentPage_13_5, A1=>layerType
   );
   ix3966 : nand02 port map ( Y=>nx3965, A0=>outMuls_13_5, A1=>nx5250);
   ix1671 : nand02 port map ( Y=>addersInputs_13_6, A0=>nx3968, A1=>nx3970);
   ix3969 : nand02 port map ( Y=>nx3968, A0=>currentPage_13_6, A1=>layerType
   );
   ix3971 : nand02 port map ( Y=>nx3970, A0=>outMuls_13_6, A1=>nx5252);
   ix1679 : nand02 port map ( Y=>addersInputs_13_7, A0=>nx3973, A1=>nx3975);
   ix3974 : nand02 port map ( Y=>nx3973, A0=>currentPage_13_7, A1=>layerType
   );
   ix3976 : nand02 port map ( Y=>nx3975, A0=>outMuls_13_7, A1=>nx5252);
   ix1687 : nand02 port map ( Y=>addersInputs_13_8, A0=>nx3978, A1=>nx3980);
   ix3979 : nand02 port map ( Y=>nx3978, A0=>currentPage_13_8, A1=>layerType
   );
   ix3981 : nand02 port map ( Y=>nx3980, A0=>outMuls_13_8, A1=>nx5252);
   ix1695 : nand02 port map ( Y=>addersInputs_13_9, A0=>nx3983, A1=>nx3985);
   ix3984 : nand02 port map ( Y=>nx3983, A0=>currentPage_13_9, A1=>layerType
   );
   ix3986 : nand02 port map ( Y=>nx3985, A0=>outMuls_13_9, A1=>nx5252);
   ix1703 : nand02 port map ( Y=>addersInputs_13_10, A0=>nx3988, A1=>nx3990
   );
   ix3989 : nand02 port map ( Y=>nx3988, A0=>currentPage_13_10, A1=>
      layerType);
   ix3991 : nand02 port map ( Y=>nx3990, A0=>outMuls_13_10, A1=>nx5252);
   ix1711 : nand02 port map ( Y=>addersInputs_13_11, A0=>nx3993, A1=>nx3995
   );
   ix3994 : nand02 port map ( Y=>nx3993, A0=>currentPage_13_11, A1=>
      layerType);
   ix3996 : nand02 port map ( Y=>nx3995, A0=>outMuls_13_11, A1=>nx5252);
   ix1719 : nand02 port map ( Y=>addersInputs_13_12, A0=>nx3998, A1=>nx4000
   );
   ix3999 : nand02 port map ( Y=>nx3998, A0=>currentPage_13_12, A1=>
      layerType);
   ix4001 : nand02 port map ( Y=>nx4000, A0=>outMuls_13_12, A1=>nx5252);
   ix1727 : nand02 port map ( Y=>addersInputs_13_13, A0=>nx4003, A1=>nx4005
   );
   ix4004 : nand02 port map ( Y=>nx4003, A0=>currentPage_13_13, A1=>
      layerType);
   ix4006 : nand02 port map ( Y=>nx4005, A0=>outMuls_13_13, A1=>nx5254);
   ix1735 : nand02 port map ( Y=>addersInputs_13_14, A0=>nx4008, A1=>nx4010
   );
   ix4009 : nand02 port map ( Y=>nx4008, A0=>currentPage_13_14, A1=>
      layerType);
   ix4011 : nand02 port map ( Y=>nx4010, A0=>outMuls_13_14, A1=>nx5254);
   ix1743 : nand02 port map ( Y=>addersInputs_13_15, A0=>nx4013, A1=>nx4015
   );
   ix4014 : nand02 port map ( Y=>nx4013, A0=>currentPage_13_15, A1=>
      layerType);
   ix4016 : nand02 port map ( Y=>nx4015, A0=>outMuls_13_15, A1=>nx5254);
   ix1751 : nand02 port map ( Y=>addersInputs_12_0, A0=>nx4018, A1=>nx4020);
   ix4019 : nand02 port map ( Y=>nx4018, A0=>currentPage_12_0, A1=>layerType
   );
   ix4021 : nand02 port map ( Y=>nx4020, A0=>outMuls_12_0, A1=>nx5254);
   ix1759 : nand02 port map ( Y=>addersInputs_12_1, A0=>nx4023, A1=>nx4025);
   ix4024 : nand02 port map ( Y=>nx4023, A0=>currentPage_12_1, A1=>layerType
   );
   ix4026 : nand02 port map ( Y=>nx4025, A0=>outMuls_12_1, A1=>nx5254);
   ix1767 : nand02 port map ( Y=>addersInputs_12_2, A0=>nx4028, A1=>nx4030);
   ix4029 : nand02 port map ( Y=>nx4028, A0=>currentPage_12_2, A1=>layerType
   );
   ix4031 : nand02 port map ( Y=>nx4030, A0=>outMuls_12_2, A1=>nx5254);
   ix1775 : nand02 port map ( Y=>addersInputs_12_3, A0=>nx4033, A1=>nx4035);
   ix4034 : nand02 port map ( Y=>nx4033, A0=>currentPage_12_3, A1=>layerType
   );
   ix4036 : nand02 port map ( Y=>nx4035, A0=>outMuls_12_3, A1=>nx5254);
   ix1783 : nand02 port map ( Y=>addersInputs_12_4, A0=>nx4038, A1=>nx4040);
   ix4039 : nand02 port map ( Y=>nx4038, A0=>currentPage_12_4, A1=>layerType
   );
   ix4041 : nand02 port map ( Y=>nx4040, A0=>outMuls_12_4, A1=>nx5256);
   ix1791 : nand02 port map ( Y=>addersInputs_12_5, A0=>nx4043, A1=>nx4045);
   ix4044 : nand02 port map ( Y=>nx4043, A0=>currentPage_12_5, A1=>layerType
   );
   ix4046 : nand02 port map ( Y=>nx4045, A0=>outMuls_12_5, A1=>nx5256);
   ix1799 : nand02 port map ( Y=>addersInputs_12_6, A0=>nx4048, A1=>nx4050);
   ix4049 : nand02 port map ( Y=>nx4048, A0=>currentPage_12_6, A1=>layerType
   );
   ix4051 : nand02 port map ( Y=>nx4050, A0=>outMuls_12_6, A1=>nx5256);
   ix1807 : nand02 port map ( Y=>addersInputs_12_7, A0=>nx4053, A1=>nx4055);
   ix4054 : nand02 port map ( Y=>nx4053, A0=>currentPage_12_7, A1=>layerType
   );
   ix4056 : nand02 port map ( Y=>nx4055, A0=>outMuls_12_7, A1=>nx5256);
   ix1815 : nand02 port map ( Y=>addersInputs_12_8, A0=>nx4058, A1=>nx4060);
   ix4059 : nand02 port map ( Y=>nx4058, A0=>currentPage_12_8, A1=>layerType
   );
   ix4061 : nand02 port map ( Y=>nx4060, A0=>outMuls_12_8, A1=>nx5256);
   ix1823 : nand02 port map ( Y=>addersInputs_12_9, A0=>nx4063, A1=>nx4065);
   ix4064 : nand02 port map ( Y=>nx4063, A0=>currentPage_12_9, A1=>layerType
   );
   ix4066 : nand02 port map ( Y=>nx4065, A0=>outMuls_12_9, A1=>nx5256);
   ix1831 : nand02 port map ( Y=>addersInputs_12_10, A0=>nx4068, A1=>nx4070
   );
   ix4069 : nand02 port map ( Y=>nx4068, A0=>currentPage_12_10, A1=>
      layerType);
   ix4071 : nand02 port map ( Y=>nx4070, A0=>outMuls_12_10, A1=>nx5256);
   ix1839 : nand02 port map ( Y=>addersInputs_12_11, A0=>nx4073, A1=>nx4075
   );
   ix4074 : nand02 port map ( Y=>nx4073, A0=>currentPage_12_11, A1=>
      layerType);
   ix4076 : nand02 port map ( Y=>nx4075, A0=>outMuls_12_11, A1=>nx5258);
   ix1847 : nand02 port map ( Y=>addersInputs_12_12, A0=>nx4078, A1=>nx4080
   );
   ix4079 : nand02 port map ( Y=>nx4078, A0=>currentPage_12_12, A1=>
      layerType);
   ix4081 : nand02 port map ( Y=>nx4080, A0=>outMuls_12_12, A1=>nx5258);
   ix1855 : nand02 port map ( Y=>addersInputs_12_13, A0=>nx4083, A1=>nx4085
   );
   ix4084 : nand02 port map ( Y=>nx4083, A0=>currentPage_12_13, A1=>
      layerType);
   ix4086 : nand02 port map ( Y=>nx4085, A0=>outMuls_12_13, A1=>nx5258);
   ix1863 : nand02 port map ( Y=>addersInputs_12_14, A0=>nx4088, A1=>nx4090
   );
   ix4089 : nand02 port map ( Y=>nx4088, A0=>currentPage_12_14, A1=>
      layerType);
   ix4091 : nand02 port map ( Y=>nx4090, A0=>outMuls_12_14, A1=>nx5258);
   ix1871 : nand02 port map ( Y=>addersInputs_12_15, A0=>nx4093, A1=>nx4095
   );
   ix4094 : nand02 port map ( Y=>nx4093, A0=>currentPage_12_15, A1=>
      layerType);
   ix4096 : nand02 port map ( Y=>nx4095, A0=>outMuls_12_15, A1=>nx5258);
   ix1879 : nand02 port map ( Y=>addersInputs_11_0, A0=>nx4098, A1=>nx4100);
   ix4099 : nand02 port map ( Y=>nx4098, A0=>currentPage_11_0, A1=>layerType
   );
   ix4101 : nand02 port map ( Y=>nx4100, A0=>outMuls_11_0, A1=>nx5258);
   ix1887 : nand02 port map ( Y=>addersInputs_11_1, A0=>nx4103, A1=>nx4105);
   ix4104 : nand02 port map ( Y=>nx4103, A0=>currentPage_11_1, A1=>layerType
   );
   ix4106 : nand02 port map ( Y=>nx4105, A0=>outMuls_11_1, A1=>nx5258);
   ix1895 : nand02 port map ( Y=>addersInputs_11_2, A0=>nx4108, A1=>nx4110);
   ix4109 : nand02 port map ( Y=>nx4108, A0=>currentPage_11_2, A1=>layerType
   );
   ix4111 : nand02 port map ( Y=>nx4110, A0=>outMuls_11_2, A1=>nx5260);
   ix1903 : nand02 port map ( Y=>addersInputs_11_3, A0=>nx4113, A1=>nx4115);
   ix4114 : nand02 port map ( Y=>nx4113, A0=>currentPage_11_3, A1=>layerType
   );
   ix4116 : nand02 port map ( Y=>nx4115, A0=>outMuls_11_3, A1=>nx5260);
   ix1911 : nand02 port map ( Y=>addersInputs_11_4, A0=>nx4118, A1=>nx4120);
   ix4119 : nand02 port map ( Y=>nx4118, A0=>currentPage_11_4, A1=>layerType
   );
   ix4121 : nand02 port map ( Y=>nx4120, A0=>outMuls_11_4, A1=>nx5260);
   ix1919 : nand02 port map ( Y=>addersInputs_11_5, A0=>nx4123, A1=>nx4125);
   ix4124 : nand02 port map ( Y=>nx4123, A0=>currentPage_11_5, A1=>layerType
   );
   ix4126 : nand02 port map ( Y=>nx4125, A0=>outMuls_11_5, A1=>nx5260);
   ix1927 : nand02 port map ( Y=>addersInputs_11_6, A0=>nx4128, A1=>nx4130);
   ix4129 : nand02 port map ( Y=>nx4128, A0=>currentPage_11_6, A1=>layerType
   );
   ix4131 : nand02 port map ( Y=>nx4130, A0=>outMuls_11_6, A1=>nx5260);
   ix1935 : nand02 port map ( Y=>addersInputs_11_7, A0=>nx4133, A1=>nx4135);
   ix4134 : nand02 port map ( Y=>nx4133, A0=>currentPage_11_7, A1=>layerType
   );
   ix4136 : nand02 port map ( Y=>nx4135, A0=>outMuls_11_7, A1=>nx5260);
   ix1943 : nand02 port map ( Y=>addersInputs_11_8, A0=>nx4138, A1=>nx4140);
   ix4139 : nand02 port map ( Y=>nx4138, A0=>currentPage_11_8, A1=>layerType
   );
   ix4141 : nand02 port map ( Y=>nx4140, A0=>outMuls_11_8, A1=>nx5260);
   ix1951 : nand02 port map ( Y=>addersInputs_11_9, A0=>nx4143, A1=>nx4145);
   ix4144 : nand02 port map ( Y=>nx4143, A0=>currentPage_11_9, A1=>layerType
   );
   ix4146 : nand02 port map ( Y=>nx4145, A0=>outMuls_11_9, A1=>nx5262);
   ix1959 : nand02 port map ( Y=>addersInputs_11_10, A0=>nx4148, A1=>nx4150
   );
   ix4149 : nand02 port map ( Y=>nx4148, A0=>currentPage_11_10, A1=>
      layerType);
   ix4151 : nand02 port map ( Y=>nx4150, A0=>outMuls_11_10, A1=>nx5262);
   ix1967 : nand02 port map ( Y=>addersInputs_11_11, A0=>nx4153, A1=>nx4155
   );
   ix4154 : nand02 port map ( Y=>nx4153, A0=>currentPage_11_11, A1=>
      layerType);
   ix4156 : nand02 port map ( Y=>nx4155, A0=>outMuls_11_11, A1=>nx5262);
   ix1975 : nand02 port map ( Y=>addersInputs_11_12, A0=>nx4158, A1=>nx4160
   );
   ix4159 : nand02 port map ( Y=>nx4158, A0=>currentPage_11_12, A1=>
      layerType);
   ix4161 : nand02 port map ( Y=>nx4160, A0=>outMuls_11_12, A1=>nx5262);
   ix1983 : nand02 port map ( Y=>addersInputs_11_13, A0=>nx4163, A1=>nx4165
   );
   ix4164 : nand02 port map ( Y=>nx4163, A0=>currentPage_11_13, A1=>
      layerType);
   ix4166 : nand02 port map ( Y=>nx4165, A0=>outMuls_11_13, A1=>nx5262);
   ix1991 : nand02 port map ( Y=>addersInputs_11_14, A0=>nx4168, A1=>nx4170
   );
   ix4169 : nand02 port map ( Y=>nx4168, A0=>currentPage_11_14, A1=>
      layerType);
   ix4171 : nand02 port map ( Y=>nx4170, A0=>outMuls_11_14, A1=>nx5262);
   ix1999 : nand02 port map ( Y=>addersInputs_11_15, A0=>nx4173, A1=>nx4175
   );
   ix4174 : nand02 port map ( Y=>nx4173, A0=>currentPage_11_15, A1=>
      layerType);
   ix4176 : nand02 port map ( Y=>nx4175, A0=>outMuls_11_15, A1=>nx5262);
   ix2007 : nand02 port map ( Y=>addersInputs_10_0, A0=>nx4178, A1=>nx4180);
   ix4179 : nand02 port map ( Y=>nx4178, A0=>currentPage_10_0, A1=>layerType
   );
   ix4181 : nand02 port map ( Y=>nx4180, A0=>outMuls_10_0, A1=>nx5264);
   ix2015 : nand02 port map ( Y=>addersInputs_10_1, A0=>nx4183, A1=>nx4185);
   ix4184 : nand02 port map ( Y=>nx4183, A0=>currentPage_10_1, A1=>layerType
   );
   ix4186 : nand02 port map ( Y=>nx4185, A0=>outMuls_10_1, A1=>nx5264);
   ix2023 : nand02 port map ( Y=>addersInputs_10_2, A0=>nx4188, A1=>nx4190);
   ix4189 : nand02 port map ( Y=>nx4188, A0=>currentPage_10_2, A1=>layerType
   );
   ix4191 : nand02 port map ( Y=>nx4190, A0=>outMuls_10_2, A1=>nx5264);
   ix2031 : nand02 port map ( Y=>addersInputs_10_3, A0=>nx4193, A1=>nx4195);
   ix4194 : nand02 port map ( Y=>nx4193, A0=>currentPage_10_3, A1=>layerType
   );
   ix4196 : nand02 port map ( Y=>nx4195, A0=>outMuls_10_3, A1=>nx5264);
   ix2039 : nand02 port map ( Y=>addersInputs_10_4, A0=>nx4198, A1=>nx4200);
   ix4199 : nand02 port map ( Y=>nx4198, A0=>currentPage_10_4, A1=>layerType
   );
   ix4201 : nand02 port map ( Y=>nx4200, A0=>outMuls_10_4, A1=>nx5264);
   ix2047 : nand02 port map ( Y=>addersInputs_10_5, A0=>nx4203, A1=>nx4205);
   ix4204 : nand02 port map ( Y=>nx4203, A0=>currentPage_10_5, A1=>layerType
   );
   ix4206 : nand02 port map ( Y=>nx4205, A0=>outMuls_10_5, A1=>nx5264);
   ix2055 : nand02 port map ( Y=>addersInputs_10_6, A0=>nx4208, A1=>nx4210);
   ix4209 : nand02 port map ( Y=>nx4208, A0=>currentPage_10_6, A1=>layerType
   );
   ix4211 : nand02 port map ( Y=>nx4210, A0=>outMuls_10_6, A1=>nx5264);
   ix2063 : nand02 port map ( Y=>addersInputs_10_7, A0=>nx4213, A1=>nx4215);
   ix4214 : nand02 port map ( Y=>nx4213, A0=>currentPage_10_7, A1=>layerType
   );
   ix4216 : nand02 port map ( Y=>nx4215, A0=>outMuls_10_7, A1=>nx5266);
   ix2071 : nand02 port map ( Y=>addersInputs_10_8, A0=>nx4218, A1=>nx4220);
   ix4219 : nand02 port map ( Y=>nx4218, A0=>currentPage_10_8, A1=>layerType
   );
   ix4221 : nand02 port map ( Y=>nx4220, A0=>outMuls_10_8, A1=>nx5266);
   ix2079 : nand02 port map ( Y=>addersInputs_10_9, A0=>nx4223, A1=>nx4225);
   ix4224 : nand02 port map ( Y=>nx4223, A0=>currentPage_10_9, A1=>layerType
   );
   ix4226 : nand02 port map ( Y=>nx4225, A0=>outMuls_10_9, A1=>nx5266);
   ix2087 : nand02 port map ( Y=>addersInputs_10_10, A0=>nx4228, A1=>nx4230
   );
   ix4229 : nand02 port map ( Y=>nx4228, A0=>currentPage_10_10, A1=>
      layerType);
   ix4231 : nand02 port map ( Y=>nx4230, A0=>outMuls_10_10, A1=>nx5266);
   ix2095 : nand02 port map ( Y=>addersInputs_10_11, A0=>nx4233, A1=>nx4235
   );
   ix4234 : nand02 port map ( Y=>nx4233, A0=>currentPage_10_11, A1=>
      layerType);
   ix4236 : nand02 port map ( Y=>nx4235, A0=>outMuls_10_11, A1=>nx5266);
   ix2103 : nand02 port map ( Y=>addersInputs_10_12, A0=>nx4238, A1=>nx4240
   );
   ix4239 : nand02 port map ( Y=>nx4238, A0=>currentPage_10_12, A1=>
      layerType);
   ix4241 : nand02 port map ( Y=>nx4240, A0=>outMuls_10_12, A1=>nx5266);
   ix2111 : nand02 port map ( Y=>addersInputs_10_13, A0=>nx4243, A1=>nx4245
   );
   ix4244 : nand02 port map ( Y=>nx4243, A0=>currentPage_10_13, A1=>
      layerType);
   ix4246 : nand02 port map ( Y=>nx4245, A0=>outMuls_10_13, A1=>nx5266);
   ix2119 : nand02 port map ( Y=>addersInputs_10_14, A0=>nx4248, A1=>nx4250
   );
   ix4249 : nand02 port map ( Y=>nx4248, A0=>currentPage_10_14, A1=>
      layerType);
   ix4251 : nand02 port map ( Y=>nx4250, A0=>outMuls_10_14, A1=>nx5268);
   ix2127 : nand02 port map ( Y=>addersInputs_10_15, A0=>nx4253, A1=>nx4255
   );
   ix4254 : nand02 port map ( Y=>nx4253, A0=>currentPage_10_15, A1=>
      layerType);
   ix4256 : nand02 port map ( Y=>nx4255, A0=>outMuls_10_15, A1=>nx5268);
   ix2135 : nand02 port map ( Y=>addersInputs_9_0, A0=>nx4258, A1=>nx4260);
   ix4259 : nand02 port map ( Y=>nx4258, A0=>currentPage_9_0, A1=>layerType
   );
   ix4261 : nand02 port map ( Y=>nx4260, A0=>outMuls_9_0, A1=>nx5268);
   ix2143 : nand02 port map ( Y=>addersInputs_9_1, A0=>nx4263, A1=>nx4265);
   ix4264 : nand02 port map ( Y=>nx4263, A0=>currentPage_9_1, A1=>layerType
   );
   ix4266 : nand02 port map ( Y=>nx4265, A0=>outMuls_9_1, A1=>nx5268);
   ix2151 : nand02 port map ( Y=>addersInputs_9_2, A0=>nx4268, A1=>nx4270);
   ix4269 : nand02 port map ( Y=>nx4268, A0=>currentPage_9_2, A1=>layerType
   );
   ix4271 : nand02 port map ( Y=>nx4270, A0=>outMuls_9_2, A1=>nx5268);
   ix2159 : nand02 port map ( Y=>addersInputs_9_3, A0=>nx4273, A1=>nx4275);
   ix4274 : nand02 port map ( Y=>nx4273, A0=>currentPage_9_3, A1=>layerType
   );
   ix4276 : nand02 port map ( Y=>nx4275, A0=>outMuls_9_3, A1=>nx5268);
   ix2167 : nand02 port map ( Y=>addersInputs_9_4, A0=>nx4278, A1=>nx4280);
   ix4279 : nand02 port map ( Y=>nx4278, A0=>currentPage_9_4, A1=>layerType
   );
   ix4281 : nand02 port map ( Y=>nx4280, A0=>outMuls_9_4, A1=>nx5268);
   ix2175 : nand02 port map ( Y=>addersInputs_9_5, A0=>nx4283, A1=>nx4285);
   ix4284 : nand02 port map ( Y=>nx4283, A0=>currentPage_9_5, A1=>layerType
   );
   ix4286 : nand02 port map ( Y=>nx4285, A0=>outMuls_9_5, A1=>nx5270);
   ix2183 : nand02 port map ( Y=>addersInputs_9_6, A0=>nx4288, A1=>nx4290);
   ix4289 : nand02 port map ( Y=>nx4288, A0=>currentPage_9_6, A1=>layerType
   );
   ix4291 : nand02 port map ( Y=>nx4290, A0=>outMuls_9_6, A1=>nx5270);
   ix2191 : nand02 port map ( Y=>addersInputs_9_7, A0=>nx4293, A1=>nx4295);
   ix4294 : nand02 port map ( Y=>nx4293, A0=>currentPage_9_7, A1=>layerType
   );
   ix4296 : nand02 port map ( Y=>nx4295, A0=>outMuls_9_7, A1=>nx5270);
   ix2199 : nand02 port map ( Y=>addersInputs_9_8, A0=>nx4298, A1=>nx4300);
   ix4299 : nand02 port map ( Y=>nx4298, A0=>currentPage_9_8, A1=>layerType
   );
   ix4301 : nand02 port map ( Y=>nx4300, A0=>outMuls_9_8, A1=>nx5270);
   ix2207 : nand02 port map ( Y=>addersInputs_9_9, A0=>nx4303, A1=>nx4305);
   ix4304 : nand02 port map ( Y=>nx4303, A0=>currentPage_9_9, A1=>layerType
   );
   ix4306 : nand02 port map ( Y=>nx4305, A0=>outMuls_9_9, A1=>nx5270);
   ix2215 : nand02 port map ( Y=>addersInputs_9_10, A0=>nx4308, A1=>nx4310);
   ix4309 : nand02 port map ( Y=>nx4308, A0=>currentPage_9_10, A1=>layerType
   );
   ix4311 : nand02 port map ( Y=>nx4310, A0=>outMuls_9_10, A1=>nx5270);
   ix2223 : nand02 port map ( Y=>addersInputs_9_11, A0=>nx4313, A1=>nx4315);
   ix4314 : nand02 port map ( Y=>nx4313, A0=>currentPage_9_11, A1=>layerType
   );
   ix4316 : nand02 port map ( Y=>nx4315, A0=>outMuls_9_11, A1=>nx5270);
   ix2231 : nand02 port map ( Y=>addersInputs_9_12, A0=>nx4318, A1=>nx4320);
   ix4319 : nand02 port map ( Y=>nx4318, A0=>currentPage_9_12, A1=>layerType
   );
   ix4321 : nand02 port map ( Y=>nx4320, A0=>outMuls_9_12, A1=>nx5272);
   ix2239 : nand02 port map ( Y=>addersInputs_9_13, A0=>nx4323, A1=>nx4325);
   ix4324 : nand02 port map ( Y=>nx4323, A0=>currentPage_9_13, A1=>layerType
   );
   ix4326 : nand02 port map ( Y=>nx4325, A0=>outMuls_9_13, A1=>nx5272);
   ix2247 : nand02 port map ( Y=>addersInputs_9_14, A0=>nx4328, A1=>nx4330);
   ix4329 : nand02 port map ( Y=>nx4328, A0=>currentPage_9_14, A1=>layerType
   );
   ix4331 : nand02 port map ( Y=>nx4330, A0=>outMuls_9_14, A1=>nx5272);
   ix2255 : nand02 port map ( Y=>addersInputs_9_15, A0=>nx4333, A1=>nx4335);
   ix4334 : nand02 port map ( Y=>nx4333, A0=>currentPage_9_15, A1=>layerType
   );
   ix4336 : nand02 port map ( Y=>nx4335, A0=>outMuls_9_15, A1=>nx5272);
   ix2263 : nand02 port map ( Y=>addersInputs_8_0, A0=>nx4338, A1=>nx4340);
   ix4339 : nand02 port map ( Y=>nx4338, A0=>currentPage_8_0, A1=>layerType
   );
   ix4341 : nand02 port map ( Y=>nx4340, A0=>outMuls_8_0, A1=>nx5272);
   ix2271 : nand02 port map ( Y=>addersInputs_8_1, A0=>nx4343, A1=>nx4345);
   ix4344 : nand02 port map ( Y=>nx4343, A0=>currentPage_8_1, A1=>layerType
   );
   ix4346 : nand02 port map ( Y=>nx4345, A0=>outMuls_8_1, A1=>nx5272);
   ix2279 : nand02 port map ( Y=>addersInputs_8_2, A0=>nx4348, A1=>nx4350);
   ix4349 : nand02 port map ( Y=>nx4348, A0=>currentPage_8_2, A1=>layerType
   );
   ix4351 : nand02 port map ( Y=>nx4350, A0=>outMuls_8_2, A1=>nx5272);
   ix2287 : nand02 port map ( Y=>addersInputs_8_3, A0=>nx4353, A1=>nx4355);
   ix4354 : nand02 port map ( Y=>nx4353, A0=>currentPage_8_3, A1=>layerType
   );
   ix4356 : nand02 port map ( Y=>nx4355, A0=>outMuls_8_3, A1=>nx5274);
   ix2295 : nand02 port map ( Y=>addersInputs_8_4, A0=>nx4358, A1=>nx4360);
   ix4359 : nand02 port map ( Y=>nx4358, A0=>currentPage_8_4, A1=>layerType
   );
   ix4361 : nand02 port map ( Y=>nx4360, A0=>outMuls_8_4, A1=>nx5274);
   ix2303 : nand02 port map ( Y=>addersInputs_8_5, A0=>nx4363, A1=>nx4365);
   ix4364 : nand02 port map ( Y=>nx4363, A0=>currentPage_8_5, A1=>layerType
   );
   ix4366 : nand02 port map ( Y=>nx4365, A0=>outMuls_8_5, A1=>nx5274);
   ix2311 : nand02 port map ( Y=>addersInputs_8_6, A0=>nx4368, A1=>nx4370);
   ix4369 : nand02 port map ( Y=>nx4368, A0=>currentPage_8_6, A1=>layerType
   );
   ix4371 : nand02 port map ( Y=>nx4370, A0=>outMuls_8_6, A1=>nx5274);
   ix2319 : nand02 port map ( Y=>addersInputs_8_7, A0=>nx4373, A1=>nx4375);
   ix4374 : nand02 port map ( Y=>nx4373, A0=>currentPage_8_7, A1=>layerType
   );
   ix4376 : nand02 port map ( Y=>nx4375, A0=>outMuls_8_7, A1=>nx5274);
   ix2327 : nand02 port map ( Y=>addersInputs_8_8, A0=>nx4378, A1=>nx4380);
   ix4379 : nand02 port map ( Y=>nx4378, A0=>currentPage_8_8, A1=>layerType
   );
   ix4381 : nand02 port map ( Y=>nx4380, A0=>outMuls_8_8, A1=>nx5274);
   ix2335 : nand02 port map ( Y=>addersInputs_8_9, A0=>nx4383, A1=>nx4385);
   ix4384 : nand02 port map ( Y=>nx4383, A0=>currentPage_8_9, A1=>layerType
   );
   ix4386 : nand02 port map ( Y=>nx4385, A0=>outMuls_8_9, A1=>nx5274);
   ix2343 : nand02 port map ( Y=>addersInputs_8_10, A0=>nx4388, A1=>nx4390);
   ix4389 : nand02 port map ( Y=>nx4388, A0=>currentPage_8_10, A1=>layerType
   );
   ix4391 : nand02 port map ( Y=>nx4390, A0=>outMuls_8_10, A1=>nx5276);
   ix2351 : nand02 port map ( Y=>addersInputs_8_11, A0=>nx4393, A1=>nx4395);
   ix4394 : nand02 port map ( Y=>nx4393, A0=>currentPage_8_11, A1=>layerType
   );
   ix4396 : nand02 port map ( Y=>nx4395, A0=>outMuls_8_11, A1=>nx5276);
   ix2359 : nand02 port map ( Y=>addersInputs_8_12, A0=>nx4398, A1=>nx4400);
   ix4399 : nand02 port map ( Y=>nx4398, A0=>currentPage_8_12, A1=>layerType
   );
   ix4401 : nand02 port map ( Y=>nx4400, A0=>outMuls_8_12, A1=>nx5276);
   ix2367 : nand02 port map ( Y=>addersInputs_8_13, A0=>nx4403, A1=>nx4405);
   ix4404 : nand02 port map ( Y=>nx4403, A0=>currentPage_8_13, A1=>layerType
   );
   ix4406 : nand02 port map ( Y=>nx4405, A0=>outMuls_8_13, A1=>nx5276);
   ix2375 : nand02 port map ( Y=>addersInputs_8_14, A0=>nx4408, A1=>nx4410);
   ix4409 : nand02 port map ( Y=>nx4408, A0=>currentPage_8_14, A1=>layerType
   );
   ix4411 : nand02 port map ( Y=>nx4410, A0=>outMuls_8_14, A1=>nx5276);
   ix2383 : nand02 port map ( Y=>addersInputs_8_15, A0=>nx4413, A1=>nx4415);
   ix4414 : nand02 port map ( Y=>nx4413, A0=>currentPage_8_15, A1=>layerType
   );
   ix4416 : nand02 port map ( Y=>nx4415, A0=>outMuls_8_15, A1=>nx5276);
   ix2391 : nand02 port map ( Y=>addersInputs_7_0, A0=>nx4418, A1=>nx4420);
   ix4419 : nand02 port map ( Y=>nx4418, A0=>currentPage_7_0, A1=>layerType
   );
   ix4421 : nand02 port map ( Y=>nx4420, A0=>outMuls_7_0, A1=>nx5276);
   ix2399 : nand02 port map ( Y=>addersInputs_7_1, A0=>nx4423, A1=>nx4425);
   ix4424 : nand02 port map ( Y=>nx4423, A0=>currentPage_7_1, A1=>layerType
   );
   ix4426 : nand02 port map ( Y=>nx4425, A0=>outMuls_7_1, A1=>nx5278);
   ix2407 : nand02 port map ( Y=>addersInputs_7_2, A0=>nx4428, A1=>nx4430);
   ix4429 : nand02 port map ( Y=>nx4428, A0=>currentPage_7_2, A1=>layerType
   );
   ix4431 : nand02 port map ( Y=>nx4430, A0=>outMuls_7_2, A1=>nx5278);
   ix2415 : nand02 port map ( Y=>addersInputs_7_3, A0=>nx4433, A1=>nx4435);
   ix4434 : nand02 port map ( Y=>nx4433, A0=>currentPage_7_3, A1=>layerType
   );
   ix4436 : nand02 port map ( Y=>nx4435, A0=>outMuls_7_3, A1=>nx5278);
   ix2423 : nand02 port map ( Y=>addersInputs_7_4, A0=>nx4438, A1=>nx4440);
   ix4439 : nand02 port map ( Y=>nx4438, A0=>currentPage_7_4, A1=>layerType
   );
   ix4441 : nand02 port map ( Y=>nx4440, A0=>outMuls_7_4, A1=>nx5278);
   ix2431 : nand02 port map ( Y=>addersInputs_7_5, A0=>nx4443, A1=>nx4445);
   ix4444 : nand02 port map ( Y=>nx4443, A0=>currentPage_7_5, A1=>layerType
   );
   ix4446 : nand02 port map ( Y=>nx4445, A0=>outMuls_7_5, A1=>nx5278);
   ix2439 : nand02 port map ( Y=>addersInputs_7_6, A0=>nx4448, A1=>nx4450);
   ix4449 : nand02 port map ( Y=>nx4448, A0=>currentPage_7_6, A1=>layerType
   );
   ix4451 : nand02 port map ( Y=>nx4450, A0=>outMuls_7_6, A1=>nx5278);
   ix2447 : nand02 port map ( Y=>addersInputs_7_7, A0=>nx4453, A1=>nx4455);
   ix4454 : nand02 port map ( Y=>nx4453, A0=>currentPage_7_7, A1=>layerType
   );
   ix4456 : nand02 port map ( Y=>nx4455, A0=>outMuls_7_7, A1=>nx5278);
   ix2455 : nand02 port map ( Y=>addersInputs_7_8, A0=>nx4458, A1=>nx4460);
   ix4459 : nand02 port map ( Y=>nx4458, A0=>currentPage_7_8, A1=>layerType
   );
   ix4461 : nand02 port map ( Y=>nx4460, A0=>outMuls_7_8, A1=>nx5280);
   ix2463 : nand02 port map ( Y=>addersInputs_7_9, A0=>nx4463, A1=>nx4465);
   ix4464 : nand02 port map ( Y=>nx4463, A0=>currentPage_7_9, A1=>layerType
   );
   ix4466 : nand02 port map ( Y=>nx4465, A0=>outMuls_7_9, A1=>nx5280);
   ix2471 : nand02 port map ( Y=>addersInputs_7_10, A0=>nx4468, A1=>nx4470);
   ix4469 : nand02 port map ( Y=>nx4468, A0=>currentPage_7_10, A1=>layerType
   );
   ix4471 : nand02 port map ( Y=>nx4470, A0=>outMuls_7_10, A1=>nx5280);
   ix2479 : nand02 port map ( Y=>addersInputs_7_11, A0=>nx4473, A1=>nx4475);
   ix4474 : nand02 port map ( Y=>nx4473, A0=>currentPage_7_11, A1=>layerType
   );
   ix4476 : nand02 port map ( Y=>nx4475, A0=>outMuls_7_11, A1=>nx5280);
   ix2487 : nand02 port map ( Y=>addersInputs_7_12, A0=>nx4478, A1=>nx4480);
   ix4479 : nand02 port map ( Y=>nx4478, A0=>currentPage_7_12, A1=>layerType
   );
   ix4481 : nand02 port map ( Y=>nx4480, A0=>outMuls_7_12, A1=>nx5280);
   ix2495 : nand02 port map ( Y=>addersInputs_7_13, A0=>nx4483, A1=>nx4485);
   ix4484 : nand02 port map ( Y=>nx4483, A0=>currentPage_7_13, A1=>layerType
   );
   ix4486 : nand02 port map ( Y=>nx4485, A0=>outMuls_7_13, A1=>nx5280);
   ix2503 : nand02 port map ( Y=>addersInputs_7_14, A0=>nx4488, A1=>nx4490);
   ix4489 : nand02 port map ( Y=>nx4488, A0=>currentPage_7_14, A1=>layerType
   );
   ix4491 : nand02 port map ( Y=>nx4490, A0=>outMuls_7_14, A1=>nx5280);
   ix2511 : nand02 port map ( Y=>addersInputs_7_15, A0=>nx4493, A1=>nx4495);
   ix4494 : nand02 port map ( Y=>nx4493, A0=>currentPage_7_15, A1=>layerType
   );
   ix4496 : nand02 port map ( Y=>nx4495, A0=>outMuls_7_15, A1=>nx5282);
   ix2519 : nand02 port map ( Y=>addersInputs_6_0, A0=>nx4498, A1=>nx4500);
   ix4499 : nand02 port map ( Y=>nx4498, A0=>currentPage_6_0, A1=>layerType
   );
   ix4501 : nand02 port map ( Y=>nx4500, A0=>outMuls_6_0, A1=>nx5282);
   ix2527 : nand02 port map ( Y=>addersInputs_6_1, A0=>nx4503, A1=>nx4505);
   ix4504 : nand02 port map ( Y=>nx4503, A0=>currentPage_6_1, A1=>layerType
   );
   ix4506 : nand02 port map ( Y=>nx4505, A0=>outMuls_6_1, A1=>nx5282);
   ix2535 : nand02 port map ( Y=>addersInputs_6_2, A0=>nx4508, A1=>nx4510);
   ix4509 : nand02 port map ( Y=>nx4508, A0=>currentPage_6_2, A1=>layerType
   );
   ix4511 : nand02 port map ( Y=>nx4510, A0=>outMuls_6_2, A1=>nx5282);
   ix2543 : nand02 port map ( Y=>addersInputs_6_3, A0=>nx4513, A1=>nx4515);
   ix4514 : nand02 port map ( Y=>nx4513, A0=>currentPage_6_3, A1=>layerType
   );
   ix4516 : nand02 port map ( Y=>nx4515, A0=>outMuls_6_3, A1=>nx5282);
   ix2551 : nand02 port map ( Y=>addersInputs_6_4, A0=>nx4518, A1=>nx4520);
   ix4519 : nand02 port map ( Y=>nx4518, A0=>currentPage_6_4, A1=>layerType
   );
   ix4521 : nand02 port map ( Y=>nx4520, A0=>outMuls_6_4, A1=>nx5282);
   ix2559 : nand02 port map ( Y=>addersInputs_6_5, A0=>nx4523, A1=>nx4525);
   ix4524 : nand02 port map ( Y=>nx4523, A0=>currentPage_6_5, A1=>layerType
   );
   ix4526 : nand02 port map ( Y=>nx4525, A0=>outMuls_6_5, A1=>nx5282);
   ix2567 : nand02 port map ( Y=>addersInputs_6_6, A0=>nx4528, A1=>nx4530);
   ix4529 : nand02 port map ( Y=>nx4528, A0=>currentPage_6_6, A1=>layerType
   );
   ix4531 : nand02 port map ( Y=>nx4530, A0=>outMuls_6_6, A1=>nx5284);
   ix2575 : nand02 port map ( Y=>addersInputs_6_7, A0=>nx4533, A1=>nx4535);
   ix4534 : nand02 port map ( Y=>nx4533, A0=>currentPage_6_7, A1=>layerType
   );
   ix4536 : nand02 port map ( Y=>nx4535, A0=>outMuls_6_7, A1=>nx5284);
   ix2583 : nand02 port map ( Y=>addersInputs_6_8, A0=>nx4538, A1=>nx4540);
   ix4539 : nand02 port map ( Y=>nx4538, A0=>currentPage_6_8, A1=>layerType
   );
   ix4541 : nand02 port map ( Y=>nx4540, A0=>outMuls_6_8, A1=>nx5284);
   ix2591 : nand02 port map ( Y=>addersInputs_6_9, A0=>nx4543, A1=>nx4545);
   ix4544 : nand02 port map ( Y=>nx4543, A0=>currentPage_6_9, A1=>layerType
   );
   ix4546 : nand02 port map ( Y=>nx4545, A0=>outMuls_6_9, A1=>nx5284);
   ix2599 : nand02 port map ( Y=>addersInputs_6_10, A0=>nx4548, A1=>nx4550);
   ix4549 : nand02 port map ( Y=>nx4548, A0=>currentPage_6_10, A1=>layerType
   );
   ix4551 : nand02 port map ( Y=>nx4550, A0=>outMuls_6_10, A1=>nx5284);
   ix2607 : nand02 port map ( Y=>addersInputs_6_11, A0=>nx4553, A1=>nx4555);
   ix4554 : nand02 port map ( Y=>nx4553, A0=>currentPage_6_11, A1=>layerType
   );
   ix4556 : nand02 port map ( Y=>nx4555, A0=>outMuls_6_11, A1=>nx5284);
   ix2615 : nand02 port map ( Y=>addersInputs_6_12, A0=>nx4558, A1=>nx4560);
   ix4559 : nand02 port map ( Y=>nx4558, A0=>currentPage_6_12, A1=>layerType
   );
   ix4561 : nand02 port map ( Y=>nx4560, A0=>outMuls_6_12, A1=>nx5284);
   ix2623 : nand02 port map ( Y=>addersInputs_6_13, A0=>nx4563, A1=>nx4565);
   ix4564 : nand02 port map ( Y=>nx4563, A0=>currentPage_6_13, A1=>layerType
   );
   ix4566 : nand02 port map ( Y=>nx4565, A0=>outMuls_6_13, A1=>nx5286);
   ix2631 : nand02 port map ( Y=>addersInputs_6_14, A0=>nx4568, A1=>nx4570);
   ix4569 : nand02 port map ( Y=>nx4568, A0=>currentPage_6_14, A1=>layerType
   );
   ix4571 : nand02 port map ( Y=>nx4570, A0=>outMuls_6_14, A1=>nx5286);
   ix2639 : nand02 port map ( Y=>addersInputs_6_15, A0=>nx4573, A1=>nx4575);
   ix4574 : nand02 port map ( Y=>nx4573, A0=>currentPage_6_15, A1=>layerType
   );
   ix4576 : nand02 port map ( Y=>nx4575, A0=>outMuls_6_15, A1=>nx5286);
   ix2647 : nand02 port map ( Y=>addersInputs_5_0, A0=>nx4578, A1=>nx4580);
   ix4579 : nand02 port map ( Y=>nx4578, A0=>currentPage_5_0, A1=>layerType
   );
   ix4581 : nand02 port map ( Y=>nx4580, A0=>outMuls_5_0, A1=>nx5286);
   ix2655 : nand02 port map ( Y=>addersInputs_5_1, A0=>nx4583, A1=>nx4585);
   ix4584 : nand02 port map ( Y=>nx4583, A0=>currentPage_5_1, A1=>layerType
   );
   ix4586 : nand02 port map ( Y=>nx4585, A0=>outMuls_5_1, A1=>nx5286);
   ix2663 : nand02 port map ( Y=>addersInputs_5_2, A0=>nx4588, A1=>nx4590);
   ix4589 : nand02 port map ( Y=>nx4588, A0=>currentPage_5_2, A1=>layerType
   );
   ix4591 : nand02 port map ( Y=>nx4590, A0=>outMuls_5_2, A1=>nx5286);
   ix2671 : nand02 port map ( Y=>addersInputs_5_3, A0=>nx4593, A1=>nx4595);
   ix4594 : nand02 port map ( Y=>nx4593, A0=>currentPage_5_3, A1=>layerType
   );
   ix4596 : nand02 port map ( Y=>nx4595, A0=>outMuls_5_3, A1=>nx5286);
   ix2679 : nand02 port map ( Y=>addersInputs_5_4, A0=>nx4598, A1=>nx4600);
   ix4599 : nand02 port map ( Y=>nx4598, A0=>currentPage_5_4, A1=>layerType
   );
   ix4601 : nand02 port map ( Y=>nx4600, A0=>outMuls_5_4, A1=>nx5288);
   ix2687 : nand02 port map ( Y=>addersInputs_5_5, A0=>nx4603, A1=>nx4605);
   ix4604 : nand02 port map ( Y=>nx4603, A0=>currentPage_5_5, A1=>layerType
   );
   ix4606 : nand02 port map ( Y=>nx4605, A0=>outMuls_5_5, A1=>nx5288);
   ix2695 : nand02 port map ( Y=>addersInputs_5_6, A0=>nx4608, A1=>nx4610);
   ix4609 : nand02 port map ( Y=>nx4608, A0=>currentPage_5_6, A1=>layerType
   );
   ix4611 : nand02 port map ( Y=>nx4610, A0=>outMuls_5_6, A1=>nx5288);
   ix2703 : nand02 port map ( Y=>addersInputs_5_7, A0=>nx4613, A1=>nx4615);
   ix4614 : nand02 port map ( Y=>nx4613, A0=>currentPage_5_7, A1=>layerType
   );
   ix4616 : nand02 port map ( Y=>nx4615, A0=>outMuls_5_7, A1=>nx5288);
   ix2711 : nand02 port map ( Y=>addersInputs_5_8, A0=>nx4618, A1=>nx4620);
   ix4619 : nand02 port map ( Y=>nx4618, A0=>currentPage_5_8, A1=>layerType
   );
   ix4621 : nand02 port map ( Y=>nx4620, A0=>outMuls_5_8, A1=>nx5288);
   ix2719 : nand02 port map ( Y=>addersInputs_5_9, A0=>nx4623, A1=>nx4625);
   ix4624 : nand02 port map ( Y=>nx4623, A0=>currentPage_5_9, A1=>layerType
   );
   ix4626 : nand02 port map ( Y=>nx4625, A0=>outMuls_5_9, A1=>nx5288);
   ix2727 : nand02 port map ( Y=>addersInputs_5_10, A0=>nx4628, A1=>nx4630);
   ix4629 : nand02 port map ( Y=>nx4628, A0=>currentPage_5_10, A1=>layerType
   );
   ix4631 : nand02 port map ( Y=>nx4630, A0=>outMuls_5_10, A1=>nx5288);
   ix2735 : nand02 port map ( Y=>addersInputs_5_11, A0=>nx4633, A1=>nx4635);
   ix4634 : nand02 port map ( Y=>nx4633, A0=>currentPage_5_11, A1=>layerType
   );
   ix4636 : nand02 port map ( Y=>nx4635, A0=>outMuls_5_11, A1=>nx5290);
   ix2743 : nand02 port map ( Y=>addersInputs_5_12, A0=>nx4638, A1=>nx4640);
   ix4639 : nand02 port map ( Y=>nx4638, A0=>currentPage_5_12, A1=>layerType
   );
   ix4641 : nand02 port map ( Y=>nx4640, A0=>outMuls_5_12, A1=>nx5290);
   ix2751 : nand02 port map ( Y=>addersInputs_5_13, A0=>nx4643, A1=>nx4645);
   ix4644 : nand02 port map ( Y=>nx4643, A0=>currentPage_5_13, A1=>layerType
   );
   ix4646 : nand02 port map ( Y=>nx4645, A0=>outMuls_5_13, A1=>nx5290);
   ix2759 : nand02 port map ( Y=>addersInputs_5_14, A0=>nx4648, A1=>nx4650);
   ix4649 : nand02 port map ( Y=>nx4648, A0=>currentPage_5_14, A1=>layerType
   );
   ix4651 : nand02 port map ( Y=>nx4650, A0=>outMuls_5_14, A1=>nx5290);
   ix2767 : nand02 port map ( Y=>addersInputs_5_15, A0=>nx4653, A1=>nx4655);
   ix4654 : nand02 port map ( Y=>nx4653, A0=>currentPage_5_15, A1=>layerType
   );
   ix4656 : nand02 port map ( Y=>nx4655, A0=>outMuls_5_15, A1=>nx5290);
   ix2775 : nand02 port map ( Y=>addersInputs_4_0, A0=>nx4658, A1=>nx4660);
   ix4659 : nand02 port map ( Y=>nx4658, A0=>currentPage_4_0, A1=>layerType
   );
   ix4661 : nand02 port map ( Y=>nx4660, A0=>outMuls_4_0, A1=>nx5290);
   ix2783 : nand02 port map ( Y=>addersInputs_4_1, A0=>nx4663, A1=>nx4665);
   ix4664 : nand02 port map ( Y=>nx4663, A0=>currentPage_4_1, A1=>layerType
   );
   ix4666 : nand02 port map ( Y=>nx4665, A0=>outMuls_4_1, A1=>nx5290);
   ix2791 : nand02 port map ( Y=>addersInputs_4_2, A0=>nx4668, A1=>nx4670);
   ix4669 : nand02 port map ( Y=>nx4668, A0=>currentPage_4_2, A1=>layerType
   );
   ix4671 : nand02 port map ( Y=>nx4670, A0=>outMuls_4_2, A1=>nx5292);
   ix2799 : nand02 port map ( Y=>addersInputs_4_3, A0=>nx4673, A1=>nx4675);
   ix4674 : nand02 port map ( Y=>nx4673, A0=>currentPage_4_3, A1=>layerType
   );
   ix4676 : nand02 port map ( Y=>nx4675, A0=>outMuls_4_3, A1=>nx5292);
   ix2807 : nand02 port map ( Y=>addersInputs_4_4, A0=>nx4678, A1=>nx4680);
   ix4679 : nand02 port map ( Y=>nx4678, A0=>currentPage_4_4, A1=>layerType
   );
   ix4681 : nand02 port map ( Y=>nx4680, A0=>outMuls_4_4, A1=>nx5292);
   ix2815 : nand02 port map ( Y=>addersInputs_4_5, A0=>nx4683, A1=>nx4685);
   ix4684 : nand02 port map ( Y=>nx4683, A0=>currentPage_4_5, A1=>layerType
   );
   ix4686 : nand02 port map ( Y=>nx4685, A0=>outMuls_4_5, A1=>nx5292);
   ix2823 : nand02 port map ( Y=>addersInputs_4_6, A0=>nx4688, A1=>nx4690);
   ix4689 : nand02 port map ( Y=>nx4688, A0=>currentPage_4_6, A1=>layerType
   );
   ix4691 : nand02 port map ( Y=>nx4690, A0=>outMuls_4_6, A1=>nx5292);
   ix2831 : nand02 port map ( Y=>addersInputs_4_7, A0=>nx4693, A1=>nx4695);
   ix4694 : nand02 port map ( Y=>nx4693, A0=>currentPage_4_7, A1=>layerType
   );
   ix4696 : nand02 port map ( Y=>nx4695, A0=>outMuls_4_7, A1=>nx5292);
   ix2839 : nand02 port map ( Y=>addersInputs_4_8, A0=>nx4698, A1=>nx4700);
   ix4699 : nand02 port map ( Y=>nx4698, A0=>currentPage_4_8, A1=>layerType
   );
   ix4701 : nand02 port map ( Y=>nx4700, A0=>outMuls_4_8, A1=>nx5292);
   ix2847 : nand02 port map ( Y=>addersInputs_4_9, A0=>nx4703, A1=>nx4705);
   ix4704 : nand02 port map ( Y=>nx4703, A0=>currentPage_4_9, A1=>layerType
   );
   ix4706 : nand02 port map ( Y=>nx4705, A0=>outMuls_4_9, A1=>nx5294);
   ix2855 : nand02 port map ( Y=>addersInputs_4_10, A0=>nx4708, A1=>nx4710);
   ix4709 : nand02 port map ( Y=>nx4708, A0=>currentPage_4_10, A1=>layerType
   );
   ix4711 : nand02 port map ( Y=>nx4710, A0=>outMuls_4_10, A1=>nx5294);
   ix2863 : nand02 port map ( Y=>addersInputs_4_11, A0=>nx4713, A1=>nx4715);
   ix4714 : nand02 port map ( Y=>nx4713, A0=>currentPage_4_11, A1=>layerType
   );
   ix4716 : nand02 port map ( Y=>nx4715, A0=>outMuls_4_11, A1=>nx5294);
   ix2871 : nand02 port map ( Y=>addersInputs_4_12, A0=>nx4718, A1=>nx4720);
   ix4719 : nand02 port map ( Y=>nx4718, A0=>currentPage_4_12, A1=>layerType
   );
   ix4721 : nand02 port map ( Y=>nx4720, A0=>outMuls_4_12, A1=>nx5294);
   ix2879 : nand02 port map ( Y=>addersInputs_4_13, A0=>nx4723, A1=>nx4725);
   ix4724 : nand02 port map ( Y=>nx4723, A0=>currentPage_4_13, A1=>layerType
   );
   ix4726 : nand02 port map ( Y=>nx4725, A0=>outMuls_4_13, A1=>nx5294);
   ix2887 : nand02 port map ( Y=>addersInputs_4_14, A0=>nx4728, A1=>nx4730);
   ix4729 : nand02 port map ( Y=>nx4728, A0=>currentPage_4_14, A1=>layerType
   );
   ix4731 : nand02 port map ( Y=>nx4730, A0=>outMuls_4_14, A1=>nx5294);
   ix2895 : nand02 port map ( Y=>addersInputs_4_15, A0=>nx4733, A1=>nx4735);
   ix4734 : nand02 port map ( Y=>nx4733, A0=>currentPage_4_15, A1=>layerType
   );
   ix4736 : nand02 port map ( Y=>nx4735, A0=>outMuls_4_15, A1=>nx5294);
   ix2903 : nand02 port map ( Y=>addersInputs_3_0, A0=>nx4738, A1=>nx4740);
   ix4739 : nand02 port map ( Y=>nx4738, A0=>currentPage_3_0, A1=>layerType
   );
   ix4741 : nand02 port map ( Y=>nx4740, A0=>outMuls_3_0, A1=>nx5296);
   ix2911 : nand02 port map ( Y=>addersInputs_3_1, A0=>nx4743, A1=>nx4745);
   ix4744 : nand02 port map ( Y=>nx4743, A0=>currentPage_3_1, A1=>layerType
   );
   ix4746 : nand02 port map ( Y=>nx4745, A0=>outMuls_3_1, A1=>nx5296);
   ix2919 : nand02 port map ( Y=>addersInputs_3_2, A0=>nx4748, A1=>nx4750);
   ix4749 : nand02 port map ( Y=>nx4748, A0=>currentPage_3_2, A1=>layerType
   );
   ix4751 : nand02 port map ( Y=>nx4750, A0=>outMuls_3_2, A1=>nx5296);
   ix2927 : nand02 port map ( Y=>addersInputs_3_3, A0=>nx4753, A1=>nx4755);
   ix4754 : nand02 port map ( Y=>nx4753, A0=>currentPage_3_3, A1=>layerType
   );
   ix4756 : nand02 port map ( Y=>nx4755, A0=>outMuls_3_3, A1=>nx5296);
   ix2935 : nand02 port map ( Y=>addersInputs_3_4, A0=>nx4758, A1=>nx4760);
   ix4759 : nand02 port map ( Y=>nx4758, A0=>currentPage_3_4, A1=>layerType
   );
   ix4761 : nand02 port map ( Y=>nx4760, A0=>outMuls_3_4, A1=>nx5296);
   ix2943 : nand02 port map ( Y=>addersInputs_3_5, A0=>nx4763, A1=>nx4765);
   ix4764 : nand02 port map ( Y=>nx4763, A0=>currentPage_3_5, A1=>layerType
   );
   ix4766 : nand02 port map ( Y=>nx4765, A0=>outMuls_3_5, A1=>nx5296);
   ix2951 : nand02 port map ( Y=>addersInputs_3_6, A0=>nx4768, A1=>nx4770);
   ix4769 : nand02 port map ( Y=>nx4768, A0=>currentPage_3_6, A1=>layerType
   );
   ix4771 : nand02 port map ( Y=>nx4770, A0=>outMuls_3_6, A1=>nx5296);
   ix2959 : nand02 port map ( Y=>addersInputs_3_7, A0=>nx4773, A1=>nx4775);
   ix4774 : nand02 port map ( Y=>nx4773, A0=>currentPage_3_7, A1=>layerType
   );
   ix4776 : nand02 port map ( Y=>nx4775, A0=>outMuls_3_7, A1=>nx5298);
   ix2967 : nand02 port map ( Y=>addersInputs_3_8, A0=>nx4778, A1=>nx4780);
   ix4779 : nand02 port map ( Y=>nx4778, A0=>currentPage_3_8, A1=>layerType
   );
   ix4781 : nand02 port map ( Y=>nx4780, A0=>outMuls_3_8, A1=>nx5298);
   ix2975 : nand02 port map ( Y=>addersInputs_3_9, A0=>nx4783, A1=>nx4785);
   ix4784 : nand02 port map ( Y=>nx4783, A0=>currentPage_3_9, A1=>layerType
   );
   ix4786 : nand02 port map ( Y=>nx4785, A0=>outMuls_3_9, A1=>nx5298);
   ix2983 : nand02 port map ( Y=>addersInputs_3_10, A0=>nx4788, A1=>nx4790);
   ix4789 : nand02 port map ( Y=>nx4788, A0=>currentPage_3_10, A1=>layerType
   );
   ix4791 : nand02 port map ( Y=>nx4790, A0=>outMuls_3_10, A1=>nx5298);
   ix2991 : nand02 port map ( Y=>addersInputs_3_11, A0=>nx4793, A1=>nx4795);
   ix4794 : nand02 port map ( Y=>nx4793, A0=>currentPage_3_11, A1=>layerType
   );
   ix4796 : nand02 port map ( Y=>nx4795, A0=>outMuls_3_11, A1=>nx5298);
   ix2999 : nand02 port map ( Y=>addersInputs_3_12, A0=>nx4798, A1=>nx4800);
   ix4799 : nand02 port map ( Y=>nx4798, A0=>currentPage_3_12, A1=>layerType
   );
   ix4801 : nand02 port map ( Y=>nx4800, A0=>outMuls_3_12, A1=>nx5298);
   ix3007 : nand02 port map ( Y=>addersInputs_3_13, A0=>nx4803, A1=>nx4805);
   ix4804 : nand02 port map ( Y=>nx4803, A0=>currentPage_3_13, A1=>layerType
   );
   ix4806 : nand02 port map ( Y=>nx4805, A0=>outMuls_3_13, A1=>nx5298);
   ix3015 : nand02 port map ( Y=>addersInputs_3_14, A0=>nx4808, A1=>nx4810);
   ix4809 : nand02 port map ( Y=>nx4808, A0=>currentPage_3_14, A1=>layerType
   );
   ix4811 : nand02 port map ( Y=>nx4810, A0=>outMuls_3_14, A1=>nx5300);
   ix3023 : nand02 port map ( Y=>addersInputs_3_15, A0=>nx4813, A1=>nx4815);
   ix4814 : nand02 port map ( Y=>nx4813, A0=>currentPage_3_15, A1=>layerType
   );
   ix4816 : nand02 port map ( Y=>nx4815, A0=>outMuls_3_15, A1=>nx5300);
   ix3031 : nand02 port map ( Y=>addersInputs_2_0, A0=>nx4818, A1=>nx4820);
   ix4819 : nand02 port map ( Y=>nx4818, A0=>currentPage_2_0, A1=>layerType
   );
   ix4821 : nand02 port map ( Y=>nx4820, A0=>outMuls_2_0, A1=>nx5300);
   ix3039 : nand02 port map ( Y=>addersInputs_2_1, A0=>nx4823, A1=>nx4825);
   ix4824 : nand02 port map ( Y=>nx4823, A0=>currentPage_2_1, A1=>layerType
   );
   ix4826 : nand02 port map ( Y=>nx4825, A0=>outMuls_2_1, A1=>nx5300);
   ix3047 : nand02 port map ( Y=>addersInputs_2_2, A0=>nx4828, A1=>nx4830);
   ix4829 : nand02 port map ( Y=>nx4828, A0=>currentPage_2_2, A1=>layerType
   );
   ix4831 : nand02 port map ( Y=>nx4830, A0=>outMuls_2_2, A1=>nx5300);
   ix3055 : nand02 port map ( Y=>addersInputs_2_3, A0=>nx4833, A1=>nx4835);
   ix4834 : nand02 port map ( Y=>nx4833, A0=>currentPage_2_3, A1=>layerType
   );
   ix4836 : nand02 port map ( Y=>nx4835, A0=>outMuls_2_3, A1=>nx5300);
   ix3063 : nand02 port map ( Y=>addersInputs_2_4, A0=>nx4838, A1=>nx4840);
   ix4839 : nand02 port map ( Y=>nx4838, A0=>currentPage_2_4, A1=>layerType
   );
   ix4841 : nand02 port map ( Y=>nx4840, A0=>outMuls_2_4, A1=>nx5300);
   ix3071 : nand02 port map ( Y=>addersInputs_2_5, A0=>nx4843, A1=>nx4845);
   ix4844 : nand02 port map ( Y=>nx4843, A0=>currentPage_2_5, A1=>layerType
   );
   ix4846 : nand02 port map ( Y=>nx4845, A0=>outMuls_2_5, A1=>nx5302);
   ix3079 : nand02 port map ( Y=>addersInputs_2_6, A0=>nx4848, A1=>nx4850);
   ix4849 : nand02 port map ( Y=>nx4848, A0=>currentPage_2_6, A1=>layerType
   );
   ix4851 : nand02 port map ( Y=>nx4850, A0=>outMuls_2_6, A1=>nx5302);
   ix3087 : nand02 port map ( Y=>addersInputs_2_7, A0=>nx4853, A1=>nx4855);
   ix4854 : nand02 port map ( Y=>nx4853, A0=>currentPage_2_7, A1=>layerType
   );
   ix4856 : nand02 port map ( Y=>nx4855, A0=>outMuls_2_7, A1=>nx5302);
   ix3095 : nand02 port map ( Y=>addersInputs_2_8, A0=>nx4858, A1=>nx4860);
   ix4859 : nand02 port map ( Y=>nx4858, A0=>currentPage_2_8, A1=>layerType
   );
   ix4861 : nand02 port map ( Y=>nx4860, A0=>outMuls_2_8, A1=>nx5302);
   ix3103 : nand02 port map ( Y=>addersInputs_2_9, A0=>nx4863, A1=>nx4865);
   ix4864 : nand02 port map ( Y=>nx4863, A0=>currentPage_2_9, A1=>layerType
   );
   ix4866 : nand02 port map ( Y=>nx4865, A0=>outMuls_2_9, A1=>nx5302);
   ix3111 : nand02 port map ( Y=>addersInputs_2_10, A0=>nx4868, A1=>nx4870);
   ix4869 : nand02 port map ( Y=>nx4868, A0=>currentPage_2_10, A1=>layerType
   );
   ix4871 : nand02 port map ( Y=>nx4870, A0=>outMuls_2_10, A1=>nx5302);
   ix3119 : nand02 port map ( Y=>addersInputs_2_11, A0=>nx4873, A1=>nx4875);
   ix4874 : nand02 port map ( Y=>nx4873, A0=>currentPage_2_11, A1=>layerType
   );
   ix4876 : nand02 port map ( Y=>nx4875, A0=>outMuls_2_11, A1=>nx5302);
   ix3127 : nand02 port map ( Y=>addersInputs_2_12, A0=>nx4878, A1=>nx4880);
   ix4879 : nand02 port map ( Y=>nx4878, A0=>currentPage_2_12, A1=>layerType
   );
   ix4881 : nand02 port map ( Y=>nx4880, A0=>outMuls_2_12, A1=>nx5304);
   ix3135 : nand02 port map ( Y=>addersInputs_2_13, A0=>nx4883, A1=>nx4885);
   ix4884 : nand02 port map ( Y=>nx4883, A0=>currentPage_2_13, A1=>layerType
   );
   ix4886 : nand02 port map ( Y=>nx4885, A0=>outMuls_2_13, A1=>nx5304);
   ix3143 : nand02 port map ( Y=>addersInputs_2_14, A0=>nx4888, A1=>nx4890);
   ix4889 : nand02 port map ( Y=>nx4888, A0=>currentPage_2_14, A1=>layerType
   );
   ix4891 : nand02 port map ( Y=>nx4890, A0=>outMuls_2_14, A1=>nx5304);
   ix3151 : nand02 port map ( Y=>addersInputs_2_15, A0=>nx4893, A1=>nx4895);
   ix4894 : nand02 port map ( Y=>nx4893, A0=>currentPage_2_15, A1=>layerType
   );
   ix4896 : nand02 port map ( Y=>nx4895, A0=>outMuls_2_15, A1=>nx5304);
   ix3159 : nand02 port map ( Y=>addersInputs_1_0, A0=>nx4898, A1=>nx4900);
   ix4899 : nand02 port map ( Y=>nx4898, A0=>currentPage_1_0, A1=>layerType
   );
   ix4901 : nand02 port map ( Y=>nx4900, A0=>outMuls_1_0, A1=>nx5304);
   ix3167 : nand02 port map ( Y=>addersInputs_1_1, A0=>nx4903, A1=>nx4905);
   ix4904 : nand02 port map ( Y=>nx4903, A0=>currentPage_1_1, A1=>layerType
   );
   ix4906 : nand02 port map ( Y=>nx4905, A0=>outMuls_1_1, A1=>nx5304);
   ix3175 : nand02 port map ( Y=>addersInputs_1_2, A0=>nx4908, A1=>nx4910);
   ix4909 : nand02 port map ( Y=>nx4908, A0=>currentPage_1_2, A1=>layerType
   );
   ix4911 : nand02 port map ( Y=>nx4910, A0=>outMuls_1_2, A1=>nx5304);
   ix3183 : nand02 port map ( Y=>addersInputs_1_3, A0=>nx4913, A1=>nx4915);
   ix4914 : nand02 port map ( Y=>nx4913, A0=>currentPage_1_3, A1=>layerType
   );
   ix4916 : nand02 port map ( Y=>nx4915, A0=>outMuls_1_3, A1=>nx5306);
   ix3191 : nand02 port map ( Y=>addersInputs_1_4, A0=>nx4918, A1=>nx4920);
   ix4919 : nand02 port map ( Y=>nx4918, A0=>currentPage_1_4, A1=>layerType
   );
   ix4921 : nand02 port map ( Y=>nx4920, A0=>outMuls_1_4, A1=>nx5306);
   ix3199 : nand02 port map ( Y=>addersInputs_1_5, A0=>nx4923, A1=>nx4925);
   ix4924 : nand02 port map ( Y=>nx4923, A0=>currentPage_1_5, A1=>layerType
   );
   ix4926 : nand02 port map ( Y=>nx4925, A0=>outMuls_1_5, A1=>nx5306);
   ix3207 : nand02 port map ( Y=>addersInputs_1_6, A0=>nx4928, A1=>nx4930);
   ix4929 : nand02 port map ( Y=>nx4928, A0=>currentPage_1_6, A1=>layerType
   );
   ix4931 : nand02 port map ( Y=>nx4930, A0=>outMuls_1_6, A1=>nx5306);
   ix3215 : nand02 port map ( Y=>addersInputs_1_7, A0=>nx4933, A1=>nx4935);
   ix4934 : nand02 port map ( Y=>nx4933, A0=>currentPage_1_7, A1=>layerType
   );
   ix4936 : nand02 port map ( Y=>nx4935, A0=>outMuls_1_7, A1=>nx5306);
   ix3223 : nand02 port map ( Y=>addersInputs_1_8, A0=>nx4938, A1=>nx4940);
   ix4939 : nand02 port map ( Y=>nx4938, A0=>currentPage_1_8, A1=>layerType
   );
   ix4941 : nand02 port map ( Y=>nx4940, A0=>outMuls_1_8, A1=>nx5306);
   ix3231 : nand02 port map ( Y=>addersInputs_1_9, A0=>nx4943, A1=>nx4945);
   ix4944 : nand02 port map ( Y=>nx4943, A0=>currentPage_1_9, A1=>layerType
   );
   ix4946 : nand02 port map ( Y=>nx4945, A0=>outMuls_1_9, A1=>nx5306);
   ix3239 : nand02 port map ( Y=>addersInputs_1_10, A0=>nx4948, A1=>nx4950);
   ix4949 : nand02 port map ( Y=>nx4948, A0=>currentPage_1_10, A1=>layerType
   );
   ix4951 : nand02 port map ( Y=>nx4950, A0=>outMuls_1_10, A1=>nx5308);
   ix3247 : nand02 port map ( Y=>addersInputs_1_11, A0=>nx4953, A1=>nx4955);
   ix4954 : nand02 port map ( Y=>nx4953, A0=>currentPage_1_11, A1=>layerType
   );
   ix4956 : nand02 port map ( Y=>nx4955, A0=>outMuls_1_11, A1=>nx5308);
   ix3255 : nand02 port map ( Y=>addersInputs_1_12, A0=>nx4958, A1=>nx4960);
   ix4959 : nand02 port map ( Y=>nx4958, A0=>currentPage_1_12, A1=>layerType
   );
   ix4961 : nand02 port map ( Y=>nx4960, A0=>outMuls_1_12, A1=>nx5308);
   ix3263 : nand02 port map ( Y=>addersInputs_1_13, A0=>nx4963, A1=>nx4965);
   ix4964 : nand02 port map ( Y=>nx4963, A0=>currentPage_1_13, A1=>layerType
   );
   ix4966 : nand02 port map ( Y=>nx4965, A0=>outMuls_1_13, A1=>nx5308);
   ix3271 : nand02 port map ( Y=>addersInputs_1_14, A0=>nx4968, A1=>nx4970);
   ix4969 : nand02 port map ( Y=>nx4968, A0=>currentPage_1_14, A1=>layerType
   );
   ix4971 : nand02 port map ( Y=>nx4970, A0=>outMuls_1_14, A1=>nx5308);
   ix3279 : nand02 port map ( Y=>addersInputs_1_15, A0=>nx4973, A1=>nx4975);
   ix4974 : nand02 port map ( Y=>nx4973, A0=>currentPage_1_15, A1=>layerType
   );
   ix4976 : nand02 port map ( Y=>nx4975, A0=>outMuls_1_15, A1=>nx5308);
   ix3287 : nand02 port map ( Y=>addersInputs_0_0, A0=>nx4978, A1=>nx4980);
   ix4979 : nand02 port map ( Y=>nx4978, A0=>currentPage_0_0, A1=>layerType
   );
   ix4981 : nand02 port map ( Y=>nx4980, A0=>outMuls_0_0, A1=>nx5308);
   ix3295 : nand02 port map ( Y=>addersInputs_0_1, A0=>nx4983, A1=>nx4985);
   ix4984 : nand02 port map ( Y=>nx4983, A0=>currentPage_0_1, A1=>layerType
   );
   ix4986 : nand02 port map ( Y=>nx4985, A0=>outMuls_0_1, A1=>nx5310);
   ix3303 : nand02 port map ( Y=>addersInputs_0_2, A0=>nx4988, A1=>nx4990);
   ix4989 : nand02 port map ( Y=>nx4988, A0=>currentPage_0_2, A1=>layerType
   );
   ix4991 : nand02 port map ( Y=>nx4990, A0=>outMuls_0_2, A1=>nx5310);
   ix3311 : nand02 port map ( Y=>addersInputs_0_3, A0=>nx4993, A1=>nx4995);
   ix4994 : nand02 port map ( Y=>nx4993, A0=>currentPage_0_3, A1=>layerType
   );
   ix4996 : nand02 port map ( Y=>nx4995, A0=>outMuls_0_3, A1=>nx5310);
   ix3319 : nand02 port map ( Y=>addersInputs_0_4, A0=>nx4998, A1=>nx5000);
   ix4999 : nand02 port map ( Y=>nx4998, A0=>currentPage_0_4, A1=>layerType
   );
   ix5001 : nand02 port map ( Y=>nx5000, A0=>outMuls_0_4, A1=>nx5310);
   ix3327 : nand02 port map ( Y=>addersInputs_0_5, A0=>nx5003, A1=>nx5005);
   ix5004 : nand02 port map ( Y=>nx5003, A0=>currentPage_0_5, A1=>layerType
   );
   ix5006 : nand02 port map ( Y=>nx5005, A0=>outMuls_0_5, A1=>nx5310);
   ix3335 : nand02 port map ( Y=>addersInputs_0_6, A0=>nx5008, A1=>nx5010);
   ix5009 : nand02 port map ( Y=>nx5008, A0=>currentPage_0_6, A1=>layerType
   );
   ix5011 : nand02 port map ( Y=>nx5010, A0=>outMuls_0_6, A1=>nx5310);
   ix3343 : nand02 port map ( Y=>addersInputs_0_7, A0=>nx5013, A1=>nx5015);
   ix5014 : nand02 port map ( Y=>nx5013, A0=>currentPage_0_7, A1=>layerType
   );
   ix5016 : nand02 port map ( Y=>nx5015, A0=>outMuls_0_7, A1=>nx5310);
   ix3351 : nand02 port map ( Y=>addersInputs_0_8, A0=>nx5018, A1=>nx5020);
   ix5019 : nand02 port map ( Y=>nx5018, A0=>currentPage_0_8, A1=>layerType
   );
   ix5021 : nand02 port map ( Y=>nx5020, A0=>outMuls_0_8, A1=>nx5312);
   ix3359 : nand02 port map ( Y=>addersInputs_0_9, A0=>nx5023, A1=>nx5025);
   ix5024 : nand02 port map ( Y=>nx5023, A0=>currentPage_0_9, A1=>layerType
   );
   ix5026 : nand02 port map ( Y=>nx5025, A0=>outMuls_0_9, A1=>nx5312);
   ix3367 : nand02 port map ( Y=>addersInputs_0_10, A0=>nx5028, A1=>nx5030);
   ix5029 : nand02 port map ( Y=>nx5028, A0=>currentPage_0_10, A1=>layerType
   );
   ix5031 : nand02 port map ( Y=>nx5030, A0=>outMuls_0_10, A1=>nx5312);
   ix3375 : nand02 port map ( Y=>addersInputs_0_11, A0=>nx5033, A1=>nx5035);
   ix5034 : nand02 port map ( Y=>nx5033, A0=>currentPage_0_11, A1=>layerType
   );
   ix5036 : nand02 port map ( Y=>nx5035, A0=>outMuls_0_11, A1=>nx5312);
   ix3383 : nand02 port map ( Y=>addersInputs_0_12, A0=>nx5038, A1=>nx5040);
   ix5039 : nand02 port map ( Y=>nx5038, A0=>currentPage_0_12, A1=>layerType
   );
   ix5041 : nand02 port map ( Y=>nx5040, A0=>outMuls_0_12, A1=>nx5312);
   ix3391 : nand02 port map ( Y=>addersInputs_0_13, A0=>nx5043, A1=>nx5045);
   ix5044 : nand02 port map ( Y=>nx5043, A0=>currentPage_0_13, A1=>layerType
   );
   ix5046 : nand02 port map ( Y=>nx5045, A0=>outMuls_0_13, A1=>nx5312);
   ix3399 : nand02 port map ( Y=>addersInputs_0_14, A0=>nx5048, A1=>nx5050);
   ix5049 : nand02 port map ( Y=>nx5048, A0=>currentPage_0_14, A1=>layerType
   );
   ix5051 : nand02 port map ( Y=>nx5050, A0=>outMuls_0_14, A1=>nx5312);
   ix3407 : nand02 port map ( Y=>addersInputs_0_15, A0=>nx5053, A1=>nx5055);
   ix5054 : nand02 port map ( Y=>nx5053, A0=>currentPage_0_15, A1=>layerType
   );
   ix5056 : nand02 port map ( Y=>nx5055, A0=>outMuls_0_15, A1=>nx5314);
   ix47 : nand04 port map ( Y=>finalSum(0), A0=>nx5058, A1=>nx5060, A2=>
      nx5063, A3=>nx5067);
   ix5059 : nand03 port map ( Y=>nx5058, A0=>addersMap_totalSum_0, A1=>
      filterType, A2=>nx5314);
   ix5061 : nand02 port map ( Y=>nx5060, A0=>addersMap_sum3Filter_0, A1=>
      nx5196);
   ix5 : nor02_2x port map ( Y=>nx4, A0=>filterType, A1=>layerType);
   ix5064 : nand03 port map ( Y=>nx5063, A0=>addersMap_sum3Filter_3, A1=>
      nx5320, A2=>layerType);
   ix5068 : nand03 port map ( Y=>nx5067, A0=>addersMap_totalSum_5, A1=>
      filterType, A2=>layerType);
   ix61 : nand04 port map ( Y=>finalSum(1), A0=>nx5070, A1=>nx5072, A2=>
      nx5074, A3=>nx5076);
   ix5071 : nand03 port map ( Y=>nx5070, A0=>addersMap_totalSum_1, A1=>
      filterType, A2=>nx5314);
   ix5073 : nand02 port map ( Y=>nx5072, A0=>addersMap_sum3Filter_1, A1=>
      nx5196);
   ix5075 : nand03 port map ( Y=>nx5074, A0=>addersMap_sum3Filter_4, A1=>
      nx5320, A2=>layerType);
   ix5077 : nand03 port map ( Y=>nx5076, A0=>addersMap_totalSum_6, A1=>
      filterType, A2=>layerType);
   ix75 : nand04 port map ( Y=>finalSum(2), A0=>nx5079, A1=>nx5081, A2=>
      nx5083, A3=>nx5085);
   ix5080 : nand03 port map ( Y=>nx5079, A0=>addersMap_totalSum_2, A1=>
      filterType, A2=>nx5314);
   ix5082 : nand02 port map ( Y=>nx5081, A0=>addersMap_sum3Filter_2, A1=>
      nx5196);
   ix5084 : nand03 port map ( Y=>nx5083, A0=>addersMap_sum3Filter_5, A1=>
      nx5320, A2=>layerType);
   ix5086 : nand03 port map ( Y=>nx5085, A0=>addersMap_totalSum_7, A1=>
      filterType, A2=>layerType);
   ix89 : nand04 port map ( Y=>finalSum(3), A0=>nx5088, A1=>nx5090, A2=>
      nx5092, A3=>nx5094);
   ix5089 : nand03 port map ( Y=>nx5088, A0=>addersMap_totalSum_3, A1=>
      filterType, A2=>nx5314);
   ix5091 : nand02 port map ( Y=>nx5090, A0=>addersMap_sum3Filter_3, A1=>
      nx5196);
   ix5093 : nand03 port map ( Y=>nx5092, A0=>addersMap_sum3Filter_6, A1=>
      nx5320, A2=>layerType);
   ix5095 : nand03 port map ( Y=>nx5094, A0=>addersMap_totalSum_8, A1=>
      filterType, A2=>layerType);
   ix103 : nand04 port map ( Y=>finalSum(4), A0=>nx5097, A1=>nx5099, A2=>
      nx5101, A3=>nx5103);
   ix5098 : nand03 port map ( Y=>nx5097, A0=>addersMap_totalSum_4, A1=>
      filterType, A2=>nx5314);
   ix5100 : nand02 port map ( Y=>nx5099, A0=>addersMap_sum3Filter_4, A1=>
      nx5196);
   ix5102 : nand03 port map ( Y=>nx5101, A0=>addersMap_sum3Filter_7, A1=>
      nx5320, A2=>layerType);
   ix5104 : nand03 port map ( Y=>nx5103, A0=>addersMap_totalSum_9, A1=>
      filterType, A2=>layerType);
   ix117 : nand04 port map ( Y=>finalSum(5), A0=>nx5106, A1=>nx5108, A2=>
      nx5110, A3=>nx5112);
   ix5107 : nand03 port map ( Y=>nx5106, A0=>addersMap_totalSum_5, A1=>
      filterType, A2=>nx5314);
   ix5109 : nand02 port map ( Y=>nx5108, A0=>addersMap_sum3Filter_5, A1=>
      nx5196);
   ix5111 : nand03 port map ( Y=>nx5110, A0=>addersMap_sum3Filter_8, A1=>
      nx5320, A2=>layerType);
   ix5113 : nand03 port map ( Y=>nx5112, A0=>addersMap_totalSum_10, A1=>
      filterType, A2=>layerType);
   ix131 : nand04 port map ( Y=>finalSum(6), A0=>nx5115, A1=>nx5117, A2=>
      nx5119, A3=>nx5121);
   ix5116 : nand03 port map ( Y=>nx5115, A0=>addersMap_totalSum_6, A1=>
      filterType, A2=>nx5316);
   ix5118 : nand02 port map ( Y=>nx5117, A0=>addersMap_sum3Filter_6, A1=>
      nx5196);
   ix5120 : nand03 port map ( Y=>nx5119, A0=>addersMap_sum3Filter_9, A1=>
      nx5320, A2=>layerType);
   ix5122 : nand03 port map ( Y=>nx5121, A0=>addersMap_totalSum_11, A1=>
      filterType, A2=>layerType);
   ix145 : nand04 port map ( Y=>finalSum(7), A0=>nx5124, A1=>nx5126, A2=>
      nx5128, A3=>nx5130);
   ix5125 : nand03 port map ( Y=>nx5124, A0=>addersMap_totalSum_7, A1=>
      filterType, A2=>nx5316);
   ix5127 : nand02 port map ( Y=>nx5126, A0=>addersMap_sum3Filter_7, A1=>
      nx5198);
   ix5129 : nand03 port map ( Y=>nx5128, A0=>addersMap_sum3Filter_10, A1=>
      nx5322, A2=>layerType);
   ix5131 : nand03 port map ( Y=>nx5130, A0=>addersMap_totalSum_12, A1=>
      filterType, A2=>layerType);
   ix159 : nand04 port map ( Y=>finalSum(8), A0=>nx5133, A1=>nx5135, A2=>
      nx5137, A3=>nx5139);
   ix5134 : nand03 port map ( Y=>nx5133, A0=>addersMap_totalSum_8, A1=>
      filterType, A2=>nx5316);
   ix5136 : nand02 port map ( Y=>nx5135, A0=>addersMap_sum3Filter_8, A1=>
      nx5198);
   ix5138 : nand03 port map ( Y=>nx5137, A0=>addersMap_sum3Filter_11, A1=>
      nx5322, A2=>layerType);
   ix5140 : nand03 port map ( Y=>nx5139, A0=>addersMap_totalSum_13, A1=>
      filterType, A2=>layerType);
   ix173 : nand04 port map ( Y=>finalSum(9), A0=>nx5142, A1=>nx5144, A2=>
      nx5146, A3=>nx5148);
   ix5143 : nand03 port map ( Y=>nx5142, A0=>addersMap_totalSum_9, A1=>
      filterType, A2=>nx5316);
   ix5145 : nand02 port map ( Y=>nx5144, A0=>addersMap_sum3Filter_9, A1=>
      nx5198);
   ix5147 : nand03 port map ( Y=>nx5146, A0=>addersMap_sum3Filter_12, A1=>
      nx5322, A2=>layerType);
   ix5149 : nand03 port map ( Y=>nx5148, A0=>addersMap_totalSum_14, A1=>
      filterType, A2=>layerType);
   ix187 : nand04 port map ( Y=>finalSum(10), A0=>nx5151, A1=>nx5153, A2=>
      nx5155, A3=>nx5157);
   ix5152 : nand03 port map ( Y=>nx5151, A0=>addersMap_totalSum_10, A1=>
      filterType, A2=>nx5316);
   ix5154 : nand02 port map ( Y=>nx5153, A0=>addersMap_sum3Filter_10, A1=>
      nx5198);
   ix5156 : nand03 port map ( Y=>nx5155, A0=>addersMap_sum3Filter_13, A1=>
      nx5322, A2=>layerType);
   ix5158 : nand03 port map ( Y=>nx5157, A0=>addersMap_totalSum_15, A1=>
      filterType, A2=>layerType);
   ix197 : nand03 port map ( Y=>finalSum(11), A0=>nx5160, A1=>nx5162, A2=>
      nx5164);
   ix5161 : nand02 port map ( Y=>nx5160, A0=>addersMap_sum3Filter_11, A1=>
      nx5198);
   ix5163 : nand03 port map ( Y=>nx5162, A0=>addersMap_sum3Filter_14, A1=>
      nx5322, A2=>layerType);
   ix5165 : nand03 port map ( Y=>nx5164, A0=>addersMap_totalSum_11, A1=>
      filterType, A2=>nx5316);
   ix207 : nand03 port map ( Y=>finalSum(12), A0=>nx5167, A1=>nx5169, A2=>
      nx5171);
   ix5168 : nand02 port map ( Y=>nx5167, A0=>addersMap_sum3Filter_12, A1=>
      nx5198);
   ix5170 : nand03 port map ( Y=>nx5169, A0=>addersMap_sum3Filter_15, A1=>
      nx5322, A2=>layerType);
   ix5172 : nand03 port map ( Y=>nx5171, A0=>addersMap_totalSum_12, A1=>
      filterType, A2=>nx5316);
   ix15 : nand02 port map ( Y=>finalSum(13), A0=>nx5174, A1=>nx5176);
   ix5175 : nand03 port map ( Y=>nx5174, A0=>addersMap_totalSum_13, A1=>
      filterType, A2=>nx5318);
   ix5177 : nand02 port map ( Y=>nx5176, A0=>addersMap_sum3Filter_13, A1=>
      nx5198);
   ix21 : nand02 port map ( Y=>finalSum(14), A0=>nx5179, A1=>nx5181);
   ix5180 : nand03 port map ( Y=>nx5179, A0=>addersMap_totalSum_14, A1=>
      filterType, A2=>nx5318);
   ix5182 : nand02 port map ( Y=>nx5181, A0=>addersMap_sum3Filter_14, A1=>
      nx4);
   ix27 : nand02 port map ( Y=>finalSum(15), A0=>nx5184, A1=>nx5186);
   ix5185 : nand03 port map ( Y=>nx5184, A0=>addersMap_totalSum_15, A1=>
      filterType, A2=>nx5318);
   ix5187 : nand02 port map ( Y=>nx5186, A0=>addersMap_sum3Filter_15, A1=>
      nx4);
   ix3481 : inv01 port map ( Y=>done, A=>nx5189);
   ix5190 : nor02_2x port map ( Y=>nx5189, A0=>layerType, A1=>doneMul);
   ix5195 : nor02_2x port map ( Y=>nx5196, A0=>filterType, A1=>layerType);
   ix5197 : nor02_2x port map ( Y=>nx5198, A0=>filterType, A1=>layerType);
   ix5199 : inv02 port map ( Y=>nx5200, A=>layerType);
   ix5201 : inv02 port map ( Y=>nx5202, A=>layerType);
   ix5203 : inv02 port map ( Y=>nx5204, A=>layerType);
   ix5205 : inv02 port map ( Y=>nx5206, A=>layerType);
   ix5207 : inv02 port map ( Y=>nx5208, A=>layerType);
   ix5209 : inv02 port map ( Y=>nx5210, A=>layerType);
   ix5211 : inv02 port map ( Y=>nx5212, A=>layerType);
   ix5213 : inv02 port map ( Y=>nx5214, A=>layerType);
   ix5215 : inv02 port map ( Y=>nx5216, A=>layerType);
   ix5217 : inv02 port map ( Y=>nx5218, A=>layerType);
   ix5219 : inv02 port map ( Y=>nx5220, A=>layerType);
   ix5221 : inv02 port map ( Y=>nx5222, A=>layerType);
   ix5223 : inv02 port map ( Y=>nx5224, A=>layerType);
   ix5225 : inv02 port map ( Y=>nx5226, A=>layerType);
   ix5227 : inv02 port map ( Y=>nx5228, A=>layerType);
   ix5229 : inv02 port map ( Y=>nx5230, A=>layerType);
   ix5231 : inv02 port map ( Y=>nx5232, A=>layerType);
   ix5233 : inv02 port map ( Y=>nx5234, A=>layerType);
   ix5235 : inv02 port map ( Y=>nx5236, A=>layerType);
   ix5237 : inv02 port map ( Y=>nx5238, A=>layerType);
   ix5239 : inv02 port map ( Y=>nx5240, A=>layerType);
   ix5241 : inv02 port map ( Y=>nx5242, A=>layerType);
   ix5243 : inv02 port map ( Y=>nx5244, A=>layerType);
   ix5245 : inv02 port map ( Y=>nx5246, A=>layerType);
   ix5247 : inv02 port map ( Y=>nx5248, A=>layerType);
   ix5249 : inv02 port map ( Y=>nx5250, A=>layerType);
   ix5251 : inv02 port map ( Y=>nx5252, A=>layerType);
   ix5253 : inv02 port map ( Y=>nx5254, A=>layerType);
   ix5255 : inv02 port map ( Y=>nx5256, A=>layerType);
   ix5257 : inv02 port map ( Y=>nx5258, A=>layerType);
   ix5259 : inv02 port map ( Y=>nx5260, A=>layerType);
   ix5261 : inv02 port map ( Y=>nx5262, A=>layerType);
   ix5263 : inv02 port map ( Y=>nx5264, A=>layerType);
   ix5265 : inv02 port map ( Y=>nx5266, A=>layerType);
   ix5267 : inv02 port map ( Y=>nx5268, A=>layerType);
   ix5269 : inv02 port map ( Y=>nx5270, A=>layerType);
   ix5271 : inv02 port map ( Y=>nx5272, A=>layerType);
   ix5273 : inv02 port map ( Y=>nx5274, A=>layerType);
   ix5275 : inv02 port map ( Y=>nx5276, A=>layerType);
   ix5277 : inv02 port map ( Y=>nx5278, A=>layerType);
   ix5279 : inv02 port map ( Y=>nx5280, A=>layerType);
   ix5281 : inv02 port map ( Y=>nx5282, A=>layerType);
   ix5283 : inv02 port map ( Y=>nx5284, A=>layerType);
   ix5285 : inv02 port map ( Y=>nx5286, A=>layerType);
   ix5287 : inv02 port map ( Y=>nx5288, A=>layerType);
   ix5289 : inv02 port map ( Y=>nx5290, A=>layerType);
   ix5291 : inv02 port map ( Y=>nx5292, A=>layerType);
   ix5293 : inv02 port map ( Y=>nx5294, A=>layerType);
   ix5295 : inv02 port map ( Y=>nx5296, A=>layerType);
   ix5297 : inv02 port map ( Y=>nx5298, A=>layerType);
   ix5299 : inv02 port map ( Y=>nx5300, A=>layerType);
   ix5301 : inv02 port map ( Y=>nx5302, A=>layerType);
   ix5303 : inv02 port map ( Y=>nx5304, A=>layerType);
   ix5305 : inv02 port map ( Y=>nx5306, A=>layerType);
   ix5307 : inv02 port map ( Y=>nx5308, A=>layerType);
   ix5309 : inv02 port map ( Y=>nx5310, A=>layerType);
   ix5311 : inv02 port map ( Y=>nx5312, A=>layerType);
   ix5313 : inv02 port map ( Y=>nx5314, A=>layerType);
   ix5315 : inv02 port map ( Y=>nx5316, A=>layerType);
   ix5317 : inv02 port map ( Y=>nx5318, A=>layerType);
   ix5319 : inv02 port map ( Y=>nx5320, A=>filterType);
   ix5321 : inv02 port map ( Y=>nx5322, A=>filterType);
   ix5327 : buf02 port map ( Y=>nx5328, A=>regFileMap_filterEnables_0);
   ix5329 : buf02 port map ( Y=>nx5330, A=>regFileMap_filterEnables_0);
   ix5331 : buf02 port map ( Y=>nx5332, A=>regFileMap_filterEnables_1);
   ix5333 : buf02 port map ( Y=>nx5334, A=>regFileMap_filterEnables_1);
   ix5335 : buf02 port map ( Y=>nx5336, A=>regFileMap_filterEnables_2);
   ix5337 : buf02 port map ( Y=>nx5338, A=>regFileMap_filterEnables_2);
   ix5339 : buf02 port map ( Y=>nx5340, A=>regFileMap_filterEnables_3);
   ix5341 : buf02 port map ( Y=>nx5342, A=>regFileMap_filterEnables_3);
   ix5343 : inv02 port map ( Y=>nx5344, A=>nx2917);
   ix5345 : inv02 port map ( Y=>nx5346, A=>nx2917);
end CNNCoresArch ;

