PACKAGE constants IS    

-- configurations
CONSTANT outputSize: integer:=0;
CONSTANT filterSize: integer:=1;
CONSTANT inputSize: integer:=2; -- height or width size of the input image
constant configCount: integer :=3;





constant addressSize: integer := 20 -- bits
constant maxImageSize: integer := 28 -- bits


END constants;