//
// Verilog description for cell CNNCores, 
// Thu Apr 11 17:37:23 2019
//
// LeonardoSpectrum Level 3, 2018a.2 
//


module CNNCores ( filterBus, windowBus, decoderRow, clk, rst, writePage1, 
                  writePage2, writeFilter, shift2To1, shift1To2, pageTurn, start, 
                  layerType, filterType, done, finalSum ) ;

    input [39:0]filterBus ;
    input [79:0]windowBus ;
    input [2:0]decoderRow ;
    input clk ;
    input rst ;
    input writePage1 ;
    input writePage2 ;
    input writeFilter ;
    input shift2To1 ;
    input shift1To2 ;
    input pageTurn ;
    input start ;
    input layerType ;
    input filterType ;
    output done ;
    output [15:0]finalSum ;

    wire currentPage_0__15, currentPage_0__14, currentPage_0__13, 
         currentPage_0__12, currentPage_0__11, currentPage_0__10, 
         currentPage_0__9, currentPage_0__8, currentPage_0__7, currentPage_0__6, 
         currentPage_0__5, currentPage_0__4, currentPage_0__3, currentPage_0__2, 
         currentPage_0__1, currentPage_0__0, currentPage_1__15, 
         currentPage_1__14, currentPage_1__13, currentPage_1__12, 
         currentPage_1__11, currentPage_1__10, currentPage_1__9, 
         currentPage_1__8, currentPage_1__7, currentPage_1__6, currentPage_1__5, 
         currentPage_1__4, currentPage_1__3, currentPage_1__2, currentPage_1__1, 
         currentPage_1__0, currentPage_2__15, currentPage_2__14, 
         currentPage_2__13, currentPage_2__12, currentPage_2__11, 
         currentPage_2__10, currentPage_2__9, currentPage_2__8, currentPage_2__7, 
         currentPage_2__6, currentPage_2__5, currentPage_2__4, currentPage_2__3, 
         currentPage_2__2, currentPage_2__1, currentPage_2__0, currentPage_3__15, 
         currentPage_3__14, currentPage_3__13, currentPage_3__12, 
         currentPage_3__11, currentPage_3__10, currentPage_3__9, 
         currentPage_3__8, currentPage_3__7, currentPage_3__6, currentPage_3__5, 
         currentPage_3__4, currentPage_3__3, currentPage_3__2, currentPage_3__1, 
         currentPage_3__0, currentPage_4__15, currentPage_4__14, 
         currentPage_4__13, currentPage_4__12, currentPage_4__11, 
         currentPage_4__10, currentPage_4__9, currentPage_4__8, currentPage_4__7, 
         currentPage_4__6, currentPage_4__5, currentPage_4__4, currentPage_4__3, 
         currentPage_4__2, currentPage_4__1, currentPage_4__0, currentPage_5__15, 
         currentPage_5__14, currentPage_5__13, currentPage_5__12, 
         currentPage_5__11, currentPage_5__10, currentPage_5__9, 
         currentPage_5__8, currentPage_5__7, currentPage_5__6, currentPage_5__5, 
         currentPage_5__4, currentPage_5__3, currentPage_5__2, currentPage_5__1, 
         currentPage_5__0, currentPage_6__15, currentPage_6__14, 
         currentPage_6__13, currentPage_6__12, currentPage_6__11, 
         currentPage_6__10, currentPage_6__9, currentPage_6__8, currentPage_6__7, 
         currentPage_6__6, currentPage_6__5, currentPage_6__4, currentPage_6__3, 
         currentPage_6__2, currentPage_6__1, currentPage_6__0, currentPage_7__15, 
         currentPage_7__14, currentPage_7__13, currentPage_7__12, 
         currentPage_7__11, currentPage_7__10, currentPage_7__9, 
         currentPage_7__8, currentPage_7__7, currentPage_7__6, currentPage_7__5, 
         currentPage_7__4, currentPage_7__3, currentPage_7__2, currentPage_7__1, 
         currentPage_7__0, currentPage_8__15, currentPage_8__14, 
         currentPage_8__13, currentPage_8__12, currentPage_8__11, 
         currentPage_8__10, currentPage_8__9, currentPage_8__8, currentPage_8__7, 
         currentPage_8__6, currentPage_8__5, currentPage_8__4, currentPage_8__3, 
         currentPage_8__2, currentPage_8__1, currentPage_8__0, currentPage_9__15, 
         currentPage_9__14, currentPage_9__13, currentPage_9__12, 
         currentPage_9__11, currentPage_9__10, currentPage_9__9, 
         currentPage_9__8, currentPage_9__7, currentPage_9__6, currentPage_9__5, 
         currentPage_9__4, currentPage_9__3, currentPage_9__2, currentPage_9__1, 
         currentPage_9__0, currentPage_10__15, currentPage_10__14, 
         currentPage_10__13, currentPage_10__12, currentPage_10__11, 
         currentPage_10__10, currentPage_10__9, currentPage_10__8, 
         currentPage_10__7, currentPage_10__6, currentPage_10__5, 
         currentPage_10__4, currentPage_10__3, currentPage_10__2, 
         currentPage_10__1, currentPage_10__0, currentPage_11__15, 
         currentPage_11__14, currentPage_11__13, currentPage_11__12, 
         currentPage_11__11, currentPage_11__10, currentPage_11__9, 
         currentPage_11__8, currentPage_11__7, currentPage_11__6, 
         currentPage_11__5, currentPage_11__4, currentPage_11__3, 
         currentPage_11__2, currentPage_11__1, currentPage_11__0, 
         currentPage_12__15, currentPage_12__14, currentPage_12__13, 
         currentPage_12__12, currentPage_12__11, currentPage_12__10, 
         currentPage_12__9, currentPage_12__8, currentPage_12__7, 
         currentPage_12__6, currentPage_12__5, currentPage_12__4, 
         currentPage_12__3, currentPage_12__2, currentPage_12__1, 
         currentPage_12__0, currentPage_13__15, currentPage_13__14, 
         currentPage_13__13, currentPage_13__12, currentPage_13__11, 
         currentPage_13__10, currentPage_13__9, currentPage_13__8, 
         currentPage_13__7, currentPage_13__6, currentPage_13__5, 
         currentPage_13__4, currentPage_13__3, currentPage_13__2, 
         currentPage_13__1, currentPage_13__0, currentPage_14__15, 
         currentPage_14__14, currentPage_14__13, currentPage_14__12, 
         currentPage_14__11, currentPage_14__10, currentPage_14__9, 
         currentPage_14__8, currentPage_14__7, currentPage_14__6, 
         currentPage_14__5, currentPage_14__4, currentPage_14__3, 
         currentPage_14__2, currentPage_14__1, currentPage_14__0, 
         currentPage_15__15, currentPage_15__14, currentPage_15__13, 
         currentPage_15__12, currentPage_15__11, currentPage_15__10, 
         currentPage_15__9, currentPage_15__8, currentPage_15__7, 
         currentPage_15__6, currentPage_15__5, currentPage_15__4, 
         currentPage_15__3, currentPage_15__2, currentPage_15__1, 
         currentPage_15__0, currentPage_16__15, currentPage_16__14, 
         currentPage_16__13, currentPage_16__12, currentPage_16__11, 
         currentPage_16__10, currentPage_16__9, currentPage_16__8, 
         currentPage_16__7, currentPage_16__6, currentPage_16__5, 
         currentPage_16__4, currentPage_16__3, currentPage_16__2, 
         currentPage_16__1, currentPage_16__0, currentPage_17__15, 
         currentPage_17__14, currentPage_17__13, currentPage_17__12, 
         currentPage_17__11, currentPage_17__10, currentPage_17__9, 
         currentPage_17__8, currentPage_17__7, currentPage_17__6, 
         currentPage_17__5, currentPage_17__4, currentPage_17__3, 
         currentPage_17__2, currentPage_17__1, currentPage_17__0, 
         currentPage_18__15, currentPage_18__14, currentPage_18__13, 
         currentPage_18__12, currentPage_18__11, currentPage_18__10, 
         currentPage_18__9, currentPage_18__8, currentPage_18__7, 
         currentPage_18__6, currentPage_18__5, currentPage_18__4, 
         currentPage_18__3, currentPage_18__2, currentPage_18__1, 
         currentPage_18__0, currentPage_19__15, currentPage_19__14, 
         currentPage_19__13, currentPage_19__12, currentPage_19__11, 
         currentPage_19__10, currentPage_19__9, currentPage_19__8, 
         currentPage_19__7, currentPage_19__6, currentPage_19__5, 
         currentPage_19__4, currentPage_19__3, currentPage_19__2, 
         currentPage_19__1, currentPage_19__0, currentPage_20__15, 
         currentPage_20__14, currentPage_20__13, currentPage_20__12, 
         currentPage_20__11, currentPage_20__10, currentPage_20__9, 
         currentPage_20__8, currentPage_20__7, currentPage_20__6, 
         currentPage_20__5, currentPage_20__4, currentPage_20__3, 
         currentPage_20__2, currentPage_20__1, currentPage_20__0, 
         currentPage_21__15, currentPage_21__14, currentPage_21__13, 
         currentPage_21__12, currentPage_21__11, currentPage_21__10, 
         currentPage_21__9, currentPage_21__8, currentPage_21__7, 
         currentPage_21__6, currentPage_21__5, currentPage_21__4, 
         currentPage_21__3, currentPage_21__2, currentPage_21__1, 
         currentPage_21__0, currentPage_22__15, currentPage_22__14, 
         currentPage_22__13, currentPage_22__12, currentPage_22__11, 
         currentPage_22__10, currentPage_22__9, currentPage_22__8, 
         currentPage_22__7, currentPage_22__6, currentPage_22__5, 
         currentPage_22__4, currentPage_22__3, currentPage_22__2, 
         currentPage_22__1, currentPage_22__0, currentPage_23__15, 
         currentPage_23__14, currentPage_23__13, currentPage_23__12, 
         currentPage_23__11, currentPage_23__10, currentPage_23__9, 
         currentPage_23__8, currentPage_23__7, currentPage_23__6, 
         currentPage_23__5, currentPage_23__4, currentPage_23__3, 
         currentPage_23__2, currentPage_23__1, currentPage_23__0, 
         currentPage_24__15, currentPage_24__14, currentPage_24__13, 
         currentPage_24__12, currentPage_24__11, currentPage_24__10, 
         currentPage_24__9, currentPage_24__8, currentPage_24__7, 
         currentPage_24__6, currentPage_24__5, currentPage_24__4, 
         currentPage_24__3, currentPage_24__2, currentPage_24__1, 
         currentPage_24__0, outMuls_0__15, outMuls_0__14, outMuls_0__13, 
         outMuls_0__12, outMuls_0__11, outMuls_0__10, outMuls_0__9, outMuls_0__8, 
         outMuls_0__7, outMuls_0__6, outMuls_0__5, outMuls_0__4, outMuls_0__3, 
         outMuls_0__2, outMuls_0__1, outMuls_0__0, outMuls_1__15, outMuls_1__14, 
         outMuls_1__13, outMuls_1__12, outMuls_1__11, outMuls_1__10, 
         outMuls_1__9, outMuls_1__8, outMuls_1__7, outMuls_1__6, outMuls_1__5, 
         outMuls_1__4, outMuls_1__3, outMuls_1__2, outMuls_1__1, outMuls_1__0, 
         outMuls_2__15, outMuls_2__14, outMuls_2__13, outMuls_2__12, 
         outMuls_2__11, outMuls_2__10, outMuls_2__9, outMuls_2__8, outMuls_2__7, 
         outMuls_2__6, outMuls_2__5, outMuls_2__4, outMuls_2__3, outMuls_2__2, 
         outMuls_2__1, outMuls_2__0, outMuls_3__15, outMuls_3__14, outMuls_3__13, 
         outMuls_3__12, outMuls_3__11, outMuls_3__10, outMuls_3__9, outMuls_3__8, 
         outMuls_3__7, outMuls_3__6, outMuls_3__5, outMuls_3__4, outMuls_3__3, 
         outMuls_3__2, outMuls_3__1, outMuls_3__0, outMuls_4__15, outMuls_4__14, 
         outMuls_4__13, outMuls_4__12, outMuls_4__11, outMuls_4__10, 
         outMuls_4__9, outMuls_4__8, outMuls_4__7, outMuls_4__6, outMuls_4__5, 
         outMuls_4__4, outMuls_4__3, outMuls_4__2, outMuls_4__1, outMuls_4__0, 
         outMuls_5__15, outMuls_5__14, outMuls_5__13, outMuls_5__12, 
         outMuls_5__11, outMuls_5__10, outMuls_5__9, outMuls_5__8, outMuls_5__7, 
         outMuls_5__6, outMuls_5__5, outMuls_5__4, outMuls_5__3, outMuls_5__2, 
         outMuls_5__1, outMuls_5__0, outMuls_6__15, outMuls_6__14, outMuls_6__13, 
         outMuls_6__12, outMuls_6__11, outMuls_6__10, outMuls_6__9, outMuls_6__8, 
         outMuls_6__7, outMuls_6__6, outMuls_6__5, outMuls_6__4, outMuls_6__3, 
         outMuls_6__2, outMuls_6__1, outMuls_6__0, outMuls_7__15, outMuls_7__14, 
         outMuls_7__13, outMuls_7__12, outMuls_7__11, outMuls_7__10, 
         outMuls_7__9, outMuls_7__8, outMuls_7__7, outMuls_7__6, outMuls_7__5, 
         outMuls_7__4, outMuls_7__3, outMuls_7__2, outMuls_7__1, outMuls_7__0, 
         outMuls_8__15, outMuls_8__14, outMuls_8__13, outMuls_8__12, 
         outMuls_8__11, outMuls_8__10, outMuls_8__9, outMuls_8__8, outMuls_8__7, 
         outMuls_8__6, outMuls_8__5, outMuls_8__4, outMuls_8__3, outMuls_8__2, 
         outMuls_8__1, outMuls_8__0, outMuls_9__15, outMuls_9__14, outMuls_9__13, 
         outMuls_9__12, outMuls_9__11, outMuls_9__10, outMuls_9__9, outMuls_9__8, 
         outMuls_9__7, outMuls_9__6, outMuls_9__5, outMuls_9__4, outMuls_9__3, 
         outMuls_9__2, outMuls_9__1, outMuls_9__0, outMuls_10__15, 
         outMuls_10__14, outMuls_10__13, outMuls_10__12, outMuls_10__11, 
         outMuls_10__10, outMuls_10__9, outMuls_10__8, outMuls_10__7, 
         outMuls_10__6, outMuls_10__5, outMuls_10__4, outMuls_10__3, 
         outMuls_10__2, outMuls_10__1, outMuls_10__0, outMuls_11__15, 
         outMuls_11__14, outMuls_11__13, outMuls_11__12, outMuls_11__11, 
         outMuls_11__10, outMuls_11__9, outMuls_11__8, outMuls_11__7, 
         outMuls_11__6, outMuls_11__5, outMuls_11__4, outMuls_11__3, 
         outMuls_11__2, outMuls_11__1, outMuls_11__0, outMuls_12__15, 
         outMuls_12__14, outMuls_12__13, outMuls_12__12, outMuls_12__11, 
         outMuls_12__10, outMuls_12__9, outMuls_12__8, outMuls_12__7, 
         outMuls_12__6, outMuls_12__5, outMuls_12__4, outMuls_12__3, 
         outMuls_12__2, outMuls_12__1, outMuls_12__0, outMuls_13__15, 
         outMuls_13__14, outMuls_13__13, outMuls_13__12, outMuls_13__11, 
         outMuls_13__10, outMuls_13__9, outMuls_13__8, outMuls_13__7, 
         outMuls_13__6, outMuls_13__5, outMuls_13__4, outMuls_13__3, 
         outMuls_13__2, outMuls_13__1, outMuls_13__0, outMuls_14__15, 
         outMuls_14__14, outMuls_14__13, outMuls_14__12, outMuls_14__11, 
         outMuls_14__10, outMuls_14__9, outMuls_14__8, outMuls_14__7, 
         outMuls_14__6, outMuls_14__5, outMuls_14__4, outMuls_14__3, 
         outMuls_14__2, outMuls_14__1, outMuls_14__0, outMuls_15__15, 
         outMuls_15__14, outMuls_15__13, outMuls_15__12, outMuls_15__11, 
         outMuls_15__10, outMuls_15__9, outMuls_15__8, outMuls_15__7, 
         outMuls_15__6, outMuls_15__5, outMuls_15__4, outMuls_15__3, 
         outMuls_15__2, outMuls_15__1, outMuls_15__0, outMuls_16__15, 
         outMuls_16__14, outMuls_16__13, outMuls_16__12, outMuls_16__11, 
         outMuls_16__10, outMuls_16__9, outMuls_16__8, outMuls_16__7, 
         outMuls_16__6, outMuls_16__5, outMuls_16__4, outMuls_16__3, 
         outMuls_16__2, outMuls_16__1, outMuls_16__0, outMuls_17__15, 
         outMuls_17__14, outMuls_17__13, outMuls_17__12, outMuls_17__11, 
         outMuls_17__10, outMuls_17__9, outMuls_17__8, outMuls_17__7, 
         outMuls_17__6, outMuls_17__5, outMuls_17__4, outMuls_17__3, 
         outMuls_17__2, outMuls_17__1, outMuls_17__0, outMuls_18__15, 
         outMuls_18__14, outMuls_18__13, outMuls_18__12, outMuls_18__11, 
         outMuls_18__10, outMuls_18__9, outMuls_18__8, outMuls_18__7, 
         outMuls_18__6, outMuls_18__5, outMuls_18__4, outMuls_18__3, 
         outMuls_18__2, outMuls_18__1, outMuls_18__0, outMuls_19__15, 
         outMuls_19__14, outMuls_19__13, outMuls_19__12, outMuls_19__11, 
         outMuls_19__10, outMuls_19__9, outMuls_19__8, outMuls_19__7, 
         outMuls_19__6, outMuls_19__5, outMuls_19__4, outMuls_19__3, 
         outMuls_19__2, outMuls_19__1, outMuls_19__0, outMuls_20__15, 
         outMuls_20__14, outMuls_20__13, outMuls_20__12, outMuls_20__11, 
         outMuls_20__10, outMuls_20__9, outMuls_20__8, outMuls_20__7, 
         outMuls_20__6, outMuls_20__5, outMuls_20__4, outMuls_20__3, 
         outMuls_20__2, outMuls_20__1, outMuls_20__0, outMuls_21__15, 
         outMuls_21__14, outMuls_21__13, outMuls_21__12, outMuls_21__11, 
         outMuls_21__10, outMuls_21__9, outMuls_21__8, outMuls_21__7, 
         outMuls_21__6, outMuls_21__5, outMuls_21__4, outMuls_21__3, 
         outMuls_21__2, outMuls_21__1, outMuls_21__0, outMuls_22__15, 
         outMuls_22__14, outMuls_22__13, outMuls_22__12, outMuls_22__11, 
         outMuls_22__10, outMuls_22__9, outMuls_22__8, outMuls_22__7, 
         outMuls_22__6, outMuls_22__5, outMuls_22__4, outMuls_22__3, 
         outMuls_22__2, outMuls_22__1, outMuls_22__0, outMuls_23__15, 
         outMuls_23__14, outMuls_23__13, outMuls_23__12, outMuls_23__11, 
         outMuls_23__10, outMuls_23__9, outMuls_23__8, outMuls_23__7, 
         outMuls_23__6, outMuls_23__5, outMuls_23__4, outMuls_23__3, 
         outMuls_23__2, outMuls_23__1, outMuls_23__0, outMuls_24__15, 
         outMuls_24__14, outMuls_24__13, outMuls_24__12, outMuls_24__11, 
         outMuls_24__10, outMuls_24__9, outMuls_24__8, outMuls_24__7, 
         outMuls_24__6, outMuls_24__5, outMuls_24__4, outMuls_24__3, 
         outMuls_24__2, outMuls_24__1, outMuls_24__0, addersInputs_0__15, 
         addersInputs_0__14, addersInputs_0__13, addersInputs_0__12, 
         addersInputs_0__11, addersInputs_0__10, addersInputs_0__9, 
         addersInputs_0__8, addersInputs_0__7, addersInputs_0__6, 
         addersInputs_0__5, addersInputs_0__4, addersInputs_0__3, 
         addersInputs_0__2, addersInputs_0__1, addersInputs_0__0, 
         addersInputs_1__15, addersInputs_1__14, addersInputs_1__13, 
         addersInputs_1__12, addersInputs_1__11, addersInputs_1__10, 
         addersInputs_1__9, addersInputs_1__8, addersInputs_1__7, 
         addersInputs_1__6, addersInputs_1__5, addersInputs_1__4, 
         addersInputs_1__3, addersInputs_1__2, addersInputs_1__1, 
         addersInputs_1__0, addersInputs_2__15, addersInputs_2__14, 
         addersInputs_2__13, addersInputs_2__12, addersInputs_2__11, 
         addersInputs_2__10, addersInputs_2__9, addersInputs_2__8, 
         addersInputs_2__7, addersInputs_2__6, addersInputs_2__5, 
         addersInputs_2__4, addersInputs_2__3, addersInputs_2__2, 
         addersInputs_2__1, addersInputs_2__0, addersInputs_3__15, 
         addersInputs_3__14, addersInputs_3__13, addersInputs_3__12, 
         addersInputs_3__11, addersInputs_3__10, addersInputs_3__9, 
         addersInputs_3__8, addersInputs_3__7, addersInputs_3__6, 
         addersInputs_3__5, addersInputs_3__4, addersInputs_3__3, 
         addersInputs_3__2, addersInputs_3__1, addersInputs_3__0, 
         addersInputs_4__15, addersInputs_4__14, addersInputs_4__13, 
         addersInputs_4__12, addersInputs_4__11, addersInputs_4__10, 
         addersInputs_4__9, addersInputs_4__8, addersInputs_4__7, 
         addersInputs_4__6, addersInputs_4__5, addersInputs_4__4, 
         addersInputs_4__3, addersInputs_4__2, addersInputs_4__1, 
         addersInputs_4__0, addersInputs_5__15, addersInputs_5__14, 
         addersInputs_5__13, addersInputs_5__12, addersInputs_5__11, 
         addersInputs_5__10, addersInputs_5__9, addersInputs_5__8, 
         addersInputs_5__7, addersInputs_5__6, addersInputs_5__5, 
         addersInputs_5__4, addersInputs_5__3, addersInputs_5__2, 
         addersInputs_5__1, addersInputs_5__0, addersInputs_6__15, 
         addersInputs_6__14, addersInputs_6__13, addersInputs_6__12, 
         addersInputs_6__11, addersInputs_6__10, addersInputs_6__9, 
         addersInputs_6__8, addersInputs_6__7, addersInputs_6__6, 
         addersInputs_6__5, addersInputs_6__4, addersInputs_6__3, 
         addersInputs_6__2, addersInputs_6__1, addersInputs_6__0, 
         addersInputs_7__15, addersInputs_7__14, addersInputs_7__13, 
         addersInputs_7__12, addersInputs_7__11, addersInputs_7__10, 
         addersInputs_7__9, addersInputs_7__8, addersInputs_7__7, 
         addersInputs_7__6, addersInputs_7__5, addersInputs_7__4, 
         addersInputs_7__3, addersInputs_7__2, addersInputs_7__1, 
         addersInputs_7__0, addersInputs_8__15, addersInputs_8__14, 
         addersInputs_8__13, addersInputs_8__12, addersInputs_8__11, 
         addersInputs_8__10, addersInputs_8__9, addersInputs_8__8, 
         addersInputs_8__7, addersInputs_8__6, addersInputs_8__5, 
         addersInputs_8__4, addersInputs_8__3, addersInputs_8__2, 
         addersInputs_8__1, addersInputs_8__0, addersInputs_9__15, 
         addersInputs_9__14, addersInputs_9__13, addersInputs_9__12, 
         addersInputs_9__11, addersInputs_9__10, addersInputs_9__9, 
         addersInputs_9__8, addersInputs_9__7, addersInputs_9__6, 
         addersInputs_9__5, addersInputs_9__4, addersInputs_9__3, 
         addersInputs_9__2, addersInputs_9__1, addersInputs_9__0, 
         addersInputs_10__15, addersInputs_10__14, addersInputs_10__13, 
         addersInputs_10__12, addersInputs_10__11, addersInputs_10__10, 
         addersInputs_10__9, addersInputs_10__8, addersInputs_10__7, 
         addersInputs_10__6, addersInputs_10__5, addersInputs_10__4, 
         addersInputs_10__3, addersInputs_10__2, addersInputs_10__1, 
         addersInputs_10__0, addersInputs_11__15, addersInputs_11__14, 
         addersInputs_11__13, addersInputs_11__12, addersInputs_11__11, 
         addersInputs_11__10, addersInputs_11__9, addersInputs_11__8, 
         addersInputs_11__7, addersInputs_11__6, addersInputs_11__5, 
         addersInputs_11__4, addersInputs_11__3, addersInputs_11__2, 
         addersInputs_11__1, addersInputs_11__0, addersInputs_12__15, 
         addersInputs_12__14, addersInputs_12__13, addersInputs_12__12, 
         addersInputs_12__11, addersInputs_12__10, addersInputs_12__9, 
         addersInputs_12__8, addersInputs_12__7, addersInputs_12__6, 
         addersInputs_12__5, addersInputs_12__4, addersInputs_12__3, 
         addersInputs_12__2, addersInputs_12__1, addersInputs_12__0, 
         addersInputs_13__15, addersInputs_13__14, addersInputs_13__13, 
         addersInputs_13__12, addersInputs_13__11, addersInputs_13__10, 
         addersInputs_13__9, addersInputs_13__8, addersInputs_13__7, 
         addersInputs_13__6, addersInputs_13__5, addersInputs_13__4, 
         addersInputs_13__3, addersInputs_13__2, addersInputs_13__1, 
         addersInputs_13__0, addersInputs_14__15, addersInputs_14__14, 
         addersInputs_14__13, addersInputs_14__12, addersInputs_14__11, 
         addersInputs_14__10, addersInputs_14__9, addersInputs_14__8, 
         addersInputs_14__7, addersInputs_14__6, addersInputs_14__5, 
         addersInputs_14__4, addersInputs_14__3, addersInputs_14__2, 
         addersInputs_14__1, addersInputs_14__0, addersInputs_15__15, 
         addersInputs_15__14, addersInputs_15__13, addersInputs_15__12, 
         addersInputs_15__11, addersInputs_15__10, addersInputs_15__9, 
         addersInputs_15__8, addersInputs_15__7, addersInputs_15__6, 
         addersInputs_15__5, addersInputs_15__4, addersInputs_15__3, 
         addersInputs_15__2, addersInputs_15__1, addersInputs_15__0, 
         addersInputs_16__15, addersInputs_16__14, addersInputs_16__13, 
         addersInputs_16__12, addersInputs_16__11, addersInputs_16__10, 
         addersInputs_16__9, addersInputs_16__8, addersInputs_16__7, 
         addersInputs_16__6, addersInputs_16__5, addersInputs_16__4, 
         addersInputs_16__3, addersInputs_16__2, addersInputs_16__1, 
         addersInputs_16__0, addersInputs_17__15, addersInputs_17__14, 
         addersInputs_17__13, addersInputs_17__12, addersInputs_17__11, 
         addersInputs_17__10, addersInputs_17__9, addersInputs_17__8, 
         addersInputs_17__7, addersInputs_17__6, addersInputs_17__5, 
         addersInputs_17__4, addersInputs_17__3, addersInputs_17__2, 
         addersInputs_17__1, addersInputs_17__0, addersInputs_18__15, 
         addersInputs_18__14, addersInputs_18__13, addersInputs_18__12, 
         addersInputs_18__11, addersInputs_18__10, addersInputs_18__9, 
         addersInputs_18__8, addersInputs_18__7, addersInputs_18__6, 
         addersInputs_18__5, addersInputs_18__4, addersInputs_18__3, 
         addersInputs_18__2, addersInputs_18__1, addersInputs_18__0, 
         addersInputs_19__15, addersInputs_19__14, addersInputs_19__13, 
         addersInputs_19__12, addersInputs_19__11, addersInputs_19__10, 
         addersInputs_19__9, addersInputs_19__8, addersInputs_19__7, 
         addersInputs_19__6, addersInputs_19__5, addersInputs_19__4, 
         addersInputs_19__3, addersInputs_19__2, addersInputs_19__1, 
         addersInputs_19__0, addersInputs_20__15, addersInputs_20__14, 
         addersInputs_20__13, addersInputs_20__12, addersInputs_20__11, 
         addersInputs_20__10, addersInputs_20__9, addersInputs_20__8, 
         addersInputs_20__7, addersInputs_20__6, addersInputs_20__5, 
         addersInputs_20__4, addersInputs_20__3, addersInputs_20__2, 
         addersInputs_20__1, addersInputs_20__0, addersInputs_21__15, 
         addersInputs_21__14, addersInputs_21__13, addersInputs_21__12, 
         addersInputs_21__11, addersInputs_21__10, addersInputs_21__9, 
         addersInputs_21__8, addersInputs_21__7, addersInputs_21__6, 
         addersInputs_21__5, addersInputs_21__4, addersInputs_21__3, 
         addersInputs_21__2, addersInputs_21__1, addersInputs_21__0, 
         addersInputs_22__15, addersInputs_22__14, addersInputs_22__13, 
         addersInputs_22__12, addersInputs_22__11, addersInputs_22__10, 
         addersInputs_22__9, addersInputs_22__8, addersInputs_22__7, 
         addersInputs_22__6, addersInputs_22__5, addersInputs_22__4, 
         addersInputs_22__3, addersInputs_22__2, addersInputs_22__1, 
         addersInputs_22__0, addersInputs_23__15, addersInputs_23__14, 
         addersInputs_23__13, addersInputs_23__12, addersInputs_23__11, 
         addersInputs_23__10, addersInputs_23__9, addersInputs_23__8, 
         addersInputs_23__7, addersInputs_23__6, addersInputs_23__5, 
         addersInputs_23__4, addersInputs_23__3, addersInputs_23__2, 
         addersInputs_23__1, addersInputs_23__0, addersInputs_24__15, 
         addersInputs_24__14, addersInputs_24__13, addersInputs_24__12, 
         addersInputs_24__11, addersInputs_24__10, addersInputs_24__9, 
         addersInputs_24__8, addersInputs_24__7, addersInputs_24__6, 
         addersInputs_24__5, addersInputs_24__4, addersInputs_24__3, 
         addersInputs_24__2, addersInputs_24__1, addersInputs_24__0, filter_0__7, 
         filter_0__6, filter_0__5, filter_0__4, filter_0__3, filter_0__2, 
         filter_0__1, filter_0__0, filter_1__7, filter_1__6, filter_1__5, 
         filter_1__4, filter_1__3, filter_1__2, filter_1__1, filter_1__0, 
         filter_2__7, filter_2__6, filter_2__5, filter_2__4, filter_2__3, 
         filter_2__2, filter_2__1, filter_2__0, filter_3__7, filter_3__6, 
         filter_3__5, filter_3__4, filter_3__3, filter_3__2, filter_3__1, 
         filter_3__0, filter_4__7, filter_4__6, filter_4__5, filter_4__4, 
         filter_4__3, filter_4__2, filter_4__1, filter_4__0, filter_5__7, 
         filter_5__6, filter_5__5, filter_5__4, filter_5__3, filter_5__2, 
         filter_5__1, filter_5__0, filter_6__7, filter_6__6, filter_6__5, 
         filter_6__4, filter_6__3, filter_6__2, filter_6__1, filter_6__0, 
         filter_7__7, filter_7__6, filter_7__5, filter_7__4, filter_7__3, 
         filter_7__2, filter_7__1, filter_7__0, filter_8__7, filter_8__6, 
         filter_8__5, filter_8__4, filter_8__3, filter_8__2, filter_8__1, 
         filter_8__0, filter_9__7, filter_9__6, filter_9__5, filter_9__4, 
         filter_9__3, filter_9__2, filter_9__1, filter_9__0, filter_10__7, 
         filter_10__6, filter_10__5, filter_10__4, filter_10__3, filter_10__2, 
         filter_10__1, filter_10__0, filter_11__7, filter_11__6, filter_11__5, 
         filter_11__4, filter_11__3, filter_11__2, filter_11__1, filter_11__0, 
         filter_12__7, filter_12__6, filter_12__5, filter_12__4, filter_12__3, 
         filter_12__2, filter_12__1, filter_12__0, filter_13__7, filter_13__6, 
         filter_13__5, filter_13__4, filter_13__3, filter_13__2, filter_13__1, 
         filter_13__0, filter_14__7, filter_14__6, filter_14__5, filter_14__4, 
         filter_14__3, filter_14__2, filter_14__1, filter_14__0, filter_15__7, 
         filter_15__6, filter_15__5, filter_15__4, filter_15__3, filter_15__2, 
         filter_15__1, filter_15__0, filter_16__7, filter_16__6, filter_16__5, 
         filter_16__4, filter_16__3, filter_16__2, filter_16__1, filter_16__0, 
         filter_17__7, filter_17__6, filter_17__5, filter_17__4, filter_17__3, 
         filter_17__2, filter_17__1, filter_17__0, filter_18__7, filter_18__6, 
         filter_18__5, filter_18__4, filter_18__3, filter_18__2, filter_18__1, 
         filter_18__0, filter_19__7, filter_19__6, filter_19__5, filter_19__4, 
         filter_19__3, filter_19__2, filter_19__1, filter_19__0, filter_20__7, 
         filter_20__6, filter_20__5, filter_20__4, filter_20__3, filter_20__2, 
         filter_20__1, filter_20__0, filter_21__7, filter_21__6, filter_21__5, 
         filter_21__4, filter_21__3, filter_21__2, filter_21__1, filter_21__0, 
         filter_22__7, filter_22__6, filter_22__5, filter_22__4, filter_22__3, 
         filter_22__2, filter_22__1, filter_22__0, filter_23__7, filter_23__6, 
         filter_23__5, filter_23__4, filter_23__3, filter_23__2, filter_23__1, 
         filter_23__0, filter_24__7, filter_24__6, filter_24__5, filter_24__4, 
         filter_24__3, filter_24__2, filter_24__1, filter_24__0, doneMul, 
         regFileMap_page1Out_5__15, regFileMap_page1Out_5__14, 
         regFileMap_page1Out_5__13, regFileMap_page1Out_5__12, 
         regFileMap_page1Out_5__11, regFileMap_page1Out_5__10, 
         regFileMap_page1Out_5__9, regFileMap_page1Out_5__8, 
         regFileMap_page1Out_5__7, regFileMap_page1Out_5__6, 
         regFileMap_page1Out_5__5, regFileMap_page1Out_5__4, 
         regFileMap_page1Out_5__3, regFileMap_page1Out_5__2, 
         regFileMap_page1Out_5__1, regFileMap_page1Out_5__0, 
         regFileMap_page1Out_6__15, regFileMap_page1Out_6__14, 
         regFileMap_page1Out_6__13, regFileMap_page1Out_6__12, 
         regFileMap_page1Out_6__11, regFileMap_page1Out_6__10, 
         regFileMap_page1Out_6__9, regFileMap_page1Out_6__8, 
         regFileMap_page1Out_6__7, regFileMap_page1Out_6__6, 
         regFileMap_page1Out_6__5, regFileMap_page1Out_6__4, 
         regFileMap_page1Out_6__3, regFileMap_page1Out_6__2, 
         regFileMap_page1Out_6__1, regFileMap_page1Out_6__0, 
         regFileMap_page1Out_7__15, regFileMap_page1Out_7__14, 
         regFileMap_page1Out_7__13, regFileMap_page1Out_7__12, 
         regFileMap_page1Out_7__11, regFileMap_page1Out_7__10, 
         regFileMap_page1Out_7__9, regFileMap_page1Out_7__8, 
         regFileMap_page1Out_7__7, regFileMap_page1Out_7__6, 
         regFileMap_page1Out_7__5, regFileMap_page1Out_7__4, 
         regFileMap_page1Out_7__3, regFileMap_page1Out_7__2, 
         regFileMap_page1Out_7__1, regFileMap_page1Out_7__0, 
         regFileMap_page1Out_8__15, regFileMap_page1Out_8__14, 
         regFileMap_page1Out_8__13, regFileMap_page1Out_8__12, 
         regFileMap_page1Out_8__11, regFileMap_page1Out_8__10, 
         regFileMap_page1Out_8__9, regFileMap_page1Out_8__8, 
         regFileMap_page1Out_8__7, regFileMap_page1Out_8__6, 
         regFileMap_page1Out_8__5, regFileMap_page1Out_8__4, 
         regFileMap_page1Out_8__3, regFileMap_page1Out_8__2, 
         regFileMap_page1Out_8__1, regFileMap_page1Out_8__0, 
         regFileMap_page1Out_9__15, regFileMap_page1Out_9__14, 
         regFileMap_page1Out_9__13, regFileMap_page1Out_9__12, 
         regFileMap_page1Out_9__11, regFileMap_page1Out_9__10, 
         regFileMap_page1Out_9__9, regFileMap_page1Out_9__8, 
         regFileMap_page1Out_9__7, regFileMap_page1Out_9__6, 
         regFileMap_page1Out_9__5, regFileMap_page1Out_9__4, 
         regFileMap_page1Out_9__3, regFileMap_page1Out_9__2, 
         regFileMap_page1Out_9__1, regFileMap_page1Out_9__0, 
         regFileMap_page1Out_10__15, regFileMap_page1Out_10__14, 
         regFileMap_page1Out_10__13, regFileMap_page1Out_10__12, 
         regFileMap_page1Out_10__11, regFileMap_page1Out_10__10, 
         regFileMap_page1Out_10__9, regFileMap_page1Out_10__8, 
         regFileMap_page1Out_10__7, regFileMap_page1Out_10__6, 
         regFileMap_page1Out_10__5, regFileMap_page1Out_10__4, 
         regFileMap_page1Out_10__3, regFileMap_page1Out_10__2, 
         regFileMap_page1Out_10__1, regFileMap_page1Out_10__0, 
         regFileMap_page1Out_11__15, regFileMap_page1Out_11__14, 
         regFileMap_page1Out_11__13, regFileMap_page1Out_11__12, 
         regFileMap_page1Out_11__11, regFileMap_page1Out_11__10, 
         regFileMap_page1Out_11__9, regFileMap_page1Out_11__8, 
         regFileMap_page1Out_11__7, regFileMap_page1Out_11__6, 
         regFileMap_page1Out_11__5, regFileMap_page1Out_11__4, 
         regFileMap_page1Out_11__3, regFileMap_page1Out_11__2, 
         regFileMap_page1Out_11__1, regFileMap_page1Out_11__0, 
         regFileMap_page1Out_12__15, regFileMap_page1Out_12__14, 
         regFileMap_page1Out_12__13, regFileMap_page1Out_12__12, 
         regFileMap_page1Out_12__11, regFileMap_page1Out_12__10, 
         regFileMap_page1Out_12__9, regFileMap_page1Out_12__8, 
         regFileMap_page1Out_12__7, regFileMap_page1Out_12__6, 
         regFileMap_page1Out_12__5, regFileMap_page1Out_12__4, 
         regFileMap_page1Out_12__3, regFileMap_page1Out_12__2, 
         regFileMap_page1Out_12__1, regFileMap_page1Out_12__0, 
         regFileMap_page1Out_13__15, regFileMap_page1Out_13__14, 
         regFileMap_page1Out_13__13, regFileMap_page1Out_13__12, 
         regFileMap_page1Out_13__11, regFileMap_page1Out_13__10, 
         regFileMap_page1Out_13__9, regFileMap_page1Out_13__8, 
         regFileMap_page1Out_13__7, regFileMap_page1Out_13__6, 
         regFileMap_page1Out_13__5, regFileMap_page1Out_13__4, 
         regFileMap_page1Out_13__3, regFileMap_page1Out_13__2, 
         regFileMap_page1Out_13__1, regFileMap_page1Out_13__0, 
         regFileMap_page1Out_14__15, regFileMap_page1Out_14__14, 
         regFileMap_page1Out_14__13, regFileMap_page1Out_14__12, 
         regFileMap_page1Out_14__11, regFileMap_page1Out_14__10, 
         regFileMap_page1Out_14__9, regFileMap_page1Out_14__8, 
         regFileMap_page1Out_14__7, regFileMap_page1Out_14__6, 
         regFileMap_page1Out_14__5, regFileMap_page1Out_14__4, 
         regFileMap_page1Out_14__3, regFileMap_page1Out_14__2, 
         regFileMap_page1Out_14__1, regFileMap_page1Out_14__0, 
         regFileMap_page1Out_15__15, regFileMap_page1Out_15__14, 
         regFileMap_page1Out_15__13, regFileMap_page1Out_15__12, 
         regFileMap_page1Out_15__11, regFileMap_page1Out_15__10, 
         regFileMap_page1Out_15__9, regFileMap_page1Out_15__8, 
         regFileMap_page1Out_15__7, regFileMap_page1Out_15__6, 
         regFileMap_page1Out_15__5, regFileMap_page1Out_15__4, 
         regFileMap_page1Out_15__3, regFileMap_page1Out_15__2, 
         regFileMap_page1Out_15__1, regFileMap_page1Out_15__0, 
         regFileMap_page1Out_16__15, regFileMap_page1Out_16__14, 
         regFileMap_page1Out_16__13, regFileMap_page1Out_16__12, 
         regFileMap_page1Out_16__11, regFileMap_page1Out_16__10, 
         regFileMap_page1Out_16__9, regFileMap_page1Out_16__8, 
         regFileMap_page1Out_16__7, regFileMap_page1Out_16__6, 
         regFileMap_page1Out_16__5, regFileMap_page1Out_16__4, 
         regFileMap_page1Out_16__3, regFileMap_page1Out_16__2, 
         regFileMap_page1Out_16__1, regFileMap_page1Out_16__0, 
         regFileMap_page1Out_17__15, regFileMap_page1Out_17__14, 
         regFileMap_page1Out_17__13, regFileMap_page1Out_17__12, 
         regFileMap_page1Out_17__11, regFileMap_page1Out_17__10, 
         regFileMap_page1Out_17__9, regFileMap_page1Out_17__8, 
         regFileMap_page1Out_17__7, regFileMap_page1Out_17__6, 
         regFileMap_page1Out_17__5, regFileMap_page1Out_17__4, 
         regFileMap_page1Out_17__3, regFileMap_page1Out_17__2, 
         regFileMap_page1Out_17__1, regFileMap_page1Out_17__0, 
         regFileMap_page1Out_18__15, regFileMap_page1Out_18__14, 
         regFileMap_page1Out_18__13, regFileMap_page1Out_18__12, 
         regFileMap_page1Out_18__11, regFileMap_page1Out_18__10, 
         regFileMap_page1Out_18__9, regFileMap_page1Out_18__8, 
         regFileMap_page1Out_18__7, regFileMap_page1Out_18__6, 
         regFileMap_page1Out_18__5, regFileMap_page1Out_18__4, 
         regFileMap_page1Out_18__3, regFileMap_page1Out_18__2, 
         regFileMap_page1Out_18__1, regFileMap_page1Out_18__0, 
         regFileMap_page1Out_19__15, regFileMap_page1Out_19__14, 
         regFileMap_page1Out_19__13, regFileMap_page1Out_19__12, 
         regFileMap_page1Out_19__11, regFileMap_page1Out_19__10, 
         regFileMap_page1Out_19__9, regFileMap_page1Out_19__8, 
         regFileMap_page1Out_19__7, regFileMap_page1Out_19__6, 
         regFileMap_page1Out_19__5, regFileMap_page1Out_19__4, 
         regFileMap_page1Out_19__3, regFileMap_page1Out_19__2, 
         regFileMap_page1Out_19__1, regFileMap_page1Out_19__0, 
         regFileMap_page1Out_20__15, regFileMap_page1Out_20__14, 
         regFileMap_page1Out_20__13, regFileMap_page1Out_20__12, 
         regFileMap_page1Out_20__11, regFileMap_page1Out_20__10, 
         regFileMap_page1Out_20__9, regFileMap_page1Out_20__8, 
         regFileMap_page1Out_20__7, regFileMap_page1Out_20__6, 
         regFileMap_page1Out_20__5, regFileMap_page1Out_20__4, 
         regFileMap_page1Out_20__3, regFileMap_page1Out_20__2, 
         regFileMap_page1Out_20__1, regFileMap_page1Out_20__0, 
         regFileMap_page1Out_21__15, regFileMap_page1Out_21__14, 
         regFileMap_page1Out_21__13, regFileMap_page1Out_21__12, 
         regFileMap_page1Out_21__11, regFileMap_page1Out_21__10, 
         regFileMap_page1Out_21__9, regFileMap_page1Out_21__8, 
         regFileMap_page1Out_21__7, regFileMap_page1Out_21__6, 
         regFileMap_page1Out_21__5, regFileMap_page1Out_21__4, 
         regFileMap_page1Out_21__3, regFileMap_page1Out_21__2, 
         regFileMap_page1Out_21__1, regFileMap_page1Out_21__0, 
         regFileMap_page1Out_22__15, regFileMap_page1Out_22__14, 
         regFileMap_page1Out_22__13, regFileMap_page1Out_22__12, 
         regFileMap_page1Out_22__11, regFileMap_page1Out_22__10, 
         regFileMap_page1Out_22__9, regFileMap_page1Out_22__8, 
         regFileMap_page1Out_22__7, regFileMap_page1Out_22__6, 
         regFileMap_page1Out_22__5, regFileMap_page1Out_22__4, 
         regFileMap_page1Out_22__3, regFileMap_page1Out_22__2, 
         regFileMap_page1Out_22__1, regFileMap_page1Out_22__0, 
         regFileMap_page1Out_23__15, regFileMap_page1Out_23__14, 
         regFileMap_page1Out_23__13, regFileMap_page1Out_23__12, 
         regFileMap_page1Out_23__11, regFileMap_page1Out_23__10, 
         regFileMap_page1Out_23__9, regFileMap_page1Out_23__8, 
         regFileMap_page1Out_23__7, regFileMap_page1Out_23__6, 
         regFileMap_page1Out_23__5, regFileMap_page1Out_23__4, 
         regFileMap_page1Out_23__3, regFileMap_page1Out_23__2, 
         regFileMap_page1Out_23__1, regFileMap_page1Out_23__0, 
         regFileMap_page1Out_24__15, regFileMap_page1Out_24__14, 
         regFileMap_page1Out_24__13, regFileMap_page1Out_24__12, 
         regFileMap_page1Out_24__11, regFileMap_page1Out_24__10, 
         regFileMap_page1Out_24__9, regFileMap_page1Out_24__8, 
         regFileMap_page1Out_24__7, regFileMap_page1Out_24__6, 
         regFileMap_page1Out_24__5, regFileMap_page1Out_24__4, 
         regFileMap_page1Out_24__3, regFileMap_page1Out_24__2, 
         regFileMap_page1Out_24__1, regFileMap_page1Out_24__0, 
         regFileMap_page2Out_5__15, regFileMap_page2Out_5__14, 
         regFileMap_page2Out_5__13, regFileMap_page2Out_5__12, 
         regFileMap_page2Out_5__11, regFileMap_page2Out_5__10, 
         regFileMap_page2Out_5__9, regFileMap_page2Out_5__8, 
         regFileMap_page2Out_5__7, regFileMap_page2Out_5__6, 
         regFileMap_page2Out_5__5, regFileMap_page2Out_5__4, 
         regFileMap_page2Out_5__3, regFileMap_page2Out_5__2, 
         regFileMap_page2Out_5__1, regFileMap_page2Out_5__0, 
         regFileMap_page2Out_6__15, regFileMap_page2Out_6__14, 
         regFileMap_page2Out_6__13, regFileMap_page2Out_6__12, 
         regFileMap_page2Out_6__11, regFileMap_page2Out_6__10, 
         regFileMap_page2Out_6__9, regFileMap_page2Out_6__8, 
         regFileMap_page2Out_6__7, regFileMap_page2Out_6__6, 
         regFileMap_page2Out_6__5, regFileMap_page2Out_6__4, 
         regFileMap_page2Out_6__3, regFileMap_page2Out_6__2, 
         regFileMap_page2Out_6__1, regFileMap_page2Out_6__0, 
         regFileMap_page2Out_7__15, regFileMap_page2Out_7__14, 
         regFileMap_page2Out_7__13, regFileMap_page2Out_7__12, 
         regFileMap_page2Out_7__11, regFileMap_page2Out_7__10, 
         regFileMap_page2Out_7__9, regFileMap_page2Out_7__8, 
         regFileMap_page2Out_7__7, regFileMap_page2Out_7__6, 
         regFileMap_page2Out_7__5, regFileMap_page2Out_7__4, 
         regFileMap_page2Out_7__3, regFileMap_page2Out_7__2, 
         regFileMap_page2Out_7__1, regFileMap_page2Out_7__0, 
         regFileMap_page2Out_8__15, regFileMap_page2Out_8__14, 
         regFileMap_page2Out_8__13, regFileMap_page2Out_8__12, 
         regFileMap_page2Out_8__11, regFileMap_page2Out_8__10, 
         regFileMap_page2Out_8__9, regFileMap_page2Out_8__8, 
         regFileMap_page2Out_8__7, regFileMap_page2Out_8__6, 
         regFileMap_page2Out_8__5, regFileMap_page2Out_8__4, 
         regFileMap_page2Out_8__3, regFileMap_page2Out_8__2, 
         regFileMap_page2Out_8__1, regFileMap_page2Out_8__0, 
         regFileMap_page2Out_9__15, regFileMap_page2Out_9__14, 
         regFileMap_page2Out_9__13, regFileMap_page2Out_9__12, 
         regFileMap_page2Out_9__11, regFileMap_page2Out_9__10, 
         regFileMap_page2Out_9__9, regFileMap_page2Out_9__8, 
         regFileMap_page2Out_9__7, regFileMap_page2Out_9__6, 
         regFileMap_page2Out_9__5, regFileMap_page2Out_9__4, 
         regFileMap_page2Out_9__3, regFileMap_page2Out_9__2, 
         regFileMap_page2Out_9__1, regFileMap_page2Out_9__0, 
         regFileMap_page2Out_10__15, regFileMap_page2Out_10__14, 
         regFileMap_page2Out_10__13, regFileMap_page2Out_10__12, 
         regFileMap_page2Out_10__11, regFileMap_page2Out_10__10, 
         regFileMap_page2Out_10__9, regFileMap_page2Out_10__8, 
         regFileMap_page2Out_10__7, regFileMap_page2Out_10__6, 
         regFileMap_page2Out_10__5, regFileMap_page2Out_10__4, 
         regFileMap_page2Out_10__3, regFileMap_page2Out_10__2, 
         regFileMap_page2Out_10__1, regFileMap_page2Out_10__0, 
         regFileMap_page2Out_11__15, regFileMap_page2Out_11__14, 
         regFileMap_page2Out_11__13, regFileMap_page2Out_11__12, 
         regFileMap_page2Out_11__11, regFileMap_page2Out_11__10, 
         regFileMap_page2Out_11__9, regFileMap_page2Out_11__8, 
         regFileMap_page2Out_11__7, regFileMap_page2Out_11__6, 
         regFileMap_page2Out_11__5, regFileMap_page2Out_11__4, 
         regFileMap_page2Out_11__3, regFileMap_page2Out_11__2, 
         regFileMap_page2Out_11__1, regFileMap_page2Out_11__0, 
         regFileMap_page2Out_12__15, regFileMap_page2Out_12__14, 
         regFileMap_page2Out_12__13, regFileMap_page2Out_12__12, 
         regFileMap_page2Out_12__11, regFileMap_page2Out_12__10, 
         regFileMap_page2Out_12__9, regFileMap_page2Out_12__8, 
         regFileMap_page2Out_12__7, regFileMap_page2Out_12__6, 
         regFileMap_page2Out_12__5, regFileMap_page2Out_12__4, 
         regFileMap_page2Out_12__3, regFileMap_page2Out_12__2, 
         regFileMap_page2Out_12__1, regFileMap_page2Out_12__0, 
         regFileMap_page2Out_13__15, regFileMap_page2Out_13__14, 
         regFileMap_page2Out_13__13, regFileMap_page2Out_13__12, 
         regFileMap_page2Out_13__11, regFileMap_page2Out_13__10, 
         regFileMap_page2Out_13__9, regFileMap_page2Out_13__8, 
         regFileMap_page2Out_13__7, regFileMap_page2Out_13__6, 
         regFileMap_page2Out_13__5, regFileMap_page2Out_13__4, 
         regFileMap_page2Out_13__3, regFileMap_page2Out_13__2, 
         regFileMap_page2Out_13__1, regFileMap_page2Out_13__0, 
         regFileMap_page2Out_14__15, regFileMap_page2Out_14__14, 
         regFileMap_page2Out_14__13, regFileMap_page2Out_14__12, 
         regFileMap_page2Out_14__11, regFileMap_page2Out_14__10, 
         regFileMap_page2Out_14__9, regFileMap_page2Out_14__8, 
         regFileMap_page2Out_14__7, regFileMap_page2Out_14__6, 
         regFileMap_page2Out_14__5, regFileMap_page2Out_14__4, 
         regFileMap_page2Out_14__3, regFileMap_page2Out_14__2, 
         regFileMap_page2Out_14__1, regFileMap_page2Out_14__0, 
         regFileMap_page2Out_15__15, regFileMap_page2Out_15__14, 
         regFileMap_page2Out_15__13, regFileMap_page2Out_15__12, 
         regFileMap_page2Out_15__11, regFileMap_page2Out_15__10, 
         regFileMap_page2Out_15__9, regFileMap_page2Out_15__8, 
         regFileMap_page2Out_15__7, regFileMap_page2Out_15__6, 
         regFileMap_page2Out_15__5, regFileMap_page2Out_15__4, 
         regFileMap_page2Out_15__3, regFileMap_page2Out_15__2, 
         regFileMap_page2Out_15__1, regFileMap_page2Out_15__0, 
         regFileMap_page2Out_16__15, regFileMap_page2Out_16__14, 
         regFileMap_page2Out_16__13, regFileMap_page2Out_16__12, 
         regFileMap_page2Out_16__11, regFileMap_page2Out_16__10, 
         regFileMap_page2Out_16__9, regFileMap_page2Out_16__8, 
         regFileMap_page2Out_16__7, regFileMap_page2Out_16__6, 
         regFileMap_page2Out_16__5, regFileMap_page2Out_16__4, 
         regFileMap_page2Out_16__3, regFileMap_page2Out_16__2, 
         regFileMap_page2Out_16__1, regFileMap_page2Out_16__0, 
         regFileMap_page2Out_17__15, regFileMap_page2Out_17__14, 
         regFileMap_page2Out_17__13, regFileMap_page2Out_17__12, 
         regFileMap_page2Out_17__11, regFileMap_page2Out_17__10, 
         regFileMap_page2Out_17__9, regFileMap_page2Out_17__8, 
         regFileMap_page2Out_17__7, regFileMap_page2Out_17__6, 
         regFileMap_page2Out_17__5, regFileMap_page2Out_17__4, 
         regFileMap_page2Out_17__3, regFileMap_page2Out_17__2, 
         regFileMap_page2Out_17__1, regFileMap_page2Out_17__0, 
         regFileMap_page2Out_18__15, regFileMap_page2Out_18__14, 
         regFileMap_page2Out_18__13, regFileMap_page2Out_18__12, 
         regFileMap_page2Out_18__11, regFileMap_page2Out_18__10, 
         regFileMap_page2Out_18__9, regFileMap_page2Out_18__8, 
         regFileMap_page2Out_18__7, regFileMap_page2Out_18__6, 
         regFileMap_page2Out_18__5, regFileMap_page2Out_18__4, 
         regFileMap_page2Out_18__3, regFileMap_page2Out_18__2, 
         regFileMap_page2Out_18__1, regFileMap_page2Out_18__0, 
         regFileMap_page2Out_19__15, regFileMap_page2Out_19__14, 
         regFileMap_page2Out_19__13, regFileMap_page2Out_19__12, 
         regFileMap_page2Out_19__11, regFileMap_page2Out_19__10, 
         regFileMap_page2Out_19__9, regFileMap_page2Out_19__8, 
         regFileMap_page2Out_19__7, regFileMap_page2Out_19__6, 
         regFileMap_page2Out_19__5, regFileMap_page2Out_19__4, 
         regFileMap_page2Out_19__3, regFileMap_page2Out_19__2, 
         regFileMap_page2Out_19__1, regFileMap_page2Out_19__0, 
         regFileMap_page2Out_20__15, regFileMap_page2Out_20__14, 
         regFileMap_page2Out_20__13, regFileMap_page2Out_20__12, 
         regFileMap_page2Out_20__11, regFileMap_page2Out_20__10, 
         regFileMap_page2Out_20__9, regFileMap_page2Out_20__8, 
         regFileMap_page2Out_20__7, regFileMap_page2Out_20__6, 
         regFileMap_page2Out_20__5, regFileMap_page2Out_20__4, 
         regFileMap_page2Out_20__3, regFileMap_page2Out_20__2, 
         regFileMap_page2Out_20__1, regFileMap_page2Out_20__0, 
         regFileMap_page2Out_21__15, regFileMap_page2Out_21__14, 
         regFileMap_page2Out_21__13, regFileMap_page2Out_21__12, 
         regFileMap_page2Out_21__11, regFileMap_page2Out_21__10, 
         regFileMap_page2Out_21__9, regFileMap_page2Out_21__8, 
         regFileMap_page2Out_21__7, regFileMap_page2Out_21__6, 
         regFileMap_page2Out_21__5, regFileMap_page2Out_21__4, 
         regFileMap_page2Out_21__3, regFileMap_page2Out_21__2, 
         regFileMap_page2Out_21__1, regFileMap_page2Out_21__0, 
         regFileMap_page2Out_22__15, regFileMap_page2Out_22__14, 
         regFileMap_page2Out_22__13, regFileMap_page2Out_22__12, 
         regFileMap_page2Out_22__11, regFileMap_page2Out_22__10, 
         regFileMap_page2Out_22__9, regFileMap_page2Out_22__8, 
         regFileMap_page2Out_22__7, regFileMap_page2Out_22__6, 
         regFileMap_page2Out_22__5, regFileMap_page2Out_22__4, 
         regFileMap_page2Out_22__3, regFileMap_page2Out_22__2, 
         regFileMap_page2Out_22__1, regFileMap_page2Out_22__0, 
         regFileMap_page2Out_23__15, regFileMap_page2Out_23__14, 
         regFileMap_page2Out_23__13, regFileMap_page2Out_23__12, 
         regFileMap_page2Out_23__11, regFileMap_page2Out_23__10, 
         regFileMap_page2Out_23__9, regFileMap_page2Out_23__8, 
         regFileMap_page2Out_23__7, regFileMap_page2Out_23__6, 
         regFileMap_page2Out_23__5, regFileMap_page2Out_23__4, 
         regFileMap_page2Out_23__3, regFileMap_page2Out_23__2, 
         regFileMap_page2Out_23__1, regFileMap_page2Out_23__0, 
         regFileMap_page2Out_24__15, regFileMap_page2Out_24__14, 
         regFileMap_page2Out_24__13, regFileMap_page2Out_24__12, 
         regFileMap_page2Out_24__11, regFileMap_page2Out_24__10, 
         regFileMap_page2Out_24__9, regFileMap_page2Out_24__8, 
         regFileMap_page2Out_24__7, regFileMap_page2Out_24__6, 
         regFileMap_page2Out_24__5, regFileMap_page2Out_24__4, 
         regFileMap_page2Out_24__3, regFileMap_page2Out_24__2, 
         regFileMap_page2Out_24__1, regFileMap_page2Out_24__0, 
         regFileMap_page1Enables_0, regFileMap_page1Enables_1, 
         regFileMap_page1Enables_2, regFileMap_page1Enables_3, 
         regFileMap_page1Enables_4, regFileMap_page2Enables_0, 
         regFileMap_page2Enables_1, regFileMap_page2Enables_2, 
         regFileMap_page2Enables_3, regFileMap_page2Enables_4, 
         regFileMap_filterEnables_0, regFileMap_filterEnables_1, 
         regFileMap_filterEnables_2, regFileMap_filterEnables_3, 
         addersMap_sum1_15, addersMap_sum1_14, addersMap_sum1_13, 
         addersMap_sum1_12, addersMap_sum1_11, addersMap_sum1_10, 
         addersMap_sum1_9, addersMap_sum1_8, addersMap_sum1_7, addersMap_sum1_6, 
         addersMap_sum1_5, addersMap_sum1_4, addersMap_sum1_3, addersMap_sum1_2, 
         addersMap_sum1_1, addersMap_sum1_0, addersMap_sum2_15, 
         addersMap_sum2_14, addersMap_sum2_13, addersMap_sum2_12, 
         addersMap_sum2_11, addersMap_sum2_10, addersMap_sum2_9, 
         addersMap_sum2_8, addersMap_sum2_7, addersMap_sum2_6, addersMap_sum2_5, 
         addersMap_sum2_4, addersMap_sum2_3, addersMap_sum2_2, addersMap_sum2_1, 
         addersMap_sum2_0, addersMap_sum3_15, addersMap_sum3_14, 
         addersMap_sum3_13, addersMap_sum3_12, addersMap_sum3_11, 
         addersMap_sum3_10, addersMap_sum3_9, addersMap_sum3_8, addersMap_sum3_7, 
         addersMap_sum3_6, addersMap_sum3_5, addersMap_sum3_4, addersMap_sum3_3, 
         addersMap_sum3_2, addersMap_sum3_1, addersMap_sum3_0, 
         addersMap_sum3Filter_15, addersMap_sum3Filter_14, 
         addersMap_sum3Filter_13, addersMap_sum3Filter_12, 
         addersMap_sum3Filter_11, addersMap_sum3Filter_10, 
         addersMap_sum3Filter_9, addersMap_sum3Filter_8, addersMap_sum3Filter_7, 
         addersMap_sum3Filter_6, addersMap_sum3Filter_5, addersMap_sum3Filter_4, 
         addersMap_sum3Filter_3, addersMap_sum3Filter_2, addersMap_sum3Filter_1, 
         addersMap_sum3Filter_0, addersMap_sum4_15, addersMap_sum4_14, 
         addersMap_sum4_13, addersMap_sum4_12, addersMap_sum4_11, 
         addersMap_sum4_10, addersMap_sum4_9, addersMap_sum4_8, addersMap_sum4_7, 
         addersMap_sum4_6, addersMap_sum4_5, addersMap_sum4_4, addersMap_sum4_3, 
         addersMap_sum4_2, addersMap_sum4_1, addersMap_sum4_0, 
         addersMap_totalSum_15, addersMap_totalSum_14, addersMap_totalSum_13, 
         addersMap_totalSum_12, addersMap_totalSum_11, addersMap_totalSum_10, 
         addersMap_totalSum_9, addersMap_totalSum_8, addersMap_totalSum_7, 
         addersMap_totalSum_6, addersMap_totalSum_5, addersMap_totalSum_4, 
         addersMap_totalSum_3, addersMap_totalSum_2, addersMap_totalSum_1, 
         addersMap_totalSum_0, addersMap_sum1Map_sum1_15__dup_0, 
         addersMap_sum1Map_sum1_14__dup_0, addersMap_sum1Map_sum1_13__dup_0, 
         addersMap_sum1Map_sum1_12__dup_0, addersMap_sum1Map_sum1_11__dup_0, 
         addersMap_sum1Map_sum1_10__dup_0, addersMap_sum1Map_sum1_9__dup_0, 
         addersMap_sum1Map_sum1_8__dup_0, addersMap_sum1Map_sum1_7__dup_0, 
         addersMap_sum1Map_sum1_6__dup_0, addersMap_sum1Map_sum1_5__dup_0, 
         addersMap_sum1Map_sum1_4__dup_0, addersMap_sum1Map_sum1_3__dup_0, 
         addersMap_sum1Map_sum1_2__dup_0, addersMap_sum1Map_sum1_1__dup_0, 
         addersMap_sum1Map_sum1_0__dup_0, addersMap_sum1Map_sum2_15__dup_0, 
         addersMap_sum1Map_sum2_14__dup_0, addersMap_sum1Map_sum2_13__dup_0, 
         addersMap_sum1Map_sum2_12__dup_0, addersMap_sum1Map_sum2_11__dup_0, 
         addersMap_sum1Map_sum2_10__dup_0, addersMap_sum1Map_sum2_9__dup_0, 
         addersMap_sum1Map_sum2_8__dup_0, addersMap_sum1Map_sum2_7__dup_0, 
         addersMap_sum1Map_sum2_6__dup_0, addersMap_sum1Map_sum2_5__dup_0, 
         addersMap_sum1Map_sum2_4__dup_0, addersMap_sum1Map_sum2_3__dup_0, 
         addersMap_sum1Map_sum2_2__dup_0, addersMap_sum1Map_sum2_1__dup_0, 
         addersMap_sum1Map_sum2_0__dup_0, addersMap_sum1Map_sum1Map_sum1_15, 
         addersMap_sum1Map_sum1Map_sum1_14, addersMap_sum1Map_sum1Map_sum1_13, 
         addersMap_sum1Map_sum1Map_sum1_12, addersMap_sum1Map_sum1Map_sum1_11, 
         addersMap_sum1Map_sum1Map_sum1_10, addersMap_sum1Map_sum1Map_sum1_9, 
         addersMap_sum1Map_sum1Map_sum1_8, addersMap_sum1Map_sum1Map_sum1_7, 
         addersMap_sum1Map_sum1Map_sum1_6, addersMap_sum1Map_sum1Map_sum1_5, 
         addersMap_sum1Map_sum1Map_sum1_4, addersMap_sum1Map_sum1Map_sum1_3, 
         addersMap_sum1Map_sum1Map_sum1_2, addersMap_sum1Map_sum1Map_sum1_1, 
         addersMap_sum1Map_sum1Map_sum1_0, addersMap_sum1Map_sum1Map_sum2_15, 
         addersMap_sum1Map_sum1Map_sum2_14, addersMap_sum1Map_sum1Map_sum2_13, 
         addersMap_sum1Map_sum1Map_sum2_12, addersMap_sum1Map_sum1Map_sum2_11, 
         addersMap_sum1Map_sum1Map_sum2_10, addersMap_sum1Map_sum1Map_sum2_9, 
         addersMap_sum1Map_sum1Map_sum2_8, addersMap_sum1Map_sum1Map_sum2_7, 
         addersMap_sum1Map_sum1Map_sum2_6, addersMap_sum1Map_sum1Map_sum2_5, 
         addersMap_sum1Map_sum1Map_sum2_4, addersMap_sum1Map_sum1Map_sum2_3, 
         addersMap_sum1Map_sum1Map_sum2_2, addersMap_sum1Map_sum1Map_sum2_1, 
         addersMap_sum1Map_sum1Map_sum2_0, addersMap_sum1Map_sum2Map_sum1_15, 
         addersMap_sum1Map_sum2Map_sum1_14, addersMap_sum1Map_sum2Map_sum1_13, 
         addersMap_sum1Map_sum2Map_sum1_12, addersMap_sum1Map_sum2Map_sum1_11, 
         addersMap_sum1Map_sum2Map_sum1_10, addersMap_sum1Map_sum2Map_sum1_9, 
         addersMap_sum1Map_sum2Map_sum1_8, addersMap_sum1Map_sum2Map_sum1_7, 
         addersMap_sum1Map_sum2Map_sum1_6, addersMap_sum1Map_sum2Map_sum1_5, 
         addersMap_sum1Map_sum2Map_sum1_4, addersMap_sum1Map_sum2Map_sum1_3, 
         addersMap_sum1Map_sum2Map_sum1_2, addersMap_sum1Map_sum2Map_sum1_1, 
         addersMap_sum1Map_sum2Map_sum1_0, addersMap_sum1Map_sum2Map_sum2_15, 
         addersMap_sum1Map_sum2Map_sum2_14, addersMap_sum1Map_sum2Map_sum2_13, 
         addersMap_sum1Map_sum2Map_sum2_12, addersMap_sum1Map_sum2Map_sum2_11, 
         addersMap_sum1Map_sum2Map_sum2_10, addersMap_sum1Map_sum2Map_sum2_9, 
         addersMap_sum1Map_sum2Map_sum2_8, addersMap_sum1Map_sum2Map_sum2_7, 
         addersMap_sum1Map_sum2Map_sum2_6, addersMap_sum1Map_sum2Map_sum2_5, 
         addersMap_sum1Map_sum2Map_sum2_4, addersMap_sum1Map_sum2Map_sum2_3, 
         addersMap_sum1Map_sum2Map_sum2_2, addersMap_sum1Map_sum2Map_sum2_1, 
         addersMap_sum1Map_sum2Map_sum2_0, addersMap_sum2Map_sum1_15__dup_0, 
         addersMap_sum2Map_sum1_14__dup_0, addersMap_sum2Map_sum1_13__dup_0, 
         addersMap_sum2Map_sum1_12__dup_0, addersMap_sum2Map_sum1_11__dup_0, 
         addersMap_sum2Map_sum1_10__dup_0, addersMap_sum2Map_sum1_9__dup_0, 
         addersMap_sum2Map_sum1_8__dup_0, addersMap_sum2Map_sum1_7__dup_0, 
         addersMap_sum2Map_sum1_6__dup_0, addersMap_sum2Map_sum1_5__dup_0, 
         addersMap_sum2Map_sum1_4__dup_0, addersMap_sum2Map_sum1_3__dup_0, 
         addersMap_sum2Map_sum1_2__dup_0, addersMap_sum2Map_sum1_1__dup_0, 
         addersMap_sum2Map_sum1_0__dup_0, addersMap_sum2Map_sum2_15__dup_0, 
         addersMap_sum2Map_sum2_14__dup_0, addersMap_sum2Map_sum2_13__dup_0, 
         addersMap_sum2Map_sum2_12__dup_0, addersMap_sum2Map_sum2_11__dup_0, 
         addersMap_sum2Map_sum2_10__dup_0, addersMap_sum2Map_sum2_9__dup_0, 
         addersMap_sum2Map_sum2_8__dup_0, addersMap_sum2Map_sum2_7__dup_0, 
         addersMap_sum2Map_sum2_6__dup_0, addersMap_sum2Map_sum2_5__dup_0, 
         addersMap_sum2Map_sum2_4__dup_0, addersMap_sum2Map_sum2_3__dup_0, 
         addersMap_sum2Map_sum2_2__dup_0, addersMap_sum2Map_sum2_1__dup_0, 
         addersMap_sum2Map_sum2_0__dup_0, addersMap_sum2Map_sum1Map_sum1_15, 
         addersMap_sum2Map_sum1Map_sum1_14, addersMap_sum2Map_sum1Map_sum1_13, 
         addersMap_sum2Map_sum1Map_sum1_12, addersMap_sum2Map_sum1Map_sum1_11, 
         addersMap_sum2Map_sum1Map_sum1_10, addersMap_sum2Map_sum1Map_sum1_9, 
         addersMap_sum2Map_sum1Map_sum1_8, addersMap_sum2Map_sum1Map_sum1_7, 
         addersMap_sum2Map_sum1Map_sum1_6, addersMap_sum2Map_sum1Map_sum1_5, 
         addersMap_sum2Map_sum1Map_sum1_4, addersMap_sum2Map_sum1Map_sum1_3, 
         addersMap_sum2Map_sum1Map_sum1_2, addersMap_sum2Map_sum1Map_sum1_1, 
         addersMap_sum2Map_sum1Map_sum1_0, addersMap_sum2Map_sum1Map_sum2_15, 
         addersMap_sum2Map_sum1Map_sum2_14, addersMap_sum2Map_sum1Map_sum2_13, 
         addersMap_sum2Map_sum1Map_sum2_12, addersMap_sum2Map_sum1Map_sum2_11, 
         addersMap_sum2Map_sum1Map_sum2_10, addersMap_sum2Map_sum1Map_sum2_9, 
         addersMap_sum2Map_sum1Map_sum2_8, addersMap_sum2Map_sum1Map_sum2_7, 
         addersMap_sum2Map_sum1Map_sum2_6, addersMap_sum2Map_sum1Map_sum2_5, 
         addersMap_sum2Map_sum1Map_sum2_4, addersMap_sum2Map_sum1Map_sum2_3, 
         addersMap_sum2Map_sum1Map_sum2_2, addersMap_sum2Map_sum1Map_sum2_1, 
         addersMap_sum2Map_sum1Map_sum2_0, addersMap_sum2Map_sum2Map_sum1_15, 
         addersMap_sum2Map_sum2Map_sum1_14, addersMap_sum2Map_sum2Map_sum1_13, 
         addersMap_sum2Map_sum2Map_sum1_12, addersMap_sum2Map_sum2Map_sum1_11, 
         addersMap_sum2Map_sum2Map_sum1_10, addersMap_sum2Map_sum2Map_sum1_9, 
         addersMap_sum2Map_sum2Map_sum1_8, addersMap_sum2Map_sum2Map_sum1_7, 
         addersMap_sum2Map_sum2Map_sum1_6, addersMap_sum2Map_sum2Map_sum1_5, 
         addersMap_sum2Map_sum2Map_sum1_4, addersMap_sum2Map_sum2Map_sum1_3, 
         addersMap_sum2Map_sum2Map_sum1_2, addersMap_sum2Map_sum2Map_sum1_1, 
         addersMap_sum2Map_sum2Map_sum1_0, addersMap_sum2Map_sum2Map_sum2_15, 
         addersMap_sum2Map_sum2Map_sum2_14, addersMap_sum2Map_sum2Map_sum2_13, 
         addersMap_sum2Map_sum2Map_sum2_12, addersMap_sum2Map_sum2Map_sum2_11, 
         addersMap_sum2Map_sum2Map_sum2_10, addersMap_sum2Map_sum2Map_sum2_9, 
         addersMap_sum2Map_sum2Map_sum2_8, addersMap_sum2Map_sum2Map_sum2_7, 
         addersMap_sum2Map_sum2Map_sum2_6, addersMap_sum2Map_sum2Map_sum2_5, 
         addersMap_sum2Map_sum2Map_sum2_4, addersMap_sum2Map_sum2Map_sum2_3, 
         addersMap_sum2Map_sum2Map_sum2_2, addersMap_sum2Map_sum2Map_sum2_1, 
         addersMap_sum2Map_sum2Map_sum2_0, addersMap_sum3Map_sum1_15, 
         addersMap_sum3Map_sum1_14, addersMap_sum3Map_sum1_13, 
         addersMap_sum3Map_sum1_12, addersMap_sum3Map_sum1_11, 
         addersMap_sum3Map_sum1_10, addersMap_sum3Map_sum1_9, 
         addersMap_sum3Map_sum1_8, addersMap_sum3Map_sum1_7, 
         addersMap_sum3Map_sum1_6, addersMap_sum3Map_sum1_5, 
         addersMap_sum3Map_sum1_4, addersMap_sum3Map_sum1_3, 
         addersMap_sum3Map_sum1_2, addersMap_sum3Map_sum1_1, 
         addersMap_sum3Map_sum1_0, addersMap_sum3Map_sum2_15, 
         addersMap_sum3Map_sum2_14, addersMap_sum3Map_sum2_13, 
         addersMap_sum3Map_sum2_12, addersMap_sum3Map_sum2_11, 
         addersMap_sum3Map_sum2_10, addersMap_sum3Map_sum2_9, 
         addersMap_sum3Map_sum2_8, addersMap_sum3Map_sum2_7, 
         addersMap_sum3Map_sum2_6, addersMap_sum3Map_sum2_5, 
         addersMap_sum3Map_sum2_4, addersMap_sum3Map_sum2_3, 
         addersMap_sum3Map_sum2_2, addersMap_sum3Map_sum2_1, 
         addersMap_sum3Map_sum2_0, addersMap_sum3Map_sum1Map_sum1_15, 
         addersMap_sum3Map_sum1Map_sum1_14, addersMap_sum3Map_sum1Map_sum1_13, 
         addersMap_sum3Map_sum1Map_sum1_12, addersMap_sum3Map_sum1Map_sum1_11, 
         addersMap_sum3Map_sum1Map_sum1_10, addersMap_sum3Map_sum1Map_sum1_9, 
         addersMap_sum3Map_sum1Map_sum1_8, addersMap_sum3Map_sum1Map_sum1_7, 
         addersMap_sum3Map_sum1Map_sum1_6, addersMap_sum3Map_sum1Map_sum1_5, 
         addersMap_sum3Map_sum1Map_sum1_4, addersMap_sum3Map_sum1Map_sum1_3, 
         addersMap_sum3Map_sum1Map_sum1_2, addersMap_sum3Map_sum1Map_sum1_1, 
         addersMap_sum3Map_sum1Map_sum1_0, addersMap_sum3Map_sum1Map_sum2_15, 
         addersMap_sum3Map_sum1Map_sum2_14, addersMap_sum3Map_sum1Map_sum2_13, 
         addersMap_sum3Map_sum1Map_sum2_12, addersMap_sum3Map_sum1Map_sum2_11, 
         addersMap_sum3Map_sum1Map_sum2_10, addersMap_sum3Map_sum1Map_sum2_9, 
         addersMap_sum3Map_sum1Map_sum2_8, addersMap_sum3Map_sum1Map_sum2_7, 
         addersMap_sum3Map_sum1Map_sum2_6, addersMap_sum3Map_sum1Map_sum2_5, 
         addersMap_sum3Map_sum1Map_sum2_4, addersMap_sum3Map_sum1Map_sum2_3, 
         addersMap_sum3Map_sum1Map_sum2_2, addersMap_sum3Map_sum1Map_sum2_1, 
         addersMap_sum3Map_sum1Map_sum2_0, addersMap_sum3Map_sum2Map_sum1_15, 
         addersMap_sum3Map_sum2Map_sum1_14, addersMap_sum3Map_sum2Map_sum1_13, 
         addersMap_sum3Map_sum2Map_sum1_12, addersMap_sum3Map_sum2Map_sum1_11, 
         addersMap_sum3Map_sum2Map_sum1_10, addersMap_sum3Map_sum2Map_sum1_9, 
         addersMap_sum3Map_sum2Map_sum1_8, addersMap_sum3Map_sum2Map_sum1_7, 
         addersMap_sum3Map_sum2Map_sum1_6, addersMap_sum3Map_sum2Map_sum1_5, 
         addersMap_sum3Map_sum2Map_sum1_4, addersMap_sum3Map_sum2Map_sum1_3, 
         addersMap_sum3Map_sum2Map_sum1_2, addersMap_sum3Map_sum2Map_sum1_1, 
         addersMap_sum3Map_sum2Map_sum1_0, addersMap_sum3Map_sum2Map_sum2_15, 
         addersMap_sum3Map_sum2Map_sum2_14, addersMap_sum3Map_sum2Map_sum2_13, 
         addersMap_sum3Map_sum2Map_sum2_12, addersMap_sum3Map_sum2Map_sum2_11, 
         addersMap_sum3Map_sum2Map_sum2_10, addersMap_sum3Map_sum2Map_sum2_9, 
         addersMap_sum3Map_sum2Map_sum2_8, addersMap_sum3Map_sum2Map_sum2_7, 
         addersMap_sum3Map_sum2Map_sum2_6, addersMap_sum3Map_sum2Map_sum2_5, 
         addersMap_sum3Map_sum2Map_sum2_4, addersMap_sum3Map_sum2Map_sum2_3, 
         addersMap_sum3Map_sum2Map_sum2_2, addersMap_sum3Map_sum2Map_sum2_1, 
         addersMap_sum3Map_sum2Map_sum2_0, outShifter_15, nx4, nx3412, nx3470, 
         nx2917, nx2923, nx2925, nx2929, nx2931, nx2935, nx2937, nx2941, nx2947, 
         nx2951, nx2959, nx2963, nx2971, nx2973, nx2979, nx2981, nx2985, nx2987, 
         nx2991, nx2993, nx2997, nx2999, nx3003, nx3005, nx3009, nx3011, nx3015, 
         nx3017, nx3021, nx3023, nx3027, nx3029, nx3033, nx3035, nx3039, nx3041, 
         nx3045, nx3047, nx3051, nx3053, nx3057, nx3059, nx3063, nx3065, nx3069, 
         nx3071, nx3075, nx3077, nx3081, nx3083, nx3087, nx3089, nx3093, nx3095, 
         nx3099, nx3101, nx3105, nx3107, nx3111, nx3113, nx3117, nx3119, nx3123, 
         nx3125, nx3129, nx3131, nx3135, nx3137, nx3141, nx3143, nx3147, nx3149, 
         nx3153, nx3155, nx3159, nx3161, nx3165, nx3167, nx3171, nx3173, nx3177, 
         nx3179, nx3183, nx3185, nx3189, nx3191, nx3195, nx3197, nx3201, nx3203, 
         nx3207, nx3209, nx3213, nx3215, nx3219, nx3221, nx3225, nx3227, nx3231, 
         nx3233, nx3237, nx3239, nx3243, nx3245, nx3249, nx3251, nx3255, nx3257, 
         nx3261, nx3263, nx3267, nx3269, nx3273, nx3275, nx3279, nx3281, nx3285, 
         nx3287, nx3291, nx3293, nx3297, nx3299, nx3303, nx3305, nx3309, nx3311, 
         nx3315, nx3317, nx3321, nx3323, nx3327, nx3329, nx3333, nx3335, nx3339, 
         nx3341, nx3345, nx3347, nx3351, nx3353, nx3357, nx3359, nx3363, nx3365, 
         nx3369, nx3371, nx3375, nx3377, nx3381, nx3383, nx3387, nx3389, nx3393, 
         nx3395, nx3399, nx3401, nx3405, nx3407, nx3411, nx3413, nx3417, nx3419, 
         nx3423, nx3425, nx3429, nx3431, nx3435, nx3437, nx3441, nx3443, nx3447, 
         nx3449, nx3453, nx3455, nx3459, nx3461, nx3465, nx3467, nx3471, nx3473, 
         nx3477, nx3479, nx3483, nx3485, nx3488, nx3490, nx3493, nx3495, nx3498, 
         nx3500, nx3503, nx3505, nx3508, nx3510, nx3513, nx3515, nx3518, nx3520, 
         nx3523, nx3525, nx3528, nx3530, nx3533, nx3535, nx3538, nx3540, nx3543, 
         nx3545, nx3548, nx3550, nx3553, nx3555, nx3558, nx3560, nx3563, nx3565, 
         nx3568, nx3570, nx3573, nx3575, nx3578, nx3580, nx3583, nx3585, nx3588, 
         nx3590, nx3593, nx3595, nx3598, nx3600, nx3603, nx3605, nx3608, nx3610, 
         nx3613, nx3615, nx3618, nx3620, nx3623, nx3625, nx3628, nx3630, nx3633, 
         nx3635, nx3638, nx3640, nx3643, nx3645, nx3648, nx3650, nx3653, nx3655, 
         nx3658, nx3660, nx3663, nx3665, nx3668, nx3670, nx3673, nx3675, nx3678, 
         nx3680, nx3683, nx3685, nx3688, nx3690, nx3693, nx3695, nx3698, nx3700, 
         nx3703, nx3705, nx3708, nx3710, nx3713, nx3715, nx3718, nx3720, nx3723, 
         nx3725, nx3728, nx3730, nx3733, nx3735, nx3738, nx3740, nx3743, nx3745, 
         nx3748, nx3750, nx3753, nx3755, nx3758, nx3760, nx3763, nx3765, nx3768, 
         nx3770, nx3773, nx3775, nx3778, nx3780, nx3783, nx3785, nx3788, nx3790, 
         nx3793, nx3795, nx3798, nx3800, nx3803, nx3805, nx3808, nx3810, nx3813, 
         nx3815, nx3818, nx3820, nx3823, nx3825, nx3828, nx3830, nx3833, nx3835, 
         nx3838, nx3840, nx3843, nx3845, nx3848, nx3850, nx3853, nx3855, nx3858, 
         nx3860, nx3863, nx3865, nx3868, nx3870, nx3873, nx3875, nx3878, nx3880, 
         nx3883, nx3885, nx3888, nx3890, nx3893, nx3895, nx3898, nx3900, nx3903, 
         nx3905, nx3908, nx3910, nx3913, nx3915, nx3918, nx3920, nx3923, nx3925, 
         nx3928, nx3930, nx3933, nx3935, nx3938, nx3940, nx3943, nx3945, nx3948, 
         nx3950, nx3953, nx3955, nx3958, nx3960, nx3963, nx3965, nx3968, nx3970, 
         nx3973, nx3975, nx3978, nx3980, nx3983, nx3985, nx3988, nx3990, nx3993, 
         nx3995, nx3998, nx4000, nx4003, nx4005, nx4008, nx4010, nx4013, nx4015, 
         nx4018, nx4020, nx4023, nx4025, nx4028, nx4030, nx4033, nx4035, nx4038, 
         nx4040, nx4043, nx4045, nx4048, nx4050, nx4053, nx4055, nx4058, nx4060, 
         nx4063, nx4065, nx4068, nx4070, nx4073, nx4075, nx4078, nx4080, nx4083, 
         nx4085, nx4088, nx4090, nx4093, nx4095, nx4098, nx4100, nx4103, nx4105, 
         nx4108, nx4110, nx4113, nx4115, nx4118, nx4120, nx4123, nx4125, nx4128, 
         nx4130, nx4133, nx4135, nx4138, nx4140, nx4143, nx4145, nx4148, nx4150, 
         nx4153, nx4155, nx4158, nx4160, nx4163, nx4165, nx4168, nx4170, nx4173, 
         nx4175, nx4178, nx4180, nx4183, nx4185, nx4188, nx4190, nx4193, nx4195, 
         nx4198, nx4200, nx4203, nx4205, nx4208, nx4210, nx4213, nx4215, nx4218, 
         nx4220, nx4223, nx4225, nx4228, nx4230, nx4233, nx4235, nx4238, nx4240, 
         nx4243, nx4245, nx4248, nx4250, nx4253, nx4255, nx4258, nx4260, nx4263, 
         nx4265, nx4268, nx4270, nx4273, nx4275, nx4278, nx4280, nx4283, nx4285, 
         nx4288, nx4290, nx4293, nx4295, nx4298, nx4300, nx4303, nx4305, nx4308, 
         nx4310, nx4313, nx4315, nx4318, nx4320, nx4323, nx4325, nx4328, nx4330, 
         nx4333, nx4335, nx4338, nx4340, nx4343, nx4345, nx4348, nx4350, nx4353, 
         nx4355, nx4358, nx4360, nx4363, nx4365, nx4368, nx4370, nx4373, nx4375, 
         nx4378, nx4380, nx4383, nx4385, nx4388, nx4390, nx4393, nx4395, nx4398, 
         nx4400, nx4403, nx4405, nx4408, nx4410, nx4413, nx4415, nx4418, nx4420, 
         nx4423, nx4425, nx4428, nx4430, nx4433, nx4435, nx4438, nx4440, nx4443, 
         nx4445, nx4448, nx4450, nx4453, nx4455, nx4458, nx4460, nx4463, nx4465, 
         nx4468, nx4470, nx4473, nx4475, nx4478, nx4480, nx4483, nx4485, nx4488, 
         nx4490, nx4493, nx4495, nx4498, nx4500, nx4503, nx4505, nx4508, nx4510, 
         nx4513, nx4515, nx4518, nx4520, nx4523, nx4525, nx4528, nx4530, nx4533, 
         nx4535, nx4538, nx4540, nx4543, nx4545, nx4548, nx4550, nx4553, nx4555, 
         nx4558, nx4560, nx4563, nx4565, nx4568, nx4570, nx4573, nx4575, nx4578, 
         nx4580, nx4583, nx4585, nx4588, nx4590, nx4593, nx4595, nx4598, nx4600, 
         nx4603, nx4605, nx4608, nx4610, nx4613, nx4615, nx4618, nx4620, nx4623, 
         nx4625, nx4628, nx4630, nx4633, nx4635, nx4638, nx4640, nx4643, nx4645, 
         nx4648, nx4650, nx4653, nx4655, nx4658, nx4660, nx4663, nx4665, nx4668, 
         nx4670, nx4673, nx4675, nx4678, nx4680, nx4683, nx4685, nx4688, nx4690, 
         nx4693, nx4695, nx4698, nx4700, nx4703, nx4705, nx4708, nx4710, nx4713, 
         nx4715, nx4718, nx4720, nx4723, nx4725, nx4728, nx4730, nx4733, nx4735, 
         nx4738, nx4740, nx4743, nx4745, nx4748, nx4750, nx4753, nx4755, nx4758, 
         nx4760, nx4763, nx4765, nx4768, nx4770, nx4773, nx4775, nx4778, nx4780, 
         nx4783, nx4785, nx4788, nx4790, nx4793, nx4795, nx4798, nx4800, nx4803, 
         nx4805, nx4808, nx4810, nx4813, nx4815, nx4818, nx4820, nx4823, nx4825, 
         nx4828, nx4830, nx4833, nx4835, nx4838, nx4840, nx4843, nx4845, nx4848, 
         nx4850, nx4853, nx4855, nx4858, nx4860, nx4863, nx4865, nx4868, nx4870, 
         nx4873, nx4875, nx4878, nx4880, nx4883, nx4885, nx4888, nx4890, nx4893, 
         nx4895, nx4898, nx4900, nx4903, nx4905, nx4908, nx4910, nx4913, nx4915, 
         nx4918, nx4920, nx4923, nx4925, nx4928, nx4930, nx4933, nx4935, nx4938, 
         nx4940, nx4943, nx4945, nx4948, nx4950, nx4953, nx4955, nx4958, nx4960, 
         nx4963, nx4965, nx4968, nx4970, nx4973, nx4975, nx4978, nx4980, nx4983, 
         nx4985, nx4988, nx4990, nx4993, nx4995, nx4998, nx5000, nx5003, nx5005, 
         nx5008, nx5010, nx5013, nx5015, nx5018, nx5020, nx5023, nx5025, nx5028, 
         nx5030, nx5033, nx5035, nx5038, nx5040, nx5043, nx5045, nx5048, nx5050, 
         nx5053, nx5055, nx5058, nx5060, nx5063, nx5067, nx5070, nx5072, nx5074, 
         nx5076, nx5079, nx5081, nx5083, nx5085, nx5088, nx5090, nx5092, nx5094, 
         nx5097, nx5099, nx5101, nx5103, nx5106, nx5108, nx5110, nx5112, nx5115, 
         nx5117, nx5119, nx5121, nx5124, nx5126, nx5128, nx5130, nx5133, nx5135, 
         nx5137, nx5139, nx5142, nx5144, nx5146, nx5148, nx5151, nx5153, nx5155, 
         nx5157, nx5160, nx5162, nx5164, nx5167, nx5169, nx5171, nx5174, nx5176, 
         nx5179, nx5181, nx5184, nx5186, nx5189, nx5196, nx5198, nx5200, nx5202, 
         nx5204, nx5206, nx5208, nx5210, nx5212, nx5214, nx5216, nx5218, nx5220, 
         nx5222, nx5224, nx5226, nx5228, nx5230, nx5232, nx5234, nx5236, nx5238, 
         nx5240, nx5242, nx5244, nx5246, nx5248, nx5250, nx5252, nx5254, nx5256, 
         nx5258, nx5260, nx5262, nx5264, nx5266, nx5268, nx5270, nx5272, nx5274, 
         nx5276, nx5278, nx5280, nx5282, nx5284, nx5286, nx5288, nx5290, nx5292, 
         nx5294, nx5296, nx5298, nx5300, nx5302, nx5304, nx5306, nx5308, nx5310, 
         nx5312, nx5314, nx5316, nx5318, nx5320, nx5322, nx5328, nx5330, nx5332, 
         nx5334, nx5336, nx5338, nx5340, nx5342, nx5344, nx5346;
    wire [184:0] \$dummy ;




    CNNMuls_25 mulsMap (.filter_24__7 (filter_0__7), .filter_24__6 (filter_0__6)
               , .filter_24__5 (filter_0__5), .filter_24__4 (filter_0__4), .filter_24__3 (
               filter_0__3), .filter_24__2 (filter_0__2), .filter_24__1 (
               filter_0__1), .filter_24__0 (filter_0__0), .filter_23__7 (
               filter_1__7), .filter_23__6 (filter_1__6), .filter_23__5 (
               filter_1__5), .filter_23__4 (filter_1__4), .filter_23__3 (
               filter_1__3), .filter_23__2 (filter_1__2), .filter_23__1 (
               filter_1__1), .filter_23__0 (filter_1__0), .filter_22__7 (
               filter_2__7), .filter_22__6 (filter_2__6), .filter_22__5 (
               filter_2__5), .filter_22__4 (filter_2__4), .filter_22__3 (
               filter_2__3), .filter_22__2 (filter_2__2), .filter_22__1 (
               filter_2__1), .filter_22__0 (filter_2__0), .filter_21__7 (
               filter_3__7), .filter_21__6 (filter_3__6), .filter_21__5 (
               filter_3__5), .filter_21__4 (filter_3__4), .filter_21__3 (
               filter_3__3), .filter_21__2 (filter_3__2), .filter_21__1 (
               filter_3__1), .filter_21__0 (filter_3__0), .filter_20__7 (
               filter_4__7), .filter_20__6 (filter_4__6), .filter_20__5 (
               filter_4__5), .filter_20__4 (filter_4__4), .filter_20__3 (
               filter_4__3), .filter_20__2 (filter_4__2), .filter_20__1 (
               filter_4__1), .filter_20__0 (filter_4__0), .filter_19__7 (
               filter_5__7), .filter_19__6 (filter_5__6), .filter_19__5 (
               filter_5__5), .filter_19__4 (filter_5__4), .filter_19__3 (
               filter_5__3), .filter_19__2 (filter_5__2), .filter_19__1 (
               filter_5__1), .filter_19__0 (filter_5__0), .filter_18__7 (
               filter_6__7), .filter_18__6 (filter_6__6), .filter_18__5 (
               filter_6__5), .filter_18__4 (filter_6__4), .filter_18__3 (
               filter_6__3), .filter_18__2 (filter_6__2), .filter_18__1 (
               filter_6__1), .filter_18__0 (filter_6__0), .filter_17__7 (
               filter_7__7), .filter_17__6 (filter_7__6), .filter_17__5 (
               filter_7__5), .filter_17__4 (filter_7__4), .filter_17__3 (
               filter_7__3), .filter_17__2 (filter_7__2), .filter_17__1 (
               filter_7__1), .filter_17__0 (filter_7__0), .filter_16__7 (
               filter_8__7), .filter_16__6 (filter_8__6), .filter_16__5 (
               filter_8__5), .filter_16__4 (filter_8__4), .filter_16__3 (
               filter_8__3), .filter_16__2 (filter_8__2), .filter_16__1 (
               filter_8__1), .filter_16__0 (filter_8__0), .filter_15__7 (
               filter_9__7), .filter_15__6 (filter_9__6), .filter_15__5 (
               filter_9__5), .filter_15__4 (filter_9__4), .filter_15__3 (
               filter_9__3), .filter_15__2 (filter_9__2), .filter_15__1 (
               filter_9__1), .filter_15__0 (filter_9__0), .filter_14__7 (
               filter_10__7), .filter_14__6 (filter_10__6), .filter_14__5 (
               filter_10__5), .filter_14__4 (filter_10__4), .filter_14__3 (
               filter_10__3), .filter_14__2 (filter_10__2), .filter_14__1 (
               filter_10__1), .filter_14__0 (filter_10__0), .filter_13__7 (
               filter_11__7), .filter_13__6 (filter_11__6), .filter_13__5 (
               filter_11__5), .filter_13__4 (filter_11__4), .filter_13__3 (
               filter_11__3), .filter_13__2 (filter_11__2), .filter_13__1 (
               filter_11__1), .filter_13__0 (filter_11__0), .filter_12__7 (
               filter_12__7), .filter_12__6 (filter_12__6), .filter_12__5 (
               filter_12__5), .filter_12__4 (filter_12__4), .filter_12__3 (
               filter_12__3), .filter_12__2 (filter_12__2), .filter_12__1 (
               filter_12__1), .filter_12__0 (filter_12__0), .filter_11__7 (
               filter_13__7), .filter_11__6 (filter_13__6), .filter_11__5 (
               filter_13__5), .filter_11__4 (filter_13__4), .filter_11__3 (
               filter_13__3), .filter_11__2 (filter_13__2), .filter_11__1 (
               filter_13__1), .filter_11__0 (filter_13__0), .filter_10__7 (
               filter_14__7), .filter_10__6 (filter_14__6), .filter_10__5 (
               filter_14__5), .filter_10__4 (filter_14__4), .filter_10__3 (
               filter_14__3), .filter_10__2 (filter_14__2), .filter_10__1 (
               filter_14__1), .filter_10__0 (filter_14__0), .filter_9__7 (
               filter_15__7), .filter_9__6 (filter_15__6), .filter_9__5 (
               filter_15__5), .filter_9__4 (filter_15__4), .filter_9__3 (
               filter_15__3), .filter_9__2 (filter_15__2), .filter_9__1 (
               filter_15__1), .filter_9__0 (filter_15__0), .filter_8__7 (
               filter_16__7), .filter_8__6 (filter_16__6), .filter_8__5 (
               filter_16__5), .filter_8__4 (filter_16__4), .filter_8__3 (
               filter_16__3), .filter_8__2 (filter_16__2), .filter_8__1 (
               filter_16__1), .filter_8__0 (filter_16__0), .filter_7__7 (
               filter_17__7), .filter_7__6 (filter_17__6), .filter_7__5 (
               filter_17__5), .filter_7__4 (filter_17__4), .filter_7__3 (
               filter_17__3), .filter_7__2 (filter_17__2), .filter_7__1 (
               filter_17__1), .filter_7__0 (filter_17__0), .filter_6__7 (
               filter_18__7), .filter_6__6 (filter_18__6), .filter_6__5 (
               filter_18__5), .filter_6__4 (filter_18__4), .filter_6__3 (
               filter_18__3), .filter_6__2 (filter_18__2), .filter_6__1 (
               filter_18__1), .filter_6__0 (filter_18__0), .filter_5__7 (
               filter_19__7), .filter_5__6 (filter_19__6), .filter_5__5 (
               filter_19__5), .filter_5__4 (filter_19__4), .filter_5__3 (
               filter_19__3), .filter_5__2 (filter_19__2), .filter_5__1 (
               filter_19__1), .filter_5__0 (filter_19__0), .filter_4__7 (
               filter_20__7), .filter_4__6 (filter_20__6), .filter_4__5 (
               filter_20__5), .filter_4__4 (filter_20__4), .filter_4__3 (
               filter_20__3), .filter_4__2 (filter_20__2), .filter_4__1 (
               filter_20__1), .filter_4__0 (filter_20__0), .filter_3__7 (
               filter_21__7), .filter_3__6 (filter_21__6), .filter_3__5 (
               filter_21__5), .filter_3__4 (filter_21__4), .filter_3__3 (
               filter_21__3), .filter_3__2 (filter_21__2), .filter_3__1 (
               filter_21__1), .filter_3__0 (filter_21__0), .filter_2__7 (
               filter_22__7), .filter_2__6 (filter_22__6), .filter_2__5 (
               filter_22__5), .filter_2__4 (filter_22__4), .filter_2__3 (
               filter_22__3), .filter_2__2 (filter_22__2), .filter_2__1 (
               filter_22__1), .filter_2__0 (filter_22__0), .filter_1__7 (
               filter_23__7), .filter_1__6 (filter_23__6), .filter_1__5 (
               filter_23__5), .filter_1__4 (filter_23__4), .filter_1__3 (
               filter_23__3), .filter_1__2 (filter_23__2), .filter_1__1 (
               filter_23__1), .filter_1__0 (filter_23__0), .filter_0__7 (
               filter_24__7), .filter_0__6 (filter_24__6), .filter_0__5 (
               filter_24__5), .filter_0__4 (filter_24__4), .filter_0__3 (
               filter_24__3), .filter_0__2 (filter_24__2), .filter_0__1 (
               filter_24__1), .filter_0__0 (filter_24__0), .window_24__15 (
               currentPage_0__15), .window_24__14 (currentPage_0__14), .window_24__13 (
               currentPage_0__13), .window_24__12 (currentPage_0__12), .window_24__11 (
               currentPage_0__11), .window_24__10 (currentPage_0__10), .window_24__9 (
               currentPage_0__9), .window_24__8 (currentPage_0__8), .window_24__7 (
               currentPage_0__7), .window_24__6 (currentPage_0__6), .window_24__5 (
               currentPage_0__5), .window_24__4 (currentPage_0__4), .window_24__3 (
               currentPage_0__3), .window_24__2 (currentPage_0__2), .window_24__1 (
               currentPage_0__1), .window_24__0 (currentPage_0__0), .window_23__15 (
               currentPage_1__15), .window_23__14 (currentPage_1__14), .window_23__13 (
               currentPage_1__13), .window_23__12 (currentPage_1__12), .window_23__11 (
               currentPage_1__11), .window_23__10 (currentPage_1__10), .window_23__9 (
               currentPage_1__9), .window_23__8 (currentPage_1__8), .window_23__7 (
               currentPage_1__7), .window_23__6 (currentPage_1__6), .window_23__5 (
               currentPage_1__5), .window_23__4 (currentPage_1__4), .window_23__3 (
               currentPage_1__3), .window_23__2 (currentPage_1__2), .window_23__1 (
               currentPage_1__1), .window_23__0 (currentPage_1__0), .window_22__15 (
               currentPage_2__15), .window_22__14 (currentPage_2__14), .window_22__13 (
               currentPage_2__13), .window_22__12 (currentPage_2__12), .window_22__11 (
               currentPage_2__11), .window_22__10 (currentPage_2__10), .window_22__9 (
               currentPage_2__9), .window_22__8 (currentPage_2__8), .window_22__7 (
               currentPage_2__7), .window_22__6 (currentPage_2__6), .window_22__5 (
               currentPage_2__5), .window_22__4 (currentPage_2__4), .window_22__3 (
               currentPage_2__3), .window_22__2 (currentPage_2__2), .window_22__1 (
               currentPage_2__1), .window_22__0 (currentPage_2__0), .window_21__15 (
               currentPage_3__15), .window_21__14 (currentPage_3__14), .window_21__13 (
               currentPage_3__13), .window_21__12 (currentPage_3__12), .window_21__11 (
               currentPage_3__11), .window_21__10 (currentPage_3__10), .window_21__9 (
               currentPage_3__9), .window_21__8 (currentPage_3__8), .window_21__7 (
               currentPage_3__7), .window_21__6 (currentPage_3__6), .window_21__5 (
               currentPage_3__5), .window_21__4 (currentPage_3__4), .window_21__3 (
               currentPage_3__3), .window_21__2 (currentPage_3__2), .window_21__1 (
               currentPage_3__1), .window_21__0 (currentPage_3__0), .window_20__15 (
               currentPage_4__15), .window_20__14 (currentPage_4__14), .window_20__13 (
               currentPage_4__13), .window_20__12 (currentPage_4__12), .window_20__11 (
               currentPage_4__11), .window_20__10 (currentPage_4__10), .window_20__9 (
               currentPage_4__9), .window_20__8 (currentPage_4__8), .window_20__7 (
               currentPage_4__7), .window_20__6 (currentPage_4__6), .window_20__5 (
               currentPage_4__5), .window_20__4 (currentPage_4__4), .window_20__3 (
               currentPage_4__3), .window_20__2 (currentPage_4__2), .window_20__1 (
               currentPage_4__1), .window_20__0 (currentPage_4__0), .window_19__15 (
               currentPage_5__15), .window_19__14 (currentPage_5__14), .window_19__13 (
               currentPage_5__13), .window_19__12 (currentPage_5__12), .window_19__11 (
               currentPage_5__11), .window_19__10 (currentPage_5__10), .window_19__9 (
               currentPage_5__9), .window_19__8 (currentPage_5__8), .window_19__7 (
               currentPage_5__7), .window_19__6 (currentPage_5__6), .window_19__5 (
               currentPage_5__5), .window_19__4 (currentPage_5__4), .window_19__3 (
               currentPage_5__3), .window_19__2 (currentPage_5__2), .window_19__1 (
               currentPage_5__1), .window_19__0 (currentPage_5__0), .window_18__15 (
               currentPage_6__15), .window_18__14 (currentPage_6__14), .window_18__13 (
               currentPage_6__13), .window_18__12 (currentPage_6__12), .window_18__11 (
               currentPage_6__11), .window_18__10 (currentPage_6__10), .window_18__9 (
               currentPage_6__9), .window_18__8 (currentPage_6__8), .window_18__7 (
               currentPage_6__7), .window_18__6 (currentPage_6__6), .window_18__5 (
               currentPage_6__5), .window_18__4 (currentPage_6__4), .window_18__3 (
               currentPage_6__3), .window_18__2 (currentPage_6__2), .window_18__1 (
               currentPage_6__1), .window_18__0 (currentPage_6__0), .window_17__15 (
               currentPage_7__15), .window_17__14 (currentPage_7__14), .window_17__13 (
               currentPage_7__13), .window_17__12 (currentPage_7__12), .window_17__11 (
               currentPage_7__11), .window_17__10 (currentPage_7__10), .window_17__9 (
               currentPage_7__9), .window_17__8 (currentPage_7__8), .window_17__7 (
               currentPage_7__7), .window_17__6 (currentPage_7__6), .window_17__5 (
               currentPage_7__5), .window_17__4 (currentPage_7__4), .window_17__3 (
               currentPage_7__3), .window_17__2 (currentPage_7__2), .window_17__1 (
               currentPage_7__1), .window_17__0 (currentPage_7__0), .window_16__15 (
               currentPage_8__15), .window_16__14 (currentPage_8__14), .window_16__13 (
               currentPage_8__13), .window_16__12 (currentPage_8__12), .window_16__11 (
               currentPage_8__11), .window_16__10 (currentPage_8__10), .window_16__9 (
               currentPage_8__9), .window_16__8 (currentPage_8__8), .window_16__7 (
               currentPage_8__7), .window_16__6 (currentPage_8__6), .window_16__5 (
               currentPage_8__5), .window_16__4 (currentPage_8__4), .window_16__3 (
               currentPage_8__3), .window_16__2 (currentPage_8__2), .window_16__1 (
               currentPage_8__1), .window_16__0 (currentPage_8__0), .window_15__15 (
               currentPage_9__15), .window_15__14 (currentPage_9__14), .window_15__13 (
               currentPage_9__13), .window_15__12 (currentPage_9__12), .window_15__11 (
               currentPage_9__11), .window_15__10 (currentPage_9__10), .window_15__9 (
               currentPage_9__9), .window_15__8 (currentPage_9__8), .window_15__7 (
               currentPage_9__7), .window_15__6 (currentPage_9__6), .window_15__5 (
               currentPage_9__5), .window_15__4 (currentPage_9__4), .window_15__3 (
               currentPage_9__3), .window_15__2 (currentPage_9__2), .window_15__1 (
               currentPage_9__1), .window_15__0 (currentPage_9__0), .window_14__15 (
               currentPage_10__15), .window_14__14 (currentPage_10__14), .window_14__13 (
               currentPage_10__13), .window_14__12 (currentPage_10__12), .window_14__11 (
               currentPage_10__11), .window_14__10 (currentPage_10__10), .window_14__9 (
               currentPage_10__9), .window_14__8 (currentPage_10__8), .window_14__7 (
               currentPage_10__7), .window_14__6 (currentPage_10__6), .window_14__5 (
               currentPage_10__5), .window_14__4 (currentPage_10__4), .window_14__3 (
               currentPage_10__3), .window_14__2 (currentPage_10__2), .window_14__1 (
               currentPage_10__1), .window_14__0 (currentPage_10__0), .window_13__15 (
               currentPage_11__15), .window_13__14 (currentPage_11__14), .window_13__13 (
               currentPage_11__13), .window_13__12 (currentPage_11__12), .window_13__11 (
               currentPage_11__11), .window_13__10 (currentPage_11__10), .window_13__9 (
               currentPage_11__9), .window_13__8 (currentPage_11__8), .window_13__7 (
               currentPage_11__7), .window_13__6 (currentPage_11__6), .window_13__5 (
               currentPage_11__5), .window_13__4 (currentPage_11__4), .window_13__3 (
               currentPage_11__3), .window_13__2 (currentPage_11__2), .window_13__1 (
               currentPage_11__1), .window_13__0 (currentPage_11__0), .window_12__15 (
               currentPage_12__15), .window_12__14 (currentPage_12__14), .window_12__13 (
               currentPage_12__13), .window_12__12 (currentPage_12__12), .window_12__11 (
               currentPage_12__11), .window_12__10 (currentPage_12__10), .window_12__9 (
               currentPage_12__9), .window_12__8 (currentPage_12__8), .window_12__7 (
               currentPage_12__7), .window_12__6 (currentPage_12__6), .window_12__5 (
               currentPage_12__5), .window_12__4 (currentPage_12__4), .window_12__3 (
               currentPage_12__3), .window_12__2 (currentPage_12__2), .window_12__1 (
               currentPage_12__1), .window_12__0 (currentPage_12__0), .window_11__15 (
               currentPage_13__15), .window_11__14 (currentPage_13__14), .window_11__13 (
               currentPage_13__13), .window_11__12 (currentPage_13__12), .window_11__11 (
               currentPage_13__11), .window_11__10 (currentPage_13__10), .window_11__9 (
               currentPage_13__9), .window_11__8 (currentPage_13__8), .window_11__7 (
               currentPage_13__7), .window_11__6 (currentPage_13__6), .window_11__5 (
               currentPage_13__5), .window_11__4 (currentPage_13__4), .window_11__3 (
               currentPage_13__3), .window_11__2 (currentPage_13__2), .window_11__1 (
               currentPage_13__1), .window_11__0 (currentPage_13__0), .window_10__15 (
               currentPage_14__15), .window_10__14 (currentPage_14__14), .window_10__13 (
               currentPage_14__13), .window_10__12 (currentPage_14__12), .window_10__11 (
               currentPage_14__11), .window_10__10 (currentPage_14__10), .window_10__9 (
               currentPage_14__9), .window_10__8 (currentPage_14__8), .window_10__7 (
               currentPage_14__7), .window_10__6 (currentPage_14__6), .window_10__5 (
               currentPage_14__5), .window_10__4 (currentPage_14__4), .window_10__3 (
               currentPage_14__3), .window_10__2 (currentPage_14__2), .window_10__1 (
               currentPage_14__1), .window_10__0 (currentPage_14__0), .window_9__15 (
               currentPage_15__15), .window_9__14 (currentPage_15__14), .window_9__13 (
               currentPage_15__13), .window_9__12 (currentPage_15__12), .window_9__11 (
               currentPage_15__11), .window_9__10 (currentPage_15__10), .window_9__9 (
               currentPage_15__9), .window_9__8 (currentPage_15__8), .window_9__7 (
               currentPage_15__7), .window_9__6 (currentPage_15__6), .window_9__5 (
               currentPage_15__5), .window_9__4 (currentPage_15__4), .window_9__3 (
               currentPage_15__3), .window_9__2 (currentPage_15__2), .window_9__1 (
               currentPage_15__1), .window_9__0 (currentPage_15__0), .window_8__15 (
               currentPage_16__15), .window_8__14 (currentPage_16__14), .window_8__13 (
               currentPage_16__13), .window_8__12 (currentPage_16__12), .window_8__11 (
               currentPage_16__11), .window_8__10 (currentPage_16__10), .window_8__9 (
               currentPage_16__9), .window_8__8 (currentPage_16__8), .window_8__7 (
               currentPage_16__7), .window_8__6 (currentPage_16__6), .window_8__5 (
               currentPage_16__5), .window_8__4 (currentPage_16__4), .window_8__3 (
               currentPage_16__3), .window_8__2 (currentPage_16__2), .window_8__1 (
               currentPage_16__1), .window_8__0 (currentPage_16__0), .window_7__15 (
               currentPage_17__15), .window_7__14 (currentPage_17__14), .window_7__13 (
               currentPage_17__13), .window_7__12 (currentPage_17__12), .window_7__11 (
               currentPage_17__11), .window_7__10 (currentPage_17__10), .window_7__9 (
               currentPage_17__9), .window_7__8 (currentPage_17__8), .window_7__7 (
               currentPage_17__7), .window_7__6 (currentPage_17__6), .window_7__5 (
               currentPage_17__5), .window_7__4 (currentPage_17__4), .window_7__3 (
               currentPage_17__3), .window_7__2 (currentPage_17__2), .window_7__1 (
               currentPage_17__1), .window_7__0 (currentPage_17__0), .window_6__15 (
               currentPage_18__15), .window_6__14 (currentPage_18__14), .window_6__13 (
               currentPage_18__13), .window_6__12 (currentPage_18__12), .window_6__11 (
               currentPage_18__11), .window_6__10 (currentPage_18__10), .window_6__9 (
               currentPage_18__9), .window_6__8 (currentPage_18__8), .window_6__7 (
               currentPage_18__7), .window_6__6 (currentPage_18__6), .window_6__5 (
               currentPage_18__5), .window_6__4 (currentPage_18__4), .window_6__3 (
               currentPage_18__3), .window_6__2 (currentPage_18__2), .window_6__1 (
               currentPage_18__1), .window_6__0 (currentPage_18__0), .window_5__15 (
               currentPage_19__15), .window_5__14 (currentPage_19__14), .window_5__13 (
               currentPage_19__13), .window_5__12 (currentPage_19__12), .window_5__11 (
               currentPage_19__11), .window_5__10 (currentPage_19__10), .window_5__9 (
               currentPage_19__9), .window_5__8 (currentPage_19__8), .window_5__7 (
               currentPage_19__7), .window_5__6 (currentPage_19__6), .window_5__5 (
               currentPage_19__5), .window_5__4 (currentPage_19__4), .window_5__3 (
               currentPage_19__3), .window_5__2 (currentPage_19__2), .window_5__1 (
               currentPage_19__1), .window_5__0 (currentPage_19__0), .window_4__15 (
               currentPage_20__15), .window_4__14 (currentPage_20__14), .window_4__13 (
               currentPage_20__13), .window_4__12 (currentPage_20__12), .window_4__11 (
               currentPage_20__11), .window_4__10 (currentPage_20__10), .window_4__9 (
               currentPage_20__9), .window_4__8 (currentPage_20__8), .window_4__7 (
               currentPage_20__7), .window_4__6 (currentPage_20__6), .window_4__5 (
               currentPage_20__5), .window_4__4 (currentPage_20__4), .window_4__3 (
               currentPage_20__3), .window_4__2 (currentPage_20__2), .window_4__1 (
               currentPage_20__1), .window_4__0 (currentPage_20__0), .window_3__15 (
               currentPage_21__15), .window_3__14 (currentPage_21__14), .window_3__13 (
               currentPage_21__13), .window_3__12 (currentPage_21__12), .window_3__11 (
               currentPage_21__11), .window_3__10 (currentPage_21__10), .window_3__9 (
               currentPage_21__9), .window_3__8 (currentPage_21__8), .window_3__7 (
               currentPage_21__7), .window_3__6 (currentPage_21__6), .window_3__5 (
               currentPage_21__5), .window_3__4 (currentPage_21__4), .window_3__3 (
               currentPage_21__3), .window_3__2 (currentPage_21__2), .window_3__1 (
               currentPage_21__1), .window_3__0 (currentPage_21__0), .window_2__15 (
               currentPage_22__15), .window_2__14 (currentPage_22__14), .window_2__13 (
               currentPage_22__13), .window_2__12 (currentPage_22__12), .window_2__11 (
               currentPage_22__11), .window_2__10 (currentPage_22__10), .window_2__9 (
               currentPage_22__9), .window_2__8 (currentPage_22__8), .window_2__7 (
               currentPage_22__7), .window_2__6 (currentPage_22__6), .window_2__5 (
               currentPage_22__5), .window_2__4 (currentPage_22__4), .window_2__3 (
               currentPage_22__3), .window_2__2 (currentPage_22__2), .window_2__1 (
               currentPage_22__1), .window_2__0 (currentPage_22__0), .window_1__15 (
               currentPage_23__15), .window_1__14 (currentPage_23__14), .window_1__13 (
               currentPage_23__13), .window_1__12 (currentPage_23__12), .window_1__11 (
               currentPage_23__11), .window_1__10 (currentPage_23__10), .window_1__9 (
               currentPage_23__9), .window_1__8 (currentPage_23__8), .window_1__7 (
               currentPage_23__7), .window_1__6 (currentPage_23__6), .window_1__5 (
               currentPage_23__5), .window_1__4 (currentPage_23__4), .window_1__3 (
               currentPage_23__3), .window_1__2 (currentPage_23__2), .window_1__1 (
               currentPage_23__1), .window_1__0 (currentPage_23__0), .window_0__15 (
               currentPage_24__15), .window_0__14 (currentPage_24__14), .window_0__13 (
               currentPage_24__13), .window_0__12 (currentPage_24__12), .window_0__11 (
               currentPage_24__11), .window_0__10 (currentPage_24__10), .window_0__9 (
               currentPage_24__9), .window_0__8 (currentPage_24__8), .window_0__7 (
               currentPage_24__7), .window_0__6 (currentPage_24__6), .window_0__5 (
               currentPage_24__5), .window_0__4 (currentPage_24__4), .window_0__3 (
               currentPage_24__3), .window_0__2 (currentPage_24__2), .window_0__1 (
               currentPage_24__1), .window_0__0 (currentPage_24__0), .outputs_24__15 (
               outMuls_0__15), .outputs_24__14 (outMuls_0__14), .outputs_24__13 (
               outMuls_0__13), .outputs_24__12 (outMuls_0__12), .outputs_24__11 (
               outMuls_0__11), .outputs_24__10 (outMuls_0__10), .outputs_24__9 (
               outMuls_0__9), .outputs_24__8 (outMuls_0__8), .outputs_24__7 (
               outMuls_0__7), .outputs_24__6 (outMuls_0__6), .outputs_24__5 (
               outMuls_0__5), .outputs_24__4 (outMuls_0__4), .outputs_24__3 (
               outMuls_0__3), .outputs_24__2 (outMuls_0__2), .outputs_24__1 (
               outMuls_0__1), .outputs_24__0 (outMuls_0__0), .outputs_23__15 (
               outMuls_1__15), .outputs_23__14 (outMuls_1__14), .outputs_23__13 (
               outMuls_1__13), .outputs_23__12 (outMuls_1__12), .outputs_23__11 (
               outMuls_1__11), .outputs_23__10 (outMuls_1__10), .outputs_23__9 (
               outMuls_1__9), .outputs_23__8 (outMuls_1__8), .outputs_23__7 (
               outMuls_1__7), .outputs_23__6 (outMuls_1__6), .outputs_23__5 (
               outMuls_1__5), .outputs_23__4 (outMuls_1__4), .outputs_23__3 (
               outMuls_1__3), .outputs_23__2 (outMuls_1__2), .outputs_23__1 (
               outMuls_1__1), .outputs_23__0 (outMuls_1__0), .outputs_22__15 (
               outMuls_2__15), .outputs_22__14 (outMuls_2__14), .outputs_22__13 (
               outMuls_2__13), .outputs_22__12 (outMuls_2__12), .outputs_22__11 (
               outMuls_2__11), .outputs_22__10 (outMuls_2__10), .outputs_22__9 (
               outMuls_2__9), .outputs_22__8 (outMuls_2__8), .outputs_22__7 (
               outMuls_2__7), .outputs_22__6 (outMuls_2__6), .outputs_22__5 (
               outMuls_2__5), .outputs_22__4 (outMuls_2__4), .outputs_22__3 (
               outMuls_2__3), .outputs_22__2 (outMuls_2__2), .outputs_22__1 (
               outMuls_2__1), .outputs_22__0 (outMuls_2__0), .outputs_21__15 (
               outMuls_3__15), .outputs_21__14 (outMuls_3__14), .outputs_21__13 (
               outMuls_3__13), .outputs_21__12 (outMuls_3__12), .outputs_21__11 (
               outMuls_3__11), .outputs_21__10 (outMuls_3__10), .outputs_21__9 (
               outMuls_3__9), .outputs_21__8 (outMuls_3__8), .outputs_21__7 (
               outMuls_3__7), .outputs_21__6 (outMuls_3__6), .outputs_21__5 (
               outMuls_3__5), .outputs_21__4 (outMuls_3__4), .outputs_21__3 (
               outMuls_3__3), .outputs_21__2 (outMuls_3__2), .outputs_21__1 (
               outMuls_3__1), .outputs_21__0 (outMuls_3__0), .outputs_20__15 (
               outMuls_4__15), .outputs_20__14 (outMuls_4__14), .outputs_20__13 (
               outMuls_4__13), .outputs_20__12 (outMuls_4__12), .outputs_20__11 (
               outMuls_4__11), .outputs_20__10 (outMuls_4__10), .outputs_20__9 (
               outMuls_4__9), .outputs_20__8 (outMuls_4__8), .outputs_20__7 (
               outMuls_4__7), .outputs_20__6 (outMuls_4__6), .outputs_20__5 (
               outMuls_4__5), .outputs_20__4 (outMuls_4__4), .outputs_20__3 (
               outMuls_4__3), .outputs_20__2 (outMuls_4__2), .outputs_20__1 (
               outMuls_4__1), .outputs_20__0 (outMuls_4__0), .outputs_19__15 (
               outMuls_5__15), .outputs_19__14 (outMuls_5__14), .outputs_19__13 (
               outMuls_5__13), .outputs_19__12 (outMuls_5__12), .outputs_19__11 (
               outMuls_5__11), .outputs_19__10 (outMuls_5__10), .outputs_19__9 (
               outMuls_5__9), .outputs_19__8 (outMuls_5__8), .outputs_19__7 (
               outMuls_5__7), .outputs_19__6 (outMuls_5__6), .outputs_19__5 (
               outMuls_5__5), .outputs_19__4 (outMuls_5__4), .outputs_19__3 (
               outMuls_5__3), .outputs_19__2 (outMuls_5__2), .outputs_19__1 (
               outMuls_5__1), .outputs_19__0 (outMuls_5__0), .outputs_18__15 (
               outMuls_6__15), .outputs_18__14 (outMuls_6__14), .outputs_18__13 (
               outMuls_6__13), .outputs_18__12 (outMuls_6__12), .outputs_18__11 (
               outMuls_6__11), .outputs_18__10 (outMuls_6__10), .outputs_18__9 (
               outMuls_6__9), .outputs_18__8 (outMuls_6__8), .outputs_18__7 (
               outMuls_6__7), .outputs_18__6 (outMuls_6__6), .outputs_18__5 (
               outMuls_6__5), .outputs_18__4 (outMuls_6__4), .outputs_18__3 (
               outMuls_6__3), .outputs_18__2 (outMuls_6__2), .outputs_18__1 (
               outMuls_6__1), .outputs_18__0 (outMuls_6__0), .outputs_17__15 (
               outMuls_7__15), .outputs_17__14 (outMuls_7__14), .outputs_17__13 (
               outMuls_7__13), .outputs_17__12 (outMuls_7__12), .outputs_17__11 (
               outMuls_7__11), .outputs_17__10 (outMuls_7__10), .outputs_17__9 (
               outMuls_7__9), .outputs_17__8 (outMuls_7__8), .outputs_17__7 (
               outMuls_7__7), .outputs_17__6 (outMuls_7__6), .outputs_17__5 (
               outMuls_7__5), .outputs_17__4 (outMuls_7__4), .outputs_17__3 (
               outMuls_7__3), .outputs_17__2 (outMuls_7__2), .outputs_17__1 (
               outMuls_7__1), .outputs_17__0 (outMuls_7__0), .outputs_16__15 (
               outMuls_8__15), .outputs_16__14 (outMuls_8__14), .outputs_16__13 (
               outMuls_8__13), .outputs_16__12 (outMuls_8__12), .outputs_16__11 (
               outMuls_8__11), .outputs_16__10 (outMuls_8__10), .outputs_16__9 (
               outMuls_8__9), .outputs_16__8 (outMuls_8__8), .outputs_16__7 (
               outMuls_8__7), .outputs_16__6 (outMuls_8__6), .outputs_16__5 (
               outMuls_8__5), .outputs_16__4 (outMuls_8__4), .outputs_16__3 (
               outMuls_8__3), .outputs_16__2 (outMuls_8__2), .outputs_16__1 (
               outMuls_8__1), .outputs_16__0 (outMuls_8__0), .outputs_15__15 (
               outMuls_9__15), .outputs_15__14 (outMuls_9__14), .outputs_15__13 (
               outMuls_9__13), .outputs_15__12 (outMuls_9__12), .outputs_15__11 (
               outMuls_9__11), .outputs_15__10 (outMuls_9__10), .outputs_15__9 (
               outMuls_9__9), .outputs_15__8 (outMuls_9__8), .outputs_15__7 (
               outMuls_9__7), .outputs_15__6 (outMuls_9__6), .outputs_15__5 (
               outMuls_9__5), .outputs_15__4 (outMuls_9__4), .outputs_15__3 (
               outMuls_9__3), .outputs_15__2 (outMuls_9__2), .outputs_15__1 (
               outMuls_9__1), .outputs_15__0 (outMuls_9__0), .outputs_14__15 (
               outMuls_10__15), .outputs_14__14 (outMuls_10__14), .outputs_14__13 (
               outMuls_10__13), .outputs_14__12 (outMuls_10__12), .outputs_14__11 (
               outMuls_10__11), .outputs_14__10 (outMuls_10__10), .outputs_14__9 (
               outMuls_10__9), .outputs_14__8 (outMuls_10__8), .outputs_14__7 (
               outMuls_10__7), .outputs_14__6 (outMuls_10__6), .outputs_14__5 (
               outMuls_10__5), .outputs_14__4 (outMuls_10__4), .outputs_14__3 (
               outMuls_10__3), .outputs_14__2 (outMuls_10__2), .outputs_14__1 (
               outMuls_10__1), .outputs_14__0 (outMuls_10__0), .outputs_13__15 (
               outMuls_11__15), .outputs_13__14 (outMuls_11__14), .outputs_13__13 (
               outMuls_11__13), .outputs_13__12 (outMuls_11__12), .outputs_13__11 (
               outMuls_11__11), .outputs_13__10 (outMuls_11__10), .outputs_13__9 (
               outMuls_11__9), .outputs_13__8 (outMuls_11__8), .outputs_13__7 (
               outMuls_11__7), .outputs_13__6 (outMuls_11__6), .outputs_13__5 (
               outMuls_11__5), .outputs_13__4 (outMuls_11__4), .outputs_13__3 (
               outMuls_11__3), .outputs_13__2 (outMuls_11__2), .outputs_13__1 (
               outMuls_11__1), .outputs_13__0 (outMuls_11__0), .outputs_12__15 (
               outMuls_12__15), .outputs_12__14 (outMuls_12__14), .outputs_12__13 (
               outMuls_12__13), .outputs_12__12 (outMuls_12__12), .outputs_12__11 (
               outMuls_12__11), .outputs_12__10 (outMuls_12__10), .outputs_12__9 (
               outMuls_12__9), .outputs_12__8 (outMuls_12__8), .outputs_12__7 (
               outMuls_12__7), .outputs_12__6 (outMuls_12__6), .outputs_12__5 (
               outMuls_12__5), .outputs_12__4 (outMuls_12__4), .outputs_12__3 (
               outMuls_12__3), .outputs_12__2 (outMuls_12__2), .outputs_12__1 (
               outMuls_12__1), .outputs_12__0 (outMuls_12__0), .outputs_11__15 (
               outMuls_13__15), .outputs_11__14 (outMuls_13__14), .outputs_11__13 (
               outMuls_13__13), .outputs_11__12 (outMuls_13__12), .outputs_11__11 (
               outMuls_13__11), .outputs_11__10 (outMuls_13__10), .outputs_11__9 (
               outMuls_13__9), .outputs_11__8 (outMuls_13__8), .outputs_11__7 (
               outMuls_13__7), .outputs_11__6 (outMuls_13__6), .outputs_11__5 (
               outMuls_13__5), .outputs_11__4 (outMuls_13__4), .outputs_11__3 (
               outMuls_13__3), .outputs_11__2 (outMuls_13__2), .outputs_11__1 (
               outMuls_13__1), .outputs_11__0 (outMuls_13__0), .outputs_10__15 (
               outMuls_14__15), .outputs_10__14 (outMuls_14__14), .outputs_10__13 (
               outMuls_14__13), .outputs_10__12 (outMuls_14__12), .outputs_10__11 (
               outMuls_14__11), .outputs_10__10 (outMuls_14__10), .outputs_10__9 (
               outMuls_14__9), .outputs_10__8 (outMuls_14__8), .outputs_10__7 (
               outMuls_14__7), .outputs_10__6 (outMuls_14__6), .outputs_10__5 (
               outMuls_14__5), .outputs_10__4 (outMuls_14__4), .outputs_10__3 (
               outMuls_14__3), .outputs_10__2 (outMuls_14__2), .outputs_10__1 (
               outMuls_14__1), .outputs_10__0 (outMuls_14__0), .outputs_9__15 (
               outMuls_15__15), .outputs_9__14 (outMuls_15__14), .outputs_9__13 (
               outMuls_15__13), .outputs_9__12 (outMuls_15__12), .outputs_9__11 (
               outMuls_15__11), .outputs_9__10 (outMuls_15__10), .outputs_9__9 (
               outMuls_15__9), .outputs_9__8 (outMuls_15__8), .outputs_9__7 (
               outMuls_15__7), .outputs_9__6 (outMuls_15__6), .outputs_9__5 (
               outMuls_15__5), .outputs_9__4 (outMuls_15__4), .outputs_9__3 (
               outMuls_15__3), .outputs_9__2 (outMuls_15__2), .outputs_9__1 (
               outMuls_15__1), .outputs_9__0 (outMuls_15__0), .outputs_8__15 (
               outMuls_16__15), .outputs_8__14 (outMuls_16__14), .outputs_8__13 (
               outMuls_16__13), .outputs_8__12 (outMuls_16__12), .outputs_8__11 (
               outMuls_16__11), .outputs_8__10 (outMuls_16__10), .outputs_8__9 (
               outMuls_16__9), .outputs_8__8 (outMuls_16__8), .outputs_8__7 (
               outMuls_16__7), .outputs_8__6 (outMuls_16__6), .outputs_8__5 (
               outMuls_16__5), .outputs_8__4 (outMuls_16__4), .outputs_8__3 (
               outMuls_16__3), .outputs_8__2 (outMuls_16__2), .outputs_8__1 (
               outMuls_16__1), .outputs_8__0 (outMuls_16__0), .outputs_7__15 (
               outMuls_17__15), .outputs_7__14 (outMuls_17__14), .outputs_7__13 (
               outMuls_17__13), .outputs_7__12 (outMuls_17__12), .outputs_7__11 (
               outMuls_17__11), .outputs_7__10 (outMuls_17__10), .outputs_7__9 (
               outMuls_17__9), .outputs_7__8 (outMuls_17__8), .outputs_7__7 (
               outMuls_17__7), .outputs_7__6 (outMuls_17__6), .outputs_7__5 (
               outMuls_17__5), .outputs_7__4 (outMuls_17__4), .outputs_7__3 (
               outMuls_17__3), .outputs_7__2 (outMuls_17__2), .outputs_7__1 (
               outMuls_17__1), .outputs_7__0 (outMuls_17__0), .outputs_6__15 (
               outMuls_18__15), .outputs_6__14 (outMuls_18__14), .outputs_6__13 (
               outMuls_18__13), .outputs_6__12 (outMuls_18__12), .outputs_6__11 (
               outMuls_18__11), .outputs_6__10 (outMuls_18__10), .outputs_6__9 (
               outMuls_18__9), .outputs_6__8 (outMuls_18__8), .outputs_6__7 (
               outMuls_18__7), .outputs_6__6 (outMuls_18__6), .outputs_6__5 (
               outMuls_18__5), .outputs_6__4 (outMuls_18__4), .outputs_6__3 (
               outMuls_18__3), .outputs_6__2 (outMuls_18__2), .outputs_6__1 (
               outMuls_18__1), .outputs_6__0 (outMuls_18__0), .outputs_5__15 (
               outMuls_19__15), .outputs_5__14 (outMuls_19__14), .outputs_5__13 (
               outMuls_19__13), .outputs_5__12 (outMuls_19__12), .outputs_5__11 (
               outMuls_19__11), .outputs_5__10 (outMuls_19__10), .outputs_5__9 (
               outMuls_19__9), .outputs_5__8 (outMuls_19__8), .outputs_5__7 (
               outMuls_19__7), .outputs_5__6 (outMuls_19__6), .outputs_5__5 (
               outMuls_19__5), .outputs_5__4 (outMuls_19__4), .outputs_5__3 (
               outMuls_19__3), .outputs_5__2 (outMuls_19__2), .outputs_5__1 (
               outMuls_19__1), .outputs_5__0 (outMuls_19__0), .outputs_4__15 (
               outMuls_20__15), .outputs_4__14 (outMuls_20__14), .outputs_4__13 (
               outMuls_20__13), .outputs_4__12 (outMuls_20__12), .outputs_4__11 (
               outMuls_20__11), .outputs_4__10 (outMuls_20__10), .outputs_4__9 (
               outMuls_20__9), .outputs_4__8 (outMuls_20__8), .outputs_4__7 (
               outMuls_20__7), .outputs_4__6 (outMuls_20__6), .outputs_4__5 (
               outMuls_20__5), .outputs_4__4 (outMuls_20__4), .outputs_4__3 (
               outMuls_20__3), .outputs_4__2 (outMuls_20__2), .outputs_4__1 (
               outMuls_20__1), .outputs_4__0 (outMuls_20__0), .outputs_3__15 (
               outMuls_21__15), .outputs_3__14 (outMuls_21__14), .outputs_3__13 (
               outMuls_21__13), .outputs_3__12 (outMuls_21__12), .outputs_3__11 (
               outMuls_21__11), .outputs_3__10 (outMuls_21__10), .outputs_3__9 (
               outMuls_21__9), .outputs_3__8 (outMuls_21__8), .outputs_3__7 (
               outMuls_21__7), .outputs_3__6 (outMuls_21__6), .outputs_3__5 (
               outMuls_21__5), .outputs_3__4 (outMuls_21__4), .outputs_3__3 (
               outMuls_21__3), .outputs_3__2 (outMuls_21__2), .outputs_3__1 (
               outMuls_21__1), .outputs_3__0 (outMuls_21__0), .outputs_2__15 (
               outMuls_22__15), .outputs_2__14 (outMuls_22__14), .outputs_2__13 (
               outMuls_22__13), .outputs_2__12 (outMuls_22__12), .outputs_2__11 (
               outMuls_22__11), .outputs_2__10 (outMuls_22__10), .outputs_2__9 (
               outMuls_22__9), .outputs_2__8 (outMuls_22__8), .outputs_2__7 (
               outMuls_22__7), .outputs_2__6 (outMuls_22__6), .outputs_2__5 (
               outMuls_22__5), .outputs_2__4 (outMuls_22__4), .outputs_2__3 (
               outMuls_22__3), .outputs_2__2 (outMuls_22__2), .outputs_2__1 (
               outMuls_22__1), .outputs_2__0 (outMuls_22__0), .outputs_1__15 (
               outMuls_23__15), .outputs_1__14 (outMuls_23__14), .outputs_1__13 (
               outMuls_23__13), .outputs_1__12 (outMuls_23__12), .outputs_1__11 (
               outMuls_23__11), .outputs_1__10 (outMuls_23__10), .outputs_1__9 (
               outMuls_23__9), .outputs_1__8 (outMuls_23__8), .outputs_1__7 (
               outMuls_23__7), .outputs_1__6 (outMuls_23__6), .outputs_1__5 (
               outMuls_23__5), .outputs_1__4 (outMuls_23__4), .outputs_1__3 (
               outMuls_23__3), .outputs_1__2 (outMuls_23__2), .outputs_1__1 (
               outMuls_23__1), .outputs_1__0 (outMuls_23__0), .outputs_0__15 (
               outMuls_24__15), .outputs_0__14 (outMuls_24__14), .outputs_0__13 (
               outMuls_24__13), .outputs_0__12 (outMuls_24__12), .outputs_0__11 (
               outMuls_24__11), .outputs_0__10 (outMuls_24__10), .outputs_0__9 (
               outMuls_24__9), .outputs_0__8 (outMuls_24__8), .outputs_0__7 (
               outMuls_24__7), .outputs_0__6 (outMuls_24__6), .outputs_0__5 (
               outMuls_24__5), .outputs_0__4 (outMuls_24__4), .outputs_0__3 (
               outMuls_24__3), .outputs_0__2 (outMuls_24__2), .outputs_0__1 (
               outMuls_24__1), .outputs_0__0 (outMuls_24__0), .clk (clk), .start (
               start), .rst (rst), .done (doneMul), .working (\$dummy [0])) ;
    RegUnit_8_16 regFileMap_loop1_0_regRowMap_loop1_0_regUnitMap (.filterBus ({
                 filterBus[7],filterBus[6],filterBus[5],filterBus[4],
                 filterBus[3],filterBus[2],filterBus[1],filterBus[0]}), .windowBus (
                 {windowBus[15],windowBus[14],windowBus[13],windowBus[12],
                 windowBus[11],windowBus[10],windowBus[9],windowBus[8],
                 windowBus[7],windowBus[6],windowBus[5],windowBus[4],
                 windowBus[3],windowBus[2],windowBus[1],windowBus[0]}), .regPage1NextUnit (
                 {regFileMap_page1Out_5__15,regFileMap_page1Out_5__14,
                 regFileMap_page1Out_5__13,regFileMap_page1Out_5__12,
                 regFileMap_page1Out_5__11,regFileMap_page1Out_5__10,
                 regFileMap_page1Out_5__9,regFileMap_page1Out_5__8,
                 regFileMap_page1Out_5__7,regFileMap_page1Out_5__6,
                 regFileMap_page1Out_5__5,regFileMap_page1Out_5__4,
                 regFileMap_page1Out_5__3,regFileMap_page1Out_5__2,
                 regFileMap_page1Out_5__1,regFileMap_page1Out_5__0}), .regPage2NextUnit (
                 {regFileMap_page2Out_5__15,regFileMap_page2Out_5__14,
                 regFileMap_page2Out_5__13,regFileMap_page2Out_5__12,
                 regFileMap_page2Out_5__11,regFileMap_page2Out_5__10,
                 regFileMap_page2Out_5__9,regFileMap_page2Out_5__8,
                 regFileMap_page2Out_5__7,regFileMap_page2Out_5__6,
                 regFileMap_page2Out_5__5,regFileMap_page2Out_5__4,
                 regFileMap_page2Out_5__3,regFileMap_page2Out_5__2,
                 regFileMap_page2Out_5__1,regFileMap_page2Out_5__0}), .clk (clk)
                 , .rst (rst), .enableRegPage1 (regFileMap_page1Enables_0), .enableRegPage2 (
                 regFileMap_page2Enables_0), .enableRegFilter (nx5328), .page1ReadBusOrPage2 (
                 shift2To1), .page2ReadBusOrPage1 (shift1To2), .pageTurn (
                 pageTurn), .outRegPage ({currentPage_0__15,currentPage_0__14,
                 currentPage_0__13,currentPage_0__12,currentPage_0__11,
                 currentPage_0__10,currentPage_0__9,currentPage_0__8,
                 currentPage_0__7,currentPage_0__6,currentPage_0__5,
                 currentPage_0__4,currentPage_0__3,currentPage_0__2,
                 currentPage_0__1,currentPage_0__0}), .outputRegPage1 ({
                 \$dummy [1],\$dummy [2],\$dummy [3],\$dummy [4],\$dummy [5],
                 \$dummy [6],\$dummy [7],\$dummy [8],\$dummy [9],\$dummy [10],
                 \$dummy [11],\$dummy [12],\$dummy [13],\$dummy [14],
                 \$dummy [15],\$dummy [16]}), .outputRegPage2 ({\$dummy [17],
                 \$dummy [18],\$dummy [19],\$dummy [20],\$dummy [21],
                 \$dummy [22],\$dummy [23],\$dummy [24],\$dummy [25],
                 \$dummy [26],\$dummy [27],\$dummy [28],\$dummy [29],
                 \$dummy [30],\$dummy [31],\$dummy [32]}), .outFilter ({
                 filter_0__7,filter_0__6,filter_0__5,filter_0__4,filter_0__3,
                 filter_0__2,filter_0__1,filter_0__0})) ;
    RegUnit_8_16 regFileMap_loop1_0_regRowMap_loop1_1_regUnitMap (.filterBus ({
                 filterBus[15],filterBus[14],filterBus[13],filterBus[12],
                 filterBus[11],filterBus[10],filterBus[9],filterBus[8]}), .windowBus (
                 {windowBus[31],windowBus[30],windowBus[29],windowBus[28],
                 windowBus[27],windowBus[26],windowBus[25],windowBus[24],
                 windowBus[23],windowBus[22],windowBus[21],windowBus[20],
                 windowBus[19],windowBus[18],windowBus[17],windowBus[16]}), .regPage1NextUnit (
                 {regFileMap_page1Out_6__15,regFileMap_page1Out_6__14,
                 regFileMap_page1Out_6__13,regFileMap_page1Out_6__12,
                 regFileMap_page1Out_6__11,regFileMap_page1Out_6__10,
                 regFileMap_page1Out_6__9,regFileMap_page1Out_6__8,
                 regFileMap_page1Out_6__7,regFileMap_page1Out_6__6,
                 regFileMap_page1Out_6__5,regFileMap_page1Out_6__4,
                 regFileMap_page1Out_6__3,regFileMap_page1Out_6__2,
                 regFileMap_page1Out_6__1,regFileMap_page1Out_6__0}), .regPage2NextUnit (
                 {regFileMap_page2Out_6__15,regFileMap_page2Out_6__14,
                 regFileMap_page2Out_6__13,regFileMap_page2Out_6__12,
                 regFileMap_page2Out_6__11,regFileMap_page2Out_6__10,
                 regFileMap_page2Out_6__9,regFileMap_page2Out_6__8,
                 regFileMap_page2Out_6__7,regFileMap_page2Out_6__6,
                 regFileMap_page2Out_6__5,regFileMap_page2Out_6__4,
                 regFileMap_page2Out_6__3,regFileMap_page2Out_6__2,
                 regFileMap_page2Out_6__1,regFileMap_page2Out_6__0}), .clk (clk)
                 , .rst (rst), .enableRegPage1 (regFileMap_page1Enables_0), .enableRegPage2 (
                 regFileMap_page2Enables_0), .enableRegFilter (nx5328), .page1ReadBusOrPage2 (
                 shift2To1), .page2ReadBusOrPage1 (shift1To2), .pageTurn (
                 pageTurn), .outRegPage ({currentPage_1__15,currentPage_1__14,
                 currentPage_1__13,currentPage_1__12,currentPage_1__11,
                 currentPage_1__10,currentPage_1__9,currentPage_1__8,
                 currentPage_1__7,currentPage_1__6,currentPage_1__5,
                 currentPage_1__4,currentPage_1__3,currentPage_1__2,
                 currentPage_1__1,currentPage_1__0}), .outputRegPage1 ({
                 \$dummy [33],\$dummy [34],\$dummy [35],\$dummy [36],
                 \$dummy [37],\$dummy [38],\$dummy [39],\$dummy [40],
                 \$dummy [41],\$dummy [42],\$dummy [43],\$dummy [44],
                 \$dummy [45],\$dummy [46],\$dummy [47],\$dummy [48]}), .outputRegPage2 (
                 {\$dummy [49],\$dummy [50],\$dummy [51],\$dummy [52],
                 \$dummy [53],\$dummy [54],\$dummy [55],\$dummy [56],
                 \$dummy [57],\$dummy [58],\$dummy [59],\$dummy [60],
                 \$dummy [61],\$dummy [62],\$dummy [63],\$dummy [64]}), .outFilter (
                 {filter_1__7,filter_1__6,filter_1__5,filter_1__4,filter_1__3,
                 filter_1__2,filter_1__1,filter_1__0})) ;
    RegUnit_8_16 regFileMap_loop1_0_regRowMap_loop1_2_regUnitMap (.filterBus ({
                 filterBus[23],filterBus[22],filterBus[21],filterBus[20],
                 filterBus[19],filterBus[18],filterBus[17],filterBus[16]}), .windowBus (
                 {windowBus[47],windowBus[46],windowBus[45],windowBus[44],
                 windowBus[43],windowBus[42],windowBus[41],windowBus[40],
                 windowBus[39],windowBus[38],windowBus[37],windowBus[36],
                 windowBus[35],windowBus[34],windowBus[33],windowBus[32]}), .regPage1NextUnit (
                 {regFileMap_page1Out_7__15,regFileMap_page1Out_7__14,
                 regFileMap_page1Out_7__13,regFileMap_page1Out_7__12,
                 regFileMap_page1Out_7__11,regFileMap_page1Out_7__10,
                 regFileMap_page1Out_7__9,regFileMap_page1Out_7__8,
                 regFileMap_page1Out_7__7,regFileMap_page1Out_7__6,
                 regFileMap_page1Out_7__5,regFileMap_page1Out_7__4,
                 regFileMap_page1Out_7__3,regFileMap_page1Out_7__2,
                 regFileMap_page1Out_7__1,regFileMap_page1Out_7__0}), .regPage2NextUnit (
                 {regFileMap_page2Out_7__15,regFileMap_page2Out_7__14,
                 regFileMap_page2Out_7__13,regFileMap_page2Out_7__12,
                 regFileMap_page2Out_7__11,regFileMap_page2Out_7__10,
                 regFileMap_page2Out_7__9,regFileMap_page2Out_7__8,
                 regFileMap_page2Out_7__7,regFileMap_page2Out_7__6,
                 regFileMap_page2Out_7__5,regFileMap_page2Out_7__4,
                 regFileMap_page2Out_7__3,regFileMap_page2Out_7__2,
                 regFileMap_page2Out_7__1,regFileMap_page2Out_7__0}), .clk (clk)
                 , .rst (rst), .enableRegPage1 (regFileMap_page1Enables_0), .enableRegPage2 (
                 regFileMap_page2Enables_0), .enableRegFilter (nx5328), .page1ReadBusOrPage2 (
                 shift2To1), .page2ReadBusOrPage1 (shift1To2), .pageTurn (
                 pageTurn), .outRegPage ({currentPage_2__15,currentPage_2__14,
                 currentPage_2__13,currentPage_2__12,currentPage_2__11,
                 currentPage_2__10,currentPage_2__9,currentPage_2__8,
                 currentPage_2__7,currentPage_2__6,currentPage_2__5,
                 currentPage_2__4,currentPage_2__3,currentPage_2__2,
                 currentPage_2__1,currentPage_2__0}), .outputRegPage1 ({
                 \$dummy [65],\$dummy [66],\$dummy [67],\$dummy [68],
                 \$dummy [69],\$dummy [70],\$dummy [71],\$dummy [72],
                 \$dummy [73],\$dummy [74],\$dummy [75],\$dummy [76],
                 \$dummy [77],\$dummy [78],\$dummy [79],\$dummy [80]}), .outputRegPage2 (
                 {\$dummy [81],\$dummy [82],\$dummy [83],\$dummy [84],
                 \$dummy [85],\$dummy [86],\$dummy [87],\$dummy [88],
                 \$dummy [89],\$dummy [90],\$dummy [91],\$dummy [92],
                 \$dummy [93],\$dummy [94],\$dummy [95],\$dummy [96]}), .outFilter (
                 {filter_2__7,filter_2__6,filter_2__5,filter_2__4,filter_2__3,
                 filter_2__2,filter_2__1,filter_2__0})) ;
    RegUnit_8_16 regFileMap_loop1_0_regRowMap_loop1_3_regUnitMap (.filterBus ({
                 filterBus[31],filterBus[30],filterBus[29],filterBus[28],
                 filterBus[27],filterBus[26],filterBus[25],filterBus[24]}), .windowBus (
                 {windowBus[63],windowBus[62],windowBus[61],windowBus[60],
                 windowBus[59],windowBus[58],windowBus[57],windowBus[56],
                 windowBus[55],windowBus[54],windowBus[53],windowBus[52],
                 windowBus[51],windowBus[50],windowBus[49],windowBus[48]}), .regPage1NextUnit (
                 {regFileMap_page1Out_8__15,regFileMap_page1Out_8__14,
                 regFileMap_page1Out_8__13,regFileMap_page1Out_8__12,
                 regFileMap_page1Out_8__11,regFileMap_page1Out_8__10,
                 regFileMap_page1Out_8__9,regFileMap_page1Out_8__8,
                 regFileMap_page1Out_8__7,regFileMap_page1Out_8__6,
                 regFileMap_page1Out_8__5,regFileMap_page1Out_8__4,
                 regFileMap_page1Out_8__3,regFileMap_page1Out_8__2,
                 regFileMap_page1Out_8__1,regFileMap_page1Out_8__0}), .regPage2NextUnit (
                 {regFileMap_page2Out_8__15,regFileMap_page2Out_8__14,
                 regFileMap_page2Out_8__13,regFileMap_page2Out_8__12,
                 regFileMap_page2Out_8__11,regFileMap_page2Out_8__10,
                 regFileMap_page2Out_8__9,regFileMap_page2Out_8__8,
                 regFileMap_page2Out_8__7,regFileMap_page2Out_8__6,
                 regFileMap_page2Out_8__5,regFileMap_page2Out_8__4,
                 regFileMap_page2Out_8__3,regFileMap_page2Out_8__2,
                 regFileMap_page2Out_8__1,regFileMap_page2Out_8__0}), .clk (clk)
                 , .rst (rst), .enableRegPage1 (regFileMap_page1Enables_0), .enableRegPage2 (
                 regFileMap_page2Enables_0), .enableRegFilter (nx5330), .page1ReadBusOrPage2 (
                 shift2To1), .page2ReadBusOrPage1 (shift1To2), .pageTurn (
                 pageTurn), .outRegPage ({currentPage_15__15,currentPage_15__14,
                 currentPage_15__13,currentPage_15__12,currentPage_15__11,
                 currentPage_15__10,currentPage_15__9,currentPage_15__8,
                 currentPage_15__7,currentPage_15__6,currentPage_15__5,
                 currentPage_15__4,currentPage_15__3,currentPage_15__2,
                 currentPage_15__1,currentPage_15__0}), .outputRegPage1 ({
                 \$dummy [97],\$dummy [98],\$dummy [99],\$dummy [100],
                 \$dummy [101],\$dummy [102],\$dummy [103],\$dummy [104],
                 \$dummy [105],\$dummy [106],\$dummy [107],\$dummy [108],
                 \$dummy [109],\$dummy [110],\$dummy [111],\$dummy [112]}), .outputRegPage2 (
                 {\$dummy [113],\$dummy [114],\$dummy [115],\$dummy [116],
                 \$dummy [117],\$dummy [118],\$dummy [119],\$dummy [120],
                 \$dummy [121],\$dummy [122],\$dummy [123],\$dummy [124],
                 \$dummy [125],\$dummy [126],\$dummy [127],\$dummy [128]}), .outFilter (
                 {filter_15__7,filter_15__6,filter_15__5,filter_15__4,
                 filter_15__3,filter_15__2,filter_15__1,filter_15__0})) ;
    RegUnit_8_16 regFileMap_loop1_0_regRowMap_loop1_4_regUnitMap (.filterBus ({
                 filterBus[39],filterBus[38],filterBus[37],filterBus[36],
                 filterBus[35],filterBus[34],filterBus[33],filterBus[32]}), .windowBus (
                 {windowBus[79],windowBus[78],windowBus[77],windowBus[76],
                 windowBus[75],windowBus[74],windowBus[73],windowBus[72],
                 windowBus[71],windowBus[70],windowBus[69],windowBus[68],
                 windowBus[67],windowBus[66],windowBus[65],windowBus[64]}), .regPage1NextUnit (
                 {regFileMap_page1Out_9__15,regFileMap_page1Out_9__14,
                 regFileMap_page1Out_9__13,regFileMap_page1Out_9__12,
                 regFileMap_page1Out_9__11,regFileMap_page1Out_9__10,
                 regFileMap_page1Out_9__9,regFileMap_page1Out_9__8,
                 regFileMap_page1Out_9__7,regFileMap_page1Out_9__6,
                 regFileMap_page1Out_9__5,regFileMap_page1Out_9__4,
                 regFileMap_page1Out_9__3,regFileMap_page1Out_9__2,
                 regFileMap_page1Out_9__1,regFileMap_page1Out_9__0}), .regPage2NextUnit (
                 {regFileMap_page2Out_9__15,regFileMap_page2Out_9__14,
                 regFileMap_page2Out_9__13,regFileMap_page2Out_9__12,
                 regFileMap_page2Out_9__11,regFileMap_page2Out_9__10,
                 regFileMap_page2Out_9__9,regFileMap_page2Out_9__8,
                 regFileMap_page2Out_9__7,regFileMap_page2Out_9__6,
                 regFileMap_page2Out_9__5,regFileMap_page2Out_9__4,
                 regFileMap_page2Out_9__3,regFileMap_page2Out_9__2,
                 regFileMap_page2Out_9__1,regFileMap_page2Out_9__0}), .clk (clk)
                 , .rst (rst), .enableRegPage1 (regFileMap_page1Enables_0), .enableRegPage2 (
                 regFileMap_page2Enables_0), .enableRegFilter (nx5330), .page1ReadBusOrPage2 (
                 shift2To1), .page2ReadBusOrPage1 (shift1To2), .pageTurn (
                 pageTurn), .outRegPage ({currentPage_16__15,currentPage_16__14,
                 currentPage_16__13,currentPage_16__12,currentPage_16__11,
                 currentPage_16__10,currentPage_16__9,currentPage_16__8,
                 currentPage_16__7,currentPage_16__6,currentPage_16__5,
                 currentPage_16__4,currentPage_16__3,currentPage_16__2,
                 currentPage_16__1,currentPage_16__0}), .outputRegPage1 ({
                 \$dummy [129],\$dummy [130],\$dummy [131],\$dummy [132],
                 \$dummy [133],\$dummy [134],\$dummy [135],\$dummy [136],
                 \$dummy [137],\$dummy [138],\$dummy [139],\$dummy [140],
                 \$dummy [141],\$dummy [142],\$dummy [143],\$dummy [144]}), .outputRegPage2 (
                 {\$dummy [145],\$dummy [146],\$dummy [147],\$dummy [148],
                 \$dummy [149],\$dummy [150],\$dummy [151],\$dummy [152],
                 \$dummy [153],\$dummy [154],\$dummy [155],\$dummy [156],
                 \$dummy [157],\$dummy [158],\$dummy [159],\$dummy [160]}), .outFilter (
                 {filter_16__7,filter_16__6,filter_16__5,filter_16__4,
                 filter_16__3,filter_16__2,filter_16__1,filter_16__0})) ;
    RegUnit_8_16_unfolded0 regFileMap_loop1_1_regRowMap_loop1_0_regUnitMap (.filterBus (
                           {filterBus[7],filterBus[6],filterBus[5],filterBus[4],
                           filterBus[3],filterBus[2],filterBus[1],filterBus[0]})
                           , .windowBus ({windowBus[15],windowBus[14],
                           windowBus[13],windowBus[12],windowBus[11],
                           windowBus[10],windowBus[9],windowBus[8],windowBus[7],
                           windowBus[6],windowBus[5],windowBus[4],windowBus[3],
                           windowBus[2],windowBus[1],windowBus[0]}), .regPage1NextUnit (
                           {regFileMap_page1Out_10__15,
                           regFileMap_page1Out_10__14,regFileMap_page1Out_10__13
                           ,regFileMap_page1Out_10__12,
                           regFileMap_page1Out_10__11,regFileMap_page1Out_10__10
                           ,regFileMap_page1Out_10__9,regFileMap_page1Out_10__8,
                           regFileMap_page1Out_10__7,regFileMap_page1Out_10__6,
                           regFileMap_page1Out_10__5,regFileMap_page1Out_10__4,
                           regFileMap_page1Out_10__3,regFileMap_page1Out_10__2,
                           regFileMap_page1Out_10__1,regFileMap_page1Out_10__0})
                           , .regPage2NextUnit ({regFileMap_page2Out_10__15,
                           regFileMap_page2Out_10__14,regFileMap_page2Out_10__13
                           ,regFileMap_page2Out_10__12,
                           regFileMap_page2Out_10__11,regFileMap_page2Out_10__10
                           ,regFileMap_page2Out_10__9,regFileMap_page2Out_10__8,
                           regFileMap_page2Out_10__7,regFileMap_page2Out_10__6,
                           regFileMap_page2Out_10__5,regFileMap_page2Out_10__4,
                           regFileMap_page2Out_10__3,regFileMap_page2Out_10__2,
                           regFileMap_page2Out_10__1,regFileMap_page2Out_10__0})
                           , .clk (clk), .rst (rst), .enableRegPage1 (
                           regFileMap_page1Enables_1), .enableRegPage2 (
                           regFileMap_page2Enables_1), .enableRegFilter (nx5332)
                           , .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           currentPage_3__15,currentPage_3__14,currentPage_3__13
                           ,currentPage_3__12,currentPage_3__11,
                           currentPage_3__10,currentPage_3__9,currentPage_3__8,
                           currentPage_3__7,currentPage_3__6,currentPage_3__5,
                           currentPage_3__4,currentPage_3__3,currentPage_3__2,
                           currentPage_3__1,currentPage_3__0}), .outputRegPage1 (
                           {regFileMap_page1Out_5__15,regFileMap_page1Out_5__14,
                           regFileMap_page1Out_5__13,regFileMap_page1Out_5__12,
                           regFileMap_page1Out_5__11,regFileMap_page1Out_5__10,
                           regFileMap_page1Out_5__9,regFileMap_page1Out_5__8,
                           regFileMap_page1Out_5__7,regFileMap_page1Out_5__6,
                           regFileMap_page1Out_5__5,regFileMap_page1Out_5__4,
                           regFileMap_page1Out_5__3,regFileMap_page1Out_5__2,
                           regFileMap_page1Out_5__1,regFileMap_page1Out_5__0}), 
                           .outputRegPage2 ({regFileMap_page2Out_5__15,
                           regFileMap_page2Out_5__14,regFileMap_page2Out_5__13,
                           regFileMap_page2Out_5__12,regFileMap_page2Out_5__11,
                           regFileMap_page2Out_5__10,regFileMap_page2Out_5__9,
                           regFileMap_page2Out_5__8,regFileMap_page2Out_5__7,
                           regFileMap_page2Out_5__6,regFileMap_page2Out_5__5,
                           regFileMap_page2Out_5__4,regFileMap_page2Out_5__3,
                           regFileMap_page2Out_5__2,regFileMap_page2Out_5__1,
                           regFileMap_page2Out_5__0}), .outFilter ({filter_3__7,
                           filter_3__6,filter_3__5,filter_3__4,filter_3__3,
                           filter_3__2,filter_3__1,filter_3__0})) ;
    RegUnit_8_16_unfolded0 regFileMap_loop1_1_regRowMap_loop1_1_regUnitMap (.filterBus (
                           {filterBus[15],filterBus[14],filterBus[13],
                           filterBus[12],filterBus[11],filterBus[10],
                           filterBus[9],filterBus[8]}), .windowBus ({
                           windowBus[31],windowBus[30],windowBus[29],
                           windowBus[28],windowBus[27],windowBus[26],
                           windowBus[25],windowBus[24],windowBus[23],
                           windowBus[22],windowBus[21],windowBus[20],
                           windowBus[19],windowBus[18],windowBus[17],
                           windowBus[16]}), .regPage1NextUnit ({
                           regFileMap_page1Out_11__15,regFileMap_page1Out_11__14
                           ,regFileMap_page1Out_11__13,
                           regFileMap_page1Out_11__12,regFileMap_page1Out_11__11
                           ,regFileMap_page1Out_11__10,regFileMap_page1Out_11__9
                           ,regFileMap_page1Out_11__8,regFileMap_page1Out_11__7,
                           regFileMap_page1Out_11__6,regFileMap_page1Out_11__5,
                           regFileMap_page1Out_11__4,regFileMap_page1Out_11__3,
                           regFileMap_page1Out_11__2,regFileMap_page1Out_11__1,
                           regFileMap_page1Out_11__0}), .regPage2NextUnit ({
                           regFileMap_page2Out_11__15,regFileMap_page2Out_11__14
                           ,regFileMap_page2Out_11__13,
                           regFileMap_page2Out_11__12,regFileMap_page2Out_11__11
                           ,regFileMap_page2Out_11__10,regFileMap_page2Out_11__9
                           ,regFileMap_page2Out_11__8,regFileMap_page2Out_11__7,
                           regFileMap_page2Out_11__6,regFileMap_page2Out_11__5,
                           regFileMap_page2Out_11__4,regFileMap_page2Out_11__3,
                           regFileMap_page2Out_11__2,regFileMap_page2Out_11__1,
                           regFileMap_page2Out_11__0}), .clk (clk), .rst (rst), 
                           .enableRegPage1 (regFileMap_page1Enables_1), .enableRegPage2 (
                           regFileMap_page2Enables_1), .enableRegFilter (nx5332)
                           , .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           currentPage_4__15,currentPage_4__14,currentPage_4__13
                           ,currentPage_4__12,currentPage_4__11,
                           currentPage_4__10,currentPage_4__9,currentPage_4__8,
                           currentPage_4__7,currentPage_4__6,currentPage_4__5,
                           currentPage_4__4,currentPage_4__3,currentPage_4__2,
                           currentPage_4__1,currentPage_4__0}), .outputRegPage1 (
                           {regFileMap_page1Out_6__15,regFileMap_page1Out_6__14,
                           regFileMap_page1Out_6__13,regFileMap_page1Out_6__12,
                           regFileMap_page1Out_6__11,regFileMap_page1Out_6__10,
                           regFileMap_page1Out_6__9,regFileMap_page1Out_6__8,
                           regFileMap_page1Out_6__7,regFileMap_page1Out_6__6,
                           regFileMap_page1Out_6__5,regFileMap_page1Out_6__4,
                           regFileMap_page1Out_6__3,regFileMap_page1Out_6__2,
                           regFileMap_page1Out_6__1,regFileMap_page1Out_6__0}), 
                           .outputRegPage2 ({regFileMap_page2Out_6__15,
                           regFileMap_page2Out_6__14,regFileMap_page2Out_6__13,
                           regFileMap_page2Out_6__12,regFileMap_page2Out_6__11,
                           regFileMap_page2Out_6__10,regFileMap_page2Out_6__9,
                           regFileMap_page2Out_6__8,regFileMap_page2Out_6__7,
                           regFileMap_page2Out_6__6,regFileMap_page2Out_6__5,
                           regFileMap_page2Out_6__4,regFileMap_page2Out_6__3,
                           regFileMap_page2Out_6__2,regFileMap_page2Out_6__1,
                           regFileMap_page2Out_6__0}), .outFilter ({filter_4__7,
                           filter_4__6,filter_4__5,filter_4__4,filter_4__3,
                           filter_4__2,filter_4__1,filter_4__0})) ;
    RegUnit_8_16_unfolded0 regFileMap_loop1_1_regRowMap_loop1_2_regUnitMap (.filterBus (
                           {filterBus[23],filterBus[22],filterBus[21],
                           filterBus[20],filterBus[19],filterBus[18],
                           filterBus[17],filterBus[16]}), .windowBus ({
                           windowBus[47],windowBus[46],windowBus[45],
                           windowBus[44],windowBus[43],windowBus[42],
                           windowBus[41],windowBus[40],windowBus[39],
                           windowBus[38],windowBus[37],windowBus[36],
                           windowBus[35],windowBus[34],windowBus[33],
                           windowBus[32]}), .regPage1NextUnit ({
                           regFileMap_page1Out_12__15,regFileMap_page1Out_12__14
                           ,regFileMap_page1Out_12__13,
                           regFileMap_page1Out_12__12,regFileMap_page1Out_12__11
                           ,regFileMap_page1Out_12__10,regFileMap_page1Out_12__9
                           ,regFileMap_page1Out_12__8,regFileMap_page1Out_12__7,
                           regFileMap_page1Out_12__6,regFileMap_page1Out_12__5,
                           regFileMap_page1Out_12__4,regFileMap_page1Out_12__3,
                           regFileMap_page1Out_12__2,regFileMap_page1Out_12__1,
                           regFileMap_page1Out_12__0}), .regPage2NextUnit ({
                           regFileMap_page2Out_12__15,regFileMap_page2Out_12__14
                           ,regFileMap_page2Out_12__13,
                           regFileMap_page2Out_12__12,regFileMap_page2Out_12__11
                           ,regFileMap_page2Out_12__10,regFileMap_page2Out_12__9
                           ,regFileMap_page2Out_12__8,regFileMap_page2Out_12__7,
                           regFileMap_page2Out_12__6,regFileMap_page2Out_12__5,
                           regFileMap_page2Out_12__4,regFileMap_page2Out_12__3,
                           regFileMap_page2Out_12__2,regFileMap_page2Out_12__1,
                           regFileMap_page2Out_12__0}), .clk (clk), .rst (rst), 
                           .enableRegPage1 (regFileMap_page1Enables_1), .enableRegPage2 (
                           regFileMap_page2Enables_1), .enableRegFilter (nx5332)
                           , .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           currentPage_5__15,currentPage_5__14,currentPage_5__13
                           ,currentPage_5__12,currentPage_5__11,
                           currentPage_5__10,currentPage_5__9,currentPage_5__8,
                           currentPage_5__7,currentPage_5__6,currentPage_5__5,
                           currentPage_5__4,currentPage_5__3,currentPage_5__2,
                           currentPage_5__1,currentPage_5__0}), .outputRegPage1 (
                           {regFileMap_page1Out_7__15,regFileMap_page1Out_7__14,
                           regFileMap_page1Out_7__13,regFileMap_page1Out_7__12,
                           regFileMap_page1Out_7__11,regFileMap_page1Out_7__10,
                           regFileMap_page1Out_7__9,regFileMap_page1Out_7__8,
                           regFileMap_page1Out_7__7,regFileMap_page1Out_7__6,
                           regFileMap_page1Out_7__5,regFileMap_page1Out_7__4,
                           regFileMap_page1Out_7__3,regFileMap_page1Out_7__2,
                           regFileMap_page1Out_7__1,regFileMap_page1Out_7__0}), 
                           .outputRegPage2 ({regFileMap_page2Out_7__15,
                           regFileMap_page2Out_7__14,regFileMap_page2Out_7__13,
                           regFileMap_page2Out_7__12,regFileMap_page2Out_7__11,
                           regFileMap_page2Out_7__10,regFileMap_page2Out_7__9,
                           regFileMap_page2Out_7__8,regFileMap_page2Out_7__7,
                           regFileMap_page2Out_7__6,regFileMap_page2Out_7__5,
                           regFileMap_page2Out_7__4,regFileMap_page2Out_7__3,
                           regFileMap_page2Out_7__2,regFileMap_page2Out_7__1,
                           regFileMap_page2Out_7__0}), .outFilter ({filter_5__7,
                           filter_5__6,filter_5__5,filter_5__4,filter_5__3,
                           filter_5__2,filter_5__1,filter_5__0})) ;
    RegUnit_8_16_unfolded0 regFileMap_loop1_1_regRowMap_loop1_3_regUnitMap (.filterBus (
                           {filterBus[31],filterBus[30],filterBus[29],
                           filterBus[28],filterBus[27],filterBus[26],
                           filterBus[25],filterBus[24]}), .windowBus ({
                           windowBus[63],windowBus[62],windowBus[61],
                           windowBus[60],windowBus[59],windowBus[58],
                           windowBus[57],windowBus[56],windowBus[55],
                           windowBus[54],windowBus[53],windowBus[52],
                           windowBus[51],windowBus[50],windowBus[49],
                           windowBus[48]}), .regPage1NextUnit ({
                           regFileMap_page1Out_13__15,regFileMap_page1Out_13__14
                           ,regFileMap_page1Out_13__13,
                           regFileMap_page1Out_13__12,regFileMap_page1Out_13__11
                           ,regFileMap_page1Out_13__10,regFileMap_page1Out_13__9
                           ,regFileMap_page1Out_13__8,regFileMap_page1Out_13__7,
                           regFileMap_page1Out_13__6,regFileMap_page1Out_13__5,
                           regFileMap_page1Out_13__4,regFileMap_page1Out_13__3,
                           regFileMap_page1Out_13__2,regFileMap_page1Out_13__1,
                           regFileMap_page1Out_13__0}), .regPage2NextUnit ({
                           regFileMap_page2Out_13__15,regFileMap_page2Out_13__14
                           ,regFileMap_page2Out_13__13,
                           regFileMap_page2Out_13__12,regFileMap_page2Out_13__11
                           ,regFileMap_page2Out_13__10,regFileMap_page2Out_13__9
                           ,regFileMap_page2Out_13__8,regFileMap_page2Out_13__7,
                           regFileMap_page2Out_13__6,regFileMap_page2Out_13__5,
                           regFileMap_page2Out_13__4,regFileMap_page2Out_13__3,
                           regFileMap_page2Out_13__2,regFileMap_page2Out_13__1,
                           regFileMap_page2Out_13__0}), .clk (clk), .rst (rst), 
                           .enableRegPage1 (regFileMap_page1Enables_1), .enableRegPage2 (
                           regFileMap_page2Enables_1), .enableRegFilter (nx5334)
                           , .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           currentPage_17__15,currentPage_17__14,
                           currentPage_17__13,currentPage_17__12,
                           currentPage_17__11,currentPage_17__10,
                           currentPage_17__9,currentPage_17__8,currentPage_17__7
                           ,currentPage_17__6,currentPage_17__5,
                           currentPage_17__4,currentPage_17__3,currentPage_17__2
                           ,currentPage_17__1,currentPage_17__0}), .outputRegPage1 (
                           {regFileMap_page1Out_8__15,regFileMap_page1Out_8__14,
                           regFileMap_page1Out_8__13,regFileMap_page1Out_8__12,
                           regFileMap_page1Out_8__11,regFileMap_page1Out_8__10,
                           regFileMap_page1Out_8__9,regFileMap_page1Out_8__8,
                           regFileMap_page1Out_8__7,regFileMap_page1Out_8__6,
                           regFileMap_page1Out_8__5,regFileMap_page1Out_8__4,
                           regFileMap_page1Out_8__3,regFileMap_page1Out_8__2,
                           regFileMap_page1Out_8__1,regFileMap_page1Out_8__0}), 
                           .outputRegPage2 ({regFileMap_page2Out_8__15,
                           regFileMap_page2Out_8__14,regFileMap_page2Out_8__13,
                           regFileMap_page2Out_8__12,regFileMap_page2Out_8__11,
                           regFileMap_page2Out_8__10,regFileMap_page2Out_8__9,
                           regFileMap_page2Out_8__8,regFileMap_page2Out_8__7,
                           regFileMap_page2Out_8__6,regFileMap_page2Out_8__5,
                           regFileMap_page2Out_8__4,regFileMap_page2Out_8__3,
                           regFileMap_page2Out_8__2,regFileMap_page2Out_8__1,
                           regFileMap_page2Out_8__0}), .outFilter ({filter_17__7
                           ,filter_17__6,filter_17__5,filter_17__4,filter_17__3,
                           filter_17__2,filter_17__1,filter_17__0})) ;
    RegUnit_8_16_unfolded0 regFileMap_loop1_1_regRowMap_loop1_4_regUnitMap (.filterBus (
                           {filterBus[39],filterBus[38],filterBus[37],
                           filterBus[36],filterBus[35],filterBus[34],
                           filterBus[33],filterBus[32]}), .windowBus ({
                           windowBus[79],windowBus[78],windowBus[77],
                           windowBus[76],windowBus[75],windowBus[74],
                           windowBus[73],windowBus[72],windowBus[71],
                           windowBus[70],windowBus[69],windowBus[68],
                           windowBus[67],windowBus[66],windowBus[65],
                           windowBus[64]}), .regPage1NextUnit ({
                           regFileMap_page1Out_14__15,regFileMap_page1Out_14__14
                           ,regFileMap_page1Out_14__13,
                           regFileMap_page1Out_14__12,regFileMap_page1Out_14__11
                           ,regFileMap_page1Out_14__10,regFileMap_page1Out_14__9
                           ,regFileMap_page1Out_14__8,regFileMap_page1Out_14__7,
                           regFileMap_page1Out_14__6,regFileMap_page1Out_14__5,
                           regFileMap_page1Out_14__4,regFileMap_page1Out_14__3,
                           regFileMap_page1Out_14__2,regFileMap_page1Out_14__1,
                           regFileMap_page1Out_14__0}), .regPage2NextUnit ({
                           regFileMap_page2Out_14__15,regFileMap_page2Out_14__14
                           ,regFileMap_page2Out_14__13,
                           regFileMap_page2Out_14__12,regFileMap_page2Out_14__11
                           ,regFileMap_page2Out_14__10,regFileMap_page2Out_14__9
                           ,regFileMap_page2Out_14__8,regFileMap_page2Out_14__7,
                           regFileMap_page2Out_14__6,regFileMap_page2Out_14__5,
                           regFileMap_page2Out_14__4,regFileMap_page2Out_14__3,
                           regFileMap_page2Out_14__2,regFileMap_page2Out_14__1,
                           regFileMap_page2Out_14__0}), .clk (clk), .rst (rst), 
                           .enableRegPage1 (regFileMap_page1Enables_1), .enableRegPage2 (
                           regFileMap_page2Enables_1), .enableRegFilter (nx5334)
                           , .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           currentPage_18__15,currentPage_18__14,
                           currentPage_18__13,currentPage_18__12,
                           currentPage_18__11,currentPage_18__10,
                           currentPage_18__9,currentPage_18__8,currentPage_18__7
                           ,currentPage_18__6,currentPage_18__5,
                           currentPage_18__4,currentPage_18__3,currentPage_18__2
                           ,currentPage_18__1,currentPage_18__0}), .outputRegPage1 (
                           {regFileMap_page1Out_9__15,regFileMap_page1Out_9__14,
                           regFileMap_page1Out_9__13,regFileMap_page1Out_9__12,
                           regFileMap_page1Out_9__11,regFileMap_page1Out_9__10,
                           regFileMap_page1Out_9__9,regFileMap_page1Out_9__8,
                           regFileMap_page1Out_9__7,regFileMap_page1Out_9__6,
                           regFileMap_page1Out_9__5,regFileMap_page1Out_9__4,
                           regFileMap_page1Out_9__3,regFileMap_page1Out_9__2,
                           regFileMap_page1Out_9__1,regFileMap_page1Out_9__0}), 
                           .outputRegPage2 ({regFileMap_page2Out_9__15,
                           regFileMap_page2Out_9__14,regFileMap_page2Out_9__13,
                           regFileMap_page2Out_9__12,regFileMap_page2Out_9__11,
                           regFileMap_page2Out_9__10,regFileMap_page2Out_9__9,
                           regFileMap_page2Out_9__8,regFileMap_page2Out_9__7,
                           regFileMap_page2Out_9__6,regFileMap_page2Out_9__5,
                           regFileMap_page2Out_9__4,regFileMap_page2Out_9__3,
                           regFileMap_page2Out_9__2,regFileMap_page2Out_9__1,
                           regFileMap_page2Out_9__0}), .outFilter ({filter_18__7
                           ,filter_18__6,filter_18__5,filter_18__4,filter_18__3,
                           filter_18__2,filter_18__1,filter_18__0})) ;
    RegUnit_8_16_unfolded0 regFileMap_loop1_2_regRowMap_loop1_0_regUnitMap (.filterBus (
                           {filterBus[7],filterBus[6],filterBus[5],filterBus[4],
                           filterBus[3],filterBus[2],filterBus[1],filterBus[0]})
                           , .windowBus ({windowBus[15],windowBus[14],
                           windowBus[13],windowBus[12],windowBus[11],
                           windowBus[10],windowBus[9],windowBus[8],windowBus[7],
                           windowBus[6],windowBus[5],windowBus[4],windowBus[3],
                           windowBus[2],windowBus[1],windowBus[0]}), .regPage1NextUnit (
                           {regFileMap_page1Out_15__15,
                           regFileMap_page1Out_15__14,regFileMap_page1Out_15__13
                           ,regFileMap_page1Out_15__12,
                           regFileMap_page1Out_15__11,regFileMap_page1Out_15__10
                           ,regFileMap_page1Out_15__9,regFileMap_page1Out_15__8,
                           regFileMap_page1Out_15__7,regFileMap_page1Out_15__6,
                           regFileMap_page1Out_15__5,regFileMap_page1Out_15__4,
                           regFileMap_page1Out_15__3,regFileMap_page1Out_15__2,
                           regFileMap_page1Out_15__1,regFileMap_page1Out_15__0})
                           , .regPage2NextUnit ({regFileMap_page2Out_15__15,
                           regFileMap_page2Out_15__14,regFileMap_page2Out_15__13
                           ,regFileMap_page2Out_15__12,
                           regFileMap_page2Out_15__11,regFileMap_page2Out_15__10
                           ,regFileMap_page2Out_15__9,regFileMap_page2Out_15__8,
                           regFileMap_page2Out_15__7,regFileMap_page2Out_15__6,
                           regFileMap_page2Out_15__5,regFileMap_page2Out_15__4,
                           regFileMap_page2Out_15__3,regFileMap_page2Out_15__2,
                           regFileMap_page2Out_15__1,regFileMap_page2Out_15__0})
                           , .clk (clk), .rst (rst), .enableRegPage1 (
                           regFileMap_page1Enables_2), .enableRegPage2 (
                           regFileMap_page2Enables_2), .enableRegFilter (nx5336)
                           , .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           currentPage_6__15,currentPage_6__14,currentPage_6__13
                           ,currentPage_6__12,currentPage_6__11,
                           currentPage_6__10,currentPage_6__9,currentPage_6__8,
                           currentPage_6__7,currentPage_6__6,currentPage_6__5,
                           currentPage_6__4,currentPage_6__3,currentPage_6__2,
                           currentPage_6__1,currentPage_6__0}), .outputRegPage1 (
                           {regFileMap_page1Out_10__15,
                           regFileMap_page1Out_10__14,regFileMap_page1Out_10__13
                           ,regFileMap_page1Out_10__12,
                           regFileMap_page1Out_10__11,regFileMap_page1Out_10__10
                           ,regFileMap_page1Out_10__9,regFileMap_page1Out_10__8,
                           regFileMap_page1Out_10__7,regFileMap_page1Out_10__6,
                           regFileMap_page1Out_10__5,regFileMap_page1Out_10__4,
                           regFileMap_page1Out_10__3,regFileMap_page1Out_10__2,
                           regFileMap_page1Out_10__1,regFileMap_page1Out_10__0})
                           , .outputRegPage2 ({regFileMap_page2Out_10__15,
                           regFileMap_page2Out_10__14,regFileMap_page2Out_10__13
                           ,regFileMap_page2Out_10__12,
                           regFileMap_page2Out_10__11,regFileMap_page2Out_10__10
                           ,regFileMap_page2Out_10__9,regFileMap_page2Out_10__8,
                           regFileMap_page2Out_10__7,regFileMap_page2Out_10__6,
                           regFileMap_page2Out_10__5,regFileMap_page2Out_10__4,
                           regFileMap_page2Out_10__3,regFileMap_page2Out_10__2,
                           regFileMap_page2Out_10__1,regFileMap_page2Out_10__0})
                           , .outFilter ({filter_6__7,filter_6__6,filter_6__5,
                           filter_6__4,filter_6__3,filter_6__2,filter_6__1,
                           filter_6__0})) ;
    RegUnit_8_16_unfolded0 regFileMap_loop1_2_regRowMap_loop1_1_regUnitMap (.filterBus (
                           {filterBus[15],filterBus[14],filterBus[13],
                           filterBus[12],filterBus[11],filterBus[10],
                           filterBus[9],filterBus[8]}), .windowBus ({
                           windowBus[31],windowBus[30],windowBus[29],
                           windowBus[28],windowBus[27],windowBus[26],
                           windowBus[25],windowBus[24],windowBus[23],
                           windowBus[22],windowBus[21],windowBus[20],
                           windowBus[19],windowBus[18],windowBus[17],
                           windowBus[16]}), .regPage1NextUnit ({
                           regFileMap_page1Out_16__15,regFileMap_page1Out_16__14
                           ,regFileMap_page1Out_16__13,
                           regFileMap_page1Out_16__12,regFileMap_page1Out_16__11
                           ,regFileMap_page1Out_16__10,regFileMap_page1Out_16__9
                           ,regFileMap_page1Out_16__8,regFileMap_page1Out_16__7,
                           regFileMap_page1Out_16__6,regFileMap_page1Out_16__5,
                           regFileMap_page1Out_16__4,regFileMap_page1Out_16__3,
                           regFileMap_page1Out_16__2,regFileMap_page1Out_16__1,
                           regFileMap_page1Out_16__0}), .regPage2NextUnit ({
                           regFileMap_page2Out_16__15,regFileMap_page2Out_16__14
                           ,regFileMap_page2Out_16__13,
                           regFileMap_page2Out_16__12,regFileMap_page2Out_16__11
                           ,regFileMap_page2Out_16__10,regFileMap_page2Out_16__9
                           ,regFileMap_page2Out_16__8,regFileMap_page2Out_16__7,
                           regFileMap_page2Out_16__6,regFileMap_page2Out_16__5,
                           regFileMap_page2Out_16__4,regFileMap_page2Out_16__3,
                           regFileMap_page2Out_16__2,regFileMap_page2Out_16__1,
                           regFileMap_page2Out_16__0}), .clk (clk), .rst (rst), 
                           .enableRegPage1 (regFileMap_page1Enables_2), .enableRegPage2 (
                           regFileMap_page2Enables_2), .enableRegFilter (nx5336)
                           , .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           currentPage_7__15,currentPage_7__14,currentPage_7__13
                           ,currentPage_7__12,currentPage_7__11,
                           currentPage_7__10,currentPage_7__9,currentPage_7__8,
                           currentPage_7__7,currentPage_7__6,currentPage_7__5,
                           currentPage_7__4,currentPage_7__3,currentPage_7__2,
                           currentPage_7__1,currentPage_7__0}), .outputRegPage1 (
                           {regFileMap_page1Out_11__15,
                           regFileMap_page1Out_11__14,regFileMap_page1Out_11__13
                           ,regFileMap_page1Out_11__12,
                           regFileMap_page1Out_11__11,regFileMap_page1Out_11__10
                           ,regFileMap_page1Out_11__9,regFileMap_page1Out_11__8,
                           regFileMap_page1Out_11__7,regFileMap_page1Out_11__6,
                           regFileMap_page1Out_11__5,regFileMap_page1Out_11__4,
                           regFileMap_page1Out_11__3,regFileMap_page1Out_11__2,
                           regFileMap_page1Out_11__1,regFileMap_page1Out_11__0})
                           , .outputRegPage2 ({regFileMap_page2Out_11__15,
                           regFileMap_page2Out_11__14,regFileMap_page2Out_11__13
                           ,regFileMap_page2Out_11__12,
                           regFileMap_page2Out_11__11,regFileMap_page2Out_11__10
                           ,regFileMap_page2Out_11__9,regFileMap_page2Out_11__8,
                           regFileMap_page2Out_11__7,regFileMap_page2Out_11__6,
                           regFileMap_page2Out_11__5,regFileMap_page2Out_11__4,
                           regFileMap_page2Out_11__3,regFileMap_page2Out_11__2,
                           regFileMap_page2Out_11__1,regFileMap_page2Out_11__0})
                           , .outFilter ({filter_7__7,filter_7__6,filter_7__5,
                           filter_7__4,filter_7__3,filter_7__2,filter_7__1,
                           filter_7__0})) ;
    RegUnit_8_16_unfolded0 regFileMap_loop1_2_regRowMap_loop1_2_regUnitMap (.filterBus (
                           {filterBus[23],filterBus[22],filterBus[21],
                           filterBus[20],filterBus[19],filterBus[18],
                           filterBus[17],filterBus[16]}), .windowBus ({
                           windowBus[47],windowBus[46],windowBus[45],
                           windowBus[44],windowBus[43],windowBus[42],
                           windowBus[41],windowBus[40],windowBus[39],
                           windowBus[38],windowBus[37],windowBus[36],
                           windowBus[35],windowBus[34],windowBus[33],
                           windowBus[32]}), .regPage1NextUnit ({
                           regFileMap_page1Out_17__15,regFileMap_page1Out_17__14
                           ,regFileMap_page1Out_17__13,
                           regFileMap_page1Out_17__12,regFileMap_page1Out_17__11
                           ,regFileMap_page1Out_17__10,regFileMap_page1Out_17__9
                           ,regFileMap_page1Out_17__8,regFileMap_page1Out_17__7,
                           regFileMap_page1Out_17__6,regFileMap_page1Out_17__5,
                           regFileMap_page1Out_17__4,regFileMap_page1Out_17__3,
                           regFileMap_page1Out_17__2,regFileMap_page1Out_17__1,
                           regFileMap_page1Out_17__0}), .regPage2NextUnit ({
                           regFileMap_page2Out_17__15,regFileMap_page2Out_17__14
                           ,regFileMap_page2Out_17__13,
                           regFileMap_page2Out_17__12,regFileMap_page2Out_17__11
                           ,regFileMap_page2Out_17__10,regFileMap_page2Out_17__9
                           ,regFileMap_page2Out_17__8,regFileMap_page2Out_17__7,
                           regFileMap_page2Out_17__6,regFileMap_page2Out_17__5,
                           regFileMap_page2Out_17__4,regFileMap_page2Out_17__3,
                           regFileMap_page2Out_17__2,regFileMap_page2Out_17__1,
                           regFileMap_page2Out_17__0}), .clk (clk), .rst (rst), 
                           .enableRegPage1 (regFileMap_page1Enables_2), .enableRegPage2 (
                           regFileMap_page2Enables_2), .enableRegFilter (nx5336)
                           , .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           currentPage_8__15,currentPage_8__14,currentPage_8__13
                           ,currentPage_8__12,currentPage_8__11,
                           currentPage_8__10,currentPage_8__9,currentPage_8__8,
                           currentPage_8__7,currentPage_8__6,currentPage_8__5,
                           currentPage_8__4,currentPage_8__3,currentPage_8__2,
                           currentPage_8__1,currentPage_8__0}), .outputRegPage1 (
                           {regFileMap_page1Out_12__15,
                           regFileMap_page1Out_12__14,regFileMap_page1Out_12__13
                           ,regFileMap_page1Out_12__12,
                           regFileMap_page1Out_12__11,regFileMap_page1Out_12__10
                           ,regFileMap_page1Out_12__9,regFileMap_page1Out_12__8,
                           regFileMap_page1Out_12__7,regFileMap_page1Out_12__6,
                           regFileMap_page1Out_12__5,regFileMap_page1Out_12__4,
                           regFileMap_page1Out_12__3,regFileMap_page1Out_12__2,
                           regFileMap_page1Out_12__1,regFileMap_page1Out_12__0})
                           , .outputRegPage2 ({regFileMap_page2Out_12__15,
                           regFileMap_page2Out_12__14,regFileMap_page2Out_12__13
                           ,regFileMap_page2Out_12__12,
                           regFileMap_page2Out_12__11,regFileMap_page2Out_12__10
                           ,regFileMap_page2Out_12__9,regFileMap_page2Out_12__8,
                           regFileMap_page2Out_12__7,regFileMap_page2Out_12__6,
                           regFileMap_page2Out_12__5,regFileMap_page2Out_12__4,
                           regFileMap_page2Out_12__3,regFileMap_page2Out_12__2,
                           regFileMap_page2Out_12__1,regFileMap_page2Out_12__0})
                           , .outFilter ({filter_8__7,filter_8__6,filter_8__5,
                           filter_8__4,filter_8__3,filter_8__2,filter_8__1,
                           filter_8__0})) ;
    RegUnit_8_16_unfolded0 regFileMap_loop1_2_regRowMap_loop1_3_regUnitMap (.filterBus (
                           {filterBus[31],filterBus[30],filterBus[29],
                           filterBus[28],filterBus[27],filterBus[26],
                           filterBus[25],filterBus[24]}), .windowBus ({
                           windowBus[63],windowBus[62],windowBus[61],
                           windowBus[60],windowBus[59],windowBus[58],
                           windowBus[57],windowBus[56],windowBus[55],
                           windowBus[54],windowBus[53],windowBus[52],
                           windowBus[51],windowBus[50],windowBus[49],
                           windowBus[48]}), .regPage1NextUnit ({
                           regFileMap_page1Out_18__15,regFileMap_page1Out_18__14
                           ,regFileMap_page1Out_18__13,
                           regFileMap_page1Out_18__12,regFileMap_page1Out_18__11
                           ,regFileMap_page1Out_18__10,regFileMap_page1Out_18__9
                           ,regFileMap_page1Out_18__8,regFileMap_page1Out_18__7,
                           regFileMap_page1Out_18__6,regFileMap_page1Out_18__5,
                           regFileMap_page1Out_18__4,regFileMap_page1Out_18__3,
                           regFileMap_page1Out_18__2,regFileMap_page1Out_18__1,
                           regFileMap_page1Out_18__0}), .regPage2NextUnit ({
                           regFileMap_page2Out_18__15,regFileMap_page2Out_18__14
                           ,regFileMap_page2Out_18__13,
                           regFileMap_page2Out_18__12,regFileMap_page2Out_18__11
                           ,regFileMap_page2Out_18__10,regFileMap_page2Out_18__9
                           ,regFileMap_page2Out_18__8,regFileMap_page2Out_18__7,
                           regFileMap_page2Out_18__6,regFileMap_page2Out_18__5,
                           regFileMap_page2Out_18__4,regFileMap_page2Out_18__3,
                           regFileMap_page2Out_18__2,regFileMap_page2Out_18__1,
                           regFileMap_page2Out_18__0}), .clk (clk), .rst (rst), 
                           .enableRegPage1 (regFileMap_page1Enables_2), .enableRegPage2 (
                           regFileMap_page2Enables_2), .enableRegFilter (nx5338)
                           , .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           currentPage_19__15,currentPage_19__14,
                           currentPage_19__13,currentPage_19__12,
                           currentPage_19__11,currentPage_19__10,
                           currentPage_19__9,currentPage_19__8,currentPage_19__7
                           ,currentPage_19__6,currentPage_19__5,
                           currentPage_19__4,currentPage_19__3,currentPage_19__2
                           ,currentPage_19__1,currentPage_19__0}), .outputRegPage1 (
                           {regFileMap_page1Out_13__15,
                           regFileMap_page1Out_13__14,regFileMap_page1Out_13__13
                           ,regFileMap_page1Out_13__12,
                           regFileMap_page1Out_13__11,regFileMap_page1Out_13__10
                           ,regFileMap_page1Out_13__9,regFileMap_page1Out_13__8,
                           regFileMap_page1Out_13__7,regFileMap_page1Out_13__6,
                           regFileMap_page1Out_13__5,regFileMap_page1Out_13__4,
                           regFileMap_page1Out_13__3,regFileMap_page1Out_13__2,
                           regFileMap_page1Out_13__1,regFileMap_page1Out_13__0})
                           , .outputRegPage2 ({regFileMap_page2Out_13__15,
                           regFileMap_page2Out_13__14,regFileMap_page2Out_13__13
                           ,regFileMap_page2Out_13__12,
                           regFileMap_page2Out_13__11,regFileMap_page2Out_13__10
                           ,regFileMap_page2Out_13__9,regFileMap_page2Out_13__8,
                           regFileMap_page2Out_13__7,regFileMap_page2Out_13__6,
                           regFileMap_page2Out_13__5,regFileMap_page2Out_13__4,
                           regFileMap_page2Out_13__3,regFileMap_page2Out_13__2,
                           regFileMap_page2Out_13__1,regFileMap_page2Out_13__0})
                           , .outFilter ({filter_19__7,filter_19__6,filter_19__5
                           ,filter_19__4,filter_19__3,filter_19__2,filter_19__1,
                           filter_19__0})) ;
    RegUnit_8_16_unfolded0 regFileMap_loop1_2_regRowMap_loop1_4_regUnitMap (.filterBus (
                           {filterBus[39],filterBus[38],filterBus[37],
                           filterBus[36],filterBus[35],filterBus[34],
                           filterBus[33],filterBus[32]}), .windowBus ({
                           windowBus[79],windowBus[78],windowBus[77],
                           windowBus[76],windowBus[75],windowBus[74],
                           windowBus[73],windowBus[72],windowBus[71],
                           windowBus[70],windowBus[69],windowBus[68],
                           windowBus[67],windowBus[66],windowBus[65],
                           windowBus[64]}), .regPage1NextUnit ({
                           regFileMap_page1Out_19__15,regFileMap_page1Out_19__14
                           ,regFileMap_page1Out_19__13,
                           regFileMap_page1Out_19__12,regFileMap_page1Out_19__11
                           ,regFileMap_page1Out_19__10,regFileMap_page1Out_19__9
                           ,regFileMap_page1Out_19__8,regFileMap_page1Out_19__7,
                           regFileMap_page1Out_19__6,regFileMap_page1Out_19__5,
                           regFileMap_page1Out_19__4,regFileMap_page1Out_19__3,
                           regFileMap_page1Out_19__2,regFileMap_page1Out_19__1,
                           regFileMap_page1Out_19__0}), .regPage2NextUnit ({
                           regFileMap_page2Out_19__15,regFileMap_page2Out_19__14
                           ,regFileMap_page2Out_19__13,
                           regFileMap_page2Out_19__12,regFileMap_page2Out_19__11
                           ,regFileMap_page2Out_19__10,regFileMap_page2Out_19__9
                           ,regFileMap_page2Out_19__8,regFileMap_page2Out_19__7,
                           regFileMap_page2Out_19__6,regFileMap_page2Out_19__5,
                           regFileMap_page2Out_19__4,regFileMap_page2Out_19__3,
                           regFileMap_page2Out_19__2,regFileMap_page2Out_19__1,
                           regFileMap_page2Out_19__0}), .clk (clk), .rst (rst), 
                           .enableRegPage1 (regFileMap_page1Enables_2), .enableRegPage2 (
                           regFileMap_page2Enables_2), .enableRegFilter (nx5338)
                           , .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           currentPage_20__15,currentPage_20__14,
                           currentPage_20__13,currentPage_20__12,
                           currentPage_20__11,currentPage_20__10,
                           currentPage_20__9,currentPage_20__8,currentPage_20__7
                           ,currentPage_20__6,currentPage_20__5,
                           currentPage_20__4,currentPage_20__3,currentPage_20__2
                           ,currentPage_20__1,currentPage_20__0}), .outputRegPage1 (
                           {regFileMap_page1Out_14__15,
                           regFileMap_page1Out_14__14,regFileMap_page1Out_14__13
                           ,regFileMap_page1Out_14__12,
                           regFileMap_page1Out_14__11,regFileMap_page1Out_14__10
                           ,regFileMap_page1Out_14__9,regFileMap_page1Out_14__8,
                           regFileMap_page1Out_14__7,regFileMap_page1Out_14__6,
                           regFileMap_page1Out_14__5,regFileMap_page1Out_14__4,
                           regFileMap_page1Out_14__3,regFileMap_page1Out_14__2,
                           regFileMap_page1Out_14__1,regFileMap_page1Out_14__0})
                           , .outputRegPage2 ({regFileMap_page2Out_14__15,
                           regFileMap_page2Out_14__14,regFileMap_page2Out_14__13
                           ,regFileMap_page2Out_14__12,
                           regFileMap_page2Out_14__11,regFileMap_page2Out_14__10
                           ,regFileMap_page2Out_14__9,regFileMap_page2Out_14__8,
                           regFileMap_page2Out_14__7,regFileMap_page2Out_14__6,
                           regFileMap_page2Out_14__5,regFileMap_page2Out_14__4,
                           regFileMap_page2Out_14__3,regFileMap_page2Out_14__2,
                           regFileMap_page2Out_14__1,regFileMap_page2Out_14__0})
                           , .outFilter ({filter_20__7,filter_20__6,filter_20__5
                           ,filter_20__4,filter_20__3,filter_20__2,filter_20__1,
                           filter_20__0})) ;
    RegUnit_8_16_unfolded0 regFileMap_loop1_3_regRowMap_loop1_0_regUnitMap (.filterBus (
                           {filterBus[7],filterBus[6],filterBus[5],filterBus[4],
                           filterBus[3],filterBus[2],filterBus[1],filterBus[0]})
                           , .windowBus ({windowBus[15],windowBus[14],
                           windowBus[13],windowBus[12],windowBus[11],
                           windowBus[10],windowBus[9],windowBus[8],windowBus[7],
                           windowBus[6],windowBus[5],windowBus[4],windowBus[3],
                           windowBus[2],windowBus[1],windowBus[0]}), .regPage1NextUnit (
                           {regFileMap_page1Out_20__15,
                           regFileMap_page1Out_20__14,regFileMap_page1Out_20__13
                           ,regFileMap_page1Out_20__12,
                           regFileMap_page1Out_20__11,regFileMap_page1Out_20__10
                           ,regFileMap_page1Out_20__9,regFileMap_page1Out_20__8,
                           regFileMap_page1Out_20__7,regFileMap_page1Out_20__6,
                           regFileMap_page1Out_20__5,regFileMap_page1Out_20__4,
                           regFileMap_page1Out_20__3,regFileMap_page1Out_20__2,
                           regFileMap_page1Out_20__1,regFileMap_page1Out_20__0})
                           , .regPage2NextUnit ({regFileMap_page2Out_20__15,
                           regFileMap_page2Out_20__14,regFileMap_page2Out_20__13
                           ,regFileMap_page2Out_20__12,
                           regFileMap_page2Out_20__11,regFileMap_page2Out_20__10
                           ,regFileMap_page2Out_20__9,regFileMap_page2Out_20__8,
                           regFileMap_page2Out_20__7,regFileMap_page2Out_20__6,
                           regFileMap_page2Out_20__5,regFileMap_page2Out_20__4,
                           regFileMap_page2Out_20__3,regFileMap_page2Out_20__2,
                           regFileMap_page2Out_20__1,regFileMap_page2Out_20__0})
                           , .clk (clk), .rst (rst), .enableRegPage1 (
                           regFileMap_page1Enables_3), .enableRegPage2 (
                           regFileMap_page2Enables_3), .enableRegFilter (nx5340)
                           , .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           currentPage_9__15,currentPage_9__14,currentPage_9__13
                           ,currentPage_9__12,currentPage_9__11,
                           currentPage_9__10,currentPage_9__9,currentPage_9__8,
                           currentPage_9__7,currentPage_9__6,currentPage_9__5,
                           currentPage_9__4,currentPage_9__3,currentPage_9__2,
                           currentPage_9__1,currentPage_9__0}), .outputRegPage1 (
                           {regFileMap_page1Out_15__15,
                           regFileMap_page1Out_15__14,regFileMap_page1Out_15__13
                           ,regFileMap_page1Out_15__12,
                           regFileMap_page1Out_15__11,regFileMap_page1Out_15__10
                           ,regFileMap_page1Out_15__9,regFileMap_page1Out_15__8,
                           regFileMap_page1Out_15__7,regFileMap_page1Out_15__6,
                           regFileMap_page1Out_15__5,regFileMap_page1Out_15__4,
                           regFileMap_page1Out_15__3,regFileMap_page1Out_15__2,
                           regFileMap_page1Out_15__1,regFileMap_page1Out_15__0})
                           , .outputRegPage2 ({regFileMap_page2Out_15__15,
                           regFileMap_page2Out_15__14,regFileMap_page2Out_15__13
                           ,regFileMap_page2Out_15__12,
                           regFileMap_page2Out_15__11,regFileMap_page2Out_15__10
                           ,regFileMap_page2Out_15__9,regFileMap_page2Out_15__8,
                           regFileMap_page2Out_15__7,regFileMap_page2Out_15__6,
                           regFileMap_page2Out_15__5,regFileMap_page2Out_15__4,
                           regFileMap_page2Out_15__3,regFileMap_page2Out_15__2,
                           regFileMap_page2Out_15__1,regFileMap_page2Out_15__0})
                           , .outFilter ({filter_9__7,filter_9__6,filter_9__5,
                           filter_9__4,filter_9__3,filter_9__2,filter_9__1,
                           filter_9__0})) ;
    RegUnit_8_16_unfolded0 regFileMap_loop1_3_regRowMap_loop1_1_regUnitMap (.filterBus (
                           {filterBus[15],filterBus[14],filterBus[13],
                           filterBus[12],filterBus[11],filterBus[10],
                           filterBus[9],filterBus[8]}), .windowBus ({
                           windowBus[31],windowBus[30],windowBus[29],
                           windowBus[28],windowBus[27],windowBus[26],
                           windowBus[25],windowBus[24],windowBus[23],
                           windowBus[22],windowBus[21],windowBus[20],
                           windowBus[19],windowBus[18],windowBus[17],
                           windowBus[16]}), .regPage1NextUnit ({
                           regFileMap_page1Out_21__15,regFileMap_page1Out_21__14
                           ,regFileMap_page1Out_21__13,
                           regFileMap_page1Out_21__12,regFileMap_page1Out_21__11
                           ,regFileMap_page1Out_21__10,regFileMap_page1Out_21__9
                           ,regFileMap_page1Out_21__8,regFileMap_page1Out_21__7,
                           regFileMap_page1Out_21__6,regFileMap_page1Out_21__5,
                           regFileMap_page1Out_21__4,regFileMap_page1Out_21__3,
                           regFileMap_page1Out_21__2,regFileMap_page1Out_21__1,
                           regFileMap_page1Out_21__0}), .regPage2NextUnit ({
                           regFileMap_page2Out_21__15,regFileMap_page2Out_21__14
                           ,regFileMap_page2Out_21__13,
                           regFileMap_page2Out_21__12,regFileMap_page2Out_21__11
                           ,regFileMap_page2Out_21__10,regFileMap_page2Out_21__9
                           ,regFileMap_page2Out_21__8,regFileMap_page2Out_21__7,
                           regFileMap_page2Out_21__6,regFileMap_page2Out_21__5,
                           regFileMap_page2Out_21__4,regFileMap_page2Out_21__3,
                           regFileMap_page2Out_21__2,regFileMap_page2Out_21__1,
                           regFileMap_page2Out_21__0}), .clk (clk), .rst (rst), 
                           .enableRegPage1 (regFileMap_page1Enables_3), .enableRegPage2 (
                           regFileMap_page2Enables_3), .enableRegFilter (nx5340)
                           , .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           currentPage_10__15,currentPage_10__14,
                           currentPage_10__13,currentPage_10__12,
                           currentPage_10__11,currentPage_10__10,
                           currentPage_10__9,currentPage_10__8,currentPage_10__7
                           ,currentPage_10__6,currentPage_10__5,
                           currentPage_10__4,currentPage_10__3,currentPage_10__2
                           ,currentPage_10__1,currentPage_10__0}), .outputRegPage1 (
                           {regFileMap_page1Out_16__15,
                           regFileMap_page1Out_16__14,regFileMap_page1Out_16__13
                           ,regFileMap_page1Out_16__12,
                           regFileMap_page1Out_16__11,regFileMap_page1Out_16__10
                           ,regFileMap_page1Out_16__9,regFileMap_page1Out_16__8,
                           regFileMap_page1Out_16__7,regFileMap_page1Out_16__6,
                           regFileMap_page1Out_16__5,regFileMap_page1Out_16__4,
                           regFileMap_page1Out_16__3,regFileMap_page1Out_16__2,
                           regFileMap_page1Out_16__1,regFileMap_page1Out_16__0})
                           , .outputRegPage2 ({regFileMap_page2Out_16__15,
                           regFileMap_page2Out_16__14,regFileMap_page2Out_16__13
                           ,regFileMap_page2Out_16__12,
                           regFileMap_page2Out_16__11,regFileMap_page2Out_16__10
                           ,regFileMap_page2Out_16__9,regFileMap_page2Out_16__8,
                           regFileMap_page2Out_16__7,regFileMap_page2Out_16__6,
                           regFileMap_page2Out_16__5,regFileMap_page2Out_16__4,
                           regFileMap_page2Out_16__3,regFileMap_page2Out_16__2,
                           regFileMap_page2Out_16__1,regFileMap_page2Out_16__0})
                           , .outFilter ({filter_10__7,filter_10__6,filter_10__5
                           ,filter_10__4,filter_10__3,filter_10__2,filter_10__1,
                           filter_10__0})) ;
    RegUnit_8_16_unfolded0 regFileMap_loop1_3_regRowMap_loop1_2_regUnitMap (.filterBus (
                           {filterBus[23],filterBus[22],filterBus[21],
                           filterBus[20],filterBus[19],filterBus[18],
                           filterBus[17],filterBus[16]}), .windowBus ({
                           windowBus[47],windowBus[46],windowBus[45],
                           windowBus[44],windowBus[43],windowBus[42],
                           windowBus[41],windowBus[40],windowBus[39],
                           windowBus[38],windowBus[37],windowBus[36],
                           windowBus[35],windowBus[34],windowBus[33],
                           windowBus[32]}), .regPage1NextUnit ({
                           regFileMap_page1Out_22__15,regFileMap_page1Out_22__14
                           ,regFileMap_page1Out_22__13,
                           regFileMap_page1Out_22__12,regFileMap_page1Out_22__11
                           ,regFileMap_page1Out_22__10,regFileMap_page1Out_22__9
                           ,regFileMap_page1Out_22__8,regFileMap_page1Out_22__7,
                           regFileMap_page1Out_22__6,regFileMap_page1Out_22__5,
                           regFileMap_page1Out_22__4,regFileMap_page1Out_22__3,
                           regFileMap_page1Out_22__2,regFileMap_page1Out_22__1,
                           regFileMap_page1Out_22__0}), .regPage2NextUnit ({
                           regFileMap_page2Out_22__15,regFileMap_page2Out_22__14
                           ,regFileMap_page2Out_22__13,
                           regFileMap_page2Out_22__12,regFileMap_page2Out_22__11
                           ,regFileMap_page2Out_22__10,regFileMap_page2Out_22__9
                           ,regFileMap_page2Out_22__8,regFileMap_page2Out_22__7,
                           regFileMap_page2Out_22__6,regFileMap_page2Out_22__5,
                           regFileMap_page2Out_22__4,regFileMap_page2Out_22__3,
                           regFileMap_page2Out_22__2,regFileMap_page2Out_22__1,
                           regFileMap_page2Out_22__0}), .clk (clk), .rst (rst), 
                           .enableRegPage1 (regFileMap_page1Enables_3), .enableRegPage2 (
                           regFileMap_page2Enables_3), .enableRegFilter (nx5340)
                           , .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           currentPage_11__15,currentPage_11__14,
                           currentPage_11__13,currentPage_11__12,
                           currentPage_11__11,currentPage_11__10,
                           currentPage_11__9,currentPage_11__8,currentPage_11__7
                           ,currentPage_11__6,currentPage_11__5,
                           currentPage_11__4,currentPage_11__3,currentPage_11__2
                           ,currentPage_11__1,currentPage_11__0}), .outputRegPage1 (
                           {regFileMap_page1Out_17__15,
                           regFileMap_page1Out_17__14,regFileMap_page1Out_17__13
                           ,regFileMap_page1Out_17__12,
                           regFileMap_page1Out_17__11,regFileMap_page1Out_17__10
                           ,regFileMap_page1Out_17__9,regFileMap_page1Out_17__8,
                           regFileMap_page1Out_17__7,regFileMap_page1Out_17__6,
                           regFileMap_page1Out_17__5,regFileMap_page1Out_17__4,
                           regFileMap_page1Out_17__3,regFileMap_page1Out_17__2,
                           regFileMap_page1Out_17__1,regFileMap_page1Out_17__0})
                           , .outputRegPage2 ({regFileMap_page2Out_17__15,
                           regFileMap_page2Out_17__14,regFileMap_page2Out_17__13
                           ,regFileMap_page2Out_17__12,
                           regFileMap_page2Out_17__11,regFileMap_page2Out_17__10
                           ,regFileMap_page2Out_17__9,regFileMap_page2Out_17__8,
                           regFileMap_page2Out_17__7,regFileMap_page2Out_17__6,
                           regFileMap_page2Out_17__5,regFileMap_page2Out_17__4,
                           regFileMap_page2Out_17__3,regFileMap_page2Out_17__2,
                           regFileMap_page2Out_17__1,regFileMap_page2Out_17__0})
                           , .outFilter ({filter_11__7,filter_11__6,filter_11__5
                           ,filter_11__4,filter_11__3,filter_11__2,filter_11__1,
                           filter_11__0})) ;
    RegUnit_8_16_unfolded0 regFileMap_loop1_3_regRowMap_loop1_3_regUnitMap (.filterBus (
                           {filterBus[31],filterBus[30],filterBus[29],
                           filterBus[28],filterBus[27],filterBus[26],
                           filterBus[25],filterBus[24]}), .windowBus ({
                           windowBus[63],windowBus[62],windowBus[61],
                           windowBus[60],windowBus[59],windowBus[58],
                           windowBus[57],windowBus[56],windowBus[55],
                           windowBus[54],windowBus[53],windowBus[52],
                           windowBus[51],windowBus[50],windowBus[49],
                           windowBus[48]}), .regPage1NextUnit ({
                           regFileMap_page1Out_23__15,regFileMap_page1Out_23__14
                           ,regFileMap_page1Out_23__13,
                           regFileMap_page1Out_23__12,regFileMap_page1Out_23__11
                           ,regFileMap_page1Out_23__10,regFileMap_page1Out_23__9
                           ,regFileMap_page1Out_23__8,regFileMap_page1Out_23__7,
                           regFileMap_page1Out_23__6,regFileMap_page1Out_23__5,
                           regFileMap_page1Out_23__4,regFileMap_page1Out_23__3,
                           regFileMap_page1Out_23__2,regFileMap_page1Out_23__1,
                           regFileMap_page1Out_23__0}), .regPage2NextUnit ({
                           regFileMap_page2Out_23__15,regFileMap_page2Out_23__14
                           ,regFileMap_page2Out_23__13,
                           regFileMap_page2Out_23__12,regFileMap_page2Out_23__11
                           ,regFileMap_page2Out_23__10,regFileMap_page2Out_23__9
                           ,regFileMap_page2Out_23__8,regFileMap_page2Out_23__7,
                           regFileMap_page2Out_23__6,regFileMap_page2Out_23__5,
                           regFileMap_page2Out_23__4,regFileMap_page2Out_23__3,
                           regFileMap_page2Out_23__2,regFileMap_page2Out_23__1,
                           regFileMap_page2Out_23__0}), .clk (clk), .rst (rst), 
                           .enableRegPage1 (regFileMap_page1Enables_3), .enableRegPage2 (
                           regFileMap_page2Enables_3), .enableRegFilter (nx5342)
                           , .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           currentPage_21__15,currentPage_21__14,
                           currentPage_21__13,currentPage_21__12,
                           currentPage_21__11,currentPage_21__10,
                           currentPage_21__9,currentPage_21__8,currentPage_21__7
                           ,currentPage_21__6,currentPage_21__5,
                           currentPage_21__4,currentPage_21__3,currentPage_21__2
                           ,currentPage_21__1,currentPage_21__0}), .outputRegPage1 (
                           {regFileMap_page1Out_18__15,
                           regFileMap_page1Out_18__14,regFileMap_page1Out_18__13
                           ,regFileMap_page1Out_18__12,
                           regFileMap_page1Out_18__11,regFileMap_page1Out_18__10
                           ,regFileMap_page1Out_18__9,regFileMap_page1Out_18__8,
                           regFileMap_page1Out_18__7,regFileMap_page1Out_18__6,
                           regFileMap_page1Out_18__5,regFileMap_page1Out_18__4,
                           regFileMap_page1Out_18__3,regFileMap_page1Out_18__2,
                           regFileMap_page1Out_18__1,regFileMap_page1Out_18__0})
                           , .outputRegPage2 ({regFileMap_page2Out_18__15,
                           regFileMap_page2Out_18__14,regFileMap_page2Out_18__13
                           ,regFileMap_page2Out_18__12,
                           regFileMap_page2Out_18__11,regFileMap_page2Out_18__10
                           ,regFileMap_page2Out_18__9,regFileMap_page2Out_18__8,
                           regFileMap_page2Out_18__7,regFileMap_page2Out_18__6,
                           regFileMap_page2Out_18__5,regFileMap_page2Out_18__4,
                           regFileMap_page2Out_18__3,regFileMap_page2Out_18__2,
                           regFileMap_page2Out_18__1,regFileMap_page2Out_18__0})
                           , .outFilter ({filter_21__7,filter_21__6,filter_21__5
                           ,filter_21__4,filter_21__3,filter_21__2,filter_21__1,
                           filter_21__0})) ;
    RegUnit_8_16_unfolded0 regFileMap_loop1_3_regRowMap_loop1_4_regUnitMap (.filterBus (
                           {filterBus[39],filterBus[38],filterBus[37],
                           filterBus[36],filterBus[35],filterBus[34],
                           filterBus[33],filterBus[32]}), .windowBus ({
                           windowBus[79],windowBus[78],windowBus[77],
                           windowBus[76],windowBus[75],windowBus[74],
                           windowBus[73],windowBus[72],windowBus[71],
                           windowBus[70],windowBus[69],windowBus[68],
                           windowBus[67],windowBus[66],windowBus[65],
                           windowBus[64]}), .regPage1NextUnit ({
                           regFileMap_page1Out_24__15,regFileMap_page1Out_24__14
                           ,regFileMap_page1Out_24__13,
                           regFileMap_page1Out_24__12,regFileMap_page1Out_24__11
                           ,regFileMap_page1Out_24__10,regFileMap_page1Out_24__9
                           ,regFileMap_page1Out_24__8,regFileMap_page1Out_24__7,
                           regFileMap_page1Out_24__6,regFileMap_page1Out_24__5,
                           regFileMap_page1Out_24__4,regFileMap_page1Out_24__3,
                           regFileMap_page1Out_24__2,regFileMap_page1Out_24__1,
                           regFileMap_page1Out_24__0}), .regPage2NextUnit ({
                           regFileMap_page2Out_24__15,regFileMap_page2Out_24__14
                           ,regFileMap_page2Out_24__13,
                           regFileMap_page2Out_24__12,regFileMap_page2Out_24__11
                           ,regFileMap_page2Out_24__10,regFileMap_page2Out_24__9
                           ,regFileMap_page2Out_24__8,regFileMap_page2Out_24__7,
                           regFileMap_page2Out_24__6,regFileMap_page2Out_24__5,
                           regFileMap_page2Out_24__4,regFileMap_page2Out_24__3,
                           regFileMap_page2Out_24__2,regFileMap_page2Out_24__1,
                           regFileMap_page2Out_24__0}), .clk (clk), .rst (rst), 
                           .enableRegPage1 (regFileMap_page1Enables_3), .enableRegPage2 (
                           regFileMap_page2Enables_3), .enableRegFilter (nx5342)
                           , .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           currentPage_22__15,currentPage_22__14,
                           currentPage_22__13,currentPage_22__12,
                           currentPage_22__11,currentPage_22__10,
                           currentPage_22__9,currentPage_22__8,currentPage_22__7
                           ,currentPage_22__6,currentPage_22__5,
                           currentPage_22__4,currentPage_22__3,currentPage_22__2
                           ,currentPage_22__1,currentPage_22__0}), .outputRegPage1 (
                           {regFileMap_page1Out_19__15,
                           regFileMap_page1Out_19__14,regFileMap_page1Out_19__13
                           ,regFileMap_page1Out_19__12,
                           regFileMap_page1Out_19__11,regFileMap_page1Out_19__10
                           ,regFileMap_page1Out_19__9,regFileMap_page1Out_19__8,
                           regFileMap_page1Out_19__7,regFileMap_page1Out_19__6,
                           regFileMap_page1Out_19__5,regFileMap_page1Out_19__4,
                           regFileMap_page1Out_19__3,regFileMap_page1Out_19__2,
                           regFileMap_page1Out_19__1,regFileMap_page1Out_19__0})
                           , .outputRegPage2 ({regFileMap_page2Out_19__15,
                           regFileMap_page2Out_19__14,regFileMap_page2Out_19__13
                           ,regFileMap_page2Out_19__12,
                           regFileMap_page2Out_19__11,regFileMap_page2Out_19__10
                           ,regFileMap_page2Out_19__9,regFileMap_page2Out_19__8,
                           regFileMap_page2Out_19__7,regFileMap_page2Out_19__6,
                           regFileMap_page2Out_19__5,regFileMap_page2Out_19__4,
                           regFileMap_page2Out_19__3,regFileMap_page2Out_19__2,
                           regFileMap_page2Out_19__1,regFileMap_page2Out_19__0})
                           , .outFilter ({filter_22__7,filter_22__6,filter_22__5
                           ,filter_22__4,filter_22__3,filter_22__2,filter_22__1,
                           filter_22__0})) ;
    RegUnit_8_16_unfolded1 regFileMap_loop1_4_regRowMap_loop1_0_regUnitMap (.filterBus (
                           {filterBus[7],filterBus[6],filterBus[5],filterBus[4],
                           filterBus[3],filterBus[2],filterBus[1],filterBus[0]})
                           , .windowBus ({windowBus[15],windowBus[14],
                           windowBus[13],windowBus[12],windowBus[11],
                           windowBus[10],windowBus[9],windowBus[8],windowBus[7],
                           windowBus[6],windowBus[5],windowBus[4],windowBus[3],
                           windowBus[2],windowBus[1],windowBus[0]}), .regPage1NextUnit (
                           {outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15}), .regPage2NextUnit ({outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15}), .clk (
                           clk), .rst (rst), .enableRegPage1 (
                           regFileMap_page1Enables_4), .enableRegPage2 (
                           regFileMap_page2Enables_4), .enableRegFilter (nx5344)
                           , .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           currentPage_12__15,currentPage_12__14,
                           currentPage_12__13,currentPage_12__12,
                           currentPage_12__11,currentPage_12__10,
                           currentPage_12__9,currentPage_12__8,currentPage_12__7
                           ,currentPage_12__6,currentPage_12__5,
                           currentPage_12__4,currentPage_12__3,currentPage_12__2
                           ,currentPage_12__1,currentPage_12__0}), .outputRegPage1 (
                           {regFileMap_page1Out_20__15,
                           regFileMap_page1Out_20__14,regFileMap_page1Out_20__13
                           ,regFileMap_page1Out_20__12,
                           regFileMap_page1Out_20__11,regFileMap_page1Out_20__10
                           ,regFileMap_page1Out_20__9,regFileMap_page1Out_20__8,
                           regFileMap_page1Out_20__7,regFileMap_page1Out_20__6,
                           regFileMap_page1Out_20__5,regFileMap_page1Out_20__4,
                           regFileMap_page1Out_20__3,regFileMap_page1Out_20__2,
                           regFileMap_page1Out_20__1,regFileMap_page1Out_20__0})
                           , .outputRegPage2 ({regFileMap_page2Out_20__15,
                           regFileMap_page2Out_20__14,regFileMap_page2Out_20__13
                           ,regFileMap_page2Out_20__12,
                           regFileMap_page2Out_20__11,regFileMap_page2Out_20__10
                           ,regFileMap_page2Out_20__9,regFileMap_page2Out_20__8,
                           regFileMap_page2Out_20__7,regFileMap_page2Out_20__6,
                           regFileMap_page2Out_20__5,regFileMap_page2Out_20__4,
                           regFileMap_page2Out_20__3,regFileMap_page2Out_20__2,
                           regFileMap_page2Out_20__1,regFileMap_page2Out_20__0})
                           , .outFilter ({filter_12__7,filter_12__6,filter_12__5
                           ,filter_12__4,filter_12__3,filter_12__2,filter_12__1,
                           filter_12__0})) ;
    RegUnit_8_16_unfolded1 regFileMap_loop1_4_regRowMap_loop1_1_regUnitMap (.filterBus (
                           {filterBus[15],filterBus[14],filterBus[13],
                           filterBus[12],filterBus[11],filterBus[10],
                           filterBus[9],filterBus[8]}), .windowBus ({
                           windowBus[31],windowBus[30],windowBus[29],
                           windowBus[28],windowBus[27],windowBus[26],
                           windowBus[25],windowBus[24],windowBus[23],
                           windowBus[22],windowBus[21],windowBus[20],
                           windowBus[19],windowBus[18],windowBus[17],
                           windowBus[16]}), .regPage1NextUnit ({outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15}), .regPage2NextUnit (
                           {outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15}), .clk (clk), .rst (rst), .enableRegPage1 (
                           regFileMap_page1Enables_4), .enableRegPage2 (
                           regFileMap_page2Enables_4), .enableRegFilter (nx5344)
                           , .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           currentPage_13__15,currentPage_13__14,
                           currentPage_13__13,currentPage_13__12,
                           currentPage_13__11,currentPage_13__10,
                           currentPage_13__9,currentPage_13__8,currentPage_13__7
                           ,currentPage_13__6,currentPage_13__5,
                           currentPage_13__4,currentPage_13__3,currentPage_13__2
                           ,currentPage_13__1,currentPage_13__0}), .outputRegPage1 (
                           {regFileMap_page1Out_21__15,
                           regFileMap_page1Out_21__14,regFileMap_page1Out_21__13
                           ,regFileMap_page1Out_21__12,
                           regFileMap_page1Out_21__11,regFileMap_page1Out_21__10
                           ,regFileMap_page1Out_21__9,regFileMap_page1Out_21__8,
                           regFileMap_page1Out_21__7,regFileMap_page1Out_21__6,
                           regFileMap_page1Out_21__5,regFileMap_page1Out_21__4,
                           regFileMap_page1Out_21__3,regFileMap_page1Out_21__2,
                           regFileMap_page1Out_21__1,regFileMap_page1Out_21__0})
                           , .outputRegPage2 ({regFileMap_page2Out_21__15,
                           regFileMap_page2Out_21__14,regFileMap_page2Out_21__13
                           ,regFileMap_page2Out_21__12,
                           regFileMap_page2Out_21__11,regFileMap_page2Out_21__10
                           ,regFileMap_page2Out_21__9,regFileMap_page2Out_21__8,
                           regFileMap_page2Out_21__7,regFileMap_page2Out_21__6,
                           regFileMap_page2Out_21__5,regFileMap_page2Out_21__4,
                           regFileMap_page2Out_21__3,regFileMap_page2Out_21__2,
                           regFileMap_page2Out_21__1,regFileMap_page2Out_21__0})
                           , .outFilter ({filter_13__7,filter_13__6,filter_13__5
                           ,filter_13__4,filter_13__3,filter_13__2,filter_13__1,
                           filter_13__0})) ;
    RegUnit_8_16_unfolded1 regFileMap_loop1_4_regRowMap_loop1_2_regUnitMap (.filterBus (
                           {filterBus[23],filterBus[22],filterBus[21],
                           filterBus[20],filterBus[19],filterBus[18],
                           filterBus[17],filterBus[16]}), .windowBus ({
                           windowBus[47],windowBus[46],windowBus[45],
                           windowBus[44],windowBus[43],windowBus[42],
                           windowBus[41],windowBus[40],windowBus[39],
                           windowBus[38],windowBus[37],windowBus[36],
                           windowBus[35],windowBus[34],windowBus[33],
                           windowBus[32]}), .regPage1NextUnit ({outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15}), .regPage2NextUnit (
                           {outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15}), .clk (clk), .rst (rst), .enableRegPage1 (
                           regFileMap_page1Enables_4), .enableRegPage2 (
                           regFileMap_page2Enables_4), .enableRegFilter (nx5344)
                           , .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           currentPage_14__15,currentPage_14__14,
                           currentPage_14__13,currentPage_14__12,
                           currentPage_14__11,currentPage_14__10,
                           currentPage_14__9,currentPage_14__8,currentPage_14__7
                           ,currentPage_14__6,currentPage_14__5,
                           currentPage_14__4,currentPage_14__3,currentPage_14__2
                           ,currentPage_14__1,currentPage_14__0}), .outputRegPage1 (
                           {regFileMap_page1Out_22__15,
                           regFileMap_page1Out_22__14,regFileMap_page1Out_22__13
                           ,regFileMap_page1Out_22__12,
                           regFileMap_page1Out_22__11,regFileMap_page1Out_22__10
                           ,regFileMap_page1Out_22__9,regFileMap_page1Out_22__8,
                           regFileMap_page1Out_22__7,regFileMap_page1Out_22__6,
                           regFileMap_page1Out_22__5,regFileMap_page1Out_22__4,
                           regFileMap_page1Out_22__3,regFileMap_page1Out_22__2,
                           regFileMap_page1Out_22__1,regFileMap_page1Out_22__0})
                           , .outputRegPage2 ({regFileMap_page2Out_22__15,
                           regFileMap_page2Out_22__14,regFileMap_page2Out_22__13
                           ,regFileMap_page2Out_22__12,
                           regFileMap_page2Out_22__11,regFileMap_page2Out_22__10
                           ,regFileMap_page2Out_22__9,regFileMap_page2Out_22__8,
                           regFileMap_page2Out_22__7,regFileMap_page2Out_22__6,
                           regFileMap_page2Out_22__5,regFileMap_page2Out_22__4,
                           regFileMap_page2Out_22__3,regFileMap_page2Out_22__2,
                           regFileMap_page2Out_22__1,regFileMap_page2Out_22__0})
                           , .outFilter ({filter_14__7,filter_14__6,filter_14__5
                           ,filter_14__4,filter_14__3,filter_14__2,filter_14__1,
                           filter_14__0})) ;
    RegUnit_8_16_unfolded1 regFileMap_loop1_4_regRowMap_loop1_3_regUnitMap (.filterBus (
                           {filterBus[31],filterBus[30],filterBus[29],
                           filterBus[28],filterBus[27],filterBus[26],
                           filterBus[25],filterBus[24]}), .windowBus ({
                           windowBus[63],windowBus[62],windowBus[61],
                           windowBus[60],windowBus[59],windowBus[58],
                           windowBus[57],windowBus[56],windowBus[55],
                           windowBus[54],windowBus[53],windowBus[52],
                           windowBus[51],windowBus[50],windowBus[49],
                           windowBus[48]}), .regPage1NextUnit ({outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15}), .regPage2NextUnit (
                           {outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15}), .clk (clk), .rst (rst), .enableRegPage1 (
                           regFileMap_page1Enables_4), .enableRegPage2 (
                           regFileMap_page2Enables_4), .enableRegFilter (nx5346)
                           , .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           currentPage_23__15,currentPage_23__14,
                           currentPage_23__13,currentPage_23__12,
                           currentPage_23__11,currentPage_23__10,
                           currentPage_23__9,currentPage_23__8,currentPage_23__7
                           ,currentPage_23__6,currentPage_23__5,
                           currentPage_23__4,currentPage_23__3,currentPage_23__2
                           ,currentPage_23__1,currentPage_23__0}), .outputRegPage1 (
                           {regFileMap_page1Out_23__15,
                           regFileMap_page1Out_23__14,regFileMap_page1Out_23__13
                           ,regFileMap_page1Out_23__12,
                           regFileMap_page1Out_23__11,regFileMap_page1Out_23__10
                           ,regFileMap_page1Out_23__9,regFileMap_page1Out_23__8,
                           regFileMap_page1Out_23__7,regFileMap_page1Out_23__6,
                           regFileMap_page1Out_23__5,regFileMap_page1Out_23__4,
                           regFileMap_page1Out_23__3,regFileMap_page1Out_23__2,
                           regFileMap_page1Out_23__1,regFileMap_page1Out_23__0})
                           , .outputRegPage2 ({regFileMap_page2Out_23__15,
                           regFileMap_page2Out_23__14,regFileMap_page2Out_23__13
                           ,regFileMap_page2Out_23__12,
                           regFileMap_page2Out_23__11,regFileMap_page2Out_23__10
                           ,regFileMap_page2Out_23__9,regFileMap_page2Out_23__8,
                           regFileMap_page2Out_23__7,regFileMap_page2Out_23__6,
                           regFileMap_page2Out_23__5,regFileMap_page2Out_23__4,
                           regFileMap_page2Out_23__3,regFileMap_page2Out_23__2,
                           regFileMap_page2Out_23__1,regFileMap_page2Out_23__0})
                           , .outFilter ({filter_23__7,filter_23__6,filter_23__5
                           ,filter_23__4,filter_23__3,filter_23__2,filter_23__1,
                           filter_23__0})) ;
    RegUnit_8_16_unfolded1 regFileMap_loop1_4_regRowMap_loop1_4_regUnitMap (.filterBus (
                           {filterBus[39],filterBus[38],filterBus[37],
                           filterBus[36],filterBus[35],filterBus[34],
                           filterBus[33],filterBus[32]}), .windowBus ({
                           windowBus[79],windowBus[78],windowBus[77],
                           windowBus[76],windowBus[75],windowBus[74],
                           windowBus[73],windowBus[72],windowBus[71],
                           windowBus[70],windowBus[69],windowBus[68],
                           windowBus[67],windowBus[66],windowBus[65],
                           windowBus[64]}), .regPage1NextUnit ({outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15}), .regPage2NextUnit (
                           {outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15,outShifter_15,outShifter_15,
                           outShifter_15}), .clk (clk), .rst (rst), .enableRegPage1 (
                           regFileMap_page1Enables_4), .enableRegPage2 (
                           regFileMap_page2Enables_4), .enableRegFilter (nx5346)
                           , .page1ReadBusOrPage2 (shift2To1), .page2ReadBusOrPage1 (
                           shift1To2), .pageTurn (pageTurn), .outRegPage ({
                           currentPage_24__15,currentPage_24__14,
                           currentPage_24__13,currentPage_24__12,
                           currentPage_24__11,currentPage_24__10,
                           currentPage_24__9,currentPage_24__8,currentPage_24__7
                           ,currentPage_24__6,currentPage_24__5,
                           currentPage_24__4,currentPage_24__3,currentPage_24__2
                           ,currentPage_24__1,currentPage_24__0}), .outputRegPage1 (
                           {regFileMap_page1Out_24__15,
                           regFileMap_page1Out_24__14,regFileMap_page1Out_24__13
                           ,regFileMap_page1Out_24__12,
                           regFileMap_page1Out_24__11,regFileMap_page1Out_24__10
                           ,regFileMap_page1Out_24__9,regFileMap_page1Out_24__8,
                           regFileMap_page1Out_24__7,regFileMap_page1Out_24__6,
                           regFileMap_page1Out_24__5,regFileMap_page1Out_24__4,
                           regFileMap_page1Out_24__3,regFileMap_page1Out_24__2,
                           regFileMap_page1Out_24__1,regFileMap_page1Out_24__0})
                           , .outputRegPage2 ({regFileMap_page2Out_24__15,
                           regFileMap_page2Out_24__14,regFileMap_page2Out_24__13
                           ,regFileMap_page2Out_24__12,
                           regFileMap_page2Out_24__11,regFileMap_page2Out_24__10
                           ,regFileMap_page2Out_24__9,regFileMap_page2Out_24__8,
                           regFileMap_page2Out_24__7,regFileMap_page2Out_24__6,
                           regFileMap_page2Out_24__5,regFileMap_page2Out_24__4,
                           regFileMap_page2Out_24__3,regFileMap_page2Out_24__2,
                           regFileMap_page2Out_24__1,regFileMap_page2Out_24__0})
                           , .outFilter ({filter_24__7,filter_24__6,filter_24__5
                           ,filter_24__4,filter_24__3,filter_24__2,filter_24__1,
                           filter_24__0})) ;
    NBitAdder_16 addersMap_sum3FilterMap (.a ({addersMap_sum1_15,
                 addersMap_sum1_14,addersMap_sum1_13,addersMap_sum1_12,
                 addersMap_sum1_11,addersMap_sum1_10,addersMap_sum1_9,
                 addersMap_sum1_8,addersMap_sum1_7,addersMap_sum1_6,
                 addersMap_sum1_5,addersMap_sum1_4,addersMap_sum1_3,
                 addersMap_sum1_2,addersMap_sum1_1,addersMap_sum1_0}), .b ({
                 addersInputs_8__15,addersInputs_8__14,addersInputs_8__13,
                 addersInputs_8__12,addersInputs_8__11,addersInputs_8__10,
                 addersInputs_8__9,addersInputs_8__8,addersInputs_8__7,
                 addersInputs_8__6,addersInputs_8__5,addersInputs_8__4,
                 addersInputs_8__3,addersInputs_8__2,addersInputs_8__1,
                 addersInputs_8__0}), .carryIn (outShifter_15), .sum ({
                 addersMap_sum3Filter_15,addersMap_sum3Filter_14,
                 addersMap_sum3Filter_13,addersMap_sum3Filter_12,
                 addersMap_sum3Filter_11,addersMap_sum3Filter_10,
                 addersMap_sum3Filter_9,addersMap_sum3Filter_8,
                 addersMap_sum3Filter_7,addersMap_sum3Filter_6,
                 addersMap_sum3Filter_5,addersMap_sum3Filter_4,
                 addersMap_sum3Filter_3,addersMap_sum3Filter_2,
                 addersMap_sum3Filter_1,addersMap_sum3Filter_0}), .carryOut (
                 \$dummy [161])) ;
    NBitAdder_16 addersMap_sumRestMap (.a ({addersMap_sum2_15,addersMap_sum2_14,
                 addersMap_sum2_13,addersMap_sum2_12,addersMap_sum2_11,
                 addersMap_sum2_10,addersMap_sum2_9,addersMap_sum2_8,
                 addersMap_sum2_7,addersMap_sum2_6,addersMap_sum2_5,
                 addersMap_sum2_4,addersMap_sum2_3,addersMap_sum2_2,
                 addersMap_sum2_1,addersMap_sum2_0}), .b ({addersMap_sum3_15,
                 addersMap_sum3_14,addersMap_sum3_13,addersMap_sum3_12,
                 addersMap_sum3_11,addersMap_sum3_10,addersMap_sum3_9,
                 addersMap_sum3_8,addersMap_sum3_7,addersMap_sum3_6,
                 addersMap_sum3_5,addersMap_sum3_4,addersMap_sum3_3,
                 addersMap_sum3_2,addersMap_sum3_1,addersMap_sum3_0}), .carryIn (
                 outShifter_15), .sum ({addersMap_sum4_15,addersMap_sum4_14,
                 addersMap_sum4_13,addersMap_sum4_12,addersMap_sum4_11,
                 addersMap_sum4_10,addersMap_sum4_9,addersMap_sum4_8,
                 addersMap_sum4_7,addersMap_sum4_6,addersMap_sum4_5,
                 addersMap_sum4_4,addersMap_sum4_3,addersMap_sum4_2,
                 addersMap_sum4_1,addersMap_sum4_0}), .carryOut (\$dummy [162])
                 ) ;
    NBitAdder_16 addersMap_sumFinalMap (.a ({addersMap_sum3Filter_15,
                 addersMap_sum3Filter_14,addersMap_sum3Filter_13,
                 addersMap_sum3Filter_12,addersMap_sum3Filter_11,
                 addersMap_sum3Filter_10,addersMap_sum3Filter_9,
                 addersMap_sum3Filter_8,addersMap_sum3Filter_7,
                 addersMap_sum3Filter_6,addersMap_sum3Filter_5,
                 addersMap_sum3Filter_4,addersMap_sum3Filter_3,
                 addersMap_sum3Filter_2,addersMap_sum3Filter_1,
                 addersMap_sum3Filter_0}), .b ({addersMap_sum4_15,
                 addersMap_sum4_14,addersMap_sum4_13,addersMap_sum4_12,
                 addersMap_sum4_11,addersMap_sum4_10,addersMap_sum4_9,
                 addersMap_sum4_8,addersMap_sum4_7,addersMap_sum4_6,
                 addersMap_sum4_5,addersMap_sum4_4,addersMap_sum4_3,
                 addersMap_sum4_2,addersMap_sum4_1,addersMap_sum4_0}), .carryIn (
                 outShifter_15), .sum ({addersMap_totalSum_15,
                 addersMap_totalSum_14,addersMap_totalSum_13,
                 addersMap_totalSum_12,addersMap_totalSum_11,
                 addersMap_totalSum_10,addersMap_totalSum_9,addersMap_totalSum_8
                 ,addersMap_totalSum_7,addersMap_totalSum_6,addersMap_totalSum_5
                 ,addersMap_totalSum_4,addersMap_totalSum_3,addersMap_totalSum_2
                 ,addersMap_totalSum_1,addersMap_totalSum_0}), .carryOut (
                 \$dummy [163])) ;
    NBitAdder_16 addersMap_sum1Map_sumFinalMap_dup_0 (.a ({
                 addersMap_sum1Map_sum1_15__dup_0,
                 addersMap_sum1Map_sum1_14__dup_0,
                 addersMap_sum1Map_sum1_13__dup_0,
                 addersMap_sum1Map_sum1_12__dup_0,
                 addersMap_sum1Map_sum1_11__dup_0,
                 addersMap_sum1Map_sum1_10__dup_0,
                 addersMap_sum1Map_sum1_9__dup_0,addersMap_sum1Map_sum1_8__dup_0
                 ,addersMap_sum1Map_sum1_7__dup_0,
                 addersMap_sum1Map_sum1_6__dup_0,addersMap_sum1Map_sum1_5__dup_0
                 ,addersMap_sum1Map_sum1_4__dup_0,
                 addersMap_sum1Map_sum1_3__dup_0,addersMap_sum1Map_sum1_2__dup_0
                 ,addersMap_sum1Map_sum1_1__dup_0,
                 addersMap_sum1Map_sum1_0__dup_0}), .b ({
                 addersMap_sum1Map_sum2_15__dup_0,
                 addersMap_sum1Map_sum2_14__dup_0,
                 addersMap_sum1Map_sum2_13__dup_0,
                 addersMap_sum1Map_sum2_12__dup_0,
                 addersMap_sum1Map_sum2_11__dup_0,
                 addersMap_sum1Map_sum2_10__dup_0,
                 addersMap_sum1Map_sum2_9__dup_0,addersMap_sum1Map_sum2_8__dup_0
                 ,addersMap_sum1Map_sum2_7__dup_0,
                 addersMap_sum1Map_sum2_6__dup_0,addersMap_sum1Map_sum2_5__dup_0
                 ,addersMap_sum1Map_sum2_4__dup_0,
                 addersMap_sum1Map_sum2_3__dup_0,addersMap_sum1Map_sum2_2__dup_0
                 ,addersMap_sum1Map_sum2_1__dup_0,
                 addersMap_sum1Map_sum2_0__dup_0}), .carryIn (outShifter_15), .sum (
                 {addersMap_sum1_15,addersMap_sum1_14,addersMap_sum1_13,
                 addersMap_sum1_12,addersMap_sum1_11,addersMap_sum1_10,
                 addersMap_sum1_9,addersMap_sum1_8,addersMap_sum1_7,
                 addersMap_sum1_6,addersMap_sum1_5,addersMap_sum1_4,
                 addersMap_sum1_3,addersMap_sum1_2,addersMap_sum1_1,
                 addersMap_sum1_0}), .carryOut (\$dummy [164])) ;
    NBitAdder_16 addersMap_sum1Map_sum1Map_sum1Map (.a ({addersInputs_0__15,
                 addersInputs_0__14,addersInputs_0__13,addersInputs_0__12,
                 addersInputs_0__11,addersInputs_0__10,addersInputs_0__9,
                 addersInputs_0__8,addersInputs_0__7,addersInputs_0__6,
                 addersInputs_0__5,addersInputs_0__4,addersInputs_0__3,
                 addersInputs_0__2,addersInputs_0__1,addersInputs_0__0}), .b ({
                 addersInputs_1__15,addersInputs_1__14,addersInputs_1__13,
                 addersInputs_1__12,addersInputs_1__11,addersInputs_1__10,
                 addersInputs_1__9,addersInputs_1__8,addersInputs_1__7,
                 addersInputs_1__6,addersInputs_1__5,addersInputs_1__4,
                 addersInputs_1__3,addersInputs_1__2,addersInputs_1__1,
                 addersInputs_1__0}), .carryIn (outShifter_15), .sum ({
                 addersMap_sum1Map_sum1Map_sum1_15,
                 addersMap_sum1Map_sum1Map_sum1_14,
                 addersMap_sum1Map_sum1Map_sum1_13,
                 addersMap_sum1Map_sum1Map_sum1_12,
                 addersMap_sum1Map_sum1Map_sum1_11,
                 addersMap_sum1Map_sum1Map_sum1_10,
                 addersMap_sum1Map_sum1Map_sum1_9,
                 addersMap_sum1Map_sum1Map_sum1_8,
                 addersMap_sum1Map_sum1Map_sum1_7,
                 addersMap_sum1Map_sum1Map_sum1_6,
                 addersMap_sum1Map_sum1Map_sum1_5,
                 addersMap_sum1Map_sum1Map_sum1_4,
                 addersMap_sum1Map_sum1Map_sum1_3,
                 addersMap_sum1Map_sum1Map_sum1_2,
                 addersMap_sum1Map_sum1Map_sum1_1,
                 addersMap_sum1Map_sum1Map_sum1_0}), .carryOut (\$dummy [165])
                 ) ;
    NBitAdder_16 addersMap_sum1Map_sum1Map_sum2Map (.a ({addersInputs_2__15,
                 addersInputs_2__14,addersInputs_2__13,addersInputs_2__12,
                 addersInputs_2__11,addersInputs_2__10,addersInputs_2__9,
                 addersInputs_2__8,addersInputs_2__7,addersInputs_2__6,
                 addersInputs_2__5,addersInputs_2__4,addersInputs_2__3,
                 addersInputs_2__2,addersInputs_2__1,addersInputs_2__0}), .b ({
                 addersInputs_3__15,addersInputs_3__14,addersInputs_3__13,
                 addersInputs_3__12,addersInputs_3__11,addersInputs_3__10,
                 addersInputs_3__9,addersInputs_3__8,addersInputs_3__7,
                 addersInputs_3__6,addersInputs_3__5,addersInputs_3__4,
                 addersInputs_3__3,addersInputs_3__2,addersInputs_3__1,
                 addersInputs_3__0}), .carryIn (outShifter_15), .sum ({
                 addersMap_sum1Map_sum1Map_sum2_15,
                 addersMap_sum1Map_sum1Map_sum2_14,
                 addersMap_sum1Map_sum1Map_sum2_13,
                 addersMap_sum1Map_sum1Map_sum2_12,
                 addersMap_sum1Map_sum1Map_sum2_11,
                 addersMap_sum1Map_sum1Map_sum2_10,
                 addersMap_sum1Map_sum1Map_sum2_9,
                 addersMap_sum1Map_sum1Map_sum2_8,
                 addersMap_sum1Map_sum1Map_sum2_7,
                 addersMap_sum1Map_sum1Map_sum2_6,
                 addersMap_sum1Map_sum1Map_sum2_5,
                 addersMap_sum1Map_sum1Map_sum2_4,
                 addersMap_sum1Map_sum1Map_sum2_3,
                 addersMap_sum1Map_sum1Map_sum2_2,
                 addersMap_sum1Map_sum1Map_sum2_1,
                 addersMap_sum1Map_sum1Map_sum2_0}), .carryOut (\$dummy [166])
                 ) ;
    NBitAdder_16 addersMap_sum1Map_sum1Map_sumFinalMap (.a ({
                 addersMap_sum1Map_sum1Map_sum1_15,
                 addersMap_sum1Map_sum1Map_sum1_14,
                 addersMap_sum1Map_sum1Map_sum1_13,
                 addersMap_sum1Map_sum1Map_sum1_12,
                 addersMap_sum1Map_sum1Map_sum1_11,
                 addersMap_sum1Map_sum1Map_sum1_10,
                 addersMap_sum1Map_sum1Map_sum1_9,
                 addersMap_sum1Map_sum1Map_sum1_8,
                 addersMap_sum1Map_sum1Map_sum1_7,
                 addersMap_sum1Map_sum1Map_sum1_6,
                 addersMap_sum1Map_sum1Map_sum1_5,
                 addersMap_sum1Map_sum1Map_sum1_4,
                 addersMap_sum1Map_sum1Map_sum1_3,
                 addersMap_sum1Map_sum1Map_sum1_2,
                 addersMap_sum1Map_sum1Map_sum1_1,
                 addersMap_sum1Map_sum1Map_sum1_0}), .b ({
                 addersMap_sum1Map_sum1Map_sum2_15,
                 addersMap_sum1Map_sum1Map_sum2_14,
                 addersMap_sum1Map_sum1Map_sum2_13,
                 addersMap_sum1Map_sum1Map_sum2_12,
                 addersMap_sum1Map_sum1Map_sum2_11,
                 addersMap_sum1Map_sum1Map_sum2_10,
                 addersMap_sum1Map_sum1Map_sum2_9,
                 addersMap_sum1Map_sum1Map_sum2_8,
                 addersMap_sum1Map_sum1Map_sum2_7,
                 addersMap_sum1Map_sum1Map_sum2_6,
                 addersMap_sum1Map_sum1Map_sum2_5,
                 addersMap_sum1Map_sum1Map_sum2_4,
                 addersMap_sum1Map_sum1Map_sum2_3,
                 addersMap_sum1Map_sum1Map_sum2_2,
                 addersMap_sum1Map_sum1Map_sum2_1,
                 addersMap_sum1Map_sum1Map_sum2_0}), .carryIn (outShifter_15), .sum (
                 {addersMap_sum1Map_sum1_15__dup_0,
                 addersMap_sum1Map_sum1_14__dup_0,
                 addersMap_sum1Map_sum1_13__dup_0,
                 addersMap_sum1Map_sum1_12__dup_0,
                 addersMap_sum1Map_sum1_11__dup_0,
                 addersMap_sum1Map_sum1_10__dup_0,
                 addersMap_sum1Map_sum1_9__dup_0,addersMap_sum1Map_sum1_8__dup_0
                 ,addersMap_sum1Map_sum1_7__dup_0,
                 addersMap_sum1Map_sum1_6__dup_0,addersMap_sum1Map_sum1_5__dup_0
                 ,addersMap_sum1Map_sum1_4__dup_0,
                 addersMap_sum1Map_sum1_3__dup_0,addersMap_sum1Map_sum1_2__dup_0
                 ,addersMap_sum1Map_sum1_1__dup_0,
                 addersMap_sum1Map_sum1_0__dup_0}), .carryOut (\$dummy [167])) ;
    NBitAdder_16 addersMap_sum1Map_sum2Map_sum1Map (.a ({addersInputs_4__15,
                 addersInputs_4__14,addersInputs_4__13,addersInputs_4__12,
                 addersInputs_4__11,addersInputs_4__10,addersInputs_4__9,
                 addersInputs_4__8,addersInputs_4__7,addersInputs_4__6,
                 addersInputs_4__5,addersInputs_4__4,addersInputs_4__3,
                 addersInputs_4__2,addersInputs_4__1,addersInputs_4__0}), .b ({
                 addersInputs_5__15,addersInputs_5__14,addersInputs_5__13,
                 addersInputs_5__12,addersInputs_5__11,addersInputs_5__10,
                 addersInputs_5__9,addersInputs_5__8,addersInputs_5__7,
                 addersInputs_5__6,addersInputs_5__5,addersInputs_5__4,
                 addersInputs_5__3,addersInputs_5__2,addersInputs_5__1,
                 addersInputs_5__0}), .carryIn (outShifter_15), .sum ({
                 addersMap_sum1Map_sum2Map_sum1_15,
                 addersMap_sum1Map_sum2Map_sum1_14,
                 addersMap_sum1Map_sum2Map_sum1_13,
                 addersMap_sum1Map_sum2Map_sum1_12,
                 addersMap_sum1Map_sum2Map_sum1_11,
                 addersMap_sum1Map_sum2Map_sum1_10,
                 addersMap_sum1Map_sum2Map_sum1_9,
                 addersMap_sum1Map_sum2Map_sum1_8,
                 addersMap_sum1Map_sum2Map_sum1_7,
                 addersMap_sum1Map_sum2Map_sum1_6,
                 addersMap_sum1Map_sum2Map_sum1_5,
                 addersMap_sum1Map_sum2Map_sum1_4,
                 addersMap_sum1Map_sum2Map_sum1_3,
                 addersMap_sum1Map_sum2Map_sum1_2,
                 addersMap_sum1Map_sum2Map_sum1_1,
                 addersMap_sum1Map_sum2Map_sum1_0}), .carryOut (\$dummy [168])
                 ) ;
    NBitAdder_16 addersMap_sum1Map_sum2Map_sum2Map (.a ({addersInputs_6__15,
                 addersInputs_6__14,addersInputs_6__13,addersInputs_6__12,
                 addersInputs_6__11,addersInputs_6__10,addersInputs_6__9,
                 addersInputs_6__8,addersInputs_6__7,addersInputs_6__6,
                 addersInputs_6__5,addersInputs_6__4,addersInputs_6__3,
                 addersInputs_6__2,addersInputs_6__1,addersInputs_6__0}), .b ({
                 addersInputs_7__15,addersInputs_7__14,addersInputs_7__13,
                 addersInputs_7__12,addersInputs_7__11,addersInputs_7__10,
                 addersInputs_7__9,addersInputs_7__8,addersInputs_7__7,
                 addersInputs_7__6,addersInputs_7__5,addersInputs_7__4,
                 addersInputs_7__3,addersInputs_7__2,addersInputs_7__1,
                 addersInputs_7__0}), .carryIn (outShifter_15), .sum ({
                 addersMap_sum1Map_sum2Map_sum2_15,
                 addersMap_sum1Map_sum2Map_sum2_14,
                 addersMap_sum1Map_sum2Map_sum2_13,
                 addersMap_sum1Map_sum2Map_sum2_12,
                 addersMap_sum1Map_sum2Map_sum2_11,
                 addersMap_sum1Map_sum2Map_sum2_10,
                 addersMap_sum1Map_sum2Map_sum2_9,
                 addersMap_sum1Map_sum2Map_sum2_8,
                 addersMap_sum1Map_sum2Map_sum2_7,
                 addersMap_sum1Map_sum2Map_sum2_6,
                 addersMap_sum1Map_sum2Map_sum2_5,
                 addersMap_sum1Map_sum2Map_sum2_4,
                 addersMap_sum1Map_sum2Map_sum2_3,
                 addersMap_sum1Map_sum2Map_sum2_2,
                 addersMap_sum1Map_sum2Map_sum2_1,
                 addersMap_sum1Map_sum2Map_sum2_0}), .carryOut (\$dummy [169])
                 ) ;
    NBitAdder_16 addersMap_sum1Map_sum2Map_sumFinalMap (.a ({
                 addersMap_sum1Map_sum2Map_sum1_15,
                 addersMap_sum1Map_sum2Map_sum1_14,
                 addersMap_sum1Map_sum2Map_sum1_13,
                 addersMap_sum1Map_sum2Map_sum1_12,
                 addersMap_sum1Map_sum2Map_sum1_11,
                 addersMap_sum1Map_sum2Map_sum1_10,
                 addersMap_sum1Map_sum2Map_sum1_9,
                 addersMap_sum1Map_sum2Map_sum1_8,
                 addersMap_sum1Map_sum2Map_sum1_7,
                 addersMap_sum1Map_sum2Map_sum1_6,
                 addersMap_sum1Map_sum2Map_sum1_5,
                 addersMap_sum1Map_sum2Map_sum1_4,
                 addersMap_sum1Map_sum2Map_sum1_3,
                 addersMap_sum1Map_sum2Map_sum1_2,
                 addersMap_sum1Map_sum2Map_sum1_1,
                 addersMap_sum1Map_sum2Map_sum1_0}), .b ({
                 addersMap_sum1Map_sum2Map_sum2_15,
                 addersMap_sum1Map_sum2Map_sum2_14,
                 addersMap_sum1Map_sum2Map_sum2_13,
                 addersMap_sum1Map_sum2Map_sum2_12,
                 addersMap_sum1Map_sum2Map_sum2_11,
                 addersMap_sum1Map_sum2Map_sum2_10,
                 addersMap_sum1Map_sum2Map_sum2_9,
                 addersMap_sum1Map_sum2Map_sum2_8,
                 addersMap_sum1Map_sum2Map_sum2_7,
                 addersMap_sum1Map_sum2Map_sum2_6,
                 addersMap_sum1Map_sum2Map_sum2_5,
                 addersMap_sum1Map_sum2Map_sum2_4,
                 addersMap_sum1Map_sum2Map_sum2_3,
                 addersMap_sum1Map_sum2Map_sum2_2,
                 addersMap_sum1Map_sum2Map_sum2_1,
                 addersMap_sum1Map_sum2Map_sum2_0}), .carryIn (outShifter_15), .sum (
                 {addersMap_sum1Map_sum2_15__dup_0,
                 addersMap_sum1Map_sum2_14__dup_0,
                 addersMap_sum1Map_sum2_13__dup_0,
                 addersMap_sum1Map_sum2_12__dup_0,
                 addersMap_sum1Map_sum2_11__dup_0,
                 addersMap_sum1Map_sum2_10__dup_0,
                 addersMap_sum1Map_sum2_9__dup_0,addersMap_sum1Map_sum2_8__dup_0
                 ,addersMap_sum1Map_sum2_7__dup_0,
                 addersMap_sum1Map_sum2_6__dup_0,addersMap_sum1Map_sum2_5__dup_0
                 ,addersMap_sum1Map_sum2_4__dup_0,
                 addersMap_sum1Map_sum2_3__dup_0,addersMap_sum1Map_sum2_2__dup_0
                 ,addersMap_sum1Map_sum2_1__dup_0,
                 addersMap_sum1Map_sum2_0__dup_0}), .carryOut (\$dummy [170])) ;
    NBitAdder_16 addersMap_sum2Map_sumFinalMap_dup_0 (.a ({
                 addersMap_sum2Map_sum1_15__dup_0,
                 addersMap_sum2Map_sum1_14__dup_0,
                 addersMap_sum2Map_sum1_13__dup_0,
                 addersMap_sum2Map_sum1_12__dup_0,
                 addersMap_sum2Map_sum1_11__dup_0,
                 addersMap_sum2Map_sum1_10__dup_0,
                 addersMap_sum2Map_sum1_9__dup_0,addersMap_sum2Map_sum1_8__dup_0
                 ,addersMap_sum2Map_sum1_7__dup_0,
                 addersMap_sum2Map_sum1_6__dup_0,addersMap_sum2Map_sum1_5__dup_0
                 ,addersMap_sum2Map_sum1_4__dup_0,
                 addersMap_sum2Map_sum1_3__dup_0,addersMap_sum2Map_sum1_2__dup_0
                 ,addersMap_sum2Map_sum1_1__dup_0,
                 addersMap_sum2Map_sum1_0__dup_0}), .b ({
                 addersMap_sum2Map_sum2_15__dup_0,
                 addersMap_sum2Map_sum2_14__dup_0,
                 addersMap_sum2Map_sum2_13__dup_0,
                 addersMap_sum2Map_sum2_12__dup_0,
                 addersMap_sum2Map_sum2_11__dup_0,
                 addersMap_sum2Map_sum2_10__dup_0,
                 addersMap_sum2Map_sum2_9__dup_0,addersMap_sum2Map_sum2_8__dup_0
                 ,addersMap_sum2Map_sum2_7__dup_0,
                 addersMap_sum2Map_sum2_6__dup_0,addersMap_sum2Map_sum2_5__dup_0
                 ,addersMap_sum2Map_sum2_4__dup_0,
                 addersMap_sum2Map_sum2_3__dup_0,addersMap_sum2Map_sum2_2__dup_0
                 ,addersMap_sum2Map_sum2_1__dup_0,
                 addersMap_sum2Map_sum2_0__dup_0}), .carryIn (outShifter_15), .sum (
                 {addersMap_sum2_15,addersMap_sum2_14,addersMap_sum2_13,
                 addersMap_sum2_12,addersMap_sum2_11,addersMap_sum2_10,
                 addersMap_sum2_9,addersMap_sum2_8,addersMap_sum2_7,
                 addersMap_sum2_6,addersMap_sum2_5,addersMap_sum2_4,
                 addersMap_sum2_3,addersMap_sum2_2,addersMap_sum2_1,
                 addersMap_sum2_0}), .carryOut (\$dummy [171])) ;
    NBitAdder_16 addersMap_sum2Map_sum1Map_sum1Map (.a ({addersInputs_9__15,
                 addersInputs_9__14,addersInputs_9__13,addersInputs_9__12,
                 addersInputs_9__11,addersInputs_9__10,addersInputs_9__9,
                 addersInputs_9__8,addersInputs_9__7,addersInputs_9__6,
                 addersInputs_9__5,addersInputs_9__4,addersInputs_9__3,
                 addersInputs_9__2,addersInputs_9__1,addersInputs_9__0}), .b ({
                 addersInputs_10__15,addersInputs_10__14,addersInputs_10__13,
                 addersInputs_10__12,addersInputs_10__11,addersInputs_10__10,
                 addersInputs_10__9,addersInputs_10__8,addersInputs_10__7,
                 addersInputs_10__6,addersInputs_10__5,addersInputs_10__4,
                 addersInputs_10__3,addersInputs_10__2,addersInputs_10__1,
                 addersInputs_10__0}), .carryIn (outShifter_15), .sum ({
                 addersMap_sum2Map_sum1Map_sum1_15,
                 addersMap_sum2Map_sum1Map_sum1_14,
                 addersMap_sum2Map_sum1Map_sum1_13,
                 addersMap_sum2Map_sum1Map_sum1_12,
                 addersMap_sum2Map_sum1Map_sum1_11,
                 addersMap_sum2Map_sum1Map_sum1_10,
                 addersMap_sum2Map_sum1Map_sum1_9,
                 addersMap_sum2Map_sum1Map_sum1_8,
                 addersMap_sum2Map_sum1Map_sum1_7,
                 addersMap_sum2Map_sum1Map_sum1_6,
                 addersMap_sum2Map_sum1Map_sum1_5,
                 addersMap_sum2Map_sum1Map_sum1_4,
                 addersMap_sum2Map_sum1Map_sum1_3,
                 addersMap_sum2Map_sum1Map_sum1_2,
                 addersMap_sum2Map_sum1Map_sum1_1,
                 addersMap_sum2Map_sum1Map_sum1_0}), .carryOut (\$dummy [172])
                 ) ;
    NBitAdder_16 addersMap_sum2Map_sum1Map_sum2Map (.a ({addersInputs_11__15,
                 addersInputs_11__14,addersInputs_11__13,addersInputs_11__12,
                 addersInputs_11__11,addersInputs_11__10,addersInputs_11__9,
                 addersInputs_11__8,addersInputs_11__7,addersInputs_11__6,
                 addersInputs_11__5,addersInputs_11__4,addersInputs_11__3,
                 addersInputs_11__2,addersInputs_11__1,addersInputs_11__0}), .b (
                 {addersInputs_12__15,addersInputs_12__14,addersInputs_12__13,
                 addersInputs_12__12,addersInputs_12__11,addersInputs_12__10,
                 addersInputs_12__9,addersInputs_12__8,addersInputs_12__7,
                 addersInputs_12__6,addersInputs_12__5,addersInputs_12__4,
                 addersInputs_12__3,addersInputs_12__2,addersInputs_12__1,
                 addersInputs_12__0}), .carryIn (outShifter_15), .sum ({
                 addersMap_sum2Map_sum1Map_sum2_15,
                 addersMap_sum2Map_sum1Map_sum2_14,
                 addersMap_sum2Map_sum1Map_sum2_13,
                 addersMap_sum2Map_sum1Map_sum2_12,
                 addersMap_sum2Map_sum1Map_sum2_11,
                 addersMap_sum2Map_sum1Map_sum2_10,
                 addersMap_sum2Map_sum1Map_sum2_9,
                 addersMap_sum2Map_sum1Map_sum2_8,
                 addersMap_sum2Map_sum1Map_sum2_7,
                 addersMap_sum2Map_sum1Map_sum2_6,
                 addersMap_sum2Map_sum1Map_sum2_5,
                 addersMap_sum2Map_sum1Map_sum2_4,
                 addersMap_sum2Map_sum1Map_sum2_3,
                 addersMap_sum2Map_sum1Map_sum2_2,
                 addersMap_sum2Map_sum1Map_sum2_1,
                 addersMap_sum2Map_sum1Map_sum2_0}), .carryOut (\$dummy [173])
                 ) ;
    NBitAdder_16 addersMap_sum2Map_sum1Map_sumFinalMap (.a ({
                 addersMap_sum2Map_sum1Map_sum1_15,
                 addersMap_sum2Map_sum1Map_sum1_14,
                 addersMap_sum2Map_sum1Map_sum1_13,
                 addersMap_sum2Map_sum1Map_sum1_12,
                 addersMap_sum2Map_sum1Map_sum1_11,
                 addersMap_sum2Map_sum1Map_sum1_10,
                 addersMap_sum2Map_sum1Map_sum1_9,
                 addersMap_sum2Map_sum1Map_sum1_8,
                 addersMap_sum2Map_sum1Map_sum1_7,
                 addersMap_sum2Map_sum1Map_sum1_6,
                 addersMap_sum2Map_sum1Map_sum1_5,
                 addersMap_sum2Map_sum1Map_sum1_4,
                 addersMap_sum2Map_sum1Map_sum1_3,
                 addersMap_sum2Map_sum1Map_sum1_2,
                 addersMap_sum2Map_sum1Map_sum1_1,
                 addersMap_sum2Map_sum1Map_sum1_0}), .b ({
                 addersMap_sum2Map_sum1Map_sum2_15,
                 addersMap_sum2Map_sum1Map_sum2_14,
                 addersMap_sum2Map_sum1Map_sum2_13,
                 addersMap_sum2Map_sum1Map_sum2_12,
                 addersMap_sum2Map_sum1Map_sum2_11,
                 addersMap_sum2Map_sum1Map_sum2_10,
                 addersMap_sum2Map_sum1Map_sum2_9,
                 addersMap_sum2Map_sum1Map_sum2_8,
                 addersMap_sum2Map_sum1Map_sum2_7,
                 addersMap_sum2Map_sum1Map_sum2_6,
                 addersMap_sum2Map_sum1Map_sum2_5,
                 addersMap_sum2Map_sum1Map_sum2_4,
                 addersMap_sum2Map_sum1Map_sum2_3,
                 addersMap_sum2Map_sum1Map_sum2_2,
                 addersMap_sum2Map_sum1Map_sum2_1,
                 addersMap_sum2Map_sum1Map_sum2_0}), .carryIn (outShifter_15), .sum (
                 {addersMap_sum2Map_sum1_15__dup_0,
                 addersMap_sum2Map_sum1_14__dup_0,
                 addersMap_sum2Map_sum1_13__dup_0,
                 addersMap_sum2Map_sum1_12__dup_0,
                 addersMap_sum2Map_sum1_11__dup_0,
                 addersMap_sum2Map_sum1_10__dup_0,
                 addersMap_sum2Map_sum1_9__dup_0,addersMap_sum2Map_sum1_8__dup_0
                 ,addersMap_sum2Map_sum1_7__dup_0,
                 addersMap_sum2Map_sum1_6__dup_0,addersMap_sum2Map_sum1_5__dup_0
                 ,addersMap_sum2Map_sum1_4__dup_0,
                 addersMap_sum2Map_sum1_3__dup_0,addersMap_sum2Map_sum1_2__dup_0
                 ,addersMap_sum2Map_sum1_1__dup_0,
                 addersMap_sum2Map_sum1_0__dup_0}), .carryOut (\$dummy [174])) ;
    NBitAdder_16 addersMap_sum2Map_sum2Map_sum1Map (.a ({addersInputs_13__15,
                 addersInputs_13__14,addersInputs_13__13,addersInputs_13__12,
                 addersInputs_13__11,addersInputs_13__10,addersInputs_13__9,
                 addersInputs_13__8,addersInputs_13__7,addersInputs_13__6,
                 addersInputs_13__5,addersInputs_13__4,addersInputs_13__3,
                 addersInputs_13__2,addersInputs_13__1,addersInputs_13__0}), .b (
                 {addersInputs_14__15,addersInputs_14__14,addersInputs_14__13,
                 addersInputs_14__12,addersInputs_14__11,addersInputs_14__10,
                 addersInputs_14__9,addersInputs_14__8,addersInputs_14__7,
                 addersInputs_14__6,addersInputs_14__5,addersInputs_14__4,
                 addersInputs_14__3,addersInputs_14__2,addersInputs_14__1,
                 addersInputs_14__0}), .carryIn (outShifter_15), .sum ({
                 addersMap_sum2Map_sum2Map_sum1_15,
                 addersMap_sum2Map_sum2Map_sum1_14,
                 addersMap_sum2Map_sum2Map_sum1_13,
                 addersMap_sum2Map_sum2Map_sum1_12,
                 addersMap_sum2Map_sum2Map_sum1_11,
                 addersMap_sum2Map_sum2Map_sum1_10,
                 addersMap_sum2Map_sum2Map_sum1_9,
                 addersMap_sum2Map_sum2Map_sum1_8,
                 addersMap_sum2Map_sum2Map_sum1_7,
                 addersMap_sum2Map_sum2Map_sum1_6,
                 addersMap_sum2Map_sum2Map_sum1_5,
                 addersMap_sum2Map_sum2Map_sum1_4,
                 addersMap_sum2Map_sum2Map_sum1_3,
                 addersMap_sum2Map_sum2Map_sum1_2,
                 addersMap_sum2Map_sum2Map_sum1_1,
                 addersMap_sum2Map_sum2Map_sum1_0}), .carryOut (\$dummy [175])
                 ) ;
    NBitAdder_16 addersMap_sum2Map_sum2Map_sum2Map (.a ({addersInputs_15__15,
                 addersInputs_15__14,addersInputs_15__13,addersInputs_15__12,
                 addersInputs_15__11,addersInputs_15__10,addersInputs_15__9,
                 addersInputs_15__8,addersInputs_15__7,addersInputs_15__6,
                 addersInputs_15__5,addersInputs_15__4,addersInputs_15__3,
                 addersInputs_15__2,addersInputs_15__1,addersInputs_15__0}), .b (
                 {addersInputs_16__15,addersInputs_16__14,addersInputs_16__13,
                 addersInputs_16__12,addersInputs_16__11,addersInputs_16__10,
                 addersInputs_16__9,addersInputs_16__8,addersInputs_16__7,
                 addersInputs_16__6,addersInputs_16__5,addersInputs_16__4,
                 addersInputs_16__3,addersInputs_16__2,addersInputs_16__1,
                 addersInputs_16__0}), .carryIn (outShifter_15), .sum ({
                 addersMap_sum2Map_sum2Map_sum2_15,
                 addersMap_sum2Map_sum2Map_sum2_14,
                 addersMap_sum2Map_sum2Map_sum2_13,
                 addersMap_sum2Map_sum2Map_sum2_12,
                 addersMap_sum2Map_sum2Map_sum2_11,
                 addersMap_sum2Map_sum2Map_sum2_10,
                 addersMap_sum2Map_sum2Map_sum2_9,
                 addersMap_sum2Map_sum2Map_sum2_8,
                 addersMap_sum2Map_sum2Map_sum2_7,
                 addersMap_sum2Map_sum2Map_sum2_6,
                 addersMap_sum2Map_sum2Map_sum2_5,
                 addersMap_sum2Map_sum2Map_sum2_4,
                 addersMap_sum2Map_sum2Map_sum2_3,
                 addersMap_sum2Map_sum2Map_sum2_2,
                 addersMap_sum2Map_sum2Map_sum2_1,
                 addersMap_sum2Map_sum2Map_sum2_0}), .carryOut (\$dummy [176])
                 ) ;
    NBitAdder_16 addersMap_sum2Map_sum2Map_sumFinalMap (.a ({
                 addersMap_sum2Map_sum2Map_sum1_15,
                 addersMap_sum2Map_sum2Map_sum1_14,
                 addersMap_sum2Map_sum2Map_sum1_13,
                 addersMap_sum2Map_sum2Map_sum1_12,
                 addersMap_sum2Map_sum2Map_sum1_11,
                 addersMap_sum2Map_sum2Map_sum1_10,
                 addersMap_sum2Map_sum2Map_sum1_9,
                 addersMap_sum2Map_sum2Map_sum1_8,
                 addersMap_sum2Map_sum2Map_sum1_7,
                 addersMap_sum2Map_sum2Map_sum1_6,
                 addersMap_sum2Map_sum2Map_sum1_5,
                 addersMap_sum2Map_sum2Map_sum1_4,
                 addersMap_sum2Map_sum2Map_sum1_3,
                 addersMap_sum2Map_sum2Map_sum1_2,
                 addersMap_sum2Map_sum2Map_sum1_1,
                 addersMap_sum2Map_sum2Map_sum1_0}), .b ({
                 addersMap_sum2Map_sum2Map_sum2_15,
                 addersMap_sum2Map_sum2Map_sum2_14,
                 addersMap_sum2Map_sum2Map_sum2_13,
                 addersMap_sum2Map_sum2Map_sum2_12,
                 addersMap_sum2Map_sum2Map_sum2_11,
                 addersMap_sum2Map_sum2Map_sum2_10,
                 addersMap_sum2Map_sum2Map_sum2_9,
                 addersMap_sum2Map_sum2Map_sum2_8,
                 addersMap_sum2Map_sum2Map_sum2_7,
                 addersMap_sum2Map_sum2Map_sum2_6,
                 addersMap_sum2Map_sum2Map_sum2_5,
                 addersMap_sum2Map_sum2Map_sum2_4,
                 addersMap_sum2Map_sum2Map_sum2_3,
                 addersMap_sum2Map_sum2Map_sum2_2,
                 addersMap_sum2Map_sum2Map_sum2_1,
                 addersMap_sum2Map_sum2Map_sum2_0}), .carryIn (outShifter_15), .sum (
                 {addersMap_sum2Map_sum2_15__dup_0,
                 addersMap_sum2Map_sum2_14__dup_0,
                 addersMap_sum2Map_sum2_13__dup_0,
                 addersMap_sum2Map_sum2_12__dup_0,
                 addersMap_sum2Map_sum2_11__dup_0,
                 addersMap_sum2Map_sum2_10__dup_0,
                 addersMap_sum2Map_sum2_9__dup_0,addersMap_sum2Map_sum2_8__dup_0
                 ,addersMap_sum2Map_sum2_7__dup_0,
                 addersMap_sum2Map_sum2_6__dup_0,addersMap_sum2Map_sum2_5__dup_0
                 ,addersMap_sum2Map_sum2_4__dup_0,
                 addersMap_sum2Map_sum2_3__dup_0,addersMap_sum2Map_sum2_2__dup_0
                 ,addersMap_sum2Map_sum2_1__dup_0,
                 addersMap_sum2Map_sum2_0__dup_0}), .carryOut (\$dummy [177])) ;
    NBitAdder_16 addersMap_sum3Map_sumFinalMap (.a ({addersMap_sum3Map_sum1_15,
                 addersMap_sum3Map_sum1_14,addersMap_sum3Map_sum1_13,
                 addersMap_sum3Map_sum1_12,addersMap_sum3Map_sum1_11,
                 addersMap_sum3Map_sum1_10,addersMap_sum3Map_sum1_9,
                 addersMap_sum3Map_sum1_8,addersMap_sum3Map_sum1_7,
                 addersMap_sum3Map_sum1_6,addersMap_sum3Map_sum1_5,
                 addersMap_sum3Map_sum1_4,addersMap_sum3Map_sum1_3,
                 addersMap_sum3Map_sum1_2,addersMap_sum3Map_sum1_1,
                 addersMap_sum3Map_sum1_0}), .b ({addersMap_sum3Map_sum2_15,
                 addersMap_sum3Map_sum2_14,addersMap_sum3Map_sum2_13,
                 addersMap_sum3Map_sum2_12,addersMap_sum3Map_sum2_11,
                 addersMap_sum3Map_sum2_10,addersMap_sum3Map_sum2_9,
                 addersMap_sum3Map_sum2_8,addersMap_sum3Map_sum2_7,
                 addersMap_sum3Map_sum2_6,addersMap_sum3Map_sum2_5,
                 addersMap_sum3Map_sum2_4,addersMap_sum3Map_sum2_3,
                 addersMap_sum3Map_sum2_2,addersMap_sum3Map_sum2_1,
                 addersMap_sum3Map_sum2_0}), .carryIn (outShifter_15), .sum ({
                 addersMap_sum3_15,addersMap_sum3_14,addersMap_sum3_13,
                 addersMap_sum3_12,addersMap_sum3_11,addersMap_sum3_10,
                 addersMap_sum3_9,addersMap_sum3_8,addersMap_sum3_7,
                 addersMap_sum3_6,addersMap_sum3_5,addersMap_sum3_4,
                 addersMap_sum3_3,addersMap_sum3_2,addersMap_sum3_1,
                 addersMap_sum3_0}), .carryOut (\$dummy [178])) ;
    NBitAdder_16 addersMap_sum3Map_sum1Map_sum1Map (.a ({addersInputs_17__15,
                 addersInputs_17__14,addersInputs_17__13,addersInputs_17__12,
                 addersInputs_17__11,addersInputs_17__10,addersInputs_17__9,
                 addersInputs_17__8,addersInputs_17__7,addersInputs_17__6,
                 addersInputs_17__5,addersInputs_17__4,addersInputs_17__3,
                 addersInputs_17__2,addersInputs_17__1,addersInputs_17__0}), .b (
                 {addersInputs_18__15,addersInputs_18__14,addersInputs_18__13,
                 addersInputs_18__12,addersInputs_18__11,addersInputs_18__10,
                 addersInputs_18__9,addersInputs_18__8,addersInputs_18__7,
                 addersInputs_18__6,addersInputs_18__5,addersInputs_18__4,
                 addersInputs_18__3,addersInputs_18__2,addersInputs_18__1,
                 addersInputs_18__0}), .carryIn (outShifter_15), .sum ({
                 addersMap_sum3Map_sum1Map_sum1_15,
                 addersMap_sum3Map_sum1Map_sum1_14,
                 addersMap_sum3Map_sum1Map_sum1_13,
                 addersMap_sum3Map_sum1Map_sum1_12,
                 addersMap_sum3Map_sum1Map_sum1_11,
                 addersMap_sum3Map_sum1Map_sum1_10,
                 addersMap_sum3Map_sum1Map_sum1_9,
                 addersMap_sum3Map_sum1Map_sum1_8,
                 addersMap_sum3Map_sum1Map_sum1_7,
                 addersMap_sum3Map_sum1Map_sum1_6,
                 addersMap_sum3Map_sum1Map_sum1_5,
                 addersMap_sum3Map_sum1Map_sum1_4,
                 addersMap_sum3Map_sum1Map_sum1_3,
                 addersMap_sum3Map_sum1Map_sum1_2,
                 addersMap_sum3Map_sum1Map_sum1_1,
                 addersMap_sum3Map_sum1Map_sum1_0}), .carryOut (\$dummy [179])
                 ) ;
    NBitAdder_16 addersMap_sum3Map_sum1Map_sum2Map (.a ({addersInputs_19__15,
                 addersInputs_19__14,addersInputs_19__13,addersInputs_19__12,
                 addersInputs_19__11,addersInputs_19__10,addersInputs_19__9,
                 addersInputs_19__8,addersInputs_19__7,addersInputs_19__6,
                 addersInputs_19__5,addersInputs_19__4,addersInputs_19__3,
                 addersInputs_19__2,addersInputs_19__1,addersInputs_19__0}), .b (
                 {addersInputs_20__15,addersInputs_20__14,addersInputs_20__13,
                 addersInputs_20__12,addersInputs_20__11,addersInputs_20__10,
                 addersInputs_20__9,addersInputs_20__8,addersInputs_20__7,
                 addersInputs_20__6,addersInputs_20__5,addersInputs_20__4,
                 addersInputs_20__3,addersInputs_20__2,addersInputs_20__1,
                 addersInputs_20__0}), .carryIn (outShifter_15), .sum ({
                 addersMap_sum3Map_sum1Map_sum2_15,
                 addersMap_sum3Map_sum1Map_sum2_14,
                 addersMap_sum3Map_sum1Map_sum2_13,
                 addersMap_sum3Map_sum1Map_sum2_12,
                 addersMap_sum3Map_sum1Map_sum2_11,
                 addersMap_sum3Map_sum1Map_sum2_10,
                 addersMap_sum3Map_sum1Map_sum2_9,
                 addersMap_sum3Map_sum1Map_sum2_8,
                 addersMap_sum3Map_sum1Map_sum2_7,
                 addersMap_sum3Map_sum1Map_sum2_6,
                 addersMap_sum3Map_sum1Map_sum2_5,
                 addersMap_sum3Map_sum1Map_sum2_4,
                 addersMap_sum3Map_sum1Map_sum2_3,
                 addersMap_sum3Map_sum1Map_sum2_2,
                 addersMap_sum3Map_sum1Map_sum2_1,
                 addersMap_sum3Map_sum1Map_sum2_0}), .carryOut (\$dummy [180])
                 ) ;
    NBitAdder_16 addersMap_sum3Map_sum1Map_sumFinalMap (.a ({
                 addersMap_sum3Map_sum1Map_sum1_15,
                 addersMap_sum3Map_sum1Map_sum1_14,
                 addersMap_sum3Map_sum1Map_sum1_13,
                 addersMap_sum3Map_sum1Map_sum1_12,
                 addersMap_sum3Map_sum1Map_sum1_11,
                 addersMap_sum3Map_sum1Map_sum1_10,
                 addersMap_sum3Map_sum1Map_sum1_9,
                 addersMap_sum3Map_sum1Map_sum1_8,
                 addersMap_sum3Map_sum1Map_sum1_7,
                 addersMap_sum3Map_sum1Map_sum1_6,
                 addersMap_sum3Map_sum1Map_sum1_5,
                 addersMap_sum3Map_sum1Map_sum1_4,
                 addersMap_sum3Map_sum1Map_sum1_3,
                 addersMap_sum3Map_sum1Map_sum1_2,
                 addersMap_sum3Map_sum1Map_sum1_1,
                 addersMap_sum3Map_sum1Map_sum1_0}), .b ({
                 addersMap_sum3Map_sum1Map_sum2_15,
                 addersMap_sum3Map_sum1Map_sum2_14,
                 addersMap_sum3Map_sum1Map_sum2_13,
                 addersMap_sum3Map_sum1Map_sum2_12,
                 addersMap_sum3Map_sum1Map_sum2_11,
                 addersMap_sum3Map_sum1Map_sum2_10,
                 addersMap_sum3Map_sum1Map_sum2_9,
                 addersMap_sum3Map_sum1Map_sum2_8,
                 addersMap_sum3Map_sum1Map_sum2_7,
                 addersMap_sum3Map_sum1Map_sum2_6,
                 addersMap_sum3Map_sum1Map_sum2_5,
                 addersMap_sum3Map_sum1Map_sum2_4,
                 addersMap_sum3Map_sum1Map_sum2_3,
                 addersMap_sum3Map_sum1Map_sum2_2,
                 addersMap_sum3Map_sum1Map_sum2_1,
                 addersMap_sum3Map_sum1Map_sum2_0}), .carryIn (outShifter_15), .sum (
                 {addersMap_sum3Map_sum1_15,addersMap_sum3Map_sum1_14,
                 addersMap_sum3Map_sum1_13,addersMap_sum3Map_sum1_12,
                 addersMap_sum3Map_sum1_11,addersMap_sum3Map_sum1_10,
                 addersMap_sum3Map_sum1_9,addersMap_sum3Map_sum1_8,
                 addersMap_sum3Map_sum1_7,addersMap_sum3Map_sum1_6,
                 addersMap_sum3Map_sum1_5,addersMap_sum3Map_sum1_4,
                 addersMap_sum3Map_sum1_3,addersMap_sum3Map_sum1_2,
                 addersMap_sum3Map_sum1_1,addersMap_sum3Map_sum1_0}), .carryOut (
                 \$dummy [181])) ;
    NBitAdder_16 addersMap_sum3Map_sum2Map_sum1Map (.a ({addersInputs_21__15,
                 addersInputs_21__14,addersInputs_21__13,addersInputs_21__12,
                 addersInputs_21__11,addersInputs_21__10,addersInputs_21__9,
                 addersInputs_21__8,addersInputs_21__7,addersInputs_21__6,
                 addersInputs_21__5,addersInputs_21__4,addersInputs_21__3,
                 addersInputs_21__2,addersInputs_21__1,addersInputs_21__0}), .b (
                 {addersInputs_22__15,addersInputs_22__14,addersInputs_22__13,
                 addersInputs_22__12,addersInputs_22__11,addersInputs_22__10,
                 addersInputs_22__9,addersInputs_22__8,addersInputs_22__7,
                 addersInputs_22__6,addersInputs_22__5,addersInputs_22__4,
                 addersInputs_22__3,addersInputs_22__2,addersInputs_22__1,
                 addersInputs_22__0}), .carryIn (outShifter_15), .sum ({
                 addersMap_sum3Map_sum2Map_sum1_15,
                 addersMap_sum3Map_sum2Map_sum1_14,
                 addersMap_sum3Map_sum2Map_sum1_13,
                 addersMap_sum3Map_sum2Map_sum1_12,
                 addersMap_sum3Map_sum2Map_sum1_11,
                 addersMap_sum3Map_sum2Map_sum1_10,
                 addersMap_sum3Map_sum2Map_sum1_9,
                 addersMap_sum3Map_sum2Map_sum1_8,
                 addersMap_sum3Map_sum2Map_sum1_7,
                 addersMap_sum3Map_sum2Map_sum1_6,
                 addersMap_sum3Map_sum2Map_sum1_5,
                 addersMap_sum3Map_sum2Map_sum1_4,
                 addersMap_sum3Map_sum2Map_sum1_3,
                 addersMap_sum3Map_sum2Map_sum1_2,
                 addersMap_sum3Map_sum2Map_sum1_1,
                 addersMap_sum3Map_sum2Map_sum1_0}), .carryOut (\$dummy [182])
                 ) ;
    NBitAdder_16 addersMap_sum3Map_sum2Map_sum2Map (.a ({addersInputs_23__15,
                 addersInputs_23__14,addersInputs_23__13,addersInputs_23__12,
                 addersInputs_23__11,addersInputs_23__10,addersInputs_23__9,
                 addersInputs_23__8,addersInputs_23__7,addersInputs_23__6,
                 addersInputs_23__5,addersInputs_23__4,addersInputs_23__3,
                 addersInputs_23__2,addersInputs_23__1,addersInputs_23__0}), .b (
                 {addersInputs_24__15,addersInputs_24__14,addersInputs_24__13,
                 addersInputs_24__12,addersInputs_24__11,addersInputs_24__10,
                 addersInputs_24__9,addersInputs_24__8,addersInputs_24__7,
                 addersInputs_24__6,addersInputs_24__5,addersInputs_24__4,
                 addersInputs_24__3,addersInputs_24__2,addersInputs_24__1,
                 addersInputs_24__0}), .carryIn (outShifter_15), .sum ({
                 addersMap_sum3Map_sum2Map_sum2_15,
                 addersMap_sum3Map_sum2Map_sum2_14,
                 addersMap_sum3Map_sum2Map_sum2_13,
                 addersMap_sum3Map_sum2Map_sum2_12,
                 addersMap_sum3Map_sum2Map_sum2_11,
                 addersMap_sum3Map_sum2Map_sum2_10,
                 addersMap_sum3Map_sum2Map_sum2_9,
                 addersMap_sum3Map_sum2Map_sum2_8,
                 addersMap_sum3Map_sum2Map_sum2_7,
                 addersMap_sum3Map_sum2Map_sum2_6,
                 addersMap_sum3Map_sum2Map_sum2_5,
                 addersMap_sum3Map_sum2Map_sum2_4,
                 addersMap_sum3Map_sum2Map_sum2_3,
                 addersMap_sum3Map_sum2Map_sum2_2,
                 addersMap_sum3Map_sum2Map_sum2_1,
                 addersMap_sum3Map_sum2Map_sum2_0}), .carryOut (\$dummy [183])
                 ) ;
    NBitAdder_16 addersMap_sum3Map_sum2Map_sumFinalMap (.a ({
                 addersMap_sum3Map_sum2Map_sum1_15,
                 addersMap_sum3Map_sum2Map_sum1_14,
                 addersMap_sum3Map_sum2Map_sum1_13,
                 addersMap_sum3Map_sum2Map_sum1_12,
                 addersMap_sum3Map_sum2Map_sum1_11,
                 addersMap_sum3Map_sum2Map_sum1_10,
                 addersMap_sum3Map_sum2Map_sum1_9,
                 addersMap_sum3Map_sum2Map_sum1_8,
                 addersMap_sum3Map_sum2Map_sum1_7,
                 addersMap_sum3Map_sum2Map_sum1_6,
                 addersMap_sum3Map_sum2Map_sum1_5,
                 addersMap_sum3Map_sum2Map_sum1_4,
                 addersMap_sum3Map_sum2Map_sum1_3,
                 addersMap_sum3Map_sum2Map_sum1_2,
                 addersMap_sum3Map_sum2Map_sum1_1,
                 addersMap_sum3Map_sum2Map_sum1_0}), .b ({
                 addersMap_sum3Map_sum2Map_sum2_15,
                 addersMap_sum3Map_sum2Map_sum2_14,
                 addersMap_sum3Map_sum2Map_sum2_13,
                 addersMap_sum3Map_sum2Map_sum2_12,
                 addersMap_sum3Map_sum2Map_sum2_11,
                 addersMap_sum3Map_sum2Map_sum2_10,
                 addersMap_sum3Map_sum2Map_sum2_9,
                 addersMap_sum3Map_sum2Map_sum2_8,
                 addersMap_sum3Map_sum2Map_sum2_7,
                 addersMap_sum3Map_sum2Map_sum2_6,
                 addersMap_sum3Map_sum2Map_sum2_5,
                 addersMap_sum3Map_sum2Map_sum2_4,
                 addersMap_sum3Map_sum2Map_sum2_3,
                 addersMap_sum3Map_sum2Map_sum2_2,
                 addersMap_sum3Map_sum2Map_sum2_1,
                 addersMap_sum3Map_sum2Map_sum2_0}), .carryIn (outShifter_15), .sum (
                 {addersMap_sum3Map_sum2_15,addersMap_sum3Map_sum2_14,
                 addersMap_sum3Map_sum2_13,addersMap_sum3Map_sum2_12,
                 addersMap_sum3Map_sum2_11,addersMap_sum3Map_sum2_10,
                 addersMap_sum3Map_sum2_9,addersMap_sum3Map_sum2_8,
                 addersMap_sum3Map_sum2_7,addersMap_sum3Map_sum2_6,
                 addersMap_sum3Map_sum2_5,addersMap_sum3Map_sum2_4,
                 addersMap_sum3Map_sum2_3,addersMap_sum3Map_sum2_2,
                 addersMap_sum3Map_sum2_1,addersMap_sum3Map_sum2_0}), .carryOut (
                 \$dummy [184])) ;
    fake_gnd ix2066 (.Y (outShifter_15)) ;
    nand03 ix2918 (.Y (nx2917), .A0 (writeFilter), .A1 (nx3412), .A2 (
           decoderRow[2])) ;
    nor02_2x ix3413 (.Y (nx3412), .A0 (decoderRow[1]), .A1 (decoderRow[0])) ;
    nor03_2x ix3437 (.Y (regFileMap_filterEnables_3), .A0 (nx2923), .A1 (
             decoderRow[2]), .A2 (nx2925)) ;
    inv02 ix2924 (.Y (nx2923), .A (writeFilter)) ;
    nand02 ix2926 (.Y (nx2925), .A0 (decoderRow[1]), .A1 (decoderRow[0])) ;
    nor03_2x ix3449 (.Y (regFileMap_filterEnables_2), .A0 (nx2923), .A1 (
             decoderRow[2]), .A2 (nx2929)) ;
    nand02 ix2930 (.Y (nx2929), .A0 (decoderRow[1]), .A1 (nx2931)) ;
    inv01 ix2932 (.Y (nx2931), .A (decoderRow[0])) ;
    nor03_2x ix3461 (.Y (regFileMap_filterEnables_1), .A0 (nx2923), .A1 (
             decoderRow[2]), .A2 (nx2935)) ;
    nand02 ix2936 (.Y (nx2935), .A0 (nx2937), .A1 (decoderRow[0])) ;
    inv01 ix2938 (.Y (nx2937), .A (decoderRow[1])) ;
    nor03_2x ix3475 (.Y (regFileMap_filterEnables_0), .A0 (nx2923), .A1 (
             decoderRow[2]), .A2 (nx2941)) ;
    inv01 ix2942 (.Y (nx2941), .A (nx3470)) ;
    nor02_2x ix3471 (.Y (nx3470), .A0 (decoderRow[1]), .A1 (decoderRow[0])) ;
    inv01 ix3425 (.Y (regFileMap_page2Enables_4), .A (nx2947)) ;
    nand03 ix2948 (.Y (nx2947), .A0 (writePage2), .A1 (nx3412), .A2 (
           decoderRow[2])) ;
    nor03_2x ix3439 (.Y (regFileMap_page2Enables_3), .A0 (nx2951), .A1 (
             decoderRow[2]), .A2 (nx2925)) ;
    inv02 ix2952 (.Y (nx2951), .A (writePage2)) ;
    nor03_2x ix3451 (.Y (regFileMap_page2Enables_2), .A0 (nx2951), .A1 (
             decoderRow[2]), .A2 (nx2929)) ;
    nor03_2x ix3463 (.Y (regFileMap_page2Enables_1), .A0 (nx2951), .A1 (
             decoderRow[2]), .A2 (nx2935)) ;
    nor03_2x ix3477 (.Y (regFileMap_page2Enables_0), .A0 (nx2951), .A1 (
             decoderRow[2]), .A2 (nx2941)) ;
    inv01 ix3427 (.Y (regFileMap_page1Enables_4), .A (nx2959)) ;
    nand03 ix2960 (.Y (nx2959), .A0 (writePage1), .A1 (nx3412), .A2 (
           decoderRow[2])) ;
    nor03_2x ix3441 (.Y (regFileMap_page1Enables_3), .A0 (nx2963), .A1 (
             decoderRow[2]), .A2 (nx2925)) ;
    inv02 ix2964 (.Y (nx2963), .A (writePage1)) ;
    nor03_2x ix3453 (.Y (regFileMap_page1Enables_2), .A0 (nx2963), .A1 (
             decoderRow[2]), .A2 (nx2929)) ;
    nor03_2x ix3465 (.Y (regFileMap_page1Enables_1), .A0 (nx2963), .A1 (
             decoderRow[2]), .A2 (nx2935)) ;
    nor03_2x ix3479 (.Y (regFileMap_page1Enables_0), .A0 (nx2963), .A1 (
             decoderRow[2]), .A2 (nx2941)) ;
    nand02 ix215 (.Y (addersInputs_24__0), .A0 (nx2971), .A1 (nx2973)) ;
    nand02 ix2972 (.Y (nx2971), .A0 (currentPage_24__0), .A1 (layerType)) ;
    nand02 ix2974 (.Y (nx2973), .A0 (outMuls_24__0), .A1 (nx5200)) ;
    nand02 ix223 (.Y (addersInputs_24__1), .A0 (nx2979), .A1 (nx2981)) ;
    nand02 ix2980 (.Y (nx2979), .A0 (currentPage_24__1), .A1 (layerType)) ;
    nand02 ix2982 (.Y (nx2981), .A0 (outMuls_24__1), .A1 (nx5200)) ;
    nand02 ix231 (.Y (addersInputs_24__2), .A0 (nx2985), .A1 (nx2987)) ;
    nand02 ix2986 (.Y (nx2985), .A0 (currentPage_24__2), .A1 (layerType)) ;
    nand02 ix2988 (.Y (nx2987), .A0 (outMuls_24__2), .A1 (nx5200)) ;
    nand02 ix239 (.Y (addersInputs_24__3), .A0 (nx2991), .A1 (nx2993)) ;
    nand02 ix2992 (.Y (nx2991), .A0 (currentPage_24__3), .A1 (layerType)) ;
    nand02 ix2994 (.Y (nx2993), .A0 (outMuls_24__3), .A1 (nx5200)) ;
    nand02 ix247 (.Y (addersInputs_24__4), .A0 (nx2997), .A1 (nx2999)) ;
    nand02 ix2998 (.Y (nx2997), .A0 (currentPage_24__4), .A1 (layerType)) ;
    nand02 ix3000 (.Y (nx2999), .A0 (outMuls_24__4), .A1 (nx5200)) ;
    nand02 ix255 (.Y (addersInputs_24__5), .A0 (nx3003), .A1 (nx3005)) ;
    nand02 ix3004 (.Y (nx3003), .A0 (currentPage_24__5), .A1 (layerType)) ;
    nand02 ix3006 (.Y (nx3005), .A0 (outMuls_24__5), .A1 (nx5200)) ;
    nand02 ix263 (.Y (addersInputs_24__6), .A0 (nx3009), .A1 (nx3011)) ;
    nand02 ix3010 (.Y (nx3009), .A0 (currentPage_24__6), .A1 (layerType)) ;
    nand02 ix3012 (.Y (nx3011), .A0 (outMuls_24__6), .A1 (nx5200)) ;
    nand02 ix271 (.Y (addersInputs_24__7), .A0 (nx3015), .A1 (nx3017)) ;
    nand02 ix3016 (.Y (nx3015), .A0 (currentPage_24__7), .A1 (layerType)) ;
    nand02 ix3018 (.Y (nx3017), .A0 (outMuls_24__7), .A1 (nx5202)) ;
    nand02 ix279 (.Y (addersInputs_24__8), .A0 (nx3021), .A1 (nx3023)) ;
    nand02 ix3022 (.Y (nx3021), .A0 (currentPage_24__8), .A1 (layerType)) ;
    nand02 ix3024 (.Y (nx3023), .A0 (outMuls_24__8), .A1 (nx5202)) ;
    nand02 ix287 (.Y (addersInputs_24__9), .A0 (nx3027), .A1 (nx3029)) ;
    nand02 ix3028 (.Y (nx3027), .A0 (currentPage_24__9), .A1 (layerType)) ;
    nand02 ix3030 (.Y (nx3029), .A0 (outMuls_24__9), .A1 (nx5202)) ;
    nand02 ix295 (.Y (addersInputs_24__10), .A0 (nx3033), .A1 (nx3035)) ;
    nand02 ix3034 (.Y (nx3033), .A0 (currentPage_24__10), .A1 (layerType)) ;
    nand02 ix3036 (.Y (nx3035), .A0 (outMuls_24__10), .A1 (nx5202)) ;
    nand02 ix303 (.Y (addersInputs_24__11), .A0 (nx3039), .A1 (nx3041)) ;
    nand02 ix3040 (.Y (nx3039), .A0 (currentPage_24__11), .A1 (layerType)) ;
    nand02 ix3042 (.Y (nx3041), .A0 (outMuls_24__11), .A1 (nx5202)) ;
    nand02 ix311 (.Y (addersInputs_24__12), .A0 (nx3045), .A1 (nx3047)) ;
    nand02 ix3046 (.Y (nx3045), .A0 (currentPage_24__12), .A1 (layerType)) ;
    nand02 ix3048 (.Y (nx3047), .A0 (outMuls_24__12), .A1 (nx5202)) ;
    nand02 ix319 (.Y (addersInputs_24__13), .A0 (nx3051), .A1 (nx3053)) ;
    nand02 ix3052 (.Y (nx3051), .A0 (currentPage_24__13), .A1 (layerType)) ;
    nand02 ix3054 (.Y (nx3053), .A0 (outMuls_24__13), .A1 (nx5202)) ;
    nand02 ix327 (.Y (addersInputs_24__14), .A0 (nx3057), .A1 (nx3059)) ;
    nand02 ix3058 (.Y (nx3057), .A0 (currentPage_24__14), .A1 (layerType)) ;
    nand02 ix3060 (.Y (nx3059), .A0 (outMuls_24__14), .A1 (nx5204)) ;
    nand02 ix335 (.Y (addersInputs_24__15), .A0 (nx3063), .A1 (nx3065)) ;
    nand02 ix3064 (.Y (nx3063), .A0 (currentPage_24__15), .A1 (layerType)) ;
    nand02 ix3066 (.Y (nx3065), .A0 (outMuls_24__15), .A1 (nx5204)) ;
    nand02 ix343 (.Y (addersInputs_23__0), .A0 (nx3069), .A1 (nx3071)) ;
    nand02 ix3070 (.Y (nx3069), .A0 (currentPage_23__0), .A1 (layerType)) ;
    nand02 ix3072 (.Y (nx3071), .A0 (outMuls_23__0), .A1 (nx5204)) ;
    nand02 ix351 (.Y (addersInputs_23__1), .A0 (nx3075), .A1 (nx3077)) ;
    nand02 ix3076 (.Y (nx3075), .A0 (currentPage_23__1), .A1 (layerType)) ;
    nand02 ix3078 (.Y (nx3077), .A0 (outMuls_23__1), .A1 (nx5204)) ;
    nand02 ix359 (.Y (addersInputs_23__2), .A0 (nx3081), .A1 (nx3083)) ;
    nand02 ix3082 (.Y (nx3081), .A0 (currentPage_23__2), .A1 (layerType)) ;
    nand02 ix3084 (.Y (nx3083), .A0 (outMuls_23__2), .A1 (nx5204)) ;
    nand02 ix367 (.Y (addersInputs_23__3), .A0 (nx3087), .A1 (nx3089)) ;
    nand02 ix3088 (.Y (nx3087), .A0 (currentPage_23__3), .A1 (layerType)) ;
    nand02 ix3090 (.Y (nx3089), .A0 (outMuls_23__3), .A1 (nx5204)) ;
    nand02 ix375 (.Y (addersInputs_23__4), .A0 (nx3093), .A1 (nx3095)) ;
    nand02 ix3094 (.Y (nx3093), .A0 (currentPage_23__4), .A1 (layerType)) ;
    nand02 ix3096 (.Y (nx3095), .A0 (outMuls_23__4), .A1 (nx5204)) ;
    nand02 ix383 (.Y (addersInputs_23__5), .A0 (nx3099), .A1 (nx3101)) ;
    nand02 ix3100 (.Y (nx3099), .A0 (currentPage_23__5), .A1 (layerType)) ;
    nand02 ix3102 (.Y (nx3101), .A0 (outMuls_23__5), .A1 (nx5206)) ;
    nand02 ix391 (.Y (addersInputs_23__6), .A0 (nx3105), .A1 (nx3107)) ;
    nand02 ix3106 (.Y (nx3105), .A0 (currentPage_23__6), .A1 (layerType)) ;
    nand02 ix3108 (.Y (nx3107), .A0 (outMuls_23__6), .A1 (nx5206)) ;
    nand02 ix399 (.Y (addersInputs_23__7), .A0 (nx3111), .A1 (nx3113)) ;
    nand02 ix3112 (.Y (nx3111), .A0 (currentPage_23__7), .A1 (layerType)) ;
    nand02 ix3114 (.Y (nx3113), .A0 (outMuls_23__7), .A1 (nx5206)) ;
    nand02 ix407 (.Y (addersInputs_23__8), .A0 (nx3117), .A1 (nx3119)) ;
    nand02 ix3118 (.Y (nx3117), .A0 (currentPage_23__8), .A1 (layerType)) ;
    nand02 ix3120 (.Y (nx3119), .A0 (outMuls_23__8), .A1 (nx5206)) ;
    nand02 ix415 (.Y (addersInputs_23__9), .A0 (nx3123), .A1 (nx3125)) ;
    nand02 ix3124 (.Y (nx3123), .A0 (currentPage_23__9), .A1 (layerType)) ;
    nand02 ix3126 (.Y (nx3125), .A0 (outMuls_23__9), .A1 (nx5206)) ;
    nand02 ix423 (.Y (addersInputs_23__10), .A0 (nx3129), .A1 (nx3131)) ;
    nand02 ix3130 (.Y (nx3129), .A0 (currentPage_23__10), .A1 (layerType)) ;
    nand02 ix3132 (.Y (nx3131), .A0 (outMuls_23__10), .A1 (nx5206)) ;
    nand02 ix431 (.Y (addersInputs_23__11), .A0 (nx3135), .A1 (nx3137)) ;
    nand02 ix3136 (.Y (nx3135), .A0 (currentPage_23__11), .A1 (layerType)) ;
    nand02 ix3138 (.Y (nx3137), .A0 (outMuls_23__11), .A1 (nx5206)) ;
    nand02 ix439 (.Y (addersInputs_23__12), .A0 (nx3141), .A1 (nx3143)) ;
    nand02 ix3142 (.Y (nx3141), .A0 (currentPage_23__12), .A1 (layerType)) ;
    nand02 ix3144 (.Y (nx3143), .A0 (outMuls_23__12), .A1 (nx5208)) ;
    nand02 ix447 (.Y (addersInputs_23__13), .A0 (nx3147), .A1 (nx3149)) ;
    nand02 ix3148 (.Y (nx3147), .A0 (currentPage_23__13), .A1 (layerType)) ;
    nand02 ix3150 (.Y (nx3149), .A0 (outMuls_23__13), .A1 (nx5208)) ;
    nand02 ix455 (.Y (addersInputs_23__14), .A0 (nx3153), .A1 (nx3155)) ;
    nand02 ix3154 (.Y (nx3153), .A0 (currentPage_23__14), .A1 (layerType)) ;
    nand02 ix3156 (.Y (nx3155), .A0 (outMuls_23__14), .A1 (nx5208)) ;
    nand02 ix463 (.Y (addersInputs_23__15), .A0 (nx3159), .A1 (nx3161)) ;
    nand02 ix3160 (.Y (nx3159), .A0 (currentPage_23__15), .A1 (layerType)) ;
    nand02 ix3162 (.Y (nx3161), .A0 (outMuls_23__15), .A1 (nx5208)) ;
    nand02 ix471 (.Y (addersInputs_22__0), .A0 (nx3165), .A1 (nx3167)) ;
    nand02 ix3166 (.Y (nx3165), .A0 (currentPage_22__0), .A1 (layerType)) ;
    nand02 ix3168 (.Y (nx3167), .A0 (outMuls_22__0), .A1 (nx5208)) ;
    nand02 ix479 (.Y (addersInputs_22__1), .A0 (nx3171), .A1 (nx3173)) ;
    nand02 ix3172 (.Y (nx3171), .A0 (currentPage_22__1), .A1 (layerType)) ;
    nand02 ix3174 (.Y (nx3173), .A0 (outMuls_22__1), .A1 (nx5208)) ;
    nand02 ix487 (.Y (addersInputs_22__2), .A0 (nx3177), .A1 (nx3179)) ;
    nand02 ix3178 (.Y (nx3177), .A0 (currentPage_22__2), .A1 (layerType)) ;
    nand02 ix3180 (.Y (nx3179), .A0 (outMuls_22__2), .A1 (nx5208)) ;
    nand02 ix495 (.Y (addersInputs_22__3), .A0 (nx3183), .A1 (nx3185)) ;
    nand02 ix3184 (.Y (nx3183), .A0 (currentPage_22__3), .A1 (layerType)) ;
    nand02 ix3186 (.Y (nx3185), .A0 (outMuls_22__3), .A1 (nx5210)) ;
    nand02 ix503 (.Y (addersInputs_22__4), .A0 (nx3189), .A1 (nx3191)) ;
    nand02 ix3190 (.Y (nx3189), .A0 (currentPage_22__4), .A1 (layerType)) ;
    nand02 ix3192 (.Y (nx3191), .A0 (outMuls_22__4), .A1 (nx5210)) ;
    nand02 ix511 (.Y (addersInputs_22__5), .A0 (nx3195), .A1 (nx3197)) ;
    nand02 ix3196 (.Y (nx3195), .A0 (currentPage_22__5), .A1 (layerType)) ;
    nand02 ix3198 (.Y (nx3197), .A0 (outMuls_22__5), .A1 (nx5210)) ;
    nand02 ix519 (.Y (addersInputs_22__6), .A0 (nx3201), .A1 (nx3203)) ;
    nand02 ix3202 (.Y (nx3201), .A0 (currentPage_22__6), .A1 (layerType)) ;
    nand02 ix3204 (.Y (nx3203), .A0 (outMuls_22__6), .A1 (nx5210)) ;
    nand02 ix527 (.Y (addersInputs_22__7), .A0 (nx3207), .A1 (nx3209)) ;
    nand02 ix3208 (.Y (nx3207), .A0 (currentPage_22__7), .A1 (layerType)) ;
    nand02 ix3210 (.Y (nx3209), .A0 (outMuls_22__7), .A1 (nx5210)) ;
    nand02 ix535 (.Y (addersInputs_22__8), .A0 (nx3213), .A1 (nx3215)) ;
    nand02 ix3214 (.Y (nx3213), .A0 (currentPage_22__8), .A1 (layerType)) ;
    nand02 ix3216 (.Y (nx3215), .A0 (outMuls_22__8), .A1 (nx5210)) ;
    nand02 ix543 (.Y (addersInputs_22__9), .A0 (nx3219), .A1 (nx3221)) ;
    nand02 ix3220 (.Y (nx3219), .A0 (currentPage_22__9), .A1 (layerType)) ;
    nand02 ix3222 (.Y (nx3221), .A0 (outMuls_22__9), .A1 (nx5210)) ;
    nand02 ix551 (.Y (addersInputs_22__10), .A0 (nx3225), .A1 (nx3227)) ;
    nand02 ix3226 (.Y (nx3225), .A0 (currentPage_22__10), .A1 (layerType)) ;
    nand02 ix3228 (.Y (nx3227), .A0 (outMuls_22__10), .A1 (nx5212)) ;
    nand02 ix559 (.Y (addersInputs_22__11), .A0 (nx3231), .A1 (nx3233)) ;
    nand02 ix3232 (.Y (nx3231), .A0 (currentPage_22__11), .A1 (layerType)) ;
    nand02 ix3234 (.Y (nx3233), .A0 (outMuls_22__11), .A1 (nx5212)) ;
    nand02 ix567 (.Y (addersInputs_22__12), .A0 (nx3237), .A1 (nx3239)) ;
    nand02 ix3238 (.Y (nx3237), .A0 (currentPage_22__12), .A1 (layerType)) ;
    nand02 ix3240 (.Y (nx3239), .A0 (outMuls_22__12), .A1 (nx5212)) ;
    nand02 ix575 (.Y (addersInputs_22__13), .A0 (nx3243), .A1 (nx3245)) ;
    nand02 ix3244 (.Y (nx3243), .A0 (currentPage_22__13), .A1 (layerType)) ;
    nand02 ix3246 (.Y (nx3245), .A0 (outMuls_22__13), .A1 (nx5212)) ;
    nand02 ix583 (.Y (addersInputs_22__14), .A0 (nx3249), .A1 (nx3251)) ;
    nand02 ix3250 (.Y (nx3249), .A0 (currentPage_22__14), .A1 (layerType)) ;
    nand02 ix3252 (.Y (nx3251), .A0 (outMuls_22__14), .A1 (nx5212)) ;
    nand02 ix591 (.Y (addersInputs_22__15), .A0 (nx3255), .A1 (nx3257)) ;
    nand02 ix3256 (.Y (nx3255), .A0 (currentPage_22__15), .A1 (layerType)) ;
    nand02 ix3258 (.Y (nx3257), .A0 (outMuls_22__15), .A1 (nx5212)) ;
    nand02 ix599 (.Y (addersInputs_21__0), .A0 (nx3261), .A1 (nx3263)) ;
    nand02 ix3262 (.Y (nx3261), .A0 (currentPage_21__0), .A1 (layerType)) ;
    nand02 ix3264 (.Y (nx3263), .A0 (outMuls_21__0), .A1 (nx5212)) ;
    nand02 ix607 (.Y (addersInputs_21__1), .A0 (nx3267), .A1 (nx3269)) ;
    nand02 ix3268 (.Y (nx3267), .A0 (currentPage_21__1), .A1 (layerType)) ;
    nand02 ix3270 (.Y (nx3269), .A0 (outMuls_21__1), .A1 (nx5214)) ;
    nand02 ix615 (.Y (addersInputs_21__2), .A0 (nx3273), .A1 (nx3275)) ;
    nand02 ix3274 (.Y (nx3273), .A0 (currentPage_21__2), .A1 (layerType)) ;
    nand02 ix3276 (.Y (nx3275), .A0 (outMuls_21__2), .A1 (nx5214)) ;
    nand02 ix623 (.Y (addersInputs_21__3), .A0 (nx3279), .A1 (nx3281)) ;
    nand02 ix3280 (.Y (nx3279), .A0 (currentPage_21__3), .A1 (layerType)) ;
    nand02 ix3282 (.Y (nx3281), .A0 (outMuls_21__3), .A1 (nx5214)) ;
    nand02 ix631 (.Y (addersInputs_21__4), .A0 (nx3285), .A1 (nx3287)) ;
    nand02 ix3286 (.Y (nx3285), .A0 (currentPage_21__4), .A1 (layerType)) ;
    nand02 ix3288 (.Y (nx3287), .A0 (outMuls_21__4), .A1 (nx5214)) ;
    nand02 ix639 (.Y (addersInputs_21__5), .A0 (nx3291), .A1 (nx3293)) ;
    nand02 ix3292 (.Y (nx3291), .A0 (currentPage_21__5), .A1 (layerType)) ;
    nand02 ix3294 (.Y (nx3293), .A0 (outMuls_21__5), .A1 (nx5214)) ;
    nand02 ix647 (.Y (addersInputs_21__6), .A0 (nx3297), .A1 (nx3299)) ;
    nand02 ix3298 (.Y (nx3297), .A0 (currentPage_21__6), .A1 (layerType)) ;
    nand02 ix3300 (.Y (nx3299), .A0 (outMuls_21__6), .A1 (nx5214)) ;
    nand02 ix655 (.Y (addersInputs_21__7), .A0 (nx3303), .A1 (nx3305)) ;
    nand02 ix3304 (.Y (nx3303), .A0 (currentPage_21__7), .A1 (layerType)) ;
    nand02 ix3306 (.Y (nx3305), .A0 (outMuls_21__7), .A1 (nx5214)) ;
    nand02 ix663 (.Y (addersInputs_21__8), .A0 (nx3309), .A1 (nx3311)) ;
    nand02 ix3310 (.Y (nx3309), .A0 (currentPage_21__8), .A1 (layerType)) ;
    nand02 ix3312 (.Y (nx3311), .A0 (outMuls_21__8), .A1 (nx5216)) ;
    nand02 ix671 (.Y (addersInputs_21__9), .A0 (nx3315), .A1 (nx3317)) ;
    nand02 ix3316 (.Y (nx3315), .A0 (currentPage_21__9), .A1 (layerType)) ;
    nand02 ix3318 (.Y (nx3317), .A0 (outMuls_21__9), .A1 (nx5216)) ;
    nand02 ix679 (.Y (addersInputs_21__10), .A0 (nx3321), .A1 (nx3323)) ;
    nand02 ix3322 (.Y (nx3321), .A0 (currentPage_21__10), .A1 (layerType)) ;
    nand02 ix3324 (.Y (nx3323), .A0 (outMuls_21__10), .A1 (nx5216)) ;
    nand02 ix687 (.Y (addersInputs_21__11), .A0 (nx3327), .A1 (nx3329)) ;
    nand02 ix3328 (.Y (nx3327), .A0 (currentPage_21__11), .A1 (layerType)) ;
    nand02 ix3330 (.Y (nx3329), .A0 (outMuls_21__11), .A1 (nx5216)) ;
    nand02 ix695 (.Y (addersInputs_21__12), .A0 (nx3333), .A1 (nx3335)) ;
    nand02 ix3334 (.Y (nx3333), .A0 (currentPage_21__12), .A1 (layerType)) ;
    nand02 ix3336 (.Y (nx3335), .A0 (outMuls_21__12), .A1 (nx5216)) ;
    nand02 ix703 (.Y (addersInputs_21__13), .A0 (nx3339), .A1 (nx3341)) ;
    nand02 ix3340 (.Y (nx3339), .A0 (currentPage_21__13), .A1 (layerType)) ;
    nand02 ix3342 (.Y (nx3341), .A0 (outMuls_21__13), .A1 (nx5216)) ;
    nand02 ix711 (.Y (addersInputs_21__14), .A0 (nx3345), .A1 (nx3347)) ;
    nand02 ix3346 (.Y (nx3345), .A0 (currentPage_21__14), .A1 (layerType)) ;
    nand02 ix3348 (.Y (nx3347), .A0 (outMuls_21__14), .A1 (nx5216)) ;
    nand02 ix719 (.Y (addersInputs_21__15), .A0 (nx3351), .A1 (nx3353)) ;
    nand02 ix3352 (.Y (nx3351), .A0 (currentPage_21__15), .A1 (layerType)) ;
    nand02 ix3354 (.Y (nx3353), .A0 (outMuls_21__15), .A1 (nx5218)) ;
    nand02 ix727 (.Y (addersInputs_20__0), .A0 (nx3357), .A1 (nx3359)) ;
    nand02 ix3358 (.Y (nx3357), .A0 (currentPage_20__0), .A1 (layerType)) ;
    nand02 ix3360 (.Y (nx3359), .A0 (outMuls_20__0), .A1 (nx5218)) ;
    nand02 ix735 (.Y (addersInputs_20__1), .A0 (nx3363), .A1 (nx3365)) ;
    nand02 ix3364 (.Y (nx3363), .A0 (currentPage_20__1), .A1 (layerType)) ;
    nand02 ix3366 (.Y (nx3365), .A0 (outMuls_20__1), .A1 (nx5218)) ;
    nand02 ix743 (.Y (addersInputs_20__2), .A0 (nx3369), .A1 (nx3371)) ;
    nand02 ix3370 (.Y (nx3369), .A0 (currentPage_20__2), .A1 (layerType)) ;
    nand02 ix3372 (.Y (nx3371), .A0 (outMuls_20__2), .A1 (nx5218)) ;
    nand02 ix751 (.Y (addersInputs_20__3), .A0 (nx3375), .A1 (nx3377)) ;
    nand02 ix3376 (.Y (nx3375), .A0 (currentPage_20__3), .A1 (layerType)) ;
    nand02 ix3378 (.Y (nx3377), .A0 (outMuls_20__3), .A1 (nx5218)) ;
    nand02 ix759 (.Y (addersInputs_20__4), .A0 (nx3381), .A1 (nx3383)) ;
    nand02 ix3382 (.Y (nx3381), .A0 (currentPage_20__4), .A1 (layerType)) ;
    nand02 ix3384 (.Y (nx3383), .A0 (outMuls_20__4), .A1 (nx5218)) ;
    nand02 ix767 (.Y (addersInputs_20__5), .A0 (nx3387), .A1 (nx3389)) ;
    nand02 ix3388 (.Y (nx3387), .A0 (currentPage_20__5), .A1 (layerType)) ;
    nand02 ix3390 (.Y (nx3389), .A0 (outMuls_20__5), .A1 (nx5218)) ;
    nand02 ix775 (.Y (addersInputs_20__6), .A0 (nx3393), .A1 (nx3395)) ;
    nand02 ix3394 (.Y (nx3393), .A0 (currentPage_20__6), .A1 (layerType)) ;
    nand02 ix3396 (.Y (nx3395), .A0 (outMuls_20__6), .A1 (nx5220)) ;
    nand02 ix783 (.Y (addersInputs_20__7), .A0 (nx3399), .A1 (nx3401)) ;
    nand02 ix3400 (.Y (nx3399), .A0 (currentPage_20__7), .A1 (layerType)) ;
    nand02 ix3402 (.Y (nx3401), .A0 (outMuls_20__7), .A1 (nx5220)) ;
    nand02 ix791 (.Y (addersInputs_20__8), .A0 (nx3405), .A1 (nx3407)) ;
    nand02 ix3406 (.Y (nx3405), .A0 (currentPage_20__8), .A1 (layerType)) ;
    nand02 ix3408 (.Y (nx3407), .A0 (outMuls_20__8), .A1 (nx5220)) ;
    nand02 ix799 (.Y (addersInputs_20__9), .A0 (nx3411), .A1 (nx3413)) ;
    nand02 ix3412 (.Y (nx3411), .A0 (currentPage_20__9), .A1 (layerType)) ;
    nand02 ix3414 (.Y (nx3413), .A0 (outMuls_20__9), .A1 (nx5220)) ;
    nand02 ix807 (.Y (addersInputs_20__10), .A0 (nx3417), .A1 (nx3419)) ;
    nand02 ix3418 (.Y (nx3417), .A0 (currentPage_20__10), .A1 (layerType)) ;
    nand02 ix3420 (.Y (nx3419), .A0 (outMuls_20__10), .A1 (nx5220)) ;
    nand02 ix815 (.Y (addersInputs_20__11), .A0 (nx3423), .A1 (nx3425)) ;
    nand02 ix3424 (.Y (nx3423), .A0 (currentPage_20__11), .A1 (layerType)) ;
    nand02 ix3426 (.Y (nx3425), .A0 (outMuls_20__11), .A1 (nx5220)) ;
    nand02 ix823 (.Y (addersInputs_20__12), .A0 (nx3429), .A1 (nx3431)) ;
    nand02 ix3430 (.Y (nx3429), .A0 (currentPage_20__12), .A1 (layerType)) ;
    nand02 ix3432 (.Y (nx3431), .A0 (outMuls_20__12), .A1 (nx5220)) ;
    nand02 ix831 (.Y (addersInputs_20__13), .A0 (nx3435), .A1 (nx3437)) ;
    nand02 ix3436 (.Y (nx3435), .A0 (currentPage_20__13), .A1 (layerType)) ;
    nand02 ix3438 (.Y (nx3437), .A0 (outMuls_20__13), .A1 (nx5222)) ;
    nand02 ix839 (.Y (addersInputs_20__14), .A0 (nx3441), .A1 (nx3443)) ;
    nand02 ix3442 (.Y (nx3441), .A0 (currentPage_20__14), .A1 (layerType)) ;
    nand02 ix3444 (.Y (nx3443), .A0 (outMuls_20__14), .A1 (nx5222)) ;
    nand02 ix847 (.Y (addersInputs_20__15), .A0 (nx3447), .A1 (nx3449)) ;
    nand02 ix3448 (.Y (nx3447), .A0 (currentPage_20__15), .A1 (layerType)) ;
    nand02 ix3450 (.Y (nx3449), .A0 (outMuls_20__15), .A1 (nx5222)) ;
    nand02 ix855 (.Y (addersInputs_19__0), .A0 (nx3453), .A1 (nx3455)) ;
    nand02 ix3454 (.Y (nx3453), .A0 (currentPage_19__0), .A1 (layerType)) ;
    nand02 ix3456 (.Y (nx3455), .A0 (outMuls_19__0), .A1 (nx5222)) ;
    nand02 ix863 (.Y (addersInputs_19__1), .A0 (nx3459), .A1 (nx3461)) ;
    nand02 ix3460 (.Y (nx3459), .A0 (currentPage_19__1), .A1 (layerType)) ;
    nand02 ix3462 (.Y (nx3461), .A0 (outMuls_19__1), .A1 (nx5222)) ;
    nand02 ix871 (.Y (addersInputs_19__2), .A0 (nx3465), .A1 (nx3467)) ;
    nand02 ix3466 (.Y (nx3465), .A0 (currentPage_19__2), .A1 (layerType)) ;
    nand02 ix3468 (.Y (nx3467), .A0 (outMuls_19__2), .A1 (nx5222)) ;
    nand02 ix879 (.Y (addersInputs_19__3), .A0 (nx3471), .A1 (nx3473)) ;
    nand02 ix3472 (.Y (nx3471), .A0 (currentPage_19__3), .A1 (layerType)) ;
    nand02 ix3474 (.Y (nx3473), .A0 (outMuls_19__3), .A1 (nx5222)) ;
    nand02 ix887 (.Y (addersInputs_19__4), .A0 (nx3477), .A1 (nx3479)) ;
    nand02 ix3478 (.Y (nx3477), .A0 (currentPage_19__4), .A1 (layerType)) ;
    nand02 ix3480 (.Y (nx3479), .A0 (outMuls_19__4), .A1 (nx5224)) ;
    nand02 ix895 (.Y (addersInputs_19__5), .A0 (nx3483), .A1 (nx3485)) ;
    nand02 ix3484 (.Y (nx3483), .A0 (currentPage_19__5), .A1 (layerType)) ;
    nand02 ix3486 (.Y (nx3485), .A0 (outMuls_19__5), .A1 (nx5224)) ;
    nand02 ix903 (.Y (addersInputs_19__6), .A0 (nx3488), .A1 (nx3490)) ;
    nand02 ix3489 (.Y (nx3488), .A0 (currentPage_19__6), .A1 (layerType)) ;
    nand02 ix3491 (.Y (nx3490), .A0 (outMuls_19__6), .A1 (nx5224)) ;
    nand02 ix911 (.Y (addersInputs_19__7), .A0 (nx3493), .A1 (nx3495)) ;
    nand02 ix3494 (.Y (nx3493), .A0 (currentPage_19__7), .A1 (layerType)) ;
    nand02 ix3496 (.Y (nx3495), .A0 (outMuls_19__7), .A1 (nx5224)) ;
    nand02 ix919 (.Y (addersInputs_19__8), .A0 (nx3498), .A1 (nx3500)) ;
    nand02 ix3499 (.Y (nx3498), .A0 (currentPage_19__8), .A1 (layerType)) ;
    nand02 ix3501 (.Y (nx3500), .A0 (outMuls_19__8), .A1 (nx5224)) ;
    nand02 ix927 (.Y (addersInputs_19__9), .A0 (nx3503), .A1 (nx3505)) ;
    nand02 ix3504 (.Y (nx3503), .A0 (currentPage_19__9), .A1 (layerType)) ;
    nand02 ix3506 (.Y (nx3505), .A0 (outMuls_19__9), .A1 (nx5224)) ;
    nand02 ix935 (.Y (addersInputs_19__10), .A0 (nx3508), .A1 (nx3510)) ;
    nand02 ix3509 (.Y (nx3508), .A0 (currentPage_19__10), .A1 (layerType)) ;
    nand02 ix3511 (.Y (nx3510), .A0 (outMuls_19__10), .A1 (nx5224)) ;
    nand02 ix943 (.Y (addersInputs_19__11), .A0 (nx3513), .A1 (nx3515)) ;
    nand02 ix3514 (.Y (nx3513), .A0 (currentPage_19__11), .A1 (layerType)) ;
    nand02 ix3516 (.Y (nx3515), .A0 (outMuls_19__11), .A1 (nx5226)) ;
    nand02 ix951 (.Y (addersInputs_19__12), .A0 (nx3518), .A1 (nx3520)) ;
    nand02 ix3519 (.Y (nx3518), .A0 (currentPage_19__12), .A1 (layerType)) ;
    nand02 ix3521 (.Y (nx3520), .A0 (outMuls_19__12), .A1 (nx5226)) ;
    nand02 ix959 (.Y (addersInputs_19__13), .A0 (nx3523), .A1 (nx3525)) ;
    nand02 ix3524 (.Y (nx3523), .A0 (currentPage_19__13), .A1 (layerType)) ;
    nand02 ix3526 (.Y (nx3525), .A0 (outMuls_19__13), .A1 (nx5226)) ;
    nand02 ix967 (.Y (addersInputs_19__14), .A0 (nx3528), .A1 (nx3530)) ;
    nand02 ix3529 (.Y (nx3528), .A0 (currentPage_19__14), .A1 (layerType)) ;
    nand02 ix3531 (.Y (nx3530), .A0 (outMuls_19__14), .A1 (nx5226)) ;
    nand02 ix975 (.Y (addersInputs_19__15), .A0 (nx3533), .A1 (nx3535)) ;
    nand02 ix3534 (.Y (nx3533), .A0 (currentPage_19__15), .A1 (layerType)) ;
    nand02 ix3536 (.Y (nx3535), .A0 (outMuls_19__15), .A1 (nx5226)) ;
    nand02 ix983 (.Y (addersInputs_18__0), .A0 (nx3538), .A1 (nx3540)) ;
    nand02 ix3539 (.Y (nx3538), .A0 (currentPage_18__0), .A1 (layerType)) ;
    nand02 ix3541 (.Y (nx3540), .A0 (outMuls_18__0), .A1 (nx5226)) ;
    nand02 ix991 (.Y (addersInputs_18__1), .A0 (nx3543), .A1 (nx3545)) ;
    nand02 ix3544 (.Y (nx3543), .A0 (currentPage_18__1), .A1 (layerType)) ;
    nand02 ix3546 (.Y (nx3545), .A0 (outMuls_18__1), .A1 (nx5226)) ;
    nand02 ix999 (.Y (addersInputs_18__2), .A0 (nx3548), .A1 (nx3550)) ;
    nand02 ix3549 (.Y (nx3548), .A0 (currentPage_18__2), .A1 (layerType)) ;
    nand02 ix3551 (.Y (nx3550), .A0 (outMuls_18__2), .A1 (nx5228)) ;
    nand02 ix1007 (.Y (addersInputs_18__3), .A0 (nx3553), .A1 (nx3555)) ;
    nand02 ix3554 (.Y (nx3553), .A0 (currentPage_18__3), .A1 (layerType)) ;
    nand02 ix3556 (.Y (nx3555), .A0 (outMuls_18__3), .A1 (nx5228)) ;
    nand02 ix1015 (.Y (addersInputs_18__4), .A0 (nx3558), .A1 (nx3560)) ;
    nand02 ix3559 (.Y (nx3558), .A0 (currentPage_18__4), .A1 (layerType)) ;
    nand02 ix3561 (.Y (nx3560), .A0 (outMuls_18__4), .A1 (nx5228)) ;
    nand02 ix1023 (.Y (addersInputs_18__5), .A0 (nx3563), .A1 (nx3565)) ;
    nand02 ix3564 (.Y (nx3563), .A0 (currentPage_18__5), .A1 (layerType)) ;
    nand02 ix3566 (.Y (nx3565), .A0 (outMuls_18__5), .A1 (nx5228)) ;
    nand02 ix1031 (.Y (addersInputs_18__6), .A0 (nx3568), .A1 (nx3570)) ;
    nand02 ix3569 (.Y (nx3568), .A0 (currentPage_18__6), .A1 (layerType)) ;
    nand02 ix3571 (.Y (nx3570), .A0 (outMuls_18__6), .A1 (nx5228)) ;
    nand02 ix1039 (.Y (addersInputs_18__7), .A0 (nx3573), .A1 (nx3575)) ;
    nand02 ix3574 (.Y (nx3573), .A0 (currentPage_18__7), .A1 (layerType)) ;
    nand02 ix3576 (.Y (nx3575), .A0 (outMuls_18__7), .A1 (nx5228)) ;
    nand02 ix1047 (.Y (addersInputs_18__8), .A0 (nx3578), .A1 (nx3580)) ;
    nand02 ix3579 (.Y (nx3578), .A0 (currentPage_18__8), .A1 (layerType)) ;
    nand02 ix3581 (.Y (nx3580), .A0 (outMuls_18__8), .A1 (nx5228)) ;
    nand02 ix1055 (.Y (addersInputs_18__9), .A0 (nx3583), .A1 (nx3585)) ;
    nand02 ix3584 (.Y (nx3583), .A0 (currentPage_18__9), .A1 (layerType)) ;
    nand02 ix3586 (.Y (nx3585), .A0 (outMuls_18__9), .A1 (nx5230)) ;
    nand02 ix1063 (.Y (addersInputs_18__10), .A0 (nx3588), .A1 (nx3590)) ;
    nand02 ix3589 (.Y (nx3588), .A0 (currentPage_18__10), .A1 (layerType)) ;
    nand02 ix3591 (.Y (nx3590), .A0 (outMuls_18__10), .A1 (nx5230)) ;
    nand02 ix1071 (.Y (addersInputs_18__11), .A0 (nx3593), .A1 (nx3595)) ;
    nand02 ix3594 (.Y (nx3593), .A0 (currentPage_18__11), .A1 (layerType)) ;
    nand02 ix3596 (.Y (nx3595), .A0 (outMuls_18__11), .A1 (nx5230)) ;
    nand02 ix1079 (.Y (addersInputs_18__12), .A0 (nx3598), .A1 (nx3600)) ;
    nand02 ix3599 (.Y (nx3598), .A0 (currentPage_18__12), .A1 (layerType)) ;
    nand02 ix3601 (.Y (nx3600), .A0 (outMuls_18__12), .A1 (nx5230)) ;
    nand02 ix1087 (.Y (addersInputs_18__13), .A0 (nx3603), .A1 (nx3605)) ;
    nand02 ix3604 (.Y (nx3603), .A0 (currentPage_18__13), .A1 (layerType)) ;
    nand02 ix3606 (.Y (nx3605), .A0 (outMuls_18__13), .A1 (nx5230)) ;
    nand02 ix1095 (.Y (addersInputs_18__14), .A0 (nx3608), .A1 (nx3610)) ;
    nand02 ix3609 (.Y (nx3608), .A0 (currentPage_18__14), .A1 (layerType)) ;
    nand02 ix3611 (.Y (nx3610), .A0 (outMuls_18__14), .A1 (nx5230)) ;
    nand02 ix1103 (.Y (addersInputs_18__15), .A0 (nx3613), .A1 (nx3615)) ;
    nand02 ix3614 (.Y (nx3613), .A0 (currentPage_18__15), .A1 (layerType)) ;
    nand02 ix3616 (.Y (nx3615), .A0 (outMuls_18__15), .A1 (nx5230)) ;
    nand02 ix1111 (.Y (addersInputs_17__0), .A0 (nx3618), .A1 (nx3620)) ;
    nand02 ix3619 (.Y (nx3618), .A0 (currentPage_17__0), .A1 (layerType)) ;
    nand02 ix3621 (.Y (nx3620), .A0 (outMuls_17__0), .A1 (nx5232)) ;
    nand02 ix1119 (.Y (addersInputs_17__1), .A0 (nx3623), .A1 (nx3625)) ;
    nand02 ix3624 (.Y (nx3623), .A0 (currentPage_17__1), .A1 (layerType)) ;
    nand02 ix3626 (.Y (nx3625), .A0 (outMuls_17__1), .A1 (nx5232)) ;
    nand02 ix1127 (.Y (addersInputs_17__2), .A0 (nx3628), .A1 (nx3630)) ;
    nand02 ix3629 (.Y (nx3628), .A0 (currentPage_17__2), .A1 (layerType)) ;
    nand02 ix3631 (.Y (nx3630), .A0 (outMuls_17__2), .A1 (nx5232)) ;
    nand02 ix1135 (.Y (addersInputs_17__3), .A0 (nx3633), .A1 (nx3635)) ;
    nand02 ix3634 (.Y (nx3633), .A0 (currentPage_17__3), .A1 (layerType)) ;
    nand02 ix3636 (.Y (nx3635), .A0 (outMuls_17__3), .A1 (nx5232)) ;
    nand02 ix1143 (.Y (addersInputs_17__4), .A0 (nx3638), .A1 (nx3640)) ;
    nand02 ix3639 (.Y (nx3638), .A0 (currentPage_17__4), .A1 (layerType)) ;
    nand02 ix3641 (.Y (nx3640), .A0 (outMuls_17__4), .A1 (nx5232)) ;
    nand02 ix1151 (.Y (addersInputs_17__5), .A0 (nx3643), .A1 (nx3645)) ;
    nand02 ix3644 (.Y (nx3643), .A0 (currentPage_17__5), .A1 (layerType)) ;
    nand02 ix3646 (.Y (nx3645), .A0 (outMuls_17__5), .A1 (nx5232)) ;
    nand02 ix1159 (.Y (addersInputs_17__6), .A0 (nx3648), .A1 (nx3650)) ;
    nand02 ix3649 (.Y (nx3648), .A0 (currentPage_17__6), .A1 (layerType)) ;
    nand02 ix3651 (.Y (nx3650), .A0 (outMuls_17__6), .A1 (nx5232)) ;
    nand02 ix1167 (.Y (addersInputs_17__7), .A0 (nx3653), .A1 (nx3655)) ;
    nand02 ix3654 (.Y (nx3653), .A0 (currentPage_17__7), .A1 (layerType)) ;
    nand02 ix3656 (.Y (nx3655), .A0 (outMuls_17__7), .A1 (nx5234)) ;
    nand02 ix1175 (.Y (addersInputs_17__8), .A0 (nx3658), .A1 (nx3660)) ;
    nand02 ix3659 (.Y (nx3658), .A0 (currentPage_17__8), .A1 (layerType)) ;
    nand02 ix3661 (.Y (nx3660), .A0 (outMuls_17__8), .A1 (nx5234)) ;
    nand02 ix1183 (.Y (addersInputs_17__9), .A0 (nx3663), .A1 (nx3665)) ;
    nand02 ix3664 (.Y (nx3663), .A0 (currentPage_17__9), .A1 (layerType)) ;
    nand02 ix3666 (.Y (nx3665), .A0 (outMuls_17__9), .A1 (nx5234)) ;
    nand02 ix1191 (.Y (addersInputs_17__10), .A0 (nx3668), .A1 (nx3670)) ;
    nand02 ix3669 (.Y (nx3668), .A0 (currentPage_17__10), .A1 (layerType)) ;
    nand02 ix3671 (.Y (nx3670), .A0 (outMuls_17__10), .A1 (nx5234)) ;
    nand02 ix1199 (.Y (addersInputs_17__11), .A0 (nx3673), .A1 (nx3675)) ;
    nand02 ix3674 (.Y (nx3673), .A0 (currentPage_17__11), .A1 (layerType)) ;
    nand02 ix3676 (.Y (nx3675), .A0 (outMuls_17__11), .A1 (nx5234)) ;
    nand02 ix1207 (.Y (addersInputs_17__12), .A0 (nx3678), .A1 (nx3680)) ;
    nand02 ix3679 (.Y (nx3678), .A0 (currentPage_17__12), .A1 (layerType)) ;
    nand02 ix3681 (.Y (nx3680), .A0 (outMuls_17__12), .A1 (nx5234)) ;
    nand02 ix1215 (.Y (addersInputs_17__13), .A0 (nx3683), .A1 (nx3685)) ;
    nand02 ix3684 (.Y (nx3683), .A0 (currentPage_17__13), .A1 (layerType)) ;
    nand02 ix3686 (.Y (nx3685), .A0 (outMuls_17__13), .A1 (nx5234)) ;
    nand02 ix1223 (.Y (addersInputs_17__14), .A0 (nx3688), .A1 (nx3690)) ;
    nand02 ix3689 (.Y (nx3688), .A0 (currentPage_17__14), .A1 (layerType)) ;
    nand02 ix3691 (.Y (nx3690), .A0 (outMuls_17__14), .A1 (nx5236)) ;
    nand02 ix1231 (.Y (addersInputs_17__15), .A0 (nx3693), .A1 (nx3695)) ;
    nand02 ix3694 (.Y (nx3693), .A0 (currentPage_17__15), .A1 (layerType)) ;
    nand02 ix3696 (.Y (nx3695), .A0 (outMuls_17__15), .A1 (nx5236)) ;
    nand02 ix1239 (.Y (addersInputs_16__0), .A0 (nx3698), .A1 (nx3700)) ;
    nand02 ix3699 (.Y (nx3698), .A0 (currentPage_16__0), .A1 (layerType)) ;
    nand02 ix3701 (.Y (nx3700), .A0 (outMuls_16__0), .A1 (nx5236)) ;
    nand02 ix1247 (.Y (addersInputs_16__1), .A0 (nx3703), .A1 (nx3705)) ;
    nand02 ix3704 (.Y (nx3703), .A0 (currentPage_16__1), .A1 (layerType)) ;
    nand02 ix3706 (.Y (nx3705), .A0 (outMuls_16__1), .A1 (nx5236)) ;
    nand02 ix1255 (.Y (addersInputs_16__2), .A0 (nx3708), .A1 (nx3710)) ;
    nand02 ix3709 (.Y (nx3708), .A0 (currentPage_16__2), .A1 (layerType)) ;
    nand02 ix3711 (.Y (nx3710), .A0 (outMuls_16__2), .A1 (nx5236)) ;
    nand02 ix1263 (.Y (addersInputs_16__3), .A0 (nx3713), .A1 (nx3715)) ;
    nand02 ix3714 (.Y (nx3713), .A0 (currentPage_16__3), .A1 (layerType)) ;
    nand02 ix3716 (.Y (nx3715), .A0 (outMuls_16__3), .A1 (nx5236)) ;
    nand02 ix1271 (.Y (addersInputs_16__4), .A0 (nx3718), .A1 (nx3720)) ;
    nand02 ix3719 (.Y (nx3718), .A0 (currentPage_16__4), .A1 (layerType)) ;
    nand02 ix3721 (.Y (nx3720), .A0 (outMuls_16__4), .A1 (nx5236)) ;
    nand02 ix1279 (.Y (addersInputs_16__5), .A0 (nx3723), .A1 (nx3725)) ;
    nand02 ix3724 (.Y (nx3723), .A0 (currentPage_16__5), .A1 (layerType)) ;
    nand02 ix3726 (.Y (nx3725), .A0 (outMuls_16__5), .A1 (nx5238)) ;
    nand02 ix1287 (.Y (addersInputs_16__6), .A0 (nx3728), .A1 (nx3730)) ;
    nand02 ix3729 (.Y (nx3728), .A0 (currentPage_16__6), .A1 (layerType)) ;
    nand02 ix3731 (.Y (nx3730), .A0 (outMuls_16__6), .A1 (nx5238)) ;
    nand02 ix1295 (.Y (addersInputs_16__7), .A0 (nx3733), .A1 (nx3735)) ;
    nand02 ix3734 (.Y (nx3733), .A0 (currentPage_16__7), .A1 (layerType)) ;
    nand02 ix3736 (.Y (nx3735), .A0 (outMuls_16__7), .A1 (nx5238)) ;
    nand02 ix1303 (.Y (addersInputs_16__8), .A0 (nx3738), .A1 (nx3740)) ;
    nand02 ix3739 (.Y (nx3738), .A0 (currentPage_16__8), .A1 (layerType)) ;
    nand02 ix3741 (.Y (nx3740), .A0 (outMuls_16__8), .A1 (nx5238)) ;
    nand02 ix1311 (.Y (addersInputs_16__9), .A0 (nx3743), .A1 (nx3745)) ;
    nand02 ix3744 (.Y (nx3743), .A0 (currentPage_16__9), .A1 (layerType)) ;
    nand02 ix3746 (.Y (nx3745), .A0 (outMuls_16__9), .A1 (nx5238)) ;
    nand02 ix1319 (.Y (addersInputs_16__10), .A0 (nx3748), .A1 (nx3750)) ;
    nand02 ix3749 (.Y (nx3748), .A0 (currentPage_16__10), .A1 (layerType)) ;
    nand02 ix3751 (.Y (nx3750), .A0 (outMuls_16__10), .A1 (nx5238)) ;
    nand02 ix1327 (.Y (addersInputs_16__11), .A0 (nx3753), .A1 (nx3755)) ;
    nand02 ix3754 (.Y (nx3753), .A0 (currentPage_16__11), .A1 (layerType)) ;
    nand02 ix3756 (.Y (nx3755), .A0 (outMuls_16__11), .A1 (nx5238)) ;
    nand02 ix1335 (.Y (addersInputs_16__12), .A0 (nx3758), .A1 (nx3760)) ;
    nand02 ix3759 (.Y (nx3758), .A0 (currentPage_16__12), .A1 (layerType)) ;
    nand02 ix3761 (.Y (nx3760), .A0 (outMuls_16__12), .A1 (nx5240)) ;
    nand02 ix1343 (.Y (addersInputs_16__13), .A0 (nx3763), .A1 (nx3765)) ;
    nand02 ix3764 (.Y (nx3763), .A0 (currentPage_16__13), .A1 (layerType)) ;
    nand02 ix3766 (.Y (nx3765), .A0 (outMuls_16__13), .A1 (nx5240)) ;
    nand02 ix1351 (.Y (addersInputs_16__14), .A0 (nx3768), .A1 (nx3770)) ;
    nand02 ix3769 (.Y (nx3768), .A0 (currentPage_16__14), .A1 (layerType)) ;
    nand02 ix3771 (.Y (nx3770), .A0 (outMuls_16__14), .A1 (nx5240)) ;
    nand02 ix1359 (.Y (addersInputs_16__15), .A0 (nx3773), .A1 (nx3775)) ;
    nand02 ix3774 (.Y (nx3773), .A0 (currentPage_16__15), .A1 (layerType)) ;
    nand02 ix3776 (.Y (nx3775), .A0 (outMuls_16__15), .A1 (nx5240)) ;
    nand02 ix1367 (.Y (addersInputs_15__0), .A0 (nx3778), .A1 (nx3780)) ;
    nand02 ix3779 (.Y (nx3778), .A0 (currentPage_15__0), .A1 (layerType)) ;
    nand02 ix3781 (.Y (nx3780), .A0 (outMuls_15__0), .A1 (nx5240)) ;
    nand02 ix1375 (.Y (addersInputs_15__1), .A0 (nx3783), .A1 (nx3785)) ;
    nand02 ix3784 (.Y (nx3783), .A0 (currentPage_15__1), .A1 (layerType)) ;
    nand02 ix3786 (.Y (nx3785), .A0 (outMuls_15__1), .A1 (nx5240)) ;
    nand02 ix1383 (.Y (addersInputs_15__2), .A0 (nx3788), .A1 (nx3790)) ;
    nand02 ix3789 (.Y (nx3788), .A0 (currentPage_15__2), .A1 (layerType)) ;
    nand02 ix3791 (.Y (nx3790), .A0 (outMuls_15__2), .A1 (nx5240)) ;
    nand02 ix1391 (.Y (addersInputs_15__3), .A0 (nx3793), .A1 (nx3795)) ;
    nand02 ix3794 (.Y (nx3793), .A0 (currentPage_15__3), .A1 (layerType)) ;
    nand02 ix3796 (.Y (nx3795), .A0 (outMuls_15__3), .A1 (nx5242)) ;
    nand02 ix1399 (.Y (addersInputs_15__4), .A0 (nx3798), .A1 (nx3800)) ;
    nand02 ix3799 (.Y (nx3798), .A0 (currentPage_15__4), .A1 (layerType)) ;
    nand02 ix3801 (.Y (nx3800), .A0 (outMuls_15__4), .A1 (nx5242)) ;
    nand02 ix1407 (.Y (addersInputs_15__5), .A0 (nx3803), .A1 (nx3805)) ;
    nand02 ix3804 (.Y (nx3803), .A0 (currentPage_15__5), .A1 (layerType)) ;
    nand02 ix3806 (.Y (nx3805), .A0 (outMuls_15__5), .A1 (nx5242)) ;
    nand02 ix1415 (.Y (addersInputs_15__6), .A0 (nx3808), .A1 (nx3810)) ;
    nand02 ix3809 (.Y (nx3808), .A0 (currentPage_15__6), .A1 (layerType)) ;
    nand02 ix3811 (.Y (nx3810), .A0 (outMuls_15__6), .A1 (nx5242)) ;
    nand02 ix1423 (.Y (addersInputs_15__7), .A0 (nx3813), .A1 (nx3815)) ;
    nand02 ix3814 (.Y (nx3813), .A0 (currentPage_15__7), .A1 (layerType)) ;
    nand02 ix3816 (.Y (nx3815), .A0 (outMuls_15__7), .A1 (nx5242)) ;
    nand02 ix1431 (.Y (addersInputs_15__8), .A0 (nx3818), .A1 (nx3820)) ;
    nand02 ix3819 (.Y (nx3818), .A0 (currentPage_15__8), .A1 (layerType)) ;
    nand02 ix3821 (.Y (nx3820), .A0 (outMuls_15__8), .A1 (nx5242)) ;
    nand02 ix1439 (.Y (addersInputs_15__9), .A0 (nx3823), .A1 (nx3825)) ;
    nand02 ix3824 (.Y (nx3823), .A0 (currentPage_15__9), .A1 (layerType)) ;
    nand02 ix3826 (.Y (nx3825), .A0 (outMuls_15__9), .A1 (nx5242)) ;
    nand02 ix1447 (.Y (addersInputs_15__10), .A0 (nx3828), .A1 (nx3830)) ;
    nand02 ix3829 (.Y (nx3828), .A0 (currentPage_15__10), .A1 (layerType)) ;
    nand02 ix3831 (.Y (nx3830), .A0 (outMuls_15__10), .A1 (nx5244)) ;
    nand02 ix1455 (.Y (addersInputs_15__11), .A0 (nx3833), .A1 (nx3835)) ;
    nand02 ix3834 (.Y (nx3833), .A0 (currentPage_15__11), .A1 (layerType)) ;
    nand02 ix3836 (.Y (nx3835), .A0 (outMuls_15__11), .A1 (nx5244)) ;
    nand02 ix1463 (.Y (addersInputs_15__12), .A0 (nx3838), .A1 (nx3840)) ;
    nand02 ix3839 (.Y (nx3838), .A0 (currentPage_15__12), .A1 (layerType)) ;
    nand02 ix3841 (.Y (nx3840), .A0 (outMuls_15__12), .A1 (nx5244)) ;
    nand02 ix1471 (.Y (addersInputs_15__13), .A0 (nx3843), .A1 (nx3845)) ;
    nand02 ix3844 (.Y (nx3843), .A0 (currentPage_15__13), .A1 (layerType)) ;
    nand02 ix3846 (.Y (nx3845), .A0 (outMuls_15__13), .A1 (nx5244)) ;
    nand02 ix1479 (.Y (addersInputs_15__14), .A0 (nx3848), .A1 (nx3850)) ;
    nand02 ix3849 (.Y (nx3848), .A0 (currentPage_15__14), .A1 (layerType)) ;
    nand02 ix3851 (.Y (nx3850), .A0 (outMuls_15__14), .A1 (nx5244)) ;
    nand02 ix1487 (.Y (addersInputs_15__15), .A0 (nx3853), .A1 (nx3855)) ;
    nand02 ix3854 (.Y (nx3853), .A0 (currentPage_15__15), .A1 (layerType)) ;
    nand02 ix3856 (.Y (nx3855), .A0 (outMuls_15__15), .A1 (nx5244)) ;
    nand02 ix1495 (.Y (addersInputs_14__0), .A0 (nx3858), .A1 (nx3860)) ;
    nand02 ix3859 (.Y (nx3858), .A0 (currentPage_14__0), .A1 (layerType)) ;
    nand02 ix3861 (.Y (nx3860), .A0 (outMuls_14__0), .A1 (nx5244)) ;
    nand02 ix1503 (.Y (addersInputs_14__1), .A0 (nx3863), .A1 (nx3865)) ;
    nand02 ix3864 (.Y (nx3863), .A0 (currentPage_14__1), .A1 (layerType)) ;
    nand02 ix3866 (.Y (nx3865), .A0 (outMuls_14__1), .A1 (nx5246)) ;
    nand02 ix1511 (.Y (addersInputs_14__2), .A0 (nx3868), .A1 (nx3870)) ;
    nand02 ix3869 (.Y (nx3868), .A0 (currentPage_14__2), .A1 (layerType)) ;
    nand02 ix3871 (.Y (nx3870), .A0 (outMuls_14__2), .A1 (nx5246)) ;
    nand02 ix1519 (.Y (addersInputs_14__3), .A0 (nx3873), .A1 (nx3875)) ;
    nand02 ix3874 (.Y (nx3873), .A0 (currentPage_14__3), .A1 (layerType)) ;
    nand02 ix3876 (.Y (nx3875), .A0 (outMuls_14__3), .A1 (nx5246)) ;
    nand02 ix1527 (.Y (addersInputs_14__4), .A0 (nx3878), .A1 (nx3880)) ;
    nand02 ix3879 (.Y (nx3878), .A0 (currentPage_14__4), .A1 (layerType)) ;
    nand02 ix3881 (.Y (nx3880), .A0 (outMuls_14__4), .A1 (nx5246)) ;
    nand02 ix1535 (.Y (addersInputs_14__5), .A0 (nx3883), .A1 (nx3885)) ;
    nand02 ix3884 (.Y (nx3883), .A0 (currentPage_14__5), .A1 (layerType)) ;
    nand02 ix3886 (.Y (nx3885), .A0 (outMuls_14__5), .A1 (nx5246)) ;
    nand02 ix1543 (.Y (addersInputs_14__6), .A0 (nx3888), .A1 (nx3890)) ;
    nand02 ix3889 (.Y (nx3888), .A0 (currentPage_14__6), .A1 (layerType)) ;
    nand02 ix3891 (.Y (nx3890), .A0 (outMuls_14__6), .A1 (nx5246)) ;
    nand02 ix1551 (.Y (addersInputs_14__7), .A0 (nx3893), .A1 (nx3895)) ;
    nand02 ix3894 (.Y (nx3893), .A0 (currentPage_14__7), .A1 (layerType)) ;
    nand02 ix3896 (.Y (nx3895), .A0 (outMuls_14__7), .A1 (nx5246)) ;
    nand02 ix1559 (.Y (addersInputs_14__8), .A0 (nx3898), .A1 (nx3900)) ;
    nand02 ix3899 (.Y (nx3898), .A0 (currentPage_14__8), .A1 (layerType)) ;
    nand02 ix3901 (.Y (nx3900), .A0 (outMuls_14__8), .A1 (nx5248)) ;
    nand02 ix1567 (.Y (addersInputs_14__9), .A0 (nx3903), .A1 (nx3905)) ;
    nand02 ix3904 (.Y (nx3903), .A0 (currentPage_14__9), .A1 (layerType)) ;
    nand02 ix3906 (.Y (nx3905), .A0 (outMuls_14__9), .A1 (nx5248)) ;
    nand02 ix1575 (.Y (addersInputs_14__10), .A0 (nx3908), .A1 (nx3910)) ;
    nand02 ix3909 (.Y (nx3908), .A0 (currentPage_14__10), .A1 (layerType)) ;
    nand02 ix3911 (.Y (nx3910), .A0 (outMuls_14__10), .A1 (nx5248)) ;
    nand02 ix1583 (.Y (addersInputs_14__11), .A0 (nx3913), .A1 (nx3915)) ;
    nand02 ix3914 (.Y (nx3913), .A0 (currentPage_14__11), .A1 (layerType)) ;
    nand02 ix3916 (.Y (nx3915), .A0 (outMuls_14__11), .A1 (nx5248)) ;
    nand02 ix1591 (.Y (addersInputs_14__12), .A0 (nx3918), .A1 (nx3920)) ;
    nand02 ix3919 (.Y (nx3918), .A0 (currentPage_14__12), .A1 (layerType)) ;
    nand02 ix3921 (.Y (nx3920), .A0 (outMuls_14__12), .A1 (nx5248)) ;
    nand02 ix1599 (.Y (addersInputs_14__13), .A0 (nx3923), .A1 (nx3925)) ;
    nand02 ix3924 (.Y (nx3923), .A0 (currentPage_14__13), .A1 (layerType)) ;
    nand02 ix3926 (.Y (nx3925), .A0 (outMuls_14__13), .A1 (nx5248)) ;
    nand02 ix1607 (.Y (addersInputs_14__14), .A0 (nx3928), .A1 (nx3930)) ;
    nand02 ix3929 (.Y (nx3928), .A0 (currentPage_14__14), .A1 (layerType)) ;
    nand02 ix3931 (.Y (nx3930), .A0 (outMuls_14__14), .A1 (nx5248)) ;
    nand02 ix1615 (.Y (addersInputs_14__15), .A0 (nx3933), .A1 (nx3935)) ;
    nand02 ix3934 (.Y (nx3933), .A0 (currentPage_14__15), .A1 (layerType)) ;
    nand02 ix3936 (.Y (nx3935), .A0 (outMuls_14__15), .A1 (nx5250)) ;
    nand02 ix1623 (.Y (addersInputs_13__0), .A0 (nx3938), .A1 (nx3940)) ;
    nand02 ix3939 (.Y (nx3938), .A0 (currentPage_13__0), .A1 (layerType)) ;
    nand02 ix3941 (.Y (nx3940), .A0 (outMuls_13__0), .A1 (nx5250)) ;
    nand02 ix1631 (.Y (addersInputs_13__1), .A0 (nx3943), .A1 (nx3945)) ;
    nand02 ix3944 (.Y (nx3943), .A0 (currentPage_13__1), .A1 (layerType)) ;
    nand02 ix3946 (.Y (nx3945), .A0 (outMuls_13__1), .A1 (nx5250)) ;
    nand02 ix1639 (.Y (addersInputs_13__2), .A0 (nx3948), .A1 (nx3950)) ;
    nand02 ix3949 (.Y (nx3948), .A0 (currentPage_13__2), .A1 (layerType)) ;
    nand02 ix3951 (.Y (nx3950), .A0 (outMuls_13__2), .A1 (nx5250)) ;
    nand02 ix1647 (.Y (addersInputs_13__3), .A0 (nx3953), .A1 (nx3955)) ;
    nand02 ix3954 (.Y (nx3953), .A0 (currentPage_13__3), .A1 (layerType)) ;
    nand02 ix3956 (.Y (nx3955), .A0 (outMuls_13__3), .A1 (nx5250)) ;
    nand02 ix1655 (.Y (addersInputs_13__4), .A0 (nx3958), .A1 (nx3960)) ;
    nand02 ix3959 (.Y (nx3958), .A0 (currentPage_13__4), .A1 (layerType)) ;
    nand02 ix3961 (.Y (nx3960), .A0 (outMuls_13__4), .A1 (nx5250)) ;
    nand02 ix1663 (.Y (addersInputs_13__5), .A0 (nx3963), .A1 (nx3965)) ;
    nand02 ix3964 (.Y (nx3963), .A0 (currentPage_13__5), .A1 (layerType)) ;
    nand02 ix3966 (.Y (nx3965), .A0 (outMuls_13__5), .A1 (nx5250)) ;
    nand02 ix1671 (.Y (addersInputs_13__6), .A0 (nx3968), .A1 (nx3970)) ;
    nand02 ix3969 (.Y (nx3968), .A0 (currentPage_13__6), .A1 (layerType)) ;
    nand02 ix3971 (.Y (nx3970), .A0 (outMuls_13__6), .A1 (nx5252)) ;
    nand02 ix1679 (.Y (addersInputs_13__7), .A0 (nx3973), .A1 (nx3975)) ;
    nand02 ix3974 (.Y (nx3973), .A0 (currentPage_13__7), .A1 (layerType)) ;
    nand02 ix3976 (.Y (nx3975), .A0 (outMuls_13__7), .A1 (nx5252)) ;
    nand02 ix1687 (.Y (addersInputs_13__8), .A0 (nx3978), .A1 (nx3980)) ;
    nand02 ix3979 (.Y (nx3978), .A0 (currentPage_13__8), .A1 (layerType)) ;
    nand02 ix3981 (.Y (nx3980), .A0 (outMuls_13__8), .A1 (nx5252)) ;
    nand02 ix1695 (.Y (addersInputs_13__9), .A0 (nx3983), .A1 (nx3985)) ;
    nand02 ix3984 (.Y (nx3983), .A0 (currentPage_13__9), .A1 (layerType)) ;
    nand02 ix3986 (.Y (nx3985), .A0 (outMuls_13__9), .A1 (nx5252)) ;
    nand02 ix1703 (.Y (addersInputs_13__10), .A0 (nx3988), .A1 (nx3990)) ;
    nand02 ix3989 (.Y (nx3988), .A0 (currentPage_13__10), .A1 (layerType)) ;
    nand02 ix3991 (.Y (nx3990), .A0 (outMuls_13__10), .A1 (nx5252)) ;
    nand02 ix1711 (.Y (addersInputs_13__11), .A0 (nx3993), .A1 (nx3995)) ;
    nand02 ix3994 (.Y (nx3993), .A0 (currentPage_13__11), .A1 (layerType)) ;
    nand02 ix3996 (.Y (nx3995), .A0 (outMuls_13__11), .A1 (nx5252)) ;
    nand02 ix1719 (.Y (addersInputs_13__12), .A0 (nx3998), .A1 (nx4000)) ;
    nand02 ix3999 (.Y (nx3998), .A0 (currentPage_13__12), .A1 (layerType)) ;
    nand02 ix4001 (.Y (nx4000), .A0 (outMuls_13__12), .A1 (nx5252)) ;
    nand02 ix1727 (.Y (addersInputs_13__13), .A0 (nx4003), .A1 (nx4005)) ;
    nand02 ix4004 (.Y (nx4003), .A0 (currentPage_13__13), .A1 (layerType)) ;
    nand02 ix4006 (.Y (nx4005), .A0 (outMuls_13__13), .A1 (nx5254)) ;
    nand02 ix1735 (.Y (addersInputs_13__14), .A0 (nx4008), .A1 (nx4010)) ;
    nand02 ix4009 (.Y (nx4008), .A0 (currentPage_13__14), .A1 (layerType)) ;
    nand02 ix4011 (.Y (nx4010), .A0 (outMuls_13__14), .A1 (nx5254)) ;
    nand02 ix1743 (.Y (addersInputs_13__15), .A0 (nx4013), .A1 (nx4015)) ;
    nand02 ix4014 (.Y (nx4013), .A0 (currentPage_13__15), .A1 (layerType)) ;
    nand02 ix4016 (.Y (nx4015), .A0 (outMuls_13__15), .A1 (nx5254)) ;
    nand02 ix1751 (.Y (addersInputs_12__0), .A0 (nx4018), .A1 (nx4020)) ;
    nand02 ix4019 (.Y (nx4018), .A0 (currentPage_12__0), .A1 (layerType)) ;
    nand02 ix4021 (.Y (nx4020), .A0 (outMuls_12__0), .A1 (nx5254)) ;
    nand02 ix1759 (.Y (addersInputs_12__1), .A0 (nx4023), .A1 (nx4025)) ;
    nand02 ix4024 (.Y (nx4023), .A0 (currentPage_12__1), .A1 (layerType)) ;
    nand02 ix4026 (.Y (nx4025), .A0 (outMuls_12__1), .A1 (nx5254)) ;
    nand02 ix1767 (.Y (addersInputs_12__2), .A0 (nx4028), .A1 (nx4030)) ;
    nand02 ix4029 (.Y (nx4028), .A0 (currentPage_12__2), .A1 (layerType)) ;
    nand02 ix4031 (.Y (nx4030), .A0 (outMuls_12__2), .A1 (nx5254)) ;
    nand02 ix1775 (.Y (addersInputs_12__3), .A0 (nx4033), .A1 (nx4035)) ;
    nand02 ix4034 (.Y (nx4033), .A0 (currentPage_12__3), .A1 (layerType)) ;
    nand02 ix4036 (.Y (nx4035), .A0 (outMuls_12__3), .A1 (nx5254)) ;
    nand02 ix1783 (.Y (addersInputs_12__4), .A0 (nx4038), .A1 (nx4040)) ;
    nand02 ix4039 (.Y (nx4038), .A0 (currentPage_12__4), .A1 (layerType)) ;
    nand02 ix4041 (.Y (nx4040), .A0 (outMuls_12__4), .A1 (nx5256)) ;
    nand02 ix1791 (.Y (addersInputs_12__5), .A0 (nx4043), .A1 (nx4045)) ;
    nand02 ix4044 (.Y (nx4043), .A0 (currentPage_12__5), .A1 (layerType)) ;
    nand02 ix4046 (.Y (nx4045), .A0 (outMuls_12__5), .A1 (nx5256)) ;
    nand02 ix1799 (.Y (addersInputs_12__6), .A0 (nx4048), .A1 (nx4050)) ;
    nand02 ix4049 (.Y (nx4048), .A0 (currentPage_12__6), .A1 (layerType)) ;
    nand02 ix4051 (.Y (nx4050), .A0 (outMuls_12__6), .A1 (nx5256)) ;
    nand02 ix1807 (.Y (addersInputs_12__7), .A0 (nx4053), .A1 (nx4055)) ;
    nand02 ix4054 (.Y (nx4053), .A0 (currentPage_12__7), .A1 (layerType)) ;
    nand02 ix4056 (.Y (nx4055), .A0 (outMuls_12__7), .A1 (nx5256)) ;
    nand02 ix1815 (.Y (addersInputs_12__8), .A0 (nx4058), .A1 (nx4060)) ;
    nand02 ix4059 (.Y (nx4058), .A0 (currentPage_12__8), .A1 (layerType)) ;
    nand02 ix4061 (.Y (nx4060), .A0 (outMuls_12__8), .A1 (nx5256)) ;
    nand02 ix1823 (.Y (addersInputs_12__9), .A0 (nx4063), .A1 (nx4065)) ;
    nand02 ix4064 (.Y (nx4063), .A0 (currentPage_12__9), .A1 (layerType)) ;
    nand02 ix4066 (.Y (nx4065), .A0 (outMuls_12__9), .A1 (nx5256)) ;
    nand02 ix1831 (.Y (addersInputs_12__10), .A0 (nx4068), .A1 (nx4070)) ;
    nand02 ix4069 (.Y (nx4068), .A0 (currentPage_12__10), .A1 (layerType)) ;
    nand02 ix4071 (.Y (nx4070), .A0 (outMuls_12__10), .A1 (nx5256)) ;
    nand02 ix1839 (.Y (addersInputs_12__11), .A0 (nx4073), .A1 (nx4075)) ;
    nand02 ix4074 (.Y (nx4073), .A0 (currentPage_12__11), .A1 (layerType)) ;
    nand02 ix4076 (.Y (nx4075), .A0 (outMuls_12__11), .A1 (nx5258)) ;
    nand02 ix1847 (.Y (addersInputs_12__12), .A0 (nx4078), .A1 (nx4080)) ;
    nand02 ix4079 (.Y (nx4078), .A0 (currentPage_12__12), .A1 (layerType)) ;
    nand02 ix4081 (.Y (nx4080), .A0 (outMuls_12__12), .A1 (nx5258)) ;
    nand02 ix1855 (.Y (addersInputs_12__13), .A0 (nx4083), .A1 (nx4085)) ;
    nand02 ix4084 (.Y (nx4083), .A0 (currentPage_12__13), .A1 (layerType)) ;
    nand02 ix4086 (.Y (nx4085), .A0 (outMuls_12__13), .A1 (nx5258)) ;
    nand02 ix1863 (.Y (addersInputs_12__14), .A0 (nx4088), .A1 (nx4090)) ;
    nand02 ix4089 (.Y (nx4088), .A0 (currentPage_12__14), .A1 (layerType)) ;
    nand02 ix4091 (.Y (nx4090), .A0 (outMuls_12__14), .A1 (nx5258)) ;
    nand02 ix1871 (.Y (addersInputs_12__15), .A0 (nx4093), .A1 (nx4095)) ;
    nand02 ix4094 (.Y (nx4093), .A0 (currentPage_12__15), .A1 (layerType)) ;
    nand02 ix4096 (.Y (nx4095), .A0 (outMuls_12__15), .A1 (nx5258)) ;
    nand02 ix1879 (.Y (addersInputs_11__0), .A0 (nx4098), .A1 (nx4100)) ;
    nand02 ix4099 (.Y (nx4098), .A0 (currentPage_11__0), .A1 (layerType)) ;
    nand02 ix4101 (.Y (nx4100), .A0 (outMuls_11__0), .A1 (nx5258)) ;
    nand02 ix1887 (.Y (addersInputs_11__1), .A0 (nx4103), .A1 (nx4105)) ;
    nand02 ix4104 (.Y (nx4103), .A0 (currentPage_11__1), .A1 (layerType)) ;
    nand02 ix4106 (.Y (nx4105), .A0 (outMuls_11__1), .A1 (nx5258)) ;
    nand02 ix1895 (.Y (addersInputs_11__2), .A0 (nx4108), .A1 (nx4110)) ;
    nand02 ix4109 (.Y (nx4108), .A0 (currentPage_11__2), .A1 (layerType)) ;
    nand02 ix4111 (.Y (nx4110), .A0 (outMuls_11__2), .A1 (nx5260)) ;
    nand02 ix1903 (.Y (addersInputs_11__3), .A0 (nx4113), .A1 (nx4115)) ;
    nand02 ix4114 (.Y (nx4113), .A0 (currentPage_11__3), .A1 (layerType)) ;
    nand02 ix4116 (.Y (nx4115), .A0 (outMuls_11__3), .A1 (nx5260)) ;
    nand02 ix1911 (.Y (addersInputs_11__4), .A0 (nx4118), .A1 (nx4120)) ;
    nand02 ix4119 (.Y (nx4118), .A0 (currentPage_11__4), .A1 (layerType)) ;
    nand02 ix4121 (.Y (nx4120), .A0 (outMuls_11__4), .A1 (nx5260)) ;
    nand02 ix1919 (.Y (addersInputs_11__5), .A0 (nx4123), .A1 (nx4125)) ;
    nand02 ix4124 (.Y (nx4123), .A0 (currentPage_11__5), .A1 (layerType)) ;
    nand02 ix4126 (.Y (nx4125), .A0 (outMuls_11__5), .A1 (nx5260)) ;
    nand02 ix1927 (.Y (addersInputs_11__6), .A0 (nx4128), .A1 (nx4130)) ;
    nand02 ix4129 (.Y (nx4128), .A0 (currentPage_11__6), .A1 (layerType)) ;
    nand02 ix4131 (.Y (nx4130), .A0 (outMuls_11__6), .A1 (nx5260)) ;
    nand02 ix1935 (.Y (addersInputs_11__7), .A0 (nx4133), .A1 (nx4135)) ;
    nand02 ix4134 (.Y (nx4133), .A0 (currentPage_11__7), .A1 (layerType)) ;
    nand02 ix4136 (.Y (nx4135), .A0 (outMuls_11__7), .A1 (nx5260)) ;
    nand02 ix1943 (.Y (addersInputs_11__8), .A0 (nx4138), .A1 (nx4140)) ;
    nand02 ix4139 (.Y (nx4138), .A0 (currentPage_11__8), .A1 (layerType)) ;
    nand02 ix4141 (.Y (nx4140), .A0 (outMuls_11__8), .A1 (nx5260)) ;
    nand02 ix1951 (.Y (addersInputs_11__9), .A0 (nx4143), .A1 (nx4145)) ;
    nand02 ix4144 (.Y (nx4143), .A0 (currentPage_11__9), .A1 (layerType)) ;
    nand02 ix4146 (.Y (nx4145), .A0 (outMuls_11__9), .A1 (nx5262)) ;
    nand02 ix1959 (.Y (addersInputs_11__10), .A0 (nx4148), .A1 (nx4150)) ;
    nand02 ix4149 (.Y (nx4148), .A0 (currentPage_11__10), .A1 (layerType)) ;
    nand02 ix4151 (.Y (nx4150), .A0 (outMuls_11__10), .A1 (nx5262)) ;
    nand02 ix1967 (.Y (addersInputs_11__11), .A0 (nx4153), .A1 (nx4155)) ;
    nand02 ix4154 (.Y (nx4153), .A0 (currentPage_11__11), .A1 (layerType)) ;
    nand02 ix4156 (.Y (nx4155), .A0 (outMuls_11__11), .A1 (nx5262)) ;
    nand02 ix1975 (.Y (addersInputs_11__12), .A0 (nx4158), .A1 (nx4160)) ;
    nand02 ix4159 (.Y (nx4158), .A0 (currentPage_11__12), .A1 (layerType)) ;
    nand02 ix4161 (.Y (nx4160), .A0 (outMuls_11__12), .A1 (nx5262)) ;
    nand02 ix1983 (.Y (addersInputs_11__13), .A0 (nx4163), .A1 (nx4165)) ;
    nand02 ix4164 (.Y (nx4163), .A0 (currentPage_11__13), .A1 (layerType)) ;
    nand02 ix4166 (.Y (nx4165), .A0 (outMuls_11__13), .A1 (nx5262)) ;
    nand02 ix1991 (.Y (addersInputs_11__14), .A0 (nx4168), .A1 (nx4170)) ;
    nand02 ix4169 (.Y (nx4168), .A0 (currentPage_11__14), .A1 (layerType)) ;
    nand02 ix4171 (.Y (nx4170), .A0 (outMuls_11__14), .A1 (nx5262)) ;
    nand02 ix1999 (.Y (addersInputs_11__15), .A0 (nx4173), .A1 (nx4175)) ;
    nand02 ix4174 (.Y (nx4173), .A0 (currentPage_11__15), .A1 (layerType)) ;
    nand02 ix4176 (.Y (nx4175), .A0 (outMuls_11__15), .A1 (nx5262)) ;
    nand02 ix2007 (.Y (addersInputs_10__0), .A0 (nx4178), .A1 (nx4180)) ;
    nand02 ix4179 (.Y (nx4178), .A0 (currentPage_10__0), .A1 (layerType)) ;
    nand02 ix4181 (.Y (nx4180), .A0 (outMuls_10__0), .A1 (nx5264)) ;
    nand02 ix2015 (.Y (addersInputs_10__1), .A0 (nx4183), .A1 (nx4185)) ;
    nand02 ix4184 (.Y (nx4183), .A0 (currentPage_10__1), .A1 (layerType)) ;
    nand02 ix4186 (.Y (nx4185), .A0 (outMuls_10__1), .A1 (nx5264)) ;
    nand02 ix2023 (.Y (addersInputs_10__2), .A0 (nx4188), .A1 (nx4190)) ;
    nand02 ix4189 (.Y (nx4188), .A0 (currentPage_10__2), .A1 (layerType)) ;
    nand02 ix4191 (.Y (nx4190), .A0 (outMuls_10__2), .A1 (nx5264)) ;
    nand02 ix2031 (.Y (addersInputs_10__3), .A0 (nx4193), .A1 (nx4195)) ;
    nand02 ix4194 (.Y (nx4193), .A0 (currentPage_10__3), .A1 (layerType)) ;
    nand02 ix4196 (.Y (nx4195), .A0 (outMuls_10__3), .A1 (nx5264)) ;
    nand02 ix2039 (.Y (addersInputs_10__4), .A0 (nx4198), .A1 (nx4200)) ;
    nand02 ix4199 (.Y (nx4198), .A0 (currentPage_10__4), .A1 (layerType)) ;
    nand02 ix4201 (.Y (nx4200), .A0 (outMuls_10__4), .A1 (nx5264)) ;
    nand02 ix2047 (.Y (addersInputs_10__5), .A0 (nx4203), .A1 (nx4205)) ;
    nand02 ix4204 (.Y (nx4203), .A0 (currentPage_10__5), .A1 (layerType)) ;
    nand02 ix4206 (.Y (nx4205), .A0 (outMuls_10__5), .A1 (nx5264)) ;
    nand02 ix2055 (.Y (addersInputs_10__6), .A0 (nx4208), .A1 (nx4210)) ;
    nand02 ix4209 (.Y (nx4208), .A0 (currentPage_10__6), .A1 (layerType)) ;
    nand02 ix4211 (.Y (nx4210), .A0 (outMuls_10__6), .A1 (nx5264)) ;
    nand02 ix2063 (.Y (addersInputs_10__7), .A0 (nx4213), .A1 (nx4215)) ;
    nand02 ix4214 (.Y (nx4213), .A0 (currentPage_10__7), .A1 (layerType)) ;
    nand02 ix4216 (.Y (nx4215), .A0 (outMuls_10__7), .A1 (nx5266)) ;
    nand02 ix2071 (.Y (addersInputs_10__8), .A0 (nx4218), .A1 (nx4220)) ;
    nand02 ix4219 (.Y (nx4218), .A0 (currentPage_10__8), .A1 (layerType)) ;
    nand02 ix4221 (.Y (nx4220), .A0 (outMuls_10__8), .A1 (nx5266)) ;
    nand02 ix2079 (.Y (addersInputs_10__9), .A0 (nx4223), .A1 (nx4225)) ;
    nand02 ix4224 (.Y (nx4223), .A0 (currentPage_10__9), .A1 (layerType)) ;
    nand02 ix4226 (.Y (nx4225), .A0 (outMuls_10__9), .A1 (nx5266)) ;
    nand02 ix2087 (.Y (addersInputs_10__10), .A0 (nx4228), .A1 (nx4230)) ;
    nand02 ix4229 (.Y (nx4228), .A0 (currentPage_10__10), .A1 (layerType)) ;
    nand02 ix4231 (.Y (nx4230), .A0 (outMuls_10__10), .A1 (nx5266)) ;
    nand02 ix2095 (.Y (addersInputs_10__11), .A0 (nx4233), .A1 (nx4235)) ;
    nand02 ix4234 (.Y (nx4233), .A0 (currentPage_10__11), .A1 (layerType)) ;
    nand02 ix4236 (.Y (nx4235), .A0 (outMuls_10__11), .A1 (nx5266)) ;
    nand02 ix2103 (.Y (addersInputs_10__12), .A0 (nx4238), .A1 (nx4240)) ;
    nand02 ix4239 (.Y (nx4238), .A0 (currentPage_10__12), .A1 (layerType)) ;
    nand02 ix4241 (.Y (nx4240), .A0 (outMuls_10__12), .A1 (nx5266)) ;
    nand02 ix2111 (.Y (addersInputs_10__13), .A0 (nx4243), .A1 (nx4245)) ;
    nand02 ix4244 (.Y (nx4243), .A0 (currentPage_10__13), .A1 (layerType)) ;
    nand02 ix4246 (.Y (nx4245), .A0 (outMuls_10__13), .A1 (nx5266)) ;
    nand02 ix2119 (.Y (addersInputs_10__14), .A0 (nx4248), .A1 (nx4250)) ;
    nand02 ix4249 (.Y (nx4248), .A0 (currentPage_10__14), .A1 (layerType)) ;
    nand02 ix4251 (.Y (nx4250), .A0 (outMuls_10__14), .A1 (nx5268)) ;
    nand02 ix2127 (.Y (addersInputs_10__15), .A0 (nx4253), .A1 (nx4255)) ;
    nand02 ix4254 (.Y (nx4253), .A0 (currentPage_10__15), .A1 (layerType)) ;
    nand02 ix4256 (.Y (nx4255), .A0 (outMuls_10__15), .A1 (nx5268)) ;
    nand02 ix2135 (.Y (addersInputs_9__0), .A0 (nx4258), .A1 (nx4260)) ;
    nand02 ix4259 (.Y (nx4258), .A0 (currentPage_9__0), .A1 (layerType)) ;
    nand02 ix4261 (.Y (nx4260), .A0 (outMuls_9__0), .A1 (nx5268)) ;
    nand02 ix2143 (.Y (addersInputs_9__1), .A0 (nx4263), .A1 (nx4265)) ;
    nand02 ix4264 (.Y (nx4263), .A0 (currentPage_9__1), .A1 (layerType)) ;
    nand02 ix4266 (.Y (nx4265), .A0 (outMuls_9__1), .A1 (nx5268)) ;
    nand02 ix2151 (.Y (addersInputs_9__2), .A0 (nx4268), .A1 (nx4270)) ;
    nand02 ix4269 (.Y (nx4268), .A0 (currentPage_9__2), .A1 (layerType)) ;
    nand02 ix4271 (.Y (nx4270), .A0 (outMuls_9__2), .A1 (nx5268)) ;
    nand02 ix2159 (.Y (addersInputs_9__3), .A0 (nx4273), .A1 (nx4275)) ;
    nand02 ix4274 (.Y (nx4273), .A0 (currentPage_9__3), .A1 (layerType)) ;
    nand02 ix4276 (.Y (nx4275), .A0 (outMuls_9__3), .A1 (nx5268)) ;
    nand02 ix2167 (.Y (addersInputs_9__4), .A0 (nx4278), .A1 (nx4280)) ;
    nand02 ix4279 (.Y (nx4278), .A0 (currentPage_9__4), .A1 (layerType)) ;
    nand02 ix4281 (.Y (nx4280), .A0 (outMuls_9__4), .A1 (nx5268)) ;
    nand02 ix2175 (.Y (addersInputs_9__5), .A0 (nx4283), .A1 (nx4285)) ;
    nand02 ix4284 (.Y (nx4283), .A0 (currentPage_9__5), .A1 (layerType)) ;
    nand02 ix4286 (.Y (nx4285), .A0 (outMuls_9__5), .A1 (nx5270)) ;
    nand02 ix2183 (.Y (addersInputs_9__6), .A0 (nx4288), .A1 (nx4290)) ;
    nand02 ix4289 (.Y (nx4288), .A0 (currentPage_9__6), .A1 (layerType)) ;
    nand02 ix4291 (.Y (nx4290), .A0 (outMuls_9__6), .A1 (nx5270)) ;
    nand02 ix2191 (.Y (addersInputs_9__7), .A0 (nx4293), .A1 (nx4295)) ;
    nand02 ix4294 (.Y (nx4293), .A0 (currentPage_9__7), .A1 (layerType)) ;
    nand02 ix4296 (.Y (nx4295), .A0 (outMuls_9__7), .A1 (nx5270)) ;
    nand02 ix2199 (.Y (addersInputs_9__8), .A0 (nx4298), .A1 (nx4300)) ;
    nand02 ix4299 (.Y (nx4298), .A0 (currentPage_9__8), .A1 (layerType)) ;
    nand02 ix4301 (.Y (nx4300), .A0 (outMuls_9__8), .A1 (nx5270)) ;
    nand02 ix2207 (.Y (addersInputs_9__9), .A0 (nx4303), .A1 (nx4305)) ;
    nand02 ix4304 (.Y (nx4303), .A0 (currentPage_9__9), .A1 (layerType)) ;
    nand02 ix4306 (.Y (nx4305), .A0 (outMuls_9__9), .A1 (nx5270)) ;
    nand02 ix2215 (.Y (addersInputs_9__10), .A0 (nx4308), .A1 (nx4310)) ;
    nand02 ix4309 (.Y (nx4308), .A0 (currentPage_9__10), .A1 (layerType)) ;
    nand02 ix4311 (.Y (nx4310), .A0 (outMuls_9__10), .A1 (nx5270)) ;
    nand02 ix2223 (.Y (addersInputs_9__11), .A0 (nx4313), .A1 (nx4315)) ;
    nand02 ix4314 (.Y (nx4313), .A0 (currentPage_9__11), .A1 (layerType)) ;
    nand02 ix4316 (.Y (nx4315), .A0 (outMuls_9__11), .A1 (nx5270)) ;
    nand02 ix2231 (.Y (addersInputs_9__12), .A0 (nx4318), .A1 (nx4320)) ;
    nand02 ix4319 (.Y (nx4318), .A0 (currentPage_9__12), .A1 (layerType)) ;
    nand02 ix4321 (.Y (nx4320), .A0 (outMuls_9__12), .A1 (nx5272)) ;
    nand02 ix2239 (.Y (addersInputs_9__13), .A0 (nx4323), .A1 (nx4325)) ;
    nand02 ix4324 (.Y (nx4323), .A0 (currentPage_9__13), .A1 (layerType)) ;
    nand02 ix4326 (.Y (nx4325), .A0 (outMuls_9__13), .A1 (nx5272)) ;
    nand02 ix2247 (.Y (addersInputs_9__14), .A0 (nx4328), .A1 (nx4330)) ;
    nand02 ix4329 (.Y (nx4328), .A0 (currentPage_9__14), .A1 (layerType)) ;
    nand02 ix4331 (.Y (nx4330), .A0 (outMuls_9__14), .A1 (nx5272)) ;
    nand02 ix2255 (.Y (addersInputs_9__15), .A0 (nx4333), .A1 (nx4335)) ;
    nand02 ix4334 (.Y (nx4333), .A0 (currentPage_9__15), .A1 (layerType)) ;
    nand02 ix4336 (.Y (nx4335), .A0 (outMuls_9__15), .A1 (nx5272)) ;
    nand02 ix2263 (.Y (addersInputs_8__0), .A0 (nx4338), .A1 (nx4340)) ;
    nand02 ix4339 (.Y (nx4338), .A0 (currentPage_8__0), .A1 (layerType)) ;
    nand02 ix4341 (.Y (nx4340), .A0 (outMuls_8__0), .A1 (nx5272)) ;
    nand02 ix2271 (.Y (addersInputs_8__1), .A0 (nx4343), .A1 (nx4345)) ;
    nand02 ix4344 (.Y (nx4343), .A0 (currentPage_8__1), .A1 (layerType)) ;
    nand02 ix4346 (.Y (nx4345), .A0 (outMuls_8__1), .A1 (nx5272)) ;
    nand02 ix2279 (.Y (addersInputs_8__2), .A0 (nx4348), .A1 (nx4350)) ;
    nand02 ix4349 (.Y (nx4348), .A0 (currentPage_8__2), .A1 (layerType)) ;
    nand02 ix4351 (.Y (nx4350), .A0 (outMuls_8__2), .A1 (nx5272)) ;
    nand02 ix2287 (.Y (addersInputs_8__3), .A0 (nx4353), .A1 (nx4355)) ;
    nand02 ix4354 (.Y (nx4353), .A0 (currentPage_8__3), .A1 (layerType)) ;
    nand02 ix4356 (.Y (nx4355), .A0 (outMuls_8__3), .A1 (nx5274)) ;
    nand02 ix2295 (.Y (addersInputs_8__4), .A0 (nx4358), .A1 (nx4360)) ;
    nand02 ix4359 (.Y (nx4358), .A0 (currentPage_8__4), .A1 (layerType)) ;
    nand02 ix4361 (.Y (nx4360), .A0 (outMuls_8__4), .A1 (nx5274)) ;
    nand02 ix2303 (.Y (addersInputs_8__5), .A0 (nx4363), .A1 (nx4365)) ;
    nand02 ix4364 (.Y (nx4363), .A0 (currentPage_8__5), .A1 (layerType)) ;
    nand02 ix4366 (.Y (nx4365), .A0 (outMuls_8__5), .A1 (nx5274)) ;
    nand02 ix2311 (.Y (addersInputs_8__6), .A0 (nx4368), .A1 (nx4370)) ;
    nand02 ix4369 (.Y (nx4368), .A0 (currentPage_8__6), .A1 (layerType)) ;
    nand02 ix4371 (.Y (nx4370), .A0 (outMuls_8__6), .A1 (nx5274)) ;
    nand02 ix2319 (.Y (addersInputs_8__7), .A0 (nx4373), .A1 (nx4375)) ;
    nand02 ix4374 (.Y (nx4373), .A0 (currentPage_8__7), .A1 (layerType)) ;
    nand02 ix4376 (.Y (nx4375), .A0 (outMuls_8__7), .A1 (nx5274)) ;
    nand02 ix2327 (.Y (addersInputs_8__8), .A0 (nx4378), .A1 (nx4380)) ;
    nand02 ix4379 (.Y (nx4378), .A0 (currentPage_8__8), .A1 (layerType)) ;
    nand02 ix4381 (.Y (nx4380), .A0 (outMuls_8__8), .A1 (nx5274)) ;
    nand02 ix2335 (.Y (addersInputs_8__9), .A0 (nx4383), .A1 (nx4385)) ;
    nand02 ix4384 (.Y (nx4383), .A0 (currentPage_8__9), .A1 (layerType)) ;
    nand02 ix4386 (.Y (nx4385), .A0 (outMuls_8__9), .A1 (nx5274)) ;
    nand02 ix2343 (.Y (addersInputs_8__10), .A0 (nx4388), .A1 (nx4390)) ;
    nand02 ix4389 (.Y (nx4388), .A0 (currentPage_8__10), .A1 (layerType)) ;
    nand02 ix4391 (.Y (nx4390), .A0 (outMuls_8__10), .A1 (nx5276)) ;
    nand02 ix2351 (.Y (addersInputs_8__11), .A0 (nx4393), .A1 (nx4395)) ;
    nand02 ix4394 (.Y (nx4393), .A0 (currentPage_8__11), .A1 (layerType)) ;
    nand02 ix4396 (.Y (nx4395), .A0 (outMuls_8__11), .A1 (nx5276)) ;
    nand02 ix2359 (.Y (addersInputs_8__12), .A0 (nx4398), .A1 (nx4400)) ;
    nand02 ix4399 (.Y (nx4398), .A0 (currentPage_8__12), .A1 (layerType)) ;
    nand02 ix4401 (.Y (nx4400), .A0 (outMuls_8__12), .A1 (nx5276)) ;
    nand02 ix2367 (.Y (addersInputs_8__13), .A0 (nx4403), .A1 (nx4405)) ;
    nand02 ix4404 (.Y (nx4403), .A0 (currentPage_8__13), .A1 (layerType)) ;
    nand02 ix4406 (.Y (nx4405), .A0 (outMuls_8__13), .A1 (nx5276)) ;
    nand02 ix2375 (.Y (addersInputs_8__14), .A0 (nx4408), .A1 (nx4410)) ;
    nand02 ix4409 (.Y (nx4408), .A0 (currentPage_8__14), .A1 (layerType)) ;
    nand02 ix4411 (.Y (nx4410), .A0 (outMuls_8__14), .A1 (nx5276)) ;
    nand02 ix2383 (.Y (addersInputs_8__15), .A0 (nx4413), .A1 (nx4415)) ;
    nand02 ix4414 (.Y (nx4413), .A0 (currentPage_8__15), .A1 (layerType)) ;
    nand02 ix4416 (.Y (nx4415), .A0 (outMuls_8__15), .A1 (nx5276)) ;
    nand02 ix2391 (.Y (addersInputs_7__0), .A0 (nx4418), .A1 (nx4420)) ;
    nand02 ix4419 (.Y (nx4418), .A0 (currentPage_7__0), .A1 (layerType)) ;
    nand02 ix4421 (.Y (nx4420), .A0 (outMuls_7__0), .A1 (nx5276)) ;
    nand02 ix2399 (.Y (addersInputs_7__1), .A0 (nx4423), .A1 (nx4425)) ;
    nand02 ix4424 (.Y (nx4423), .A0 (currentPage_7__1), .A1 (layerType)) ;
    nand02 ix4426 (.Y (nx4425), .A0 (outMuls_7__1), .A1 (nx5278)) ;
    nand02 ix2407 (.Y (addersInputs_7__2), .A0 (nx4428), .A1 (nx4430)) ;
    nand02 ix4429 (.Y (nx4428), .A0 (currentPage_7__2), .A1 (layerType)) ;
    nand02 ix4431 (.Y (nx4430), .A0 (outMuls_7__2), .A1 (nx5278)) ;
    nand02 ix2415 (.Y (addersInputs_7__3), .A0 (nx4433), .A1 (nx4435)) ;
    nand02 ix4434 (.Y (nx4433), .A0 (currentPage_7__3), .A1 (layerType)) ;
    nand02 ix4436 (.Y (nx4435), .A0 (outMuls_7__3), .A1 (nx5278)) ;
    nand02 ix2423 (.Y (addersInputs_7__4), .A0 (nx4438), .A1 (nx4440)) ;
    nand02 ix4439 (.Y (nx4438), .A0 (currentPage_7__4), .A1 (layerType)) ;
    nand02 ix4441 (.Y (nx4440), .A0 (outMuls_7__4), .A1 (nx5278)) ;
    nand02 ix2431 (.Y (addersInputs_7__5), .A0 (nx4443), .A1 (nx4445)) ;
    nand02 ix4444 (.Y (nx4443), .A0 (currentPage_7__5), .A1 (layerType)) ;
    nand02 ix4446 (.Y (nx4445), .A0 (outMuls_7__5), .A1 (nx5278)) ;
    nand02 ix2439 (.Y (addersInputs_7__6), .A0 (nx4448), .A1 (nx4450)) ;
    nand02 ix4449 (.Y (nx4448), .A0 (currentPage_7__6), .A1 (layerType)) ;
    nand02 ix4451 (.Y (nx4450), .A0 (outMuls_7__6), .A1 (nx5278)) ;
    nand02 ix2447 (.Y (addersInputs_7__7), .A0 (nx4453), .A1 (nx4455)) ;
    nand02 ix4454 (.Y (nx4453), .A0 (currentPage_7__7), .A1 (layerType)) ;
    nand02 ix4456 (.Y (nx4455), .A0 (outMuls_7__7), .A1 (nx5278)) ;
    nand02 ix2455 (.Y (addersInputs_7__8), .A0 (nx4458), .A1 (nx4460)) ;
    nand02 ix4459 (.Y (nx4458), .A0 (currentPage_7__8), .A1 (layerType)) ;
    nand02 ix4461 (.Y (nx4460), .A0 (outMuls_7__8), .A1 (nx5280)) ;
    nand02 ix2463 (.Y (addersInputs_7__9), .A0 (nx4463), .A1 (nx4465)) ;
    nand02 ix4464 (.Y (nx4463), .A0 (currentPage_7__9), .A1 (layerType)) ;
    nand02 ix4466 (.Y (nx4465), .A0 (outMuls_7__9), .A1 (nx5280)) ;
    nand02 ix2471 (.Y (addersInputs_7__10), .A0 (nx4468), .A1 (nx4470)) ;
    nand02 ix4469 (.Y (nx4468), .A0 (currentPage_7__10), .A1 (layerType)) ;
    nand02 ix4471 (.Y (nx4470), .A0 (outMuls_7__10), .A1 (nx5280)) ;
    nand02 ix2479 (.Y (addersInputs_7__11), .A0 (nx4473), .A1 (nx4475)) ;
    nand02 ix4474 (.Y (nx4473), .A0 (currentPage_7__11), .A1 (layerType)) ;
    nand02 ix4476 (.Y (nx4475), .A0 (outMuls_7__11), .A1 (nx5280)) ;
    nand02 ix2487 (.Y (addersInputs_7__12), .A0 (nx4478), .A1 (nx4480)) ;
    nand02 ix4479 (.Y (nx4478), .A0 (currentPage_7__12), .A1 (layerType)) ;
    nand02 ix4481 (.Y (nx4480), .A0 (outMuls_7__12), .A1 (nx5280)) ;
    nand02 ix2495 (.Y (addersInputs_7__13), .A0 (nx4483), .A1 (nx4485)) ;
    nand02 ix4484 (.Y (nx4483), .A0 (currentPage_7__13), .A1 (layerType)) ;
    nand02 ix4486 (.Y (nx4485), .A0 (outMuls_7__13), .A1 (nx5280)) ;
    nand02 ix2503 (.Y (addersInputs_7__14), .A0 (nx4488), .A1 (nx4490)) ;
    nand02 ix4489 (.Y (nx4488), .A0 (currentPage_7__14), .A1 (layerType)) ;
    nand02 ix4491 (.Y (nx4490), .A0 (outMuls_7__14), .A1 (nx5280)) ;
    nand02 ix2511 (.Y (addersInputs_7__15), .A0 (nx4493), .A1 (nx4495)) ;
    nand02 ix4494 (.Y (nx4493), .A0 (currentPage_7__15), .A1 (layerType)) ;
    nand02 ix4496 (.Y (nx4495), .A0 (outMuls_7__15), .A1 (nx5282)) ;
    nand02 ix2519 (.Y (addersInputs_6__0), .A0 (nx4498), .A1 (nx4500)) ;
    nand02 ix4499 (.Y (nx4498), .A0 (currentPage_6__0), .A1 (layerType)) ;
    nand02 ix4501 (.Y (nx4500), .A0 (outMuls_6__0), .A1 (nx5282)) ;
    nand02 ix2527 (.Y (addersInputs_6__1), .A0 (nx4503), .A1 (nx4505)) ;
    nand02 ix4504 (.Y (nx4503), .A0 (currentPage_6__1), .A1 (layerType)) ;
    nand02 ix4506 (.Y (nx4505), .A0 (outMuls_6__1), .A1 (nx5282)) ;
    nand02 ix2535 (.Y (addersInputs_6__2), .A0 (nx4508), .A1 (nx4510)) ;
    nand02 ix4509 (.Y (nx4508), .A0 (currentPage_6__2), .A1 (layerType)) ;
    nand02 ix4511 (.Y (nx4510), .A0 (outMuls_6__2), .A1 (nx5282)) ;
    nand02 ix2543 (.Y (addersInputs_6__3), .A0 (nx4513), .A1 (nx4515)) ;
    nand02 ix4514 (.Y (nx4513), .A0 (currentPage_6__3), .A1 (layerType)) ;
    nand02 ix4516 (.Y (nx4515), .A0 (outMuls_6__3), .A1 (nx5282)) ;
    nand02 ix2551 (.Y (addersInputs_6__4), .A0 (nx4518), .A1 (nx4520)) ;
    nand02 ix4519 (.Y (nx4518), .A0 (currentPage_6__4), .A1 (layerType)) ;
    nand02 ix4521 (.Y (nx4520), .A0 (outMuls_6__4), .A1 (nx5282)) ;
    nand02 ix2559 (.Y (addersInputs_6__5), .A0 (nx4523), .A1 (nx4525)) ;
    nand02 ix4524 (.Y (nx4523), .A0 (currentPage_6__5), .A1 (layerType)) ;
    nand02 ix4526 (.Y (nx4525), .A0 (outMuls_6__5), .A1 (nx5282)) ;
    nand02 ix2567 (.Y (addersInputs_6__6), .A0 (nx4528), .A1 (nx4530)) ;
    nand02 ix4529 (.Y (nx4528), .A0 (currentPage_6__6), .A1 (layerType)) ;
    nand02 ix4531 (.Y (nx4530), .A0 (outMuls_6__6), .A1 (nx5284)) ;
    nand02 ix2575 (.Y (addersInputs_6__7), .A0 (nx4533), .A1 (nx4535)) ;
    nand02 ix4534 (.Y (nx4533), .A0 (currentPage_6__7), .A1 (layerType)) ;
    nand02 ix4536 (.Y (nx4535), .A0 (outMuls_6__7), .A1 (nx5284)) ;
    nand02 ix2583 (.Y (addersInputs_6__8), .A0 (nx4538), .A1 (nx4540)) ;
    nand02 ix4539 (.Y (nx4538), .A0 (currentPage_6__8), .A1 (layerType)) ;
    nand02 ix4541 (.Y (nx4540), .A0 (outMuls_6__8), .A1 (nx5284)) ;
    nand02 ix2591 (.Y (addersInputs_6__9), .A0 (nx4543), .A1 (nx4545)) ;
    nand02 ix4544 (.Y (nx4543), .A0 (currentPage_6__9), .A1 (layerType)) ;
    nand02 ix4546 (.Y (nx4545), .A0 (outMuls_6__9), .A1 (nx5284)) ;
    nand02 ix2599 (.Y (addersInputs_6__10), .A0 (nx4548), .A1 (nx4550)) ;
    nand02 ix4549 (.Y (nx4548), .A0 (currentPage_6__10), .A1 (layerType)) ;
    nand02 ix4551 (.Y (nx4550), .A0 (outMuls_6__10), .A1 (nx5284)) ;
    nand02 ix2607 (.Y (addersInputs_6__11), .A0 (nx4553), .A1 (nx4555)) ;
    nand02 ix4554 (.Y (nx4553), .A0 (currentPage_6__11), .A1 (layerType)) ;
    nand02 ix4556 (.Y (nx4555), .A0 (outMuls_6__11), .A1 (nx5284)) ;
    nand02 ix2615 (.Y (addersInputs_6__12), .A0 (nx4558), .A1 (nx4560)) ;
    nand02 ix4559 (.Y (nx4558), .A0 (currentPage_6__12), .A1 (layerType)) ;
    nand02 ix4561 (.Y (nx4560), .A0 (outMuls_6__12), .A1 (nx5284)) ;
    nand02 ix2623 (.Y (addersInputs_6__13), .A0 (nx4563), .A1 (nx4565)) ;
    nand02 ix4564 (.Y (nx4563), .A0 (currentPage_6__13), .A1 (layerType)) ;
    nand02 ix4566 (.Y (nx4565), .A0 (outMuls_6__13), .A1 (nx5286)) ;
    nand02 ix2631 (.Y (addersInputs_6__14), .A0 (nx4568), .A1 (nx4570)) ;
    nand02 ix4569 (.Y (nx4568), .A0 (currentPage_6__14), .A1 (layerType)) ;
    nand02 ix4571 (.Y (nx4570), .A0 (outMuls_6__14), .A1 (nx5286)) ;
    nand02 ix2639 (.Y (addersInputs_6__15), .A0 (nx4573), .A1 (nx4575)) ;
    nand02 ix4574 (.Y (nx4573), .A0 (currentPage_6__15), .A1 (layerType)) ;
    nand02 ix4576 (.Y (nx4575), .A0 (outMuls_6__15), .A1 (nx5286)) ;
    nand02 ix2647 (.Y (addersInputs_5__0), .A0 (nx4578), .A1 (nx4580)) ;
    nand02 ix4579 (.Y (nx4578), .A0 (currentPage_5__0), .A1 (layerType)) ;
    nand02 ix4581 (.Y (nx4580), .A0 (outMuls_5__0), .A1 (nx5286)) ;
    nand02 ix2655 (.Y (addersInputs_5__1), .A0 (nx4583), .A1 (nx4585)) ;
    nand02 ix4584 (.Y (nx4583), .A0 (currentPage_5__1), .A1 (layerType)) ;
    nand02 ix4586 (.Y (nx4585), .A0 (outMuls_5__1), .A1 (nx5286)) ;
    nand02 ix2663 (.Y (addersInputs_5__2), .A0 (nx4588), .A1 (nx4590)) ;
    nand02 ix4589 (.Y (nx4588), .A0 (currentPage_5__2), .A1 (layerType)) ;
    nand02 ix4591 (.Y (nx4590), .A0 (outMuls_5__2), .A1 (nx5286)) ;
    nand02 ix2671 (.Y (addersInputs_5__3), .A0 (nx4593), .A1 (nx4595)) ;
    nand02 ix4594 (.Y (nx4593), .A0 (currentPage_5__3), .A1 (layerType)) ;
    nand02 ix4596 (.Y (nx4595), .A0 (outMuls_5__3), .A1 (nx5286)) ;
    nand02 ix2679 (.Y (addersInputs_5__4), .A0 (nx4598), .A1 (nx4600)) ;
    nand02 ix4599 (.Y (nx4598), .A0 (currentPage_5__4), .A1 (layerType)) ;
    nand02 ix4601 (.Y (nx4600), .A0 (outMuls_5__4), .A1 (nx5288)) ;
    nand02 ix2687 (.Y (addersInputs_5__5), .A0 (nx4603), .A1 (nx4605)) ;
    nand02 ix4604 (.Y (nx4603), .A0 (currentPage_5__5), .A1 (layerType)) ;
    nand02 ix4606 (.Y (nx4605), .A0 (outMuls_5__5), .A1 (nx5288)) ;
    nand02 ix2695 (.Y (addersInputs_5__6), .A0 (nx4608), .A1 (nx4610)) ;
    nand02 ix4609 (.Y (nx4608), .A0 (currentPage_5__6), .A1 (layerType)) ;
    nand02 ix4611 (.Y (nx4610), .A0 (outMuls_5__6), .A1 (nx5288)) ;
    nand02 ix2703 (.Y (addersInputs_5__7), .A0 (nx4613), .A1 (nx4615)) ;
    nand02 ix4614 (.Y (nx4613), .A0 (currentPage_5__7), .A1 (layerType)) ;
    nand02 ix4616 (.Y (nx4615), .A0 (outMuls_5__7), .A1 (nx5288)) ;
    nand02 ix2711 (.Y (addersInputs_5__8), .A0 (nx4618), .A1 (nx4620)) ;
    nand02 ix4619 (.Y (nx4618), .A0 (currentPage_5__8), .A1 (layerType)) ;
    nand02 ix4621 (.Y (nx4620), .A0 (outMuls_5__8), .A1 (nx5288)) ;
    nand02 ix2719 (.Y (addersInputs_5__9), .A0 (nx4623), .A1 (nx4625)) ;
    nand02 ix4624 (.Y (nx4623), .A0 (currentPage_5__9), .A1 (layerType)) ;
    nand02 ix4626 (.Y (nx4625), .A0 (outMuls_5__9), .A1 (nx5288)) ;
    nand02 ix2727 (.Y (addersInputs_5__10), .A0 (nx4628), .A1 (nx4630)) ;
    nand02 ix4629 (.Y (nx4628), .A0 (currentPage_5__10), .A1 (layerType)) ;
    nand02 ix4631 (.Y (nx4630), .A0 (outMuls_5__10), .A1 (nx5288)) ;
    nand02 ix2735 (.Y (addersInputs_5__11), .A0 (nx4633), .A1 (nx4635)) ;
    nand02 ix4634 (.Y (nx4633), .A0 (currentPage_5__11), .A1 (layerType)) ;
    nand02 ix4636 (.Y (nx4635), .A0 (outMuls_5__11), .A1 (nx5290)) ;
    nand02 ix2743 (.Y (addersInputs_5__12), .A0 (nx4638), .A1 (nx4640)) ;
    nand02 ix4639 (.Y (nx4638), .A0 (currentPage_5__12), .A1 (layerType)) ;
    nand02 ix4641 (.Y (nx4640), .A0 (outMuls_5__12), .A1 (nx5290)) ;
    nand02 ix2751 (.Y (addersInputs_5__13), .A0 (nx4643), .A1 (nx4645)) ;
    nand02 ix4644 (.Y (nx4643), .A0 (currentPage_5__13), .A1 (layerType)) ;
    nand02 ix4646 (.Y (nx4645), .A0 (outMuls_5__13), .A1 (nx5290)) ;
    nand02 ix2759 (.Y (addersInputs_5__14), .A0 (nx4648), .A1 (nx4650)) ;
    nand02 ix4649 (.Y (nx4648), .A0 (currentPage_5__14), .A1 (layerType)) ;
    nand02 ix4651 (.Y (nx4650), .A0 (outMuls_5__14), .A1 (nx5290)) ;
    nand02 ix2767 (.Y (addersInputs_5__15), .A0 (nx4653), .A1 (nx4655)) ;
    nand02 ix4654 (.Y (nx4653), .A0 (currentPage_5__15), .A1 (layerType)) ;
    nand02 ix4656 (.Y (nx4655), .A0 (outMuls_5__15), .A1 (nx5290)) ;
    nand02 ix2775 (.Y (addersInputs_4__0), .A0 (nx4658), .A1 (nx4660)) ;
    nand02 ix4659 (.Y (nx4658), .A0 (currentPage_4__0), .A1 (layerType)) ;
    nand02 ix4661 (.Y (nx4660), .A0 (outMuls_4__0), .A1 (nx5290)) ;
    nand02 ix2783 (.Y (addersInputs_4__1), .A0 (nx4663), .A1 (nx4665)) ;
    nand02 ix4664 (.Y (nx4663), .A0 (currentPage_4__1), .A1 (layerType)) ;
    nand02 ix4666 (.Y (nx4665), .A0 (outMuls_4__1), .A1 (nx5290)) ;
    nand02 ix2791 (.Y (addersInputs_4__2), .A0 (nx4668), .A1 (nx4670)) ;
    nand02 ix4669 (.Y (nx4668), .A0 (currentPage_4__2), .A1 (layerType)) ;
    nand02 ix4671 (.Y (nx4670), .A0 (outMuls_4__2), .A1 (nx5292)) ;
    nand02 ix2799 (.Y (addersInputs_4__3), .A0 (nx4673), .A1 (nx4675)) ;
    nand02 ix4674 (.Y (nx4673), .A0 (currentPage_4__3), .A1 (layerType)) ;
    nand02 ix4676 (.Y (nx4675), .A0 (outMuls_4__3), .A1 (nx5292)) ;
    nand02 ix2807 (.Y (addersInputs_4__4), .A0 (nx4678), .A1 (nx4680)) ;
    nand02 ix4679 (.Y (nx4678), .A0 (currentPage_4__4), .A1 (layerType)) ;
    nand02 ix4681 (.Y (nx4680), .A0 (outMuls_4__4), .A1 (nx5292)) ;
    nand02 ix2815 (.Y (addersInputs_4__5), .A0 (nx4683), .A1 (nx4685)) ;
    nand02 ix4684 (.Y (nx4683), .A0 (currentPage_4__5), .A1 (layerType)) ;
    nand02 ix4686 (.Y (nx4685), .A0 (outMuls_4__5), .A1 (nx5292)) ;
    nand02 ix2823 (.Y (addersInputs_4__6), .A0 (nx4688), .A1 (nx4690)) ;
    nand02 ix4689 (.Y (nx4688), .A0 (currentPage_4__6), .A1 (layerType)) ;
    nand02 ix4691 (.Y (nx4690), .A0 (outMuls_4__6), .A1 (nx5292)) ;
    nand02 ix2831 (.Y (addersInputs_4__7), .A0 (nx4693), .A1 (nx4695)) ;
    nand02 ix4694 (.Y (nx4693), .A0 (currentPage_4__7), .A1 (layerType)) ;
    nand02 ix4696 (.Y (nx4695), .A0 (outMuls_4__7), .A1 (nx5292)) ;
    nand02 ix2839 (.Y (addersInputs_4__8), .A0 (nx4698), .A1 (nx4700)) ;
    nand02 ix4699 (.Y (nx4698), .A0 (currentPage_4__8), .A1 (layerType)) ;
    nand02 ix4701 (.Y (nx4700), .A0 (outMuls_4__8), .A1 (nx5292)) ;
    nand02 ix2847 (.Y (addersInputs_4__9), .A0 (nx4703), .A1 (nx4705)) ;
    nand02 ix4704 (.Y (nx4703), .A0 (currentPage_4__9), .A1 (layerType)) ;
    nand02 ix4706 (.Y (nx4705), .A0 (outMuls_4__9), .A1 (nx5294)) ;
    nand02 ix2855 (.Y (addersInputs_4__10), .A0 (nx4708), .A1 (nx4710)) ;
    nand02 ix4709 (.Y (nx4708), .A0 (currentPage_4__10), .A1 (layerType)) ;
    nand02 ix4711 (.Y (nx4710), .A0 (outMuls_4__10), .A1 (nx5294)) ;
    nand02 ix2863 (.Y (addersInputs_4__11), .A0 (nx4713), .A1 (nx4715)) ;
    nand02 ix4714 (.Y (nx4713), .A0 (currentPage_4__11), .A1 (layerType)) ;
    nand02 ix4716 (.Y (nx4715), .A0 (outMuls_4__11), .A1 (nx5294)) ;
    nand02 ix2871 (.Y (addersInputs_4__12), .A0 (nx4718), .A1 (nx4720)) ;
    nand02 ix4719 (.Y (nx4718), .A0 (currentPage_4__12), .A1 (layerType)) ;
    nand02 ix4721 (.Y (nx4720), .A0 (outMuls_4__12), .A1 (nx5294)) ;
    nand02 ix2879 (.Y (addersInputs_4__13), .A0 (nx4723), .A1 (nx4725)) ;
    nand02 ix4724 (.Y (nx4723), .A0 (currentPage_4__13), .A1 (layerType)) ;
    nand02 ix4726 (.Y (nx4725), .A0 (outMuls_4__13), .A1 (nx5294)) ;
    nand02 ix2887 (.Y (addersInputs_4__14), .A0 (nx4728), .A1 (nx4730)) ;
    nand02 ix4729 (.Y (nx4728), .A0 (currentPage_4__14), .A1 (layerType)) ;
    nand02 ix4731 (.Y (nx4730), .A0 (outMuls_4__14), .A1 (nx5294)) ;
    nand02 ix2895 (.Y (addersInputs_4__15), .A0 (nx4733), .A1 (nx4735)) ;
    nand02 ix4734 (.Y (nx4733), .A0 (currentPage_4__15), .A1 (layerType)) ;
    nand02 ix4736 (.Y (nx4735), .A0 (outMuls_4__15), .A1 (nx5294)) ;
    nand02 ix2903 (.Y (addersInputs_3__0), .A0 (nx4738), .A1 (nx4740)) ;
    nand02 ix4739 (.Y (nx4738), .A0 (currentPage_3__0), .A1 (layerType)) ;
    nand02 ix4741 (.Y (nx4740), .A0 (outMuls_3__0), .A1 (nx5296)) ;
    nand02 ix2911 (.Y (addersInputs_3__1), .A0 (nx4743), .A1 (nx4745)) ;
    nand02 ix4744 (.Y (nx4743), .A0 (currentPage_3__1), .A1 (layerType)) ;
    nand02 ix4746 (.Y (nx4745), .A0 (outMuls_3__1), .A1 (nx5296)) ;
    nand02 ix2919 (.Y (addersInputs_3__2), .A0 (nx4748), .A1 (nx4750)) ;
    nand02 ix4749 (.Y (nx4748), .A0 (currentPage_3__2), .A1 (layerType)) ;
    nand02 ix4751 (.Y (nx4750), .A0 (outMuls_3__2), .A1 (nx5296)) ;
    nand02 ix2927 (.Y (addersInputs_3__3), .A0 (nx4753), .A1 (nx4755)) ;
    nand02 ix4754 (.Y (nx4753), .A0 (currentPage_3__3), .A1 (layerType)) ;
    nand02 ix4756 (.Y (nx4755), .A0 (outMuls_3__3), .A1 (nx5296)) ;
    nand02 ix2935 (.Y (addersInputs_3__4), .A0 (nx4758), .A1 (nx4760)) ;
    nand02 ix4759 (.Y (nx4758), .A0 (currentPage_3__4), .A1 (layerType)) ;
    nand02 ix4761 (.Y (nx4760), .A0 (outMuls_3__4), .A1 (nx5296)) ;
    nand02 ix2943 (.Y (addersInputs_3__5), .A0 (nx4763), .A1 (nx4765)) ;
    nand02 ix4764 (.Y (nx4763), .A0 (currentPage_3__5), .A1 (layerType)) ;
    nand02 ix4766 (.Y (nx4765), .A0 (outMuls_3__5), .A1 (nx5296)) ;
    nand02 ix2951 (.Y (addersInputs_3__6), .A0 (nx4768), .A1 (nx4770)) ;
    nand02 ix4769 (.Y (nx4768), .A0 (currentPage_3__6), .A1 (layerType)) ;
    nand02 ix4771 (.Y (nx4770), .A0 (outMuls_3__6), .A1 (nx5296)) ;
    nand02 ix2959 (.Y (addersInputs_3__7), .A0 (nx4773), .A1 (nx4775)) ;
    nand02 ix4774 (.Y (nx4773), .A0 (currentPage_3__7), .A1 (layerType)) ;
    nand02 ix4776 (.Y (nx4775), .A0 (outMuls_3__7), .A1 (nx5298)) ;
    nand02 ix2967 (.Y (addersInputs_3__8), .A0 (nx4778), .A1 (nx4780)) ;
    nand02 ix4779 (.Y (nx4778), .A0 (currentPage_3__8), .A1 (layerType)) ;
    nand02 ix4781 (.Y (nx4780), .A0 (outMuls_3__8), .A1 (nx5298)) ;
    nand02 ix2975 (.Y (addersInputs_3__9), .A0 (nx4783), .A1 (nx4785)) ;
    nand02 ix4784 (.Y (nx4783), .A0 (currentPage_3__9), .A1 (layerType)) ;
    nand02 ix4786 (.Y (nx4785), .A0 (outMuls_3__9), .A1 (nx5298)) ;
    nand02 ix2983 (.Y (addersInputs_3__10), .A0 (nx4788), .A1 (nx4790)) ;
    nand02 ix4789 (.Y (nx4788), .A0 (currentPage_3__10), .A1 (layerType)) ;
    nand02 ix4791 (.Y (nx4790), .A0 (outMuls_3__10), .A1 (nx5298)) ;
    nand02 ix2991 (.Y (addersInputs_3__11), .A0 (nx4793), .A1 (nx4795)) ;
    nand02 ix4794 (.Y (nx4793), .A0 (currentPage_3__11), .A1 (layerType)) ;
    nand02 ix4796 (.Y (nx4795), .A0 (outMuls_3__11), .A1 (nx5298)) ;
    nand02 ix2999 (.Y (addersInputs_3__12), .A0 (nx4798), .A1 (nx4800)) ;
    nand02 ix4799 (.Y (nx4798), .A0 (currentPage_3__12), .A1 (layerType)) ;
    nand02 ix4801 (.Y (nx4800), .A0 (outMuls_3__12), .A1 (nx5298)) ;
    nand02 ix3007 (.Y (addersInputs_3__13), .A0 (nx4803), .A1 (nx4805)) ;
    nand02 ix4804 (.Y (nx4803), .A0 (currentPage_3__13), .A1 (layerType)) ;
    nand02 ix4806 (.Y (nx4805), .A0 (outMuls_3__13), .A1 (nx5298)) ;
    nand02 ix3015 (.Y (addersInputs_3__14), .A0 (nx4808), .A1 (nx4810)) ;
    nand02 ix4809 (.Y (nx4808), .A0 (currentPage_3__14), .A1 (layerType)) ;
    nand02 ix4811 (.Y (nx4810), .A0 (outMuls_3__14), .A1 (nx5300)) ;
    nand02 ix3023 (.Y (addersInputs_3__15), .A0 (nx4813), .A1 (nx4815)) ;
    nand02 ix4814 (.Y (nx4813), .A0 (currentPage_3__15), .A1 (layerType)) ;
    nand02 ix4816 (.Y (nx4815), .A0 (outMuls_3__15), .A1 (nx5300)) ;
    nand02 ix3031 (.Y (addersInputs_2__0), .A0 (nx4818), .A1 (nx4820)) ;
    nand02 ix4819 (.Y (nx4818), .A0 (currentPage_2__0), .A1 (layerType)) ;
    nand02 ix4821 (.Y (nx4820), .A0 (outMuls_2__0), .A1 (nx5300)) ;
    nand02 ix3039 (.Y (addersInputs_2__1), .A0 (nx4823), .A1 (nx4825)) ;
    nand02 ix4824 (.Y (nx4823), .A0 (currentPage_2__1), .A1 (layerType)) ;
    nand02 ix4826 (.Y (nx4825), .A0 (outMuls_2__1), .A1 (nx5300)) ;
    nand02 ix3047 (.Y (addersInputs_2__2), .A0 (nx4828), .A1 (nx4830)) ;
    nand02 ix4829 (.Y (nx4828), .A0 (currentPage_2__2), .A1 (layerType)) ;
    nand02 ix4831 (.Y (nx4830), .A0 (outMuls_2__2), .A1 (nx5300)) ;
    nand02 ix3055 (.Y (addersInputs_2__3), .A0 (nx4833), .A1 (nx4835)) ;
    nand02 ix4834 (.Y (nx4833), .A0 (currentPage_2__3), .A1 (layerType)) ;
    nand02 ix4836 (.Y (nx4835), .A0 (outMuls_2__3), .A1 (nx5300)) ;
    nand02 ix3063 (.Y (addersInputs_2__4), .A0 (nx4838), .A1 (nx4840)) ;
    nand02 ix4839 (.Y (nx4838), .A0 (currentPage_2__4), .A1 (layerType)) ;
    nand02 ix4841 (.Y (nx4840), .A0 (outMuls_2__4), .A1 (nx5300)) ;
    nand02 ix3071 (.Y (addersInputs_2__5), .A0 (nx4843), .A1 (nx4845)) ;
    nand02 ix4844 (.Y (nx4843), .A0 (currentPage_2__5), .A1 (layerType)) ;
    nand02 ix4846 (.Y (nx4845), .A0 (outMuls_2__5), .A1 (nx5302)) ;
    nand02 ix3079 (.Y (addersInputs_2__6), .A0 (nx4848), .A1 (nx4850)) ;
    nand02 ix4849 (.Y (nx4848), .A0 (currentPage_2__6), .A1 (layerType)) ;
    nand02 ix4851 (.Y (nx4850), .A0 (outMuls_2__6), .A1 (nx5302)) ;
    nand02 ix3087 (.Y (addersInputs_2__7), .A0 (nx4853), .A1 (nx4855)) ;
    nand02 ix4854 (.Y (nx4853), .A0 (currentPage_2__7), .A1 (layerType)) ;
    nand02 ix4856 (.Y (nx4855), .A0 (outMuls_2__7), .A1 (nx5302)) ;
    nand02 ix3095 (.Y (addersInputs_2__8), .A0 (nx4858), .A1 (nx4860)) ;
    nand02 ix4859 (.Y (nx4858), .A0 (currentPage_2__8), .A1 (layerType)) ;
    nand02 ix4861 (.Y (nx4860), .A0 (outMuls_2__8), .A1 (nx5302)) ;
    nand02 ix3103 (.Y (addersInputs_2__9), .A0 (nx4863), .A1 (nx4865)) ;
    nand02 ix4864 (.Y (nx4863), .A0 (currentPage_2__9), .A1 (layerType)) ;
    nand02 ix4866 (.Y (nx4865), .A0 (outMuls_2__9), .A1 (nx5302)) ;
    nand02 ix3111 (.Y (addersInputs_2__10), .A0 (nx4868), .A1 (nx4870)) ;
    nand02 ix4869 (.Y (nx4868), .A0 (currentPage_2__10), .A1 (layerType)) ;
    nand02 ix4871 (.Y (nx4870), .A0 (outMuls_2__10), .A1 (nx5302)) ;
    nand02 ix3119 (.Y (addersInputs_2__11), .A0 (nx4873), .A1 (nx4875)) ;
    nand02 ix4874 (.Y (nx4873), .A0 (currentPage_2__11), .A1 (layerType)) ;
    nand02 ix4876 (.Y (nx4875), .A0 (outMuls_2__11), .A1 (nx5302)) ;
    nand02 ix3127 (.Y (addersInputs_2__12), .A0 (nx4878), .A1 (nx4880)) ;
    nand02 ix4879 (.Y (nx4878), .A0 (currentPage_2__12), .A1 (layerType)) ;
    nand02 ix4881 (.Y (nx4880), .A0 (outMuls_2__12), .A1 (nx5304)) ;
    nand02 ix3135 (.Y (addersInputs_2__13), .A0 (nx4883), .A1 (nx4885)) ;
    nand02 ix4884 (.Y (nx4883), .A0 (currentPage_2__13), .A1 (layerType)) ;
    nand02 ix4886 (.Y (nx4885), .A0 (outMuls_2__13), .A1 (nx5304)) ;
    nand02 ix3143 (.Y (addersInputs_2__14), .A0 (nx4888), .A1 (nx4890)) ;
    nand02 ix4889 (.Y (nx4888), .A0 (currentPage_2__14), .A1 (layerType)) ;
    nand02 ix4891 (.Y (nx4890), .A0 (outMuls_2__14), .A1 (nx5304)) ;
    nand02 ix3151 (.Y (addersInputs_2__15), .A0 (nx4893), .A1 (nx4895)) ;
    nand02 ix4894 (.Y (nx4893), .A0 (currentPage_2__15), .A1 (layerType)) ;
    nand02 ix4896 (.Y (nx4895), .A0 (outMuls_2__15), .A1 (nx5304)) ;
    nand02 ix3159 (.Y (addersInputs_1__0), .A0 (nx4898), .A1 (nx4900)) ;
    nand02 ix4899 (.Y (nx4898), .A0 (currentPage_1__0), .A1 (layerType)) ;
    nand02 ix4901 (.Y (nx4900), .A0 (outMuls_1__0), .A1 (nx5304)) ;
    nand02 ix3167 (.Y (addersInputs_1__1), .A0 (nx4903), .A1 (nx4905)) ;
    nand02 ix4904 (.Y (nx4903), .A0 (currentPage_1__1), .A1 (layerType)) ;
    nand02 ix4906 (.Y (nx4905), .A0 (outMuls_1__1), .A1 (nx5304)) ;
    nand02 ix3175 (.Y (addersInputs_1__2), .A0 (nx4908), .A1 (nx4910)) ;
    nand02 ix4909 (.Y (nx4908), .A0 (currentPage_1__2), .A1 (layerType)) ;
    nand02 ix4911 (.Y (nx4910), .A0 (outMuls_1__2), .A1 (nx5304)) ;
    nand02 ix3183 (.Y (addersInputs_1__3), .A0 (nx4913), .A1 (nx4915)) ;
    nand02 ix4914 (.Y (nx4913), .A0 (currentPage_1__3), .A1 (layerType)) ;
    nand02 ix4916 (.Y (nx4915), .A0 (outMuls_1__3), .A1 (nx5306)) ;
    nand02 ix3191 (.Y (addersInputs_1__4), .A0 (nx4918), .A1 (nx4920)) ;
    nand02 ix4919 (.Y (nx4918), .A0 (currentPage_1__4), .A1 (layerType)) ;
    nand02 ix4921 (.Y (nx4920), .A0 (outMuls_1__4), .A1 (nx5306)) ;
    nand02 ix3199 (.Y (addersInputs_1__5), .A0 (nx4923), .A1 (nx4925)) ;
    nand02 ix4924 (.Y (nx4923), .A0 (currentPage_1__5), .A1 (layerType)) ;
    nand02 ix4926 (.Y (nx4925), .A0 (outMuls_1__5), .A1 (nx5306)) ;
    nand02 ix3207 (.Y (addersInputs_1__6), .A0 (nx4928), .A1 (nx4930)) ;
    nand02 ix4929 (.Y (nx4928), .A0 (currentPage_1__6), .A1 (layerType)) ;
    nand02 ix4931 (.Y (nx4930), .A0 (outMuls_1__6), .A1 (nx5306)) ;
    nand02 ix3215 (.Y (addersInputs_1__7), .A0 (nx4933), .A1 (nx4935)) ;
    nand02 ix4934 (.Y (nx4933), .A0 (currentPage_1__7), .A1 (layerType)) ;
    nand02 ix4936 (.Y (nx4935), .A0 (outMuls_1__7), .A1 (nx5306)) ;
    nand02 ix3223 (.Y (addersInputs_1__8), .A0 (nx4938), .A1 (nx4940)) ;
    nand02 ix4939 (.Y (nx4938), .A0 (currentPage_1__8), .A1 (layerType)) ;
    nand02 ix4941 (.Y (nx4940), .A0 (outMuls_1__8), .A1 (nx5306)) ;
    nand02 ix3231 (.Y (addersInputs_1__9), .A0 (nx4943), .A1 (nx4945)) ;
    nand02 ix4944 (.Y (nx4943), .A0 (currentPage_1__9), .A1 (layerType)) ;
    nand02 ix4946 (.Y (nx4945), .A0 (outMuls_1__9), .A1 (nx5306)) ;
    nand02 ix3239 (.Y (addersInputs_1__10), .A0 (nx4948), .A1 (nx4950)) ;
    nand02 ix4949 (.Y (nx4948), .A0 (currentPage_1__10), .A1 (layerType)) ;
    nand02 ix4951 (.Y (nx4950), .A0 (outMuls_1__10), .A1 (nx5308)) ;
    nand02 ix3247 (.Y (addersInputs_1__11), .A0 (nx4953), .A1 (nx4955)) ;
    nand02 ix4954 (.Y (nx4953), .A0 (currentPage_1__11), .A1 (layerType)) ;
    nand02 ix4956 (.Y (nx4955), .A0 (outMuls_1__11), .A1 (nx5308)) ;
    nand02 ix3255 (.Y (addersInputs_1__12), .A0 (nx4958), .A1 (nx4960)) ;
    nand02 ix4959 (.Y (nx4958), .A0 (currentPage_1__12), .A1 (layerType)) ;
    nand02 ix4961 (.Y (nx4960), .A0 (outMuls_1__12), .A1 (nx5308)) ;
    nand02 ix3263 (.Y (addersInputs_1__13), .A0 (nx4963), .A1 (nx4965)) ;
    nand02 ix4964 (.Y (nx4963), .A0 (currentPage_1__13), .A1 (layerType)) ;
    nand02 ix4966 (.Y (nx4965), .A0 (outMuls_1__13), .A1 (nx5308)) ;
    nand02 ix3271 (.Y (addersInputs_1__14), .A0 (nx4968), .A1 (nx4970)) ;
    nand02 ix4969 (.Y (nx4968), .A0 (currentPage_1__14), .A1 (layerType)) ;
    nand02 ix4971 (.Y (nx4970), .A0 (outMuls_1__14), .A1 (nx5308)) ;
    nand02 ix3279 (.Y (addersInputs_1__15), .A0 (nx4973), .A1 (nx4975)) ;
    nand02 ix4974 (.Y (nx4973), .A0 (currentPage_1__15), .A1 (layerType)) ;
    nand02 ix4976 (.Y (nx4975), .A0 (outMuls_1__15), .A1 (nx5308)) ;
    nand02 ix3287 (.Y (addersInputs_0__0), .A0 (nx4978), .A1 (nx4980)) ;
    nand02 ix4979 (.Y (nx4978), .A0 (currentPage_0__0), .A1 (layerType)) ;
    nand02 ix4981 (.Y (nx4980), .A0 (outMuls_0__0), .A1 (nx5308)) ;
    nand02 ix3295 (.Y (addersInputs_0__1), .A0 (nx4983), .A1 (nx4985)) ;
    nand02 ix4984 (.Y (nx4983), .A0 (currentPage_0__1), .A1 (layerType)) ;
    nand02 ix4986 (.Y (nx4985), .A0 (outMuls_0__1), .A1 (nx5310)) ;
    nand02 ix3303 (.Y (addersInputs_0__2), .A0 (nx4988), .A1 (nx4990)) ;
    nand02 ix4989 (.Y (nx4988), .A0 (currentPage_0__2), .A1 (layerType)) ;
    nand02 ix4991 (.Y (nx4990), .A0 (outMuls_0__2), .A1 (nx5310)) ;
    nand02 ix3311 (.Y (addersInputs_0__3), .A0 (nx4993), .A1 (nx4995)) ;
    nand02 ix4994 (.Y (nx4993), .A0 (currentPage_0__3), .A1 (layerType)) ;
    nand02 ix4996 (.Y (nx4995), .A0 (outMuls_0__3), .A1 (nx5310)) ;
    nand02 ix3319 (.Y (addersInputs_0__4), .A0 (nx4998), .A1 (nx5000)) ;
    nand02 ix4999 (.Y (nx4998), .A0 (currentPage_0__4), .A1 (layerType)) ;
    nand02 ix5001 (.Y (nx5000), .A0 (outMuls_0__4), .A1 (nx5310)) ;
    nand02 ix3327 (.Y (addersInputs_0__5), .A0 (nx5003), .A1 (nx5005)) ;
    nand02 ix5004 (.Y (nx5003), .A0 (currentPage_0__5), .A1 (layerType)) ;
    nand02 ix5006 (.Y (nx5005), .A0 (outMuls_0__5), .A1 (nx5310)) ;
    nand02 ix3335 (.Y (addersInputs_0__6), .A0 (nx5008), .A1 (nx5010)) ;
    nand02 ix5009 (.Y (nx5008), .A0 (currentPage_0__6), .A1 (layerType)) ;
    nand02 ix5011 (.Y (nx5010), .A0 (outMuls_0__6), .A1 (nx5310)) ;
    nand02 ix3343 (.Y (addersInputs_0__7), .A0 (nx5013), .A1 (nx5015)) ;
    nand02 ix5014 (.Y (nx5013), .A0 (currentPage_0__7), .A1 (layerType)) ;
    nand02 ix5016 (.Y (nx5015), .A0 (outMuls_0__7), .A1 (nx5310)) ;
    nand02 ix3351 (.Y (addersInputs_0__8), .A0 (nx5018), .A1 (nx5020)) ;
    nand02 ix5019 (.Y (nx5018), .A0 (currentPage_0__8), .A1 (layerType)) ;
    nand02 ix5021 (.Y (nx5020), .A0 (outMuls_0__8), .A1 (nx5312)) ;
    nand02 ix3359 (.Y (addersInputs_0__9), .A0 (nx5023), .A1 (nx5025)) ;
    nand02 ix5024 (.Y (nx5023), .A0 (currentPage_0__9), .A1 (layerType)) ;
    nand02 ix5026 (.Y (nx5025), .A0 (outMuls_0__9), .A1 (nx5312)) ;
    nand02 ix3367 (.Y (addersInputs_0__10), .A0 (nx5028), .A1 (nx5030)) ;
    nand02 ix5029 (.Y (nx5028), .A0 (currentPage_0__10), .A1 (layerType)) ;
    nand02 ix5031 (.Y (nx5030), .A0 (outMuls_0__10), .A1 (nx5312)) ;
    nand02 ix3375 (.Y (addersInputs_0__11), .A0 (nx5033), .A1 (nx5035)) ;
    nand02 ix5034 (.Y (nx5033), .A0 (currentPage_0__11), .A1 (layerType)) ;
    nand02 ix5036 (.Y (nx5035), .A0 (outMuls_0__11), .A1 (nx5312)) ;
    nand02 ix3383 (.Y (addersInputs_0__12), .A0 (nx5038), .A1 (nx5040)) ;
    nand02 ix5039 (.Y (nx5038), .A0 (currentPage_0__12), .A1 (layerType)) ;
    nand02 ix5041 (.Y (nx5040), .A0 (outMuls_0__12), .A1 (nx5312)) ;
    nand02 ix3391 (.Y (addersInputs_0__13), .A0 (nx5043), .A1 (nx5045)) ;
    nand02 ix5044 (.Y (nx5043), .A0 (currentPage_0__13), .A1 (layerType)) ;
    nand02 ix5046 (.Y (nx5045), .A0 (outMuls_0__13), .A1 (nx5312)) ;
    nand02 ix3399 (.Y (addersInputs_0__14), .A0 (nx5048), .A1 (nx5050)) ;
    nand02 ix5049 (.Y (nx5048), .A0 (currentPage_0__14), .A1 (layerType)) ;
    nand02 ix5051 (.Y (nx5050), .A0 (outMuls_0__14), .A1 (nx5312)) ;
    nand02 ix3407 (.Y (addersInputs_0__15), .A0 (nx5053), .A1 (nx5055)) ;
    nand02 ix5054 (.Y (nx5053), .A0 (currentPage_0__15), .A1 (layerType)) ;
    nand02 ix5056 (.Y (nx5055), .A0 (outMuls_0__15), .A1 (nx5314)) ;
    nand04 ix47 (.Y (finalSum[0]), .A0 (nx5058), .A1 (nx5060), .A2 (nx5063), .A3 (
           nx5067)) ;
    nand03 ix5059 (.Y (nx5058), .A0 (addersMap_totalSum_0), .A1 (filterType), .A2 (
           nx5314)) ;
    nand02 ix5061 (.Y (nx5060), .A0 (addersMap_sum3Filter_0), .A1 (nx5196)) ;
    nor02_2x ix5 (.Y (nx4), .A0 (filterType), .A1 (layerType)) ;
    nand03 ix5064 (.Y (nx5063), .A0 (addersMap_sum3Filter_3), .A1 (nx5320), .A2 (
           layerType)) ;
    nand03 ix5068 (.Y (nx5067), .A0 (addersMap_totalSum_5), .A1 (filterType), .A2 (
           layerType)) ;
    nand04 ix61 (.Y (finalSum[1]), .A0 (nx5070), .A1 (nx5072), .A2 (nx5074), .A3 (
           nx5076)) ;
    nand03 ix5071 (.Y (nx5070), .A0 (addersMap_totalSum_1), .A1 (filterType), .A2 (
           nx5314)) ;
    nand02 ix5073 (.Y (nx5072), .A0 (addersMap_sum3Filter_1), .A1 (nx5196)) ;
    nand03 ix5075 (.Y (nx5074), .A0 (addersMap_sum3Filter_4), .A1 (nx5320), .A2 (
           layerType)) ;
    nand03 ix5077 (.Y (nx5076), .A0 (addersMap_totalSum_6), .A1 (filterType), .A2 (
           layerType)) ;
    nand04 ix75 (.Y (finalSum[2]), .A0 (nx5079), .A1 (nx5081), .A2 (nx5083), .A3 (
           nx5085)) ;
    nand03 ix5080 (.Y (nx5079), .A0 (addersMap_totalSum_2), .A1 (filterType), .A2 (
           nx5314)) ;
    nand02 ix5082 (.Y (nx5081), .A0 (addersMap_sum3Filter_2), .A1 (nx5196)) ;
    nand03 ix5084 (.Y (nx5083), .A0 (addersMap_sum3Filter_5), .A1 (nx5320), .A2 (
           layerType)) ;
    nand03 ix5086 (.Y (nx5085), .A0 (addersMap_totalSum_7), .A1 (filterType), .A2 (
           layerType)) ;
    nand04 ix89 (.Y (finalSum[3]), .A0 (nx5088), .A1 (nx5090), .A2 (nx5092), .A3 (
           nx5094)) ;
    nand03 ix5089 (.Y (nx5088), .A0 (addersMap_totalSum_3), .A1 (filterType), .A2 (
           nx5314)) ;
    nand02 ix5091 (.Y (nx5090), .A0 (addersMap_sum3Filter_3), .A1 (nx5196)) ;
    nand03 ix5093 (.Y (nx5092), .A0 (addersMap_sum3Filter_6), .A1 (nx5320), .A2 (
           layerType)) ;
    nand03 ix5095 (.Y (nx5094), .A0 (addersMap_totalSum_8), .A1 (filterType), .A2 (
           layerType)) ;
    nand04 ix103 (.Y (finalSum[4]), .A0 (nx5097), .A1 (nx5099), .A2 (nx5101), .A3 (
           nx5103)) ;
    nand03 ix5098 (.Y (nx5097), .A0 (addersMap_totalSum_4), .A1 (filterType), .A2 (
           nx5314)) ;
    nand02 ix5100 (.Y (nx5099), .A0 (addersMap_sum3Filter_4), .A1 (nx5196)) ;
    nand03 ix5102 (.Y (nx5101), .A0 (addersMap_sum3Filter_7), .A1 (nx5320), .A2 (
           layerType)) ;
    nand03 ix5104 (.Y (nx5103), .A0 (addersMap_totalSum_9), .A1 (filterType), .A2 (
           layerType)) ;
    nand04 ix117 (.Y (finalSum[5]), .A0 (nx5106), .A1 (nx5108), .A2 (nx5110), .A3 (
           nx5112)) ;
    nand03 ix5107 (.Y (nx5106), .A0 (addersMap_totalSum_5), .A1 (filterType), .A2 (
           nx5314)) ;
    nand02 ix5109 (.Y (nx5108), .A0 (addersMap_sum3Filter_5), .A1 (nx5196)) ;
    nand03 ix5111 (.Y (nx5110), .A0 (addersMap_sum3Filter_8), .A1 (nx5320), .A2 (
           layerType)) ;
    nand03 ix5113 (.Y (nx5112), .A0 (addersMap_totalSum_10), .A1 (filterType), .A2 (
           layerType)) ;
    nand04 ix131 (.Y (finalSum[6]), .A0 (nx5115), .A1 (nx5117), .A2 (nx5119), .A3 (
           nx5121)) ;
    nand03 ix5116 (.Y (nx5115), .A0 (addersMap_totalSum_6), .A1 (filterType), .A2 (
           nx5316)) ;
    nand02 ix5118 (.Y (nx5117), .A0 (addersMap_sum3Filter_6), .A1 (nx5196)) ;
    nand03 ix5120 (.Y (nx5119), .A0 (addersMap_sum3Filter_9), .A1 (nx5320), .A2 (
           layerType)) ;
    nand03 ix5122 (.Y (nx5121), .A0 (addersMap_totalSum_11), .A1 (filterType), .A2 (
           layerType)) ;
    nand04 ix145 (.Y (finalSum[7]), .A0 (nx5124), .A1 (nx5126), .A2 (nx5128), .A3 (
           nx5130)) ;
    nand03 ix5125 (.Y (nx5124), .A0 (addersMap_totalSum_7), .A1 (filterType), .A2 (
           nx5316)) ;
    nand02 ix5127 (.Y (nx5126), .A0 (addersMap_sum3Filter_7), .A1 (nx5198)) ;
    nand03 ix5129 (.Y (nx5128), .A0 (addersMap_sum3Filter_10), .A1 (nx5322), .A2 (
           layerType)) ;
    nand03 ix5131 (.Y (nx5130), .A0 (addersMap_totalSum_12), .A1 (filterType), .A2 (
           layerType)) ;
    nand04 ix159 (.Y (finalSum[8]), .A0 (nx5133), .A1 (nx5135), .A2 (nx5137), .A3 (
           nx5139)) ;
    nand03 ix5134 (.Y (nx5133), .A0 (addersMap_totalSum_8), .A1 (filterType), .A2 (
           nx5316)) ;
    nand02 ix5136 (.Y (nx5135), .A0 (addersMap_sum3Filter_8), .A1 (nx5198)) ;
    nand03 ix5138 (.Y (nx5137), .A0 (addersMap_sum3Filter_11), .A1 (nx5322), .A2 (
           layerType)) ;
    nand03 ix5140 (.Y (nx5139), .A0 (addersMap_totalSum_13), .A1 (filterType), .A2 (
           layerType)) ;
    nand04 ix173 (.Y (finalSum[9]), .A0 (nx5142), .A1 (nx5144), .A2 (nx5146), .A3 (
           nx5148)) ;
    nand03 ix5143 (.Y (nx5142), .A0 (addersMap_totalSum_9), .A1 (filterType), .A2 (
           nx5316)) ;
    nand02 ix5145 (.Y (nx5144), .A0 (addersMap_sum3Filter_9), .A1 (nx5198)) ;
    nand03 ix5147 (.Y (nx5146), .A0 (addersMap_sum3Filter_12), .A1 (nx5322), .A2 (
           layerType)) ;
    nand03 ix5149 (.Y (nx5148), .A0 (addersMap_totalSum_14), .A1 (filterType), .A2 (
           layerType)) ;
    nand04 ix187 (.Y (finalSum[10]), .A0 (nx5151), .A1 (nx5153), .A2 (nx5155), .A3 (
           nx5157)) ;
    nand03 ix5152 (.Y (nx5151), .A0 (addersMap_totalSum_10), .A1 (filterType), .A2 (
           nx5316)) ;
    nand02 ix5154 (.Y (nx5153), .A0 (addersMap_sum3Filter_10), .A1 (nx5198)) ;
    nand03 ix5156 (.Y (nx5155), .A0 (addersMap_sum3Filter_13), .A1 (nx5322), .A2 (
           layerType)) ;
    nand03 ix5158 (.Y (nx5157), .A0 (addersMap_totalSum_15), .A1 (filterType), .A2 (
           layerType)) ;
    nand03 ix197 (.Y (finalSum[11]), .A0 (nx5160), .A1 (nx5162), .A2 (nx5164)) ;
    nand02 ix5161 (.Y (nx5160), .A0 (addersMap_sum3Filter_11), .A1 (nx5198)) ;
    nand03 ix5163 (.Y (nx5162), .A0 (addersMap_sum3Filter_14), .A1 (nx5322), .A2 (
           layerType)) ;
    nand03 ix5165 (.Y (nx5164), .A0 (addersMap_totalSum_11), .A1 (filterType), .A2 (
           nx5316)) ;
    nand03 ix207 (.Y (finalSum[12]), .A0 (nx5167), .A1 (nx5169), .A2 (nx5171)) ;
    nand02 ix5168 (.Y (nx5167), .A0 (addersMap_sum3Filter_12), .A1 (nx5198)) ;
    nand03 ix5170 (.Y (nx5169), .A0 (addersMap_sum3Filter_15), .A1 (nx5322), .A2 (
           layerType)) ;
    nand03 ix5172 (.Y (nx5171), .A0 (addersMap_totalSum_12), .A1 (filterType), .A2 (
           nx5316)) ;
    nand02 ix15 (.Y (finalSum[13]), .A0 (nx5174), .A1 (nx5176)) ;
    nand03 ix5175 (.Y (nx5174), .A0 (addersMap_totalSum_13), .A1 (filterType), .A2 (
           nx5318)) ;
    nand02 ix5177 (.Y (nx5176), .A0 (addersMap_sum3Filter_13), .A1 (nx5198)) ;
    nand02 ix21 (.Y (finalSum[14]), .A0 (nx5179), .A1 (nx5181)) ;
    nand03 ix5180 (.Y (nx5179), .A0 (addersMap_totalSum_14), .A1 (filterType), .A2 (
           nx5318)) ;
    nand02 ix5182 (.Y (nx5181), .A0 (addersMap_sum3Filter_14), .A1 (nx4)) ;
    nand02 ix27 (.Y (finalSum[15]), .A0 (nx5184), .A1 (nx5186)) ;
    nand03 ix5185 (.Y (nx5184), .A0 (addersMap_totalSum_15), .A1 (filterType), .A2 (
           nx5318)) ;
    nand02 ix5187 (.Y (nx5186), .A0 (addersMap_sum3Filter_15), .A1 (nx4)) ;
    inv01 ix3481 (.Y (done), .A (nx5189)) ;
    nor02_2x ix5190 (.Y (nx5189), .A0 (layerType), .A1 (doneMul)) ;
    nor02_2x ix5195 (.Y (nx5196), .A0 (filterType), .A1 (layerType)) ;
    nor02_2x ix5197 (.Y (nx5198), .A0 (filterType), .A1 (layerType)) ;
    inv02 ix5199 (.Y (nx5200), .A (layerType)) ;
    inv02 ix5201 (.Y (nx5202), .A (layerType)) ;
    inv02 ix5203 (.Y (nx5204), .A (layerType)) ;
    inv02 ix5205 (.Y (nx5206), .A (layerType)) ;
    inv02 ix5207 (.Y (nx5208), .A (layerType)) ;
    inv02 ix5209 (.Y (nx5210), .A (layerType)) ;
    inv02 ix5211 (.Y (nx5212), .A (layerType)) ;
    inv02 ix5213 (.Y (nx5214), .A (layerType)) ;
    inv02 ix5215 (.Y (nx5216), .A (layerType)) ;
    inv02 ix5217 (.Y (nx5218), .A (layerType)) ;
    inv02 ix5219 (.Y (nx5220), .A (layerType)) ;
    inv02 ix5221 (.Y (nx5222), .A (layerType)) ;
    inv02 ix5223 (.Y (nx5224), .A (layerType)) ;
    inv02 ix5225 (.Y (nx5226), .A (layerType)) ;
    inv02 ix5227 (.Y (nx5228), .A (layerType)) ;
    inv02 ix5229 (.Y (nx5230), .A (layerType)) ;
    inv02 ix5231 (.Y (nx5232), .A (layerType)) ;
    inv02 ix5233 (.Y (nx5234), .A (layerType)) ;
    inv02 ix5235 (.Y (nx5236), .A (layerType)) ;
    inv02 ix5237 (.Y (nx5238), .A (layerType)) ;
    inv02 ix5239 (.Y (nx5240), .A (layerType)) ;
    inv02 ix5241 (.Y (nx5242), .A (layerType)) ;
    inv02 ix5243 (.Y (nx5244), .A (layerType)) ;
    inv02 ix5245 (.Y (nx5246), .A (layerType)) ;
    inv02 ix5247 (.Y (nx5248), .A (layerType)) ;
    inv02 ix5249 (.Y (nx5250), .A (layerType)) ;
    inv02 ix5251 (.Y (nx5252), .A (layerType)) ;
    inv02 ix5253 (.Y (nx5254), .A (layerType)) ;
    inv02 ix5255 (.Y (nx5256), .A (layerType)) ;
    inv02 ix5257 (.Y (nx5258), .A (layerType)) ;
    inv02 ix5259 (.Y (nx5260), .A (layerType)) ;
    inv02 ix5261 (.Y (nx5262), .A (layerType)) ;
    inv02 ix5263 (.Y (nx5264), .A (layerType)) ;
    inv02 ix5265 (.Y (nx5266), .A (layerType)) ;
    inv02 ix5267 (.Y (nx5268), .A (layerType)) ;
    inv02 ix5269 (.Y (nx5270), .A (layerType)) ;
    inv02 ix5271 (.Y (nx5272), .A (layerType)) ;
    inv02 ix5273 (.Y (nx5274), .A (layerType)) ;
    inv02 ix5275 (.Y (nx5276), .A (layerType)) ;
    inv02 ix5277 (.Y (nx5278), .A (layerType)) ;
    inv02 ix5279 (.Y (nx5280), .A (layerType)) ;
    inv02 ix5281 (.Y (nx5282), .A (layerType)) ;
    inv02 ix5283 (.Y (nx5284), .A (layerType)) ;
    inv02 ix5285 (.Y (nx5286), .A (layerType)) ;
    inv02 ix5287 (.Y (nx5288), .A (layerType)) ;
    inv02 ix5289 (.Y (nx5290), .A (layerType)) ;
    inv02 ix5291 (.Y (nx5292), .A (layerType)) ;
    inv02 ix5293 (.Y (nx5294), .A (layerType)) ;
    inv02 ix5295 (.Y (nx5296), .A (layerType)) ;
    inv02 ix5297 (.Y (nx5298), .A (layerType)) ;
    inv02 ix5299 (.Y (nx5300), .A (layerType)) ;
    inv02 ix5301 (.Y (nx5302), .A (layerType)) ;
    inv02 ix5303 (.Y (nx5304), .A (layerType)) ;
    inv02 ix5305 (.Y (nx5306), .A (layerType)) ;
    inv02 ix5307 (.Y (nx5308), .A (layerType)) ;
    inv02 ix5309 (.Y (nx5310), .A (layerType)) ;
    inv02 ix5311 (.Y (nx5312), .A (layerType)) ;
    inv02 ix5313 (.Y (nx5314), .A (layerType)) ;
    inv02 ix5315 (.Y (nx5316), .A (layerType)) ;
    inv02 ix5317 (.Y (nx5318), .A (layerType)) ;
    inv02 ix5319 (.Y (nx5320), .A (filterType)) ;
    inv02 ix5321 (.Y (nx5322), .A (filterType)) ;
    buf02 ix5327 (.Y (nx5328), .A (regFileMap_filterEnables_0)) ;
    buf02 ix5329 (.Y (nx5330), .A (regFileMap_filterEnables_0)) ;
    buf02 ix5331 (.Y (nx5332), .A (regFileMap_filterEnables_1)) ;
    buf02 ix5333 (.Y (nx5334), .A (regFileMap_filterEnables_1)) ;
    buf02 ix5335 (.Y (nx5336), .A (regFileMap_filterEnables_2)) ;
    buf02 ix5337 (.Y (nx5338), .A (regFileMap_filterEnables_2)) ;
    buf02 ix5339 (.Y (nx5340), .A (regFileMap_filterEnables_3)) ;
    buf02 ix5341 (.Y (nx5342), .A (regFileMap_filterEnables_3)) ;
    inv02 ix5343 (.Y (nx5344), .A (nx2917)) ;
    inv02 ix5345 (.Y (nx5346), .A (nx2917)) ;
endmodule


module NBitAdder_16 ( a, b, carryIn, sum, carryOut ) ;

    input [15:0]a ;
    input [15:0]b ;
    input carryIn ;
    output [15:0]sum ;
    output carryOut ;

    wire nx2, nx8, nx10, nx18, nx24, nx26, nx34, nx40, nx42, nx50, nx56, nx58, 
         nx66, nx72, nx74, nx82, nx88, nx90, nx98, nx104, nx106, nx114, nx85, 
         nx89, nx93, nx99, nx101, nx103, nx107, nx111, nx115, nx121, nx123, 
         nx125, nx129, nx133, nx137, nx143, nx145, nx147, nx151, nx154, nx157, 
         nx161, nx163, nx165, nx168, nx171, nx174, nx178, nx180, nx182, nx185, 
         nx188, nx191, nx195, nx197, nx199, nx202, nx205, nx208, nx212, nx214, 
         nx216, nx219, nx222, nx225;



    fake_gnd ix42 (.Y (carryOut)) ;
    xnor2 ix151 (.Y (sum[0]), .A0 (b[0]), .A1 (nx85)) ;
    inv01 ix86 (.Y (nx85), .A (a[0])) ;
    xnor2 ix145 (.Y (sum[1]), .A0 (nx89), .A1 (nx2)) ;
    nand02 ix90 (.Y (nx89), .A0 (b[0]), .A1 (a[0])) ;
    xnor2 ix3 (.Y (nx2), .A0 (a[1]), .A1 (nx93)) ;
    inv01 ix94 (.Y (nx93), .A (b[1])) ;
    xnor2 ix143 (.Y (sum[2]), .A0 (nx8), .A1 (nx103)) ;
    oai22 ix9 (.Y (nx8), .A0 (nx89), .A1 (nx99), .B0 (nx93), .B1 (nx101)) ;
    xnor2 ix100 (.Y (nx99), .A0 (a[1]), .A1 (b[1])) ;
    inv01 ix102 (.Y (nx101), .A (a[1])) ;
    xnor2 ix104 (.Y (nx103), .A0 (a[2]), .A1 (b[2])) ;
    xnor2 ix141 (.Y (sum[3]), .A0 (nx107), .A1 (nx18)) ;
    aoi22 ix108 (.Y (nx107), .A0 (b[2]), .A1 (a[2]), .B0 (nx8), .B1 (nx10)) ;
    xnor2 ix11 (.Y (nx10), .A0 (a[2]), .A1 (nx111)) ;
    inv01 ix112 (.Y (nx111), .A (b[2])) ;
    xnor2 ix19 (.Y (nx18), .A0 (a[3]), .A1 (nx115)) ;
    inv01 ix116 (.Y (nx115), .A (b[3])) ;
    xnor2 ix139 (.Y (sum[4]), .A0 (nx24), .A1 (nx125)) ;
    oai21 ix25 (.Y (nx24), .A0 (nx107), .A1 (nx121), .B0 (nx123)) ;
    xnor2 ix122 (.Y (nx121), .A0 (a[3]), .A1 (b[3])) ;
    nand02 ix124 (.Y (nx123), .A0 (b[3]), .A1 (a[3])) ;
    xnor2 ix126 (.Y (nx125), .A0 (a[4]), .A1 (b[4])) ;
    xnor2 ix137 (.Y (sum[5]), .A0 (nx129), .A1 (nx34)) ;
    aoi22 ix130 (.Y (nx129), .A0 (b[4]), .A1 (a[4]), .B0 (nx24), .B1 (nx26)) ;
    xnor2 ix27 (.Y (nx26), .A0 (a[4]), .A1 (nx133)) ;
    inv01 ix134 (.Y (nx133), .A (b[4])) ;
    xnor2 ix35 (.Y (nx34), .A0 (a[5]), .A1 (nx137)) ;
    inv01 ix138 (.Y (nx137), .A (b[5])) ;
    xnor2 ix135 (.Y (sum[6]), .A0 (nx40), .A1 (nx147)) ;
    oai21 ix41 (.Y (nx40), .A0 (nx129), .A1 (nx143), .B0 (nx145)) ;
    xnor2 ix144 (.Y (nx143), .A0 (a[5]), .A1 (b[5])) ;
    nand02 ix146 (.Y (nx145), .A0 (b[5]), .A1 (a[5])) ;
    xnor2 ix148 (.Y (nx147), .A0 (a[6]), .A1 (b[6])) ;
    xnor2 ix133 (.Y (sum[7]), .A0 (nx151), .A1 (nx50)) ;
    aoi22 ix152 (.Y (nx151), .A0 (b[6]), .A1 (a[6]), .B0 (nx40), .B1 (nx42)) ;
    xnor2 ix43 (.Y (nx42), .A0 (a[6]), .A1 (nx154)) ;
    inv01 ix155 (.Y (nx154), .A (b[6])) ;
    xnor2 ix51 (.Y (nx50), .A0 (a[7]), .A1 (nx157)) ;
    inv01 ix158 (.Y (nx157), .A (b[7])) ;
    xnor2 ix131 (.Y (sum[8]), .A0 (nx56), .A1 (nx165)) ;
    oai21 ix57 (.Y (nx56), .A0 (nx151), .A1 (nx161), .B0 (nx163)) ;
    xnor2 ix162 (.Y (nx161), .A0 (a[7]), .A1 (b[7])) ;
    nand02 ix164 (.Y (nx163), .A0 (b[7]), .A1 (a[7])) ;
    xnor2 ix166 (.Y (nx165), .A0 (a[8]), .A1 (b[8])) ;
    xnor2 ix129 (.Y (sum[9]), .A0 (nx168), .A1 (nx66)) ;
    aoi22 ix169 (.Y (nx168), .A0 (b[8]), .A1 (a[8]), .B0 (nx56), .B1 (nx58)) ;
    xnor2 ix59 (.Y (nx58), .A0 (a[8]), .A1 (nx171)) ;
    inv01 ix172 (.Y (nx171), .A (b[8])) ;
    xnor2 ix67 (.Y (nx66), .A0 (a[9]), .A1 (nx174)) ;
    inv01 ix175 (.Y (nx174), .A (b[9])) ;
    xnor2 ix127 (.Y (sum[10]), .A0 (nx72), .A1 (nx182)) ;
    oai21 ix73 (.Y (nx72), .A0 (nx168), .A1 (nx178), .B0 (nx180)) ;
    xnor2 ix179 (.Y (nx178), .A0 (a[9]), .A1 (b[9])) ;
    nand02 ix181 (.Y (nx180), .A0 (b[9]), .A1 (a[9])) ;
    xnor2 ix183 (.Y (nx182), .A0 (a[10]), .A1 (b[10])) ;
    xnor2 ix125 (.Y (sum[11]), .A0 (nx185), .A1 (nx82)) ;
    aoi22 ix186 (.Y (nx185), .A0 (b[10]), .A1 (a[10]), .B0 (nx72), .B1 (nx74)) ;
    xnor2 ix75 (.Y (nx74), .A0 (a[10]), .A1 (nx188)) ;
    inv01 ix189 (.Y (nx188), .A (b[10])) ;
    xnor2 ix83 (.Y (nx82), .A0 (a[11]), .A1 (nx191)) ;
    inv01 ix192 (.Y (nx191), .A (b[11])) ;
    xnor2 ix123 (.Y (sum[12]), .A0 (nx88), .A1 (nx199)) ;
    oai21 ix89 (.Y (nx88), .A0 (nx185), .A1 (nx195), .B0 (nx197)) ;
    xnor2 ix196 (.Y (nx195), .A0 (a[11]), .A1 (b[11])) ;
    nand02 ix198 (.Y (nx197), .A0 (b[11]), .A1 (a[11])) ;
    xnor2 ix200 (.Y (nx199), .A0 (a[12]), .A1 (b[12])) ;
    xnor2 ix121 (.Y (sum[13]), .A0 (nx202), .A1 (nx98)) ;
    aoi22 ix203 (.Y (nx202), .A0 (b[12]), .A1 (a[12]), .B0 (nx88), .B1 (nx90)) ;
    xnor2 ix91 (.Y (nx90), .A0 (a[12]), .A1 (nx205)) ;
    inv01 ix206 (.Y (nx205), .A (b[12])) ;
    xnor2 ix99 (.Y (nx98), .A0 (a[13]), .A1 (nx208)) ;
    inv01 ix209 (.Y (nx208), .A (b[13])) ;
    xnor2 ix119 (.Y (sum[14]), .A0 (nx104), .A1 (nx216)) ;
    oai21 ix105 (.Y (nx104), .A0 (nx202), .A1 (nx212), .B0 (nx214)) ;
    xnor2 ix213 (.Y (nx212), .A0 (a[13]), .A1 (b[13])) ;
    nand02 ix215 (.Y (nx214), .A0 (b[13]), .A1 (a[13])) ;
    xnor2 ix217 (.Y (nx216), .A0 (a[14]), .A1 (b[14])) ;
    xnor2 ix117 (.Y (sum[15]), .A0 (nx219), .A1 (nx114)) ;
    aoi22 ix220 (.Y (nx219), .A0 (b[14]), .A1 (a[14]), .B0 (nx104), .B1 (nx106)
          ) ;
    xnor2 ix107 (.Y (nx106), .A0 (a[14]), .A1 (nx222)) ;
    inv01 ix223 (.Y (nx222), .A (b[14])) ;
    xnor2 ix115 (.Y (nx114), .A0 (a[15]), .A1 (nx225)) ;
    inv01 ix226 (.Y (nx225), .A (b[15])) ;
endmodule


module RegUnit_8_16_unfolded1 ( filterBus, windowBus, regPage1NextUnit, 
                                regPage2NextUnit, clk, rst, enableRegPage1, 
                                enableRegPage2, enableRegFilter, 
                                page1ReadBusOrPage2, page2ReadBusOrPage1, 
                                pageTurn, outRegPage, outputRegPage1, 
                                outputRegPage2, outFilter ) ;

    input [7:0]filterBus ;
    input [15:0]windowBus ;
    input [15:0]regPage1NextUnit ;
    input [15:0]regPage2NextUnit ;
    input clk ;
    input rst ;
    input enableRegPage1 ;
    input enableRegPage2 ;
    input enableRegFilter ;
    input page1ReadBusOrPage2 ;
    input page2ReadBusOrPage1 ;
    input pageTurn ;
    output [15:0]outRegPage ;
    output [15:0]outputRegPage1 ;
    output [15:0]outputRegPage2 ;
    output [7:0]outFilter ;

    wire nx133, nx143, nx153, nx163, nx173, nx183, nx193, nx203, nx213, nx223, 
         nx233, nx243, nx253, nx263, nx273, nx283, nx293, nx303, nx313, nx323, 
         nx333, nx343, nx353, nx363, nx373, nx383, nx393, nx403, nx413, nx423, 
         nx433, nx443, nx453, nx463, nx473, nx483, nx493, nx503, nx513, nx523, 
         nx535, nx539, nx544, nx546, nx551, nx553, nx558, nx560, nx565, nx567, 
         nx572, nx574, nx579, nx581, nx586, nx588, nx593, nx595, nx597, nx599, 
         nx601, nx604, nx606, nx608, nx611, nx613, nx615, nx618, nx620, nx622, 
         nx625, nx627, nx629, nx632, nx634, nx636, nx639, nx641, nx643, nx646, 
         nx648, nx650, nx653, nx655, nx657, nx660, nx662, nx664, nx667, nx669, 
         nx671, nx674, nx676, nx678, nx681, nx683, nx685, nx688, nx690, nx692, 
         nx695, nx697, nx699, nx702, nx704, nx706, nx709, nx711, nx713, nx715, 
         nx717, nx720, nx722, nx724, nx727, nx729, nx731, nx734, nx736, nx738, 
         nx741, nx743, nx745, nx748, nx750, nx752, nx755, nx757, nx759, nx762, 
         nx764, nx766, nx769, nx771, nx773, nx776, nx778, nx780, nx783, nx785, 
         nx787, nx790, nx792, nx794, nx797, nx799, nx801, nx804, nx806, nx808, 
         nx811, nx813, nx815, nx818, nx820, nx822, nx846, nx848, nx850, nx852, 
         nx854, nx856, nx858, nx860, nx862, nx868, nx870, nx872, nx874, nx876, 
         nx878, nx880, nx882, nx884, nx886, nx888, nx890;
    wire [7:0] \$dummy ;




    dffr regFilterMap_reg_Q_0 (.Q (outFilter[0]), .QB (\$dummy [0]), .D (nx453)
         , .CLK (clk), .R (rst)) ;
    nand02 ix454 (.Y (nx453), .A0 (nx535), .A1 (nx539)) ;
    nand02 ix536 (.Y (nx535), .A0 (outFilter[0]), .A1 (nx888)) ;
    nand02 ix540 (.Y (nx539), .A0 (filterBus[0]), .A1 (nx884)) ;
    dffr regFilterMap_reg_Q_1 (.Q (outFilter[1]), .QB (\$dummy [1]), .D (nx463)
         , .CLK (clk), .R (rst)) ;
    nand02 ix464 (.Y (nx463), .A0 (nx544), .A1 (nx546)) ;
    nand02 ix545 (.Y (nx544), .A0 (outFilter[1]), .A1 (nx888)) ;
    nand02 ix547 (.Y (nx546), .A0 (filterBus[1]), .A1 (nx884)) ;
    dffr regFilterMap_reg_Q_2 (.Q (outFilter[2]), .QB (\$dummy [2]), .D (nx473)
         , .CLK (clk), .R (rst)) ;
    nand02 ix474 (.Y (nx473), .A0 (nx551), .A1 (nx553)) ;
    nand02 ix552 (.Y (nx551), .A0 (outFilter[2]), .A1 (nx888)) ;
    nand02 ix554 (.Y (nx553), .A0 (filterBus[2]), .A1 (nx884)) ;
    dffr regFilterMap_reg_Q_3 (.Q (outFilter[3]), .QB (\$dummy [3]), .D (nx483)
         , .CLK (clk), .R (rst)) ;
    nand02 ix484 (.Y (nx483), .A0 (nx558), .A1 (nx560)) ;
    nand02 ix559 (.Y (nx558), .A0 (outFilter[3]), .A1 (nx888)) ;
    nand02 ix561 (.Y (nx560), .A0 (filterBus[3]), .A1 (nx884)) ;
    dffr regFilterMap_reg_Q_4 (.Q (outFilter[4]), .QB (\$dummy [4]), .D (nx493)
         , .CLK (clk), .R (rst)) ;
    nand02 ix494 (.Y (nx493), .A0 (nx565), .A1 (nx567)) ;
    nand02 ix566 (.Y (nx565), .A0 (outFilter[4]), .A1 (nx888)) ;
    nand02 ix568 (.Y (nx567), .A0 (filterBus[4]), .A1 (nx884)) ;
    dffr regFilterMap_reg_Q_5 (.Q (outFilter[5]), .QB (\$dummy [5]), .D (nx503)
         , .CLK (clk), .R (rst)) ;
    nand02 ix504 (.Y (nx503), .A0 (nx572), .A1 (nx574)) ;
    nand02 ix573 (.Y (nx572), .A0 (outFilter[5]), .A1 (nx888)) ;
    nand02 ix575 (.Y (nx574), .A0 (filterBus[5]), .A1 (nx884)) ;
    dffr regFilterMap_reg_Q_6 (.Q (outFilter[6]), .QB (\$dummy [6]), .D (nx513)
         , .CLK (clk), .R (rst)) ;
    nand02 ix514 (.Y (nx513), .A0 (nx579), .A1 (nx581)) ;
    nand02 ix580 (.Y (nx579), .A0 (outFilter[6]), .A1 (nx888)) ;
    nand02 ix582 (.Y (nx581), .A0 (filterBus[6]), .A1 (nx884)) ;
    dffr regFilterMap_reg_Q_7 (.Q (outFilter[7]), .QB (\$dummy [7]), .D (nx523)
         , .CLK (clk), .R (rst)) ;
    nand02 ix524 (.Y (nx523), .A0 (nx586), .A1 (nx588)) ;
    nand02 ix587 (.Y (nx586), .A0 (outFilter[7]), .A1 (nx846)) ;
    nand02 ix589 (.Y (nx588), .A0 (filterBus[7]), .A1 (nx886)) ;
    dffr regPage2Map_reg_Q_0 (.Q (outputRegPage2[0]), .QB (nx601), .D (nx143), .CLK (
         clk), .R (rst)) ;
    nand02 ix144 (.Y (nx143), .A0 (nx593), .A1 (nx597)) ;
    nand02 ix594 (.Y (nx593), .A0 (outputRegPage2[0]), .A1 (nx848)) ;
    nor02_2x ix596 (.Y (nx595), .A0 (nx878), .A1 (page2ReadBusOrPage1)) ;
    nand03 ix598 (.Y (nx597), .A0 (windowBus[0]), .A1 (nx852), .A2 (nx878)) ;
    inv01 ix600 (.Y (nx599), .A (page2ReadBusOrPage1)) ;
    dffr regPage2Map_reg_Q_1 (.Q (outputRegPage2[1]), .QB (nx608), .D (nx163), .CLK (
         clk), .R (rst)) ;
    nand02 ix164 (.Y (nx163), .A0 (nx604), .A1 (nx606)) ;
    nand02 ix605 (.Y (nx604), .A0 (outputRegPage2[1]), .A1 (nx848)) ;
    nand03 ix607 (.Y (nx606), .A0 (windowBus[1]), .A1 (nx852), .A2 (nx878)) ;
    dffr regPage2Map_reg_Q_2 (.Q (outputRegPage2[2]), .QB (nx615), .D (nx183), .CLK (
         clk), .R (rst)) ;
    nand02 ix184 (.Y (nx183), .A0 (nx611), .A1 (nx613)) ;
    nand02 ix612 (.Y (nx611), .A0 (outputRegPage2[2]), .A1 (nx848)) ;
    nand03 ix614 (.Y (nx613), .A0 (windowBus[2]), .A1 (nx852), .A2 (nx878)) ;
    dffr regPage2Map_reg_Q_3 (.Q (outputRegPage2[3]), .QB (nx622), .D (nx203), .CLK (
         clk), .R (rst)) ;
    nand02 ix204 (.Y (nx203), .A0 (nx618), .A1 (nx620)) ;
    nand02 ix619 (.Y (nx618), .A0 (outputRegPage2[3]), .A1 (nx848)) ;
    nand03 ix621 (.Y (nx620), .A0 (windowBus[3]), .A1 (nx852), .A2 (nx878)) ;
    dffr regPage2Map_reg_Q_4 (.Q (outputRegPage2[4]), .QB (nx629), .D (nx223), .CLK (
         clk), .R (rst)) ;
    nand02 ix224 (.Y (nx223), .A0 (nx625), .A1 (nx627)) ;
    nand02 ix626 (.Y (nx625), .A0 (outputRegPage2[4]), .A1 (nx848)) ;
    nand03 ix628 (.Y (nx627), .A0 (windowBus[4]), .A1 (nx852), .A2 (nx878)) ;
    dffr regPage2Map_reg_Q_5 (.Q (outputRegPage2[5]), .QB (nx636), .D (nx243), .CLK (
         clk), .R (rst)) ;
    nand02 ix244 (.Y (nx243), .A0 (nx632), .A1 (nx634)) ;
    nand02 ix633 (.Y (nx632), .A0 (outputRegPage2[5]), .A1 (nx848)) ;
    nand03 ix635 (.Y (nx634), .A0 (windowBus[5]), .A1 (nx852), .A2 (nx878)) ;
    dffr regPage2Map_reg_Q_6 (.Q (outputRegPage2[6]), .QB (nx643), .D (nx263), .CLK (
         clk), .R (rst)) ;
    nand02 ix264 (.Y (nx263), .A0 (nx639), .A1 (nx641)) ;
    nand02 ix640 (.Y (nx639), .A0 (outputRegPage2[6]), .A1 (nx848)) ;
    nand03 ix642 (.Y (nx641), .A0 (windowBus[6]), .A1 (nx854), .A2 (nx880)) ;
    dffr regPage2Map_reg_Q_7 (.Q (outputRegPage2[7]), .QB (nx650), .D (nx283), .CLK (
         clk), .R (rst)) ;
    nand02 ix284 (.Y (nx283), .A0 (nx646), .A1 (nx648)) ;
    nand02 ix647 (.Y (nx646), .A0 (outputRegPage2[7]), .A1 (nx850)) ;
    nand03 ix649 (.Y (nx648), .A0 (windowBus[7]), .A1 (nx854), .A2 (nx880)) ;
    dffr regPage2Map_reg_Q_8 (.Q (outputRegPage2[8]), .QB (nx657), .D (nx303), .CLK (
         clk), .R (rst)) ;
    nand02 ix304 (.Y (nx303), .A0 (nx653), .A1 (nx655)) ;
    nand02 ix654 (.Y (nx653), .A0 (outputRegPage2[8]), .A1 (nx850)) ;
    nand03 ix656 (.Y (nx655), .A0 (windowBus[8]), .A1 (nx854), .A2 (nx880)) ;
    dffr regPage2Map_reg_Q_9 (.Q (outputRegPage2[9]), .QB (nx664), .D (nx323), .CLK (
         clk), .R (rst)) ;
    nand02 ix324 (.Y (nx323), .A0 (nx660), .A1 (nx662)) ;
    nand02 ix661 (.Y (nx660), .A0 (outputRegPage2[9]), .A1 (nx850)) ;
    nand03 ix663 (.Y (nx662), .A0 (windowBus[9]), .A1 (nx854), .A2 (nx880)) ;
    dffr regPage2Map_reg_Q_10 (.Q (outputRegPage2[10]), .QB (nx671), .D (nx343)
         , .CLK (clk), .R (rst)) ;
    nand02 ix344 (.Y (nx343), .A0 (nx667), .A1 (nx669)) ;
    nand02 ix668 (.Y (nx667), .A0 (outputRegPage2[10]), .A1 (nx850)) ;
    nand03 ix670 (.Y (nx669), .A0 (windowBus[10]), .A1 (nx854), .A2 (nx880)) ;
    dffr regPage2Map_reg_Q_11 (.Q (outputRegPage2[11]), .QB (nx678), .D (nx363)
         , .CLK (clk), .R (rst)) ;
    nand02 ix364 (.Y (nx363), .A0 (nx674), .A1 (nx676)) ;
    nand02 ix675 (.Y (nx674), .A0 (outputRegPage2[11]), .A1 (nx850)) ;
    nand03 ix677 (.Y (nx676), .A0 (windowBus[11]), .A1 (nx854), .A2 (nx880)) ;
    dffr regPage2Map_reg_Q_12 (.Q (outputRegPage2[12]), .QB (nx685), .D (nx383)
         , .CLK (clk), .R (rst)) ;
    nand02 ix384 (.Y (nx383), .A0 (nx681), .A1 (nx683)) ;
    nand02 ix682 (.Y (nx681), .A0 (outputRegPage2[12]), .A1 (nx850)) ;
    nand03 ix684 (.Y (nx683), .A0 (windowBus[12]), .A1 (nx599), .A2 (nx880)) ;
    dffr regPage2Map_reg_Q_13 (.Q (outputRegPage2[13]), .QB (nx692), .D (nx403)
         , .CLK (clk), .R (rst)) ;
    nand02 ix404 (.Y (nx403), .A0 (nx688), .A1 (nx690)) ;
    nand02 ix689 (.Y (nx688), .A0 (outputRegPage2[13]), .A1 (nx850)) ;
    nand03 ix691 (.Y (nx690), .A0 (windowBus[13]), .A1 (nx599), .A2 (nx882)) ;
    dffr regPage2Map_reg_Q_14 (.Q (outputRegPage2[14]), .QB (nx699), .D (nx423)
         , .CLK (clk), .R (rst)) ;
    nand02 ix424 (.Y (nx423), .A0 (nx695), .A1 (nx697)) ;
    nand02 ix696 (.Y (nx695), .A0 (outputRegPage2[14]), .A1 (nx595)) ;
    nand03 ix698 (.Y (nx697), .A0 (windowBus[14]), .A1 (nx599), .A2 (nx882)) ;
    dffr regPage2Map_reg_Q_15 (.Q (outputRegPage2[15]), .QB (nx706), .D (nx443)
         , .CLK (clk), .R (rst)) ;
    nand02 ix444 (.Y (nx443), .A0 (nx702), .A1 (nx704)) ;
    nand02 ix703 (.Y (nx702), .A0 (outputRegPage2[15]), .A1 (nx595)) ;
    nand03 ix705 (.Y (nx704), .A0 (windowBus[15]), .A1 (nx599), .A2 (nx882)) ;
    dffr regPage1Map_reg_Q_0 (.Q (outputRegPage1[0]), .QB (nx717), .D (nx133), .CLK (
         clk), .R (rst)) ;
    nand02 ix134 (.Y (nx133), .A0 (nx709), .A1 (nx713)) ;
    nand02 ix710 (.Y (nx709), .A0 (outputRegPage1[0]), .A1 (nx856)) ;
    nor02_2x ix712 (.Y (nx711), .A0 (nx870), .A1 (page1ReadBusOrPage2)) ;
    nand03 ix714 (.Y (nx713), .A0 (windowBus[0]), .A1 (nx860), .A2 (nx870)) ;
    inv01 ix716 (.Y (nx715), .A (page1ReadBusOrPage2)) ;
    dffr regPage1Map_reg_Q_1 (.Q (outputRegPage1[1]), .QB (nx724), .D (nx153), .CLK (
         clk), .R (rst)) ;
    nand02 ix154 (.Y (nx153), .A0 (nx720), .A1 (nx722)) ;
    nand02 ix721 (.Y (nx720), .A0 (outputRegPage1[1]), .A1 (nx856)) ;
    nand03 ix723 (.Y (nx722), .A0 (windowBus[1]), .A1 (nx860), .A2 (nx870)) ;
    dffr regPage1Map_reg_Q_2 (.Q (outputRegPage1[2]), .QB (nx731), .D (nx173), .CLK (
         clk), .R (rst)) ;
    nand02 ix174 (.Y (nx173), .A0 (nx727), .A1 (nx729)) ;
    nand02 ix728 (.Y (nx727), .A0 (outputRegPage1[2]), .A1 (nx856)) ;
    nand03 ix730 (.Y (nx729), .A0 (windowBus[2]), .A1 (nx860), .A2 (nx870)) ;
    dffr regPage1Map_reg_Q_3 (.Q (outputRegPage1[3]), .QB (nx738), .D (nx193), .CLK (
         clk), .R (rst)) ;
    nand02 ix194 (.Y (nx193), .A0 (nx734), .A1 (nx736)) ;
    nand02 ix735 (.Y (nx734), .A0 (outputRegPage1[3]), .A1 (nx856)) ;
    nand03 ix737 (.Y (nx736), .A0 (windowBus[3]), .A1 (nx860), .A2 (nx870)) ;
    dffr regPage1Map_reg_Q_4 (.Q (outputRegPage1[4]), .QB (nx745), .D (nx213), .CLK (
         clk), .R (rst)) ;
    nand02 ix214 (.Y (nx213), .A0 (nx741), .A1 (nx743)) ;
    nand02 ix742 (.Y (nx741), .A0 (outputRegPage1[4]), .A1 (nx856)) ;
    nand03 ix744 (.Y (nx743), .A0 (windowBus[4]), .A1 (nx860), .A2 (nx870)) ;
    dffr regPage1Map_reg_Q_5 (.Q (outputRegPage1[5]), .QB (nx752), .D (nx233), .CLK (
         clk), .R (rst)) ;
    nand02 ix234 (.Y (nx233), .A0 (nx748), .A1 (nx750)) ;
    nand02 ix749 (.Y (nx748), .A0 (outputRegPage1[5]), .A1 (nx856)) ;
    nand03 ix751 (.Y (nx750), .A0 (windowBus[5]), .A1 (nx860), .A2 (nx870)) ;
    dffr regPage1Map_reg_Q_6 (.Q (outputRegPage1[6]), .QB (nx759), .D (nx253), .CLK (
         clk), .R (rst)) ;
    nand02 ix254 (.Y (nx253), .A0 (nx755), .A1 (nx757)) ;
    nand02 ix756 (.Y (nx755), .A0 (outputRegPage1[6]), .A1 (nx856)) ;
    nand03 ix758 (.Y (nx757), .A0 (windowBus[6]), .A1 (nx862), .A2 (nx872)) ;
    dffr regPage1Map_reg_Q_7 (.Q (outputRegPage1[7]), .QB (nx766), .D (nx273), .CLK (
         clk), .R (rst)) ;
    nand02 ix274 (.Y (nx273), .A0 (nx762), .A1 (nx764)) ;
    nand02 ix763 (.Y (nx762), .A0 (outputRegPage1[7]), .A1 (nx858)) ;
    nand03 ix765 (.Y (nx764), .A0 (windowBus[7]), .A1 (nx862), .A2 (nx872)) ;
    dffr regPage1Map_reg_Q_8 (.Q (outputRegPage1[8]), .QB (nx773), .D (nx293), .CLK (
         clk), .R (rst)) ;
    nand02 ix294 (.Y (nx293), .A0 (nx769), .A1 (nx771)) ;
    nand02 ix770 (.Y (nx769), .A0 (outputRegPage1[8]), .A1 (nx858)) ;
    nand03 ix772 (.Y (nx771), .A0 (windowBus[8]), .A1 (nx862), .A2 (nx872)) ;
    dffr regPage1Map_reg_Q_9 (.Q (outputRegPage1[9]), .QB (nx780), .D (nx313), .CLK (
         clk), .R (rst)) ;
    nand02 ix314 (.Y (nx313), .A0 (nx776), .A1 (nx778)) ;
    nand02 ix777 (.Y (nx776), .A0 (outputRegPage1[9]), .A1 (nx858)) ;
    nand03 ix779 (.Y (nx778), .A0 (windowBus[9]), .A1 (nx862), .A2 (nx872)) ;
    dffr regPage1Map_reg_Q_10 (.Q (outputRegPage1[10]), .QB (nx787), .D (nx333)
         , .CLK (clk), .R (rst)) ;
    nand02 ix334 (.Y (nx333), .A0 (nx783), .A1 (nx785)) ;
    nand02 ix784 (.Y (nx783), .A0 (outputRegPage1[10]), .A1 (nx858)) ;
    nand03 ix786 (.Y (nx785), .A0 (windowBus[10]), .A1 (nx862), .A2 (nx872)) ;
    dffr regPage1Map_reg_Q_11 (.Q (outputRegPage1[11]), .QB (nx794), .D (nx353)
         , .CLK (clk), .R (rst)) ;
    nand02 ix354 (.Y (nx353), .A0 (nx790), .A1 (nx792)) ;
    nand02 ix791 (.Y (nx790), .A0 (outputRegPage1[11]), .A1 (nx858)) ;
    nand03 ix793 (.Y (nx792), .A0 (windowBus[11]), .A1 (nx862), .A2 (nx872)) ;
    dffr regPage1Map_reg_Q_12 (.Q (outputRegPage1[12]), .QB (nx801), .D (nx373)
         , .CLK (clk), .R (rst)) ;
    nand02 ix374 (.Y (nx373), .A0 (nx797), .A1 (nx799)) ;
    nand02 ix798 (.Y (nx797), .A0 (outputRegPage1[12]), .A1 (nx858)) ;
    nand03 ix800 (.Y (nx799), .A0 (windowBus[12]), .A1 (nx715), .A2 (nx872)) ;
    dffr regPage1Map_reg_Q_13 (.Q (outputRegPage1[13]), .QB (nx808), .D (nx393)
         , .CLK (clk), .R (rst)) ;
    nand02 ix394 (.Y (nx393), .A0 (nx804), .A1 (nx806)) ;
    nand02 ix805 (.Y (nx804), .A0 (outputRegPage1[13]), .A1 (nx858)) ;
    nand03 ix807 (.Y (nx806), .A0 (windowBus[13]), .A1 (nx715), .A2 (nx874)) ;
    dffr regPage1Map_reg_Q_14 (.Q (outputRegPage1[14]), .QB (nx815), .D (nx413)
         , .CLK (clk), .R (rst)) ;
    nand02 ix414 (.Y (nx413), .A0 (nx811), .A1 (nx813)) ;
    nand02 ix812 (.Y (nx811), .A0 (outputRegPage1[14]), .A1 (nx711)) ;
    nand03 ix814 (.Y (nx813), .A0 (windowBus[14]), .A1 (nx715), .A2 (nx874)) ;
    dffr regPage1Map_reg_Q_15 (.Q (outputRegPage1[15]), .QB (nx822), .D (nx433)
         , .CLK (clk), .R (rst)) ;
    nand02 ix434 (.Y (nx433), .A0 (nx818), .A1 (nx820)) ;
    nand02 ix819 (.Y (nx818), .A0 (outputRegPage1[15]), .A1 (nx711)) ;
    nand03 ix821 (.Y (nx820), .A0 (windowBus[15]), .A1 (nx715), .A2 (nx874)) ;
    mux21 ix25 (.Y (outRegPage[0]), .A0 (nx717), .A1 (nx601), .S0 (pageTurn)) ;
    mux21 ix45 (.Y (outRegPage[1]), .A0 (nx724), .A1 (nx608), .S0 (pageTurn)) ;
    mux21 ix65 (.Y (outRegPage[2]), .A0 (nx731), .A1 (nx615), .S0 (pageTurn)) ;
    mux21 ix85 (.Y (outRegPage[3]), .A0 (nx738), .A1 (nx622), .S0 (pageTurn)) ;
    mux21 ix105 (.Y (outRegPage[4]), .A0 (nx745), .A1 (nx629), .S0 (pageTurn)) ;
    mux21 ix125 (.Y (outRegPage[5]), .A0 (nx752), .A1 (nx636), .S0 (pageTurn)) ;
    mux21 ix145 (.Y (outRegPage[6]), .A0 (nx759), .A1 (nx643), .S0 (pageTurn)) ;
    mux21 ix165 (.Y (outRegPage[7]), .A0 (nx766), .A1 (nx650), .S0 (pageTurn)) ;
    mux21 ix185 (.Y (outRegPage[8]), .A0 (nx773), .A1 (nx657), .S0 (pageTurn)) ;
    mux21 ix205 (.Y (outRegPage[9]), .A0 (nx780), .A1 (nx664), .S0 (pageTurn)) ;
    mux21 ix225 (.Y (outRegPage[10]), .A0 (nx787), .A1 (nx671), .S0 (pageTurn)
          ) ;
    mux21 ix245 (.Y (outRegPage[11]), .A0 (nx794), .A1 (nx678), .S0 (pageTurn)
          ) ;
    mux21 ix265 (.Y (outRegPage[12]), .A0 (nx801), .A1 (nx685), .S0 (pageTurn)
          ) ;
    mux21 ix285 (.Y (outRegPage[13]), .A0 (nx808), .A1 (nx692), .S0 (pageTurn)
          ) ;
    mux21 ix305 (.Y (outRegPage[14]), .A0 (nx815), .A1 (nx699), .S0 (pageTurn)
          ) ;
    mux21 ix325 (.Y (outRegPage[15]), .A0 (nx822), .A1 (nx706), .S0 (pageTurn)
          ) ;
    inv01 ix845 (.Y (nx846), .A (nx886)) ;
    nor02_2x ix847 (.Y (nx848), .A0 (nx882), .A1 (page2ReadBusOrPage1)) ;
    nor02_2x ix849 (.Y (nx850), .A0 (nx882), .A1 (page2ReadBusOrPage1)) ;
    inv01 ix851 (.Y (nx852), .A (page2ReadBusOrPage1)) ;
    inv01 ix853 (.Y (nx854), .A (page2ReadBusOrPage1)) ;
    nor02_2x ix855 (.Y (nx856), .A0 (nx874), .A1 (page1ReadBusOrPage2)) ;
    nor02_2x ix857 (.Y (nx858), .A0 (nx874), .A1 (page1ReadBusOrPage2)) ;
    inv01 ix859 (.Y (nx860), .A (page1ReadBusOrPage2)) ;
    inv01 ix861 (.Y (nx862), .A (page1ReadBusOrPage2)) ;
    inv01 ix867 (.Y (nx868), .A (enableRegPage1)) ;
    inv02 ix869 (.Y (nx870), .A (nx868)) ;
    inv02 ix871 (.Y (nx872), .A (nx868)) ;
    inv02 ix873 (.Y (nx874), .A (nx868)) ;
    inv01 ix875 (.Y (nx876), .A (enableRegPage2)) ;
    inv02 ix877 (.Y (nx878), .A (nx876)) ;
    inv02 ix879 (.Y (nx880), .A (nx876)) ;
    inv02 ix881 (.Y (nx882), .A (nx876)) ;
    inv02 ix883 (.Y (nx884), .A (nx890)) ;
    inv02 ix885 (.Y (nx886), .A (nx890)) ;
    inv02 ix887 (.Y (nx888), .A (enableRegFilter)) ;
    inv02 ix889 (.Y (nx890), .A (enableRegFilter)) ;
endmodule


module RegUnit_8_16_unfolded0 ( filterBus, windowBus, regPage1NextUnit, 
                                regPage2NextUnit, clk, rst, enableRegPage1, 
                                enableRegPage2, enableRegFilter, 
                                page1ReadBusOrPage2, page2ReadBusOrPage1, 
                                pageTurn, outRegPage, outputRegPage1, 
                                outputRegPage2, outFilter ) ;

    input [7:0]filterBus ;
    input [15:0]windowBus ;
    input [15:0]regPage1NextUnit ;
    input [15:0]regPage2NextUnit ;
    input clk ;
    input rst ;
    input enableRegPage1 ;
    input enableRegPage2 ;
    input enableRegFilter ;
    input page1ReadBusOrPage2 ;
    input page2ReadBusOrPage1 ;
    input pageTurn ;
    output [15:0]outRegPage ;
    output [15:0]outputRegPage1 ;
    output [15:0]outputRegPage2 ;
    output [7:0]outFilter ;

    wire nx345, nx355, nx365, nx375, nx385, nx395, nx405, nx415, nx425, nx435, 
         nx445, nx455, nx465, nx475, nx485, nx495, nx505, nx515, nx525, nx535, 
         nx545, nx555, nx565, nx575, nx585, nx595, nx605, nx615, nx625, nx635, 
         nx645, nx655, nx665, nx675, nx685, nx695, nx705, nx715, nx725, nx735, 
         nx747, nx751, nx756, nx758, nx763, nx765, nx770, nx772, nx777, nx779, 
         nx784, nx786, nx791, nx793, nx798, nx800, nx805, nx807, nx809, nx811, 
         nx814, nx816, nx818, nx821, nx823, nx825, nx828, nx830, nx832, nx835, 
         nx837, nx839, nx842, nx844, nx846, nx849, nx851, nx853, nx856, nx858, 
         nx860, nx863, nx865, nx867, nx870, nx872, nx874, nx877, nx879, nx881, 
         nx884, nx886, nx888, nx891, nx893, nx895, nx898, nx900, nx902, nx905, 
         nx907, nx909, nx912, nx914, nx916, nx919, nx921, nx923, nx925, nx928, 
         nx930, nx932, nx935, nx937, nx939, nx942, nx944, nx946, nx949, nx951, 
         nx953, nx956, nx958, nx960, nx963, nx965, nx967, nx970, nx972, nx974, 
         nx977, nx979, nx981, nx984, nx986, nx988, nx991, nx993, nx995, nx998, 
         nx1000, nx1002, nx1005, nx1007, nx1009, nx1012, nx1014, nx1016, nx1019, 
         nx1021, nx1023, nx1026, nx1028, nx1030, nx1054, nx1056, nx1058, nx1060, 
         nx1062, nx1064, nx1066, nx1068, nx1070, nx1072, nx1074, nx1076, nx1078, 
         nx1084, nx1086, nx1088, nx1090;
    wire [7:0] \$dummy ;




    dffr regFilterMap_reg_Q_0 (.Q (outFilter[0]), .QB (\$dummy [0]), .D (nx665)
         , .CLK (clk), .R (rst)) ;
    nand02 ix666 (.Y (nx665), .A0 (nx747), .A1 (nx751)) ;
    nand02 ix748 (.Y (nx747), .A0 (outFilter[0]), .A1 (nx1088)) ;
    nand02 ix752 (.Y (nx751), .A0 (filterBus[0]), .A1 (nx1084)) ;
    dffr regFilterMap_reg_Q_1 (.Q (outFilter[1]), .QB (\$dummy [1]), .D (nx675)
         , .CLK (clk), .R (rst)) ;
    nand02 ix676 (.Y (nx675), .A0 (nx756), .A1 (nx758)) ;
    nand02 ix757 (.Y (nx756), .A0 (outFilter[1]), .A1 (nx1088)) ;
    nand02 ix759 (.Y (nx758), .A0 (filterBus[1]), .A1 (nx1084)) ;
    dffr regFilterMap_reg_Q_2 (.Q (outFilter[2]), .QB (\$dummy [2]), .D (nx685)
         , .CLK (clk), .R (rst)) ;
    nand02 ix686 (.Y (nx685), .A0 (nx763), .A1 (nx765)) ;
    nand02 ix764 (.Y (nx763), .A0 (outFilter[2]), .A1 (nx1088)) ;
    nand02 ix766 (.Y (nx765), .A0 (filterBus[2]), .A1 (nx1084)) ;
    dffr regFilterMap_reg_Q_3 (.Q (outFilter[3]), .QB (\$dummy [3]), .D (nx695)
         , .CLK (clk), .R (rst)) ;
    nand02 ix696 (.Y (nx695), .A0 (nx770), .A1 (nx772)) ;
    nand02 ix771 (.Y (nx770), .A0 (outFilter[3]), .A1 (nx1088)) ;
    nand02 ix773 (.Y (nx772), .A0 (filterBus[3]), .A1 (nx1084)) ;
    dffr regFilterMap_reg_Q_4 (.Q (outFilter[4]), .QB (\$dummy [4]), .D (nx705)
         , .CLK (clk), .R (rst)) ;
    nand02 ix706 (.Y (nx705), .A0 (nx777), .A1 (nx779)) ;
    nand02 ix778 (.Y (nx777), .A0 (outFilter[4]), .A1 (nx1088)) ;
    nand02 ix780 (.Y (nx779), .A0 (filterBus[4]), .A1 (nx1084)) ;
    dffr regFilterMap_reg_Q_5 (.Q (outFilter[5]), .QB (\$dummy [5]), .D (nx715)
         , .CLK (clk), .R (rst)) ;
    nand02 ix716 (.Y (nx715), .A0 (nx784), .A1 (nx786)) ;
    nand02 ix785 (.Y (nx784), .A0 (outFilter[5]), .A1 (nx1088)) ;
    nand02 ix787 (.Y (nx786), .A0 (filterBus[5]), .A1 (nx1084)) ;
    dffr regFilterMap_reg_Q_6 (.Q (outFilter[6]), .QB (\$dummy [6]), .D (nx725)
         , .CLK (clk), .R (rst)) ;
    nand02 ix726 (.Y (nx725), .A0 (nx791), .A1 (nx793)) ;
    nand02 ix792 (.Y (nx791), .A0 (outFilter[6]), .A1 (nx1088)) ;
    nand02 ix794 (.Y (nx793), .A0 (filterBus[6]), .A1 (nx1084)) ;
    dffr regFilterMap_reg_Q_7 (.Q (outFilter[7]), .QB (\$dummy [7]), .D (nx735)
         , .CLK (clk), .R (rst)) ;
    nand02 ix736 (.Y (nx735), .A0 (nx798), .A1 (nx800)) ;
    nand02 ix799 (.Y (nx798), .A0 (outFilter[7]), .A1 (nx1054)) ;
    nand02 ix801 (.Y (nx800), .A0 (filterBus[7]), .A1 (nx1086)) ;
    dffr regPage2Map_reg_Q_0 (.Q (outputRegPage2[0]), .QB (nx811), .D (nx355), .CLK (
         clk), .R (rst)) ;
    oai21 ix356 (.Y (nx355), .A0 (nx805), .A1 (nx1058), .B0 (nx809)) ;
    mux21 ix806 (.Y (nx805), .A0 (windowBus[0]), .A1 (regPage1NextUnit[0]), .S0 (
          page2ReadBusOrPage1)) ;
    nor02_2x ix808 (.Y (nx807), .A0 (enableRegPage2), .A1 (page2ReadBusOrPage1)
             ) ;
    nand02 ix810 (.Y (nx809), .A0 (outputRegPage2[0]), .A1 (nx1058)) ;
    dffr regPage2Map_reg_Q_1 (.Q (outputRegPage2[1]), .QB (nx818), .D (nx375), .CLK (
         clk), .R (rst)) ;
    oai21 ix376 (.Y (nx375), .A0 (nx814), .A1 (nx1058), .B0 (nx816)) ;
    mux21 ix815 (.Y (nx814), .A0 (windowBus[1]), .A1 (regPage1NextUnit[1]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix817 (.Y (nx816), .A0 (outputRegPage2[1]), .A1 (nx1058)) ;
    dffr regPage2Map_reg_Q_2 (.Q (outputRegPage2[2]), .QB (nx825), .D (nx395), .CLK (
         clk), .R (rst)) ;
    oai21 ix396 (.Y (nx395), .A0 (nx821), .A1 (nx1058), .B0 (nx823)) ;
    mux21 ix822 (.Y (nx821), .A0 (windowBus[2]), .A1 (regPage1NextUnit[2]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix824 (.Y (nx823), .A0 (outputRegPage2[2]), .A1 (nx1058)) ;
    dffr regPage2Map_reg_Q_3 (.Q (outputRegPage2[3]), .QB (nx832), .D (nx415), .CLK (
         clk), .R (rst)) ;
    oai21 ix416 (.Y (nx415), .A0 (nx828), .A1 (nx1058), .B0 (nx830)) ;
    mux21 ix829 (.Y (nx828), .A0 (windowBus[3]), .A1 (regPage1NextUnit[3]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix831 (.Y (nx830), .A0 (outputRegPage2[3]), .A1 (nx1060)) ;
    dffr regPage2Map_reg_Q_4 (.Q (outputRegPage2[4]), .QB (nx839), .D (nx435), .CLK (
         clk), .R (rst)) ;
    oai21 ix436 (.Y (nx435), .A0 (nx835), .A1 (nx1060), .B0 (nx837)) ;
    mux21 ix836 (.Y (nx835), .A0 (windowBus[4]), .A1 (regPage1NextUnit[4]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix838 (.Y (nx837), .A0 (outputRegPage2[4]), .A1 (nx1060)) ;
    dffr regPage2Map_reg_Q_5 (.Q (outputRegPage2[5]), .QB (nx846), .D (nx455), .CLK (
         clk), .R (rst)) ;
    oai21 ix456 (.Y (nx455), .A0 (nx842), .A1 (nx1060), .B0 (nx844)) ;
    mux21 ix843 (.Y (nx842), .A0 (windowBus[5]), .A1 (regPage1NextUnit[5]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix845 (.Y (nx844), .A0 (outputRegPage2[5]), .A1 (nx1060)) ;
    dffr regPage2Map_reg_Q_6 (.Q (outputRegPage2[6]), .QB (nx853), .D (nx475), .CLK (
         clk), .R (rst)) ;
    oai21 ix476 (.Y (nx475), .A0 (nx849), .A1 (nx1060), .B0 (nx851)) ;
    mux21 ix850 (.Y (nx849), .A0 (windowBus[6]), .A1 (regPage1NextUnit[6]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix852 (.Y (nx851), .A0 (outputRegPage2[6]), .A1 (nx1060)) ;
    dffr regPage2Map_reg_Q_7 (.Q (outputRegPage2[7]), .QB (nx860), .D (nx495), .CLK (
         clk), .R (rst)) ;
    oai21 ix496 (.Y (nx495), .A0 (nx856), .A1 (nx1062), .B0 (nx858)) ;
    mux21 ix857 (.Y (nx856), .A0 (windowBus[7]), .A1 (regPage1NextUnit[7]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix859 (.Y (nx858), .A0 (outputRegPage2[7]), .A1 (nx1062)) ;
    dffr regPage2Map_reg_Q_8 (.Q (outputRegPage2[8]), .QB (nx867), .D (nx515), .CLK (
         clk), .R (rst)) ;
    oai21 ix516 (.Y (nx515), .A0 (nx863), .A1 (nx1062), .B0 (nx865)) ;
    mux21 ix864 (.Y (nx863), .A0 (windowBus[8]), .A1 (regPage1NextUnit[8]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix866 (.Y (nx865), .A0 (outputRegPage2[8]), .A1 (nx1062)) ;
    dffr regPage2Map_reg_Q_9 (.Q (outputRegPage2[9]), .QB (nx874), .D (nx535), .CLK (
         clk), .R (rst)) ;
    oai21 ix536 (.Y (nx535), .A0 (nx870), .A1 (nx1062), .B0 (nx872)) ;
    mux21 ix871 (.Y (nx870), .A0 (windowBus[9]), .A1 (regPage1NextUnit[9]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix873 (.Y (nx872), .A0 (outputRegPage2[9]), .A1 (nx1062)) ;
    dffr regPage2Map_reg_Q_10 (.Q (outputRegPage2[10]), .QB (nx881), .D (nx555)
         , .CLK (clk), .R (rst)) ;
    oai21 ix556 (.Y (nx555), .A0 (nx877), .A1 (nx1062), .B0 (nx879)) ;
    mux21 ix878 (.Y (nx877), .A0 (windowBus[10]), .A1 (regPage1NextUnit[10]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix880 (.Y (nx879), .A0 (outputRegPage2[10]), .A1 (nx1064)) ;
    dffr regPage2Map_reg_Q_11 (.Q (outputRegPage2[11]), .QB (nx888), .D (nx575)
         , .CLK (clk), .R (rst)) ;
    oai21 ix576 (.Y (nx575), .A0 (nx884), .A1 (nx1064), .B0 (nx886)) ;
    mux21 ix885 (.Y (nx884), .A0 (windowBus[11]), .A1 (regPage1NextUnit[11]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix887 (.Y (nx886), .A0 (outputRegPage2[11]), .A1 (nx1064)) ;
    dffr regPage2Map_reg_Q_12 (.Q (outputRegPage2[12]), .QB (nx895), .D (nx595)
         , .CLK (clk), .R (rst)) ;
    oai21 ix596 (.Y (nx595), .A0 (nx891), .A1 (nx1064), .B0 (nx893)) ;
    mux21 ix892 (.Y (nx891), .A0 (windowBus[12]), .A1 (regPage1NextUnit[12]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix894 (.Y (nx893), .A0 (outputRegPage2[12]), .A1 (nx1064)) ;
    dffr regPage2Map_reg_Q_13 (.Q (outputRegPage2[13]), .QB (nx902), .D (nx615)
         , .CLK (clk), .R (rst)) ;
    oai21 ix616 (.Y (nx615), .A0 (nx898), .A1 (nx1064), .B0 (nx900)) ;
    mux21 ix899 (.Y (nx898), .A0 (windowBus[13]), .A1 (regPage1NextUnit[13]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix901 (.Y (nx900), .A0 (outputRegPage2[13]), .A1 (nx1064)) ;
    dffr regPage2Map_reg_Q_14 (.Q (outputRegPage2[14]), .QB (nx909), .D (nx635)
         , .CLK (clk), .R (rst)) ;
    oai21 ix636 (.Y (nx635), .A0 (nx905), .A1 (nx1066), .B0 (nx907)) ;
    mux21 ix906 (.Y (nx905), .A0 (windowBus[14]), .A1 (regPage1NextUnit[14]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix908 (.Y (nx907), .A0 (outputRegPage2[14]), .A1 (nx1066)) ;
    dffr regPage2Map_reg_Q_15 (.Q (outputRegPage2[15]), .QB (nx916), .D (nx655)
         , .CLK (clk), .R (rst)) ;
    oai21 ix656 (.Y (nx655), .A0 (nx912), .A1 (nx1066), .B0 (nx914)) ;
    mux21 ix913 (.Y (nx912), .A0 (windowBus[15]), .A1 (regPage1NextUnit[15]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix915 (.Y (nx914), .A0 (outputRegPage2[15]), .A1 (nx1066)) ;
    dffr regPage1Map_reg_Q_0 (.Q (outputRegPage1[0]), .QB (nx925), .D (nx345), .CLK (
         clk), .R (rst)) ;
    oai21 ix346 (.Y (nx345), .A0 (nx919), .A1 (nx1070), .B0 (nx923)) ;
    mux21 ix920 (.Y (nx919), .A0 (windowBus[0]), .A1 (regPage2NextUnit[0]), .S0 (
          page1ReadBusOrPage2)) ;
    nor02_2x ix922 (.Y (nx921), .A0 (enableRegPage1), .A1 (page1ReadBusOrPage2)
             ) ;
    nand02 ix924 (.Y (nx923), .A0 (outputRegPage1[0]), .A1 (nx1070)) ;
    dffr regPage1Map_reg_Q_1 (.Q (outputRegPage1[1]), .QB (nx932), .D (nx365), .CLK (
         clk), .R (rst)) ;
    oai21 ix366 (.Y (nx365), .A0 (nx928), .A1 (nx1070), .B0 (nx930)) ;
    mux21 ix929 (.Y (nx928), .A0 (windowBus[1]), .A1 (regPage2NextUnit[1]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix931 (.Y (nx930), .A0 (outputRegPage1[1]), .A1 (nx1070)) ;
    dffr regPage1Map_reg_Q_2 (.Q (outputRegPage1[2]), .QB (nx939), .D (nx385), .CLK (
         clk), .R (rst)) ;
    oai21 ix386 (.Y (nx385), .A0 (nx935), .A1 (nx1070), .B0 (nx937)) ;
    mux21 ix936 (.Y (nx935), .A0 (windowBus[2]), .A1 (regPage2NextUnit[2]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix938 (.Y (nx937), .A0 (outputRegPage1[2]), .A1 (nx1070)) ;
    dffr regPage1Map_reg_Q_3 (.Q (outputRegPage1[3]), .QB (nx946), .D (nx405), .CLK (
         clk), .R (rst)) ;
    oai21 ix406 (.Y (nx405), .A0 (nx942), .A1 (nx1070), .B0 (nx944)) ;
    mux21 ix943 (.Y (nx942), .A0 (windowBus[3]), .A1 (regPage2NextUnit[3]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix945 (.Y (nx944), .A0 (outputRegPage1[3]), .A1 (nx1072)) ;
    dffr regPage1Map_reg_Q_4 (.Q (outputRegPage1[4]), .QB (nx953), .D (nx425), .CLK (
         clk), .R (rst)) ;
    oai21 ix426 (.Y (nx425), .A0 (nx949), .A1 (nx1072), .B0 (nx951)) ;
    mux21 ix950 (.Y (nx949), .A0 (windowBus[4]), .A1 (regPage2NextUnit[4]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix952 (.Y (nx951), .A0 (outputRegPage1[4]), .A1 (nx1072)) ;
    dffr regPage1Map_reg_Q_5 (.Q (outputRegPage1[5]), .QB (nx960), .D (nx445), .CLK (
         clk), .R (rst)) ;
    oai21 ix446 (.Y (nx445), .A0 (nx956), .A1 (nx1072), .B0 (nx958)) ;
    mux21 ix957 (.Y (nx956), .A0 (windowBus[5]), .A1 (regPage2NextUnit[5]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix959 (.Y (nx958), .A0 (outputRegPage1[5]), .A1 (nx1072)) ;
    dffr regPage1Map_reg_Q_6 (.Q (outputRegPage1[6]), .QB (nx967), .D (nx465), .CLK (
         clk), .R (rst)) ;
    oai21 ix466 (.Y (nx465), .A0 (nx963), .A1 (nx1072), .B0 (nx965)) ;
    mux21 ix964 (.Y (nx963), .A0 (windowBus[6]), .A1 (regPage2NextUnit[6]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix966 (.Y (nx965), .A0 (outputRegPage1[6]), .A1 (nx1072)) ;
    dffr regPage1Map_reg_Q_7 (.Q (outputRegPage1[7]), .QB (nx974), .D (nx485), .CLK (
         clk), .R (rst)) ;
    oai21 ix486 (.Y (nx485), .A0 (nx970), .A1 (nx1074), .B0 (nx972)) ;
    mux21 ix971 (.Y (nx970), .A0 (windowBus[7]), .A1 (regPage2NextUnit[7]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix973 (.Y (nx972), .A0 (outputRegPage1[7]), .A1 (nx1074)) ;
    dffr regPage1Map_reg_Q_8 (.Q (outputRegPage1[8]), .QB (nx981), .D (nx505), .CLK (
         clk), .R (rst)) ;
    oai21 ix506 (.Y (nx505), .A0 (nx977), .A1 (nx1074), .B0 (nx979)) ;
    mux21 ix978 (.Y (nx977), .A0 (windowBus[8]), .A1 (regPage2NextUnit[8]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix980 (.Y (nx979), .A0 (outputRegPage1[8]), .A1 (nx1074)) ;
    dffr regPage1Map_reg_Q_9 (.Q (outputRegPage1[9]), .QB (nx988), .D (nx525), .CLK (
         clk), .R (rst)) ;
    oai21 ix526 (.Y (nx525), .A0 (nx984), .A1 (nx1074), .B0 (nx986)) ;
    mux21 ix985 (.Y (nx984), .A0 (windowBus[9]), .A1 (regPage2NextUnit[9]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix987 (.Y (nx986), .A0 (outputRegPage1[9]), .A1 (nx1074)) ;
    dffr regPage1Map_reg_Q_10 (.Q (outputRegPage1[10]), .QB (nx995), .D (nx545)
         , .CLK (clk), .R (rst)) ;
    oai21 ix546 (.Y (nx545), .A0 (nx991), .A1 (nx1074), .B0 (nx993)) ;
    mux21 ix992 (.Y (nx991), .A0 (windowBus[10]), .A1 (regPage2NextUnit[10]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix994 (.Y (nx993), .A0 (outputRegPage1[10]), .A1 (nx1076)) ;
    dffr regPage1Map_reg_Q_11 (.Q (outputRegPage1[11]), .QB (nx1002), .D (nx565)
         , .CLK (clk), .R (rst)) ;
    oai21 ix566 (.Y (nx565), .A0 (nx998), .A1 (nx1076), .B0 (nx1000)) ;
    mux21 ix999 (.Y (nx998), .A0 (windowBus[11]), .A1 (regPage2NextUnit[11]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix1001 (.Y (nx1000), .A0 (outputRegPage1[11]), .A1 (nx1076)) ;
    dffr regPage1Map_reg_Q_12 (.Q (outputRegPage1[12]), .QB (nx1009), .D (nx585)
         , .CLK (clk), .R (rst)) ;
    oai21 ix586 (.Y (nx585), .A0 (nx1005), .A1 (nx1076), .B0 (nx1007)) ;
    mux21 ix1006 (.Y (nx1005), .A0 (windowBus[12]), .A1 (regPage2NextUnit[12]), 
          .S0 (page1ReadBusOrPage2)) ;
    nand02 ix1008 (.Y (nx1007), .A0 (outputRegPage1[12]), .A1 (nx1076)) ;
    dffr regPage1Map_reg_Q_13 (.Q (outputRegPage1[13]), .QB (nx1016), .D (nx605)
         , .CLK (clk), .R (rst)) ;
    oai21 ix606 (.Y (nx605), .A0 (nx1012), .A1 (nx1076), .B0 (nx1014)) ;
    mux21 ix1013 (.Y (nx1012), .A0 (windowBus[13]), .A1 (regPage2NextUnit[13]), 
          .S0 (page1ReadBusOrPage2)) ;
    nand02 ix1015 (.Y (nx1014), .A0 (outputRegPage1[13]), .A1 (nx1076)) ;
    dffr regPage1Map_reg_Q_14 (.Q (outputRegPage1[14]), .QB (nx1023), .D (nx625)
         , .CLK (clk), .R (rst)) ;
    oai21 ix626 (.Y (nx625), .A0 (nx1019), .A1 (nx1078), .B0 (nx1021)) ;
    mux21 ix1020 (.Y (nx1019), .A0 (windowBus[14]), .A1 (regPage2NextUnit[14]), 
          .S0 (page1ReadBusOrPage2)) ;
    nand02 ix1022 (.Y (nx1021), .A0 (outputRegPage1[14]), .A1 (nx1078)) ;
    dffr regPage1Map_reg_Q_15 (.Q (outputRegPage1[15]), .QB (nx1030), .D (nx645)
         , .CLK (clk), .R (rst)) ;
    oai21 ix646 (.Y (nx645), .A0 (nx1026), .A1 (nx1078), .B0 (nx1028)) ;
    mux21 ix1027 (.Y (nx1026), .A0 (windowBus[15]), .A1 (regPage2NextUnit[15]), 
          .S0 (page1ReadBusOrPage2)) ;
    nand02 ix1029 (.Y (nx1028), .A0 (outputRegPage1[15]), .A1 (nx1078)) ;
    mux21 ix33 (.Y (outRegPage[0]), .A0 (nx925), .A1 (nx811), .S0 (pageTurn)) ;
    mux21 ix61 (.Y (outRegPage[1]), .A0 (nx932), .A1 (nx818), .S0 (pageTurn)) ;
    mux21 ix89 (.Y (outRegPage[2]), .A0 (nx939), .A1 (nx825), .S0 (pageTurn)) ;
    mux21 ix117 (.Y (outRegPage[3]), .A0 (nx946), .A1 (nx832), .S0 (pageTurn)) ;
    mux21 ix145 (.Y (outRegPage[4]), .A0 (nx953), .A1 (nx839), .S0 (pageTurn)) ;
    mux21 ix173 (.Y (outRegPage[5]), .A0 (nx960), .A1 (nx846), .S0 (pageTurn)) ;
    mux21 ix201 (.Y (outRegPage[6]), .A0 (nx967), .A1 (nx853), .S0 (pageTurn)) ;
    mux21 ix229 (.Y (outRegPage[7]), .A0 (nx974), .A1 (nx860), .S0 (pageTurn)) ;
    mux21 ix257 (.Y (outRegPage[8]), .A0 (nx981), .A1 (nx867), .S0 (pageTurn)) ;
    mux21 ix285 (.Y (outRegPage[9]), .A0 (nx988), .A1 (nx874), .S0 (pageTurn)) ;
    mux21 ix313 (.Y (outRegPage[10]), .A0 (nx995), .A1 (nx881), .S0 (pageTurn)
          ) ;
    mux21 ix341 (.Y (outRegPage[11]), .A0 (nx1002), .A1 (nx888), .S0 (pageTurn)
          ) ;
    mux21 ix369 (.Y (outRegPage[12]), .A0 (nx1009), .A1 (nx895), .S0 (pageTurn)
          ) ;
    mux21 ix397 (.Y (outRegPage[13]), .A0 (nx1016), .A1 (nx902), .S0 (pageTurn)
          ) ;
    mux21 ix425 (.Y (outRegPage[14]), .A0 (nx1023), .A1 (nx909), .S0 (pageTurn)
          ) ;
    mux21 ix453 (.Y (outRegPage[15]), .A0 (nx1030), .A1 (nx916), .S0 (pageTurn)
          ) ;
    inv01 ix1053 (.Y (nx1054), .A (nx1086)) ;
    inv01 ix1055 (.Y (nx1056), .A (nx807)) ;
    inv02 ix1057 (.Y (nx1058), .A (nx1056)) ;
    inv02 ix1059 (.Y (nx1060), .A (nx1056)) ;
    inv02 ix1061 (.Y (nx1062), .A (nx1056)) ;
    inv02 ix1063 (.Y (nx1064), .A (nx1056)) ;
    inv02 ix1065 (.Y (nx1066), .A (nx1056)) ;
    inv01 ix1067 (.Y (nx1068), .A (nx921)) ;
    inv02 ix1069 (.Y (nx1070), .A (nx1068)) ;
    inv02 ix1071 (.Y (nx1072), .A (nx1068)) ;
    inv02 ix1073 (.Y (nx1074), .A (nx1068)) ;
    inv02 ix1075 (.Y (nx1076), .A (nx1068)) ;
    inv02 ix1077 (.Y (nx1078), .A (nx1068)) ;
    inv02 ix1083 (.Y (nx1084), .A (nx1090)) ;
    inv02 ix1085 (.Y (nx1086), .A (nx1090)) ;
    inv02 ix1087 (.Y (nx1088), .A (enableRegFilter)) ;
    inv02 ix1089 (.Y (nx1090), .A (enableRegFilter)) ;
endmodule


module RegUnit_8_16 ( filterBus, windowBus, regPage1NextUnit, regPage2NextUnit, 
                      clk, rst, enableRegPage1, enableRegPage2, enableRegFilter, 
                      page1ReadBusOrPage2, page2ReadBusOrPage1, pageTurn, 
                      outRegPage, outputRegPage1, outputRegPage2, outFilter ) ;

    input [7:0]filterBus ;
    input [15:0]windowBus ;
    input [15:0]regPage1NextUnit ;
    input [15:0]regPage2NextUnit ;
    input clk ;
    input rst ;
    input enableRegPage1 ;
    input enableRegPage2 ;
    input enableRegFilter ;
    input page1ReadBusOrPage2 ;
    input page2ReadBusOrPage1 ;
    input pageTurn ;
    output [15:0]outRegPage ;
    output [15:0]outputRegPage1 ;
    output [15:0]outputRegPage2 ;
    output [7:0]outFilter ;

    wire outputRegPage1_0_rename, outputRegPage2_0_rename, 
         outputRegPage1_1_rename, outputRegPage2_1_rename, 
         outputRegPage1_2_rename, outputRegPage2_2_rename, 
         outputRegPage1_3_rename, outputRegPage2_3_rename, 
         outputRegPage1_4_rename, outputRegPage2_4_rename, 
         outputRegPage1_5_rename, outputRegPage2_5_rename, 
         outputRegPage1_6_rename, outputRegPage2_6_rename, 
         outputRegPage1_7_rename, outputRegPage2_7_rename, 
         outputRegPage1_8_rename, outputRegPage2_8_rename, 
         outputRegPage1_9_rename, outputRegPage2_9_rename, 
         outputRegPage1_10_rename, outputRegPage2_10_rename, 
         outputRegPage1_11_rename, outputRegPage2_11_rename, 
         outputRegPage1_12_rename, outputRegPage2_12_rename, 
         outputRegPage1_13_rename, outputRegPage2_13_rename, 
         outputRegPage1_14_rename, outputRegPage2_14_rename, 
         outputRegPage1_15_rename, outputRegPage2_15_rename, nx133, nx143, nx153, 
         nx163, nx173, nx183, nx193, nx203, nx213, nx223, nx233, nx243, nx253, 
         nx263, nx273, nx283, nx293, nx303, nx313, nx323, nx333, nx343, nx353, 
         nx363, nx373, nx383, nx393, nx403, nx413, nx423, nx433, nx443, nx453, 
         nx463, nx473, nx483, nx493, nx503, nx513, nx523, nx535, nx539, nx544, 
         nx546, nx551, nx553, nx558, nx560, nx565, nx567, nx572, nx574, nx579, 
         nx581, nx586, nx588, nx592, nx595, nx597, nx599, nx602, nx605, nx607, 
         nx609, nx613, nx616, nx618, nx621, nx624, nx626, nx630, nx633, nx635, 
         nx638, nx641, nx643, nx647, nx650, nx652, nx655, nx658, nx660, nx664, 
         nx667, nx669, nx672, nx675, nx677, nx681, nx684, nx686, nx689, nx692, 
         nx694, nx698, nx701, nx703, nx706, nx709, nx711, nx715, nx718, nx720, 
         nx723, nx726, nx728, nx732, nx735, nx737, nx740, nx743, nx745, nx749, 
         nx752, nx754, nx757, nx760, nx762, nx766, nx769, nx771, nx774, nx777, 
         nx779, nx783, nx786, nx788, nx791, nx794, nx796, nx800, nx803, nx805, 
         nx808, nx811, nx813, nx817, nx820, nx822, nx825, nx828, nx830, nx834, 
         nx837, nx839, nx842, nx845, nx847, nx851, nx854, nx856, nx859, nx862, 
         nx864, nx874, nx876, nx878, nx880, nx882, nx884, nx886, nx888, nx890, 
         nx892, nx894, nx896, nx898, nx904, nx906, nx908, nx910;
    wire [7:0] \$dummy ;




    assign outputRegPage1[14] = outputRegPage1[15] ;
    assign outputRegPage1[13] = outputRegPage1[15] ;
    assign outputRegPage1[12] = outputRegPage1[15] ;
    assign outputRegPage1[11] = outputRegPage1[15] ;
    assign outputRegPage1[10] = outputRegPage1[15] ;
    assign outputRegPage1[9] = outputRegPage1[15] ;
    assign outputRegPage1[8] = outputRegPage1[15] ;
    assign outputRegPage1[7] = outputRegPage1[15] ;
    assign outputRegPage1[6] = outputRegPage1[15] ;
    assign outputRegPage1[5] = outputRegPage1[15] ;
    assign outputRegPage1[4] = outputRegPage1[15] ;
    assign outputRegPage1[3] = outputRegPage1[15] ;
    assign outputRegPage1[2] = outputRegPage1[15] ;
    assign outputRegPage1[1] = outputRegPage1[15] ;
    assign outputRegPage1[0] = outputRegPage1[15] ;
    assign outputRegPage2[15] = outputRegPage1[15] ;
    assign outputRegPage2[14] = outputRegPage1[15] ;
    assign outputRegPage2[13] = outputRegPage1[15] ;
    assign outputRegPage2[12] = outputRegPage1[15] ;
    assign outputRegPage2[11] = outputRegPage1[15] ;
    assign outputRegPage2[10] = outputRegPage1[15] ;
    assign outputRegPage2[9] = outputRegPage1[15] ;
    assign outputRegPage2[8] = outputRegPage1[15] ;
    assign outputRegPage2[7] = outputRegPage1[15] ;
    assign outputRegPage2[6] = outputRegPage1[15] ;
    assign outputRegPage2[5] = outputRegPage1[15] ;
    assign outputRegPage2[4] = outputRegPage1[15] ;
    assign outputRegPage2[3] = outputRegPage1[15] ;
    assign outputRegPage2[2] = outputRegPage1[15] ;
    assign outputRegPage2[1] = outputRegPage1[15] ;
    assign outputRegPage2[0] = outputRegPage1[15] ;
    fake_gnd ix54 (.Y (outputRegPage1[15])) ;
    dffr regFilterMap_reg_Q_0 (.Q (outFilter[0]), .QB (\$dummy [0]), .D (nx453)
         , .CLK (clk), .R (rst)) ;
    nand02 ix454 (.Y (nx453), .A0 (nx535), .A1 (nx539)) ;
    nand02 ix536 (.Y (nx535), .A0 (outFilter[0]), .A1 (nx908)) ;
    nand02 ix540 (.Y (nx539), .A0 (filterBus[0]), .A1 (nx904)) ;
    dffr regFilterMap_reg_Q_1 (.Q (outFilter[1]), .QB (\$dummy [1]), .D (nx463)
         , .CLK (clk), .R (rst)) ;
    nand02 ix464 (.Y (nx463), .A0 (nx544), .A1 (nx546)) ;
    nand02 ix545 (.Y (nx544), .A0 (outFilter[1]), .A1 (nx908)) ;
    nand02 ix547 (.Y (nx546), .A0 (filterBus[1]), .A1 (nx904)) ;
    dffr regFilterMap_reg_Q_2 (.Q (outFilter[2]), .QB (\$dummy [2]), .D (nx473)
         , .CLK (clk), .R (rst)) ;
    nand02 ix474 (.Y (nx473), .A0 (nx551), .A1 (nx553)) ;
    nand02 ix552 (.Y (nx551), .A0 (outFilter[2]), .A1 (nx908)) ;
    nand02 ix554 (.Y (nx553), .A0 (filterBus[2]), .A1 (nx904)) ;
    dffr regFilterMap_reg_Q_3 (.Q (outFilter[3]), .QB (\$dummy [3]), .D (nx483)
         , .CLK (clk), .R (rst)) ;
    nand02 ix484 (.Y (nx483), .A0 (nx558), .A1 (nx560)) ;
    nand02 ix559 (.Y (nx558), .A0 (outFilter[3]), .A1 (nx908)) ;
    nand02 ix561 (.Y (nx560), .A0 (filterBus[3]), .A1 (nx904)) ;
    dffr regFilterMap_reg_Q_4 (.Q (outFilter[4]), .QB (\$dummy [4]), .D (nx493)
         , .CLK (clk), .R (rst)) ;
    nand02 ix494 (.Y (nx493), .A0 (nx565), .A1 (nx567)) ;
    nand02 ix566 (.Y (nx565), .A0 (outFilter[4]), .A1 (nx908)) ;
    nand02 ix568 (.Y (nx567), .A0 (filterBus[4]), .A1 (nx904)) ;
    dffr regFilterMap_reg_Q_5 (.Q (outFilter[5]), .QB (\$dummy [5]), .D (nx503)
         , .CLK (clk), .R (rst)) ;
    nand02 ix504 (.Y (nx503), .A0 (nx572), .A1 (nx574)) ;
    nand02 ix573 (.Y (nx572), .A0 (outFilter[5]), .A1 (nx908)) ;
    nand02 ix575 (.Y (nx574), .A0 (filterBus[5]), .A1 (nx904)) ;
    dffr regFilterMap_reg_Q_6 (.Q (outFilter[6]), .QB (\$dummy [6]), .D (nx513)
         , .CLK (clk), .R (rst)) ;
    nand02 ix514 (.Y (nx513), .A0 (nx579), .A1 (nx581)) ;
    nand02 ix580 (.Y (nx579), .A0 (outFilter[6]), .A1 (nx908)) ;
    nand02 ix582 (.Y (nx581), .A0 (filterBus[6]), .A1 (nx904)) ;
    dffr regFilterMap_reg_Q_7 (.Q (outFilter[7]), .QB (\$dummy [7]), .D (nx523)
         , .CLK (clk), .R (rst)) ;
    nand02 ix524 (.Y (nx523), .A0 (nx586), .A1 (nx588)) ;
    nand02 ix587 (.Y (nx586), .A0 (outFilter[7]), .A1 (nx874)) ;
    nand02 ix589 (.Y (nx588), .A0 (filterBus[7]), .A1 (nx906)) ;
    mux21 ix33 (.Y (outRegPage[0]), .A0 (nx592), .A1 (nx602), .S0 (pageTurn)) ;
    oai21 ix134 (.Y (nx133), .A0 (nx595), .A1 (nx878), .B0 (nx599)) ;
    mux21 ix596 (.Y (nx595), .A0 (windowBus[0]), .A1 (regPage2NextUnit[0]), .S0 (
          page1ReadBusOrPage2)) ;
    nor02_2x ix598 (.Y (nx597), .A0 (enableRegPage1), .A1 (page1ReadBusOrPage2)
             ) ;
    nand02 ix600 (.Y (nx599), .A0 (outputRegPage1_0_rename), .A1 (nx878)) ;
    dffr regPage1Map_reg_Q_0 (.Q (outputRegPage1_0_rename), .QB (nx592), .D (
         nx133), .CLK (clk), .R (rst)) ;
    oai21 ix144 (.Y (nx143), .A0 (nx605), .A1 (nx890), .B0 (nx609)) ;
    mux21 ix606 (.Y (nx605), .A0 (windowBus[0]), .A1 (regPage1NextUnit[0]), .S0 (
          page2ReadBusOrPage1)) ;
    nor02_2x ix608 (.Y (nx607), .A0 (enableRegPage2), .A1 (page2ReadBusOrPage1)
             ) ;
    nand02 ix610 (.Y (nx609), .A0 (outputRegPage2_0_rename), .A1 (nx890)) ;
    dffr regPage2Map_reg_Q_0 (.Q (outputRegPage2_0_rename), .QB (nx602), .D (
         nx143), .CLK (clk), .R (rst)) ;
    mux21 ix61 (.Y (outRegPage[1]), .A0 (nx613), .A1 (nx621), .S0 (pageTurn)) ;
    oai21 ix154 (.Y (nx153), .A0 (nx616), .A1 (nx878), .B0 (nx618)) ;
    mux21 ix617 (.Y (nx616), .A0 (windowBus[1]), .A1 (regPage2NextUnit[1]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix619 (.Y (nx618), .A0 (outputRegPage1_1_rename), .A1 (nx878)) ;
    dffr regPage1Map_reg_Q_1 (.Q (outputRegPage1_1_rename), .QB (nx613), .D (
         nx153), .CLK (clk), .R (rst)) ;
    oai21 ix164 (.Y (nx163), .A0 (nx624), .A1 (nx890), .B0 (nx626)) ;
    mux21 ix625 (.Y (nx624), .A0 (windowBus[1]), .A1 (regPage1NextUnit[1]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix627 (.Y (nx626), .A0 (outputRegPage2_1_rename), .A1 (nx890)) ;
    dffr regPage2Map_reg_Q_1 (.Q (outputRegPage2_1_rename), .QB (nx621), .D (
         nx163), .CLK (clk), .R (rst)) ;
    mux21 ix89 (.Y (outRegPage[2]), .A0 (nx630), .A1 (nx638), .S0 (pageTurn)) ;
    oai21 ix174 (.Y (nx173), .A0 (nx633), .A1 (nx878), .B0 (nx635)) ;
    mux21 ix634 (.Y (nx633), .A0 (windowBus[2]), .A1 (regPage2NextUnit[2]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix636 (.Y (nx635), .A0 (outputRegPage1_2_rename), .A1 (nx878)) ;
    dffr regPage1Map_reg_Q_2 (.Q (outputRegPage1_2_rename), .QB (nx630), .D (
         nx173), .CLK (clk), .R (rst)) ;
    oai21 ix184 (.Y (nx183), .A0 (nx641), .A1 (nx890), .B0 (nx643)) ;
    mux21 ix642 (.Y (nx641), .A0 (windowBus[2]), .A1 (regPage1NextUnit[2]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix644 (.Y (nx643), .A0 (outputRegPage2_2_rename), .A1 (nx890)) ;
    dffr regPage2Map_reg_Q_2 (.Q (outputRegPage2_2_rename), .QB (nx638), .D (
         nx183), .CLK (clk), .R (rst)) ;
    mux21 ix117 (.Y (outRegPage[3]), .A0 (nx647), .A1 (nx655), .S0 (pageTurn)) ;
    oai21 ix194 (.Y (nx193), .A0 (nx650), .A1 (nx878), .B0 (nx652)) ;
    mux21 ix651 (.Y (nx650), .A0 (windowBus[3]), .A1 (regPage2NextUnit[3]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix653 (.Y (nx652), .A0 (outputRegPage1_3_rename), .A1 (nx880)) ;
    dffr regPage1Map_reg_Q_3 (.Q (outputRegPage1_3_rename), .QB (nx647), .D (
         nx193), .CLK (clk), .R (rst)) ;
    oai21 ix204 (.Y (nx203), .A0 (nx658), .A1 (nx890), .B0 (nx660)) ;
    mux21 ix659 (.Y (nx658), .A0 (windowBus[3]), .A1 (regPage1NextUnit[3]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix661 (.Y (nx660), .A0 (outputRegPage2_3_rename), .A1 (nx892)) ;
    dffr regPage2Map_reg_Q_3 (.Q (outputRegPage2_3_rename), .QB (nx655), .D (
         nx203), .CLK (clk), .R (rst)) ;
    mux21 ix145 (.Y (outRegPage[4]), .A0 (nx664), .A1 (nx672), .S0 (pageTurn)) ;
    oai21 ix214 (.Y (nx213), .A0 (nx667), .A1 (nx880), .B0 (nx669)) ;
    mux21 ix668 (.Y (nx667), .A0 (windowBus[4]), .A1 (regPage2NextUnit[4]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix670 (.Y (nx669), .A0 (outputRegPage1_4_rename), .A1 (nx880)) ;
    dffr regPage1Map_reg_Q_4 (.Q (outputRegPage1_4_rename), .QB (nx664), .D (
         nx213), .CLK (clk), .R (rst)) ;
    oai21 ix224 (.Y (nx223), .A0 (nx675), .A1 (nx892), .B0 (nx677)) ;
    mux21 ix676 (.Y (nx675), .A0 (windowBus[4]), .A1 (regPage1NextUnit[4]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix678 (.Y (nx677), .A0 (outputRegPage2_4_rename), .A1 (nx892)) ;
    dffr regPage2Map_reg_Q_4 (.Q (outputRegPage2_4_rename), .QB (nx672), .D (
         nx223), .CLK (clk), .R (rst)) ;
    mux21 ix173 (.Y (outRegPage[5]), .A0 (nx681), .A1 (nx689), .S0 (pageTurn)) ;
    oai21 ix234 (.Y (nx233), .A0 (nx684), .A1 (nx880), .B0 (nx686)) ;
    mux21 ix685 (.Y (nx684), .A0 (windowBus[5]), .A1 (regPage2NextUnit[5]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix687 (.Y (nx686), .A0 (outputRegPage1_5_rename), .A1 (nx880)) ;
    dffr regPage1Map_reg_Q_5 (.Q (outputRegPage1_5_rename), .QB (nx681), .D (
         nx233), .CLK (clk), .R (rst)) ;
    oai21 ix244 (.Y (nx243), .A0 (nx692), .A1 (nx892), .B0 (nx694)) ;
    mux21 ix693 (.Y (nx692), .A0 (windowBus[5]), .A1 (regPage1NextUnit[5]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix695 (.Y (nx694), .A0 (outputRegPage2_5_rename), .A1 (nx892)) ;
    dffr regPage2Map_reg_Q_5 (.Q (outputRegPage2_5_rename), .QB (nx689), .D (
         nx243), .CLK (clk), .R (rst)) ;
    mux21 ix201 (.Y (outRegPage[6]), .A0 (nx698), .A1 (nx706), .S0 (pageTurn)) ;
    oai21 ix254 (.Y (nx253), .A0 (nx701), .A1 (nx880), .B0 (nx703)) ;
    mux21 ix702 (.Y (nx701), .A0 (windowBus[6]), .A1 (regPage2NextUnit[6]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix704 (.Y (nx703), .A0 (outputRegPage1_6_rename), .A1 (nx880)) ;
    dffr regPage1Map_reg_Q_6 (.Q (outputRegPage1_6_rename), .QB (nx698), .D (
         nx253), .CLK (clk), .R (rst)) ;
    oai21 ix264 (.Y (nx263), .A0 (nx709), .A1 (nx892), .B0 (nx711)) ;
    mux21 ix710 (.Y (nx709), .A0 (windowBus[6]), .A1 (regPage1NextUnit[6]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix712 (.Y (nx711), .A0 (outputRegPage2_6_rename), .A1 (nx892)) ;
    dffr regPage2Map_reg_Q_6 (.Q (outputRegPage2_6_rename), .QB (nx706), .D (
         nx263), .CLK (clk), .R (rst)) ;
    mux21 ix229 (.Y (outRegPage[7]), .A0 (nx715), .A1 (nx723), .S0 (pageTurn)) ;
    oai21 ix274 (.Y (nx273), .A0 (nx718), .A1 (nx882), .B0 (nx720)) ;
    mux21 ix719 (.Y (nx718), .A0 (windowBus[7]), .A1 (regPage2NextUnit[7]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix721 (.Y (nx720), .A0 (outputRegPage1_7_rename), .A1 (nx882)) ;
    dffr regPage1Map_reg_Q_7 (.Q (outputRegPage1_7_rename), .QB (nx715), .D (
         nx273), .CLK (clk), .R (rst)) ;
    oai21 ix284 (.Y (nx283), .A0 (nx726), .A1 (nx894), .B0 (nx728)) ;
    mux21 ix727 (.Y (nx726), .A0 (windowBus[7]), .A1 (regPage1NextUnit[7]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix729 (.Y (nx728), .A0 (outputRegPage2_7_rename), .A1 (nx894)) ;
    dffr regPage2Map_reg_Q_7 (.Q (outputRegPage2_7_rename), .QB (nx723), .D (
         nx283), .CLK (clk), .R (rst)) ;
    mux21 ix257 (.Y (outRegPage[8]), .A0 (nx732), .A1 (nx740), .S0 (pageTurn)) ;
    oai21 ix294 (.Y (nx293), .A0 (nx735), .A1 (nx882), .B0 (nx737)) ;
    mux21 ix736 (.Y (nx735), .A0 (windowBus[8]), .A1 (regPage2NextUnit[8]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix738 (.Y (nx737), .A0 (outputRegPage1_8_rename), .A1 (nx882)) ;
    dffr regPage1Map_reg_Q_8 (.Q (outputRegPage1_8_rename), .QB (nx732), .D (
         nx293), .CLK (clk), .R (rst)) ;
    oai21 ix304 (.Y (nx303), .A0 (nx743), .A1 (nx894), .B0 (nx745)) ;
    mux21 ix744 (.Y (nx743), .A0 (windowBus[8]), .A1 (regPage1NextUnit[8]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix746 (.Y (nx745), .A0 (outputRegPage2_8_rename), .A1 (nx894)) ;
    dffr regPage2Map_reg_Q_8 (.Q (outputRegPage2_8_rename), .QB (nx740), .D (
         nx303), .CLK (clk), .R (rst)) ;
    mux21 ix285 (.Y (outRegPage[9]), .A0 (nx749), .A1 (nx757), .S0 (pageTurn)) ;
    oai21 ix314 (.Y (nx313), .A0 (nx752), .A1 (nx882), .B0 (nx754)) ;
    mux21 ix753 (.Y (nx752), .A0 (windowBus[9]), .A1 (regPage2NextUnit[9]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix755 (.Y (nx754), .A0 (outputRegPage1_9_rename), .A1 (nx882)) ;
    dffr regPage1Map_reg_Q_9 (.Q (outputRegPage1_9_rename), .QB (nx749), .D (
         nx313), .CLK (clk), .R (rst)) ;
    oai21 ix324 (.Y (nx323), .A0 (nx760), .A1 (nx894), .B0 (nx762)) ;
    mux21 ix761 (.Y (nx760), .A0 (windowBus[9]), .A1 (regPage1NextUnit[9]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix763 (.Y (nx762), .A0 (outputRegPage2_9_rename), .A1 (nx894)) ;
    dffr regPage2Map_reg_Q_9 (.Q (outputRegPage2_9_rename), .QB (nx757), .D (
         nx323), .CLK (clk), .R (rst)) ;
    mux21 ix313 (.Y (outRegPage[10]), .A0 (nx766), .A1 (nx774), .S0 (pageTurn)
          ) ;
    oai21 ix334 (.Y (nx333), .A0 (nx769), .A1 (nx882), .B0 (nx771)) ;
    mux21 ix770 (.Y (nx769), .A0 (windowBus[10]), .A1 (regPage2NextUnit[10]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix772 (.Y (nx771), .A0 (outputRegPage1_10_rename), .A1 (nx884)) ;
    dffr regPage1Map_reg_Q_10 (.Q (outputRegPage1_10_rename), .QB (nx766), .D (
         nx333), .CLK (clk), .R (rst)) ;
    oai21 ix344 (.Y (nx343), .A0 (nx777), .A1 (nx894), .B0 (nx779)) ;
    mux21 ix778 (.Y (nx777), .A0 (windowBus[10]), .A1 (regPage1NextUnit[10]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix780 (.Y (nx779), .A0 (outputRegPage2_10_rename), .A1 (nx896)) ;
    dffr regPage2Map_reg_Q_10 (.Q (outputRegPage2_10_rename), .QB (nx774), .D (
         nx343), .CLK (clk), .R (rst)) ;
    mux21 ix341 (.Y (outRegPage[11]), .A0 (nx783), .A1 (nx791), .S0 (pageTurn)
          ) ;
    oai21 ix354 (.Y (nx353), .A0 (nx786), .A1 (nx884), .B0 (nx788)) ;
    mux21 ix787 (.Y (nx786), .A0 (windowBus[11]), .A1 (regPage2NextUnit[11]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix789 (.Y (nx788), .A0 (outputRegPage1_11_rename), .A1 (nx884)) ;
    dffr regPage1Map_reg_Q_11 (.Q (outputRegPage1_11_rename), .QB (nx783), .D (
         nx353), .CLK (clk), .R (rst)) ;
    oai21 ix364 (.Y (nx363), .A0 (nx794), .A1 (nx896), .B0 (nx796)) ;
    mux21 ix795 (.Y (nx794), .A0 (windowBus[11]), .A1 (regPage1NextUnit[11]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix797 (.Y (nx796), .A0 (outputRegPage2_11_rename), .A1 (nx896)) ;
    dffr regPage2Map_reg_Q_11 (.Q (outputRegPage2_11_rename), .QB (nx791), .D (
         nx363), .CLK (clk), .R (rst)) ;
    mux21 ix369 (.Y (outRegPage[12]), .A0 (nx800), .A1 (nx808), .S0 (pageTurn)
          ) ;
    oai21 ix374 (.Y (nx373), .A0 (nx803), .A1 (nx884), .B0 (nx805)) ;
    mux21 ix804 (.Y (nx803), .A0 (windowBus[12]), .A1 (regPage2NextUnit[12]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix806 (.Y (nx805), .A0 (outputRegPage1_12_rename), .A1 (nx884)) ;
    dffr regPage1Map_reg_Q_12 (.Q (outputRegPage1_12_rename), .QB (nx800), .D (
         nx373), .CLK (clk), .R (rst)) ;
    oai21 ix384 (.Y (nx383), .A0 (nx811), .A1 (nx896), .B0 (nx813)) ;
    mux21 ix812 (.Y (nx811), .A0 (windowBus[12]), .A1 (regPage1NextUnit[12]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix814 (.Y (nx813), .A0 (outputRegPage2_12_rename), .A1 (nx896)) ;
    dffr regPage2Map_reg_Q_12 (.Q (outputRegPage2_12_rename), .QB (nx808), .D (
         nx383), .CLK (clk), .R (rst)) ;
    mux21 ix397 (.Y (outRegPage[13]), .A0 (nx817), .A1 (nx825), .S0 (pageTurn)
          ) ;
    oai21 ix394 (.Y (nx393), .A0 (nx820), .A1 (nx884), .B0 (nx822)) ;
    mux21 ix821 (.Y (nx820), .A0 (windowBus[13]), .A1 (regPage2NextUnit[13]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix823 (.Y (nx822), .A0 (outputRegPage1_13_rename), .A1 (nx884)) ;
    dffr regPage1Map_reg_Q_13 (.Q (outputRegPage1_13_rename), .QB (nx817), .D (
         nx393), .CLK (clk), .R (rst)) ;
    oai21 ix404 (.Y (nx403), .A0 (nx828), .A1 (nx896), .B0 (nx830)) ;
    mux21 ix829 (.Y (nx828), .A0 (windowBus[13]), .A1 (regPage1NextUnit[13]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix831 (.Y (nx830), .A0 (outputRegPage2_13_rename), .A1 (nx896)) ;
    dffr regPage2Map_reg_Q_13 (.Q (outputRegPage2_13_rename), .QB (nx825), .D (
         nx403), .CLK (clk), .R (rst)) ;
    mux21 ix425 (.Y (outRegPage[14]), .A0 (nx834), .A1 (nx842), .S0 (pageTurn)
          ) ;
    oai21 ix414 (.Y (nx413), .A0 (nx837), .A1 (nx886), .B0 (nx839)) ;
    mux21 ix838 (.Y (nx837), .A0 (windowBus[14]), .A1 (regPage2NextUnit[14]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix840 (.Y (nx839), .A0 (outputRegPage1_14_rename), .A1 (nx886)) ;
    dffr regPage1Map_reg_Q_14 (.Q (outputRegPage1_14_rename), .QB (nx834), .D (
         nx413), .CLK (clk), .R (rst)) ;
    oai21 ix424 (.Y (nx423), .A0 (nx845), .A1 (nx898), .B0 (nx847)) ;
    mux21 ix846 (.Y (nx845), .A0 (windowBus[14]), .A1 (regPage1NextUnit[14]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix848 (.Y (nx847), .A0 (outputRegPage2_14_rename), .A1 (nx898)) ;
    dffr regPage2Map_reg_Q_14 (.Q (outputRegPage2_14_rename), .QB (nx842), .D (
         nx423), .CLK (clk), .R (rst)) ;
    mux21 ix453 (.Y (outRegPage[15]), .A0 (nx851), .A1 (nx859), .S0 (pageTurn)
          ) ;
    oai21 ix434 (.Y (nx433), .A0 (nx854), .A1 (nx886), .B0 (nx856)) ;
    mux21 ix855 (.Y (nx854), .A0 (windowBus[15]), .A1 (regPage2NextUnit[15]), .S0 (
          page1ReadBusOrPage2)) ;
    nand02 ix857 (.Y (nx856), .A0 (outputRegPage1_15_rename), .A1 (nx886)) ;
    dffr regPage1Map_reg_Q_15 (.Q (outputRegPage1_15_rename), .QB (nx851), .D (
         nx433), .CLK (clk), .R (rst)) ;
    oai21 ix444 (.Y (nx443), .A0 (nx862), .A1 (nx898), .B0 (nx864)) ;
    mux21 ix863 (.Y (nx862), .A0 (windowBus[15]), .A1 (regPage1NextUnit[15]), .S0 (
          page2ReadBusOrPage1)) ;
    nand02 ix865 (.Y (nx864), .A0 (outputRegPage2_15_rename), .A1 (nx898)) ;
    dffr regPage2Map_reg_Q_15 (.Q (outputRegPage2_15_rename), .QB (nx859), .D (
         nx443), .CLK (clk), .R (rst)) ;
    inv01 ix873 (.Y (nx874), .A (nx906)) ;
    inv01 ix875 (.Y (nx876), .A (nx597)) ;
    inv02 ix877 (.Y (nx878), .A (nx876)) ;
    inv02 ix879 (.Y (nx880), .A (nx876)) ;
    inv02 ix881 (.Y (nx882), .A (nx876)) ;
    inv02 ix883 (.Y (nx884), .A (nx876)) ;
    inv02 ix885 (.Y (nx886), .A (nx876)) ;
    inv01 ix887 (.Y (nx888), .A (nx607)) ;
    inv02 ix889 (.Y (nx890), .A (nx888)) ;
    inv02 ix891 (.Y (nx892), .A (nx888)) ;
    inv02 ix893 (.Y (nx894), .A (nx888)) ;
    inv02 ix895 (.Y (nx896), .A (nx888)) ;
    inv02 ix897 (.Y (nx898), .A (nx888)) ;
    inv02 ix903 (.Y (nx904), .A (nx910)) ;
    inv02 ix905 (.Y (nx906), .A (nx910)) ;
    inv02 ix907 (.Y (nx908), .A (enableRegFilter)) ;
    inv02 ix909 (.Y (nx910), .A (enableRegFilter)) ;
endmodule


module CNNMuls_25 ( filter_24__7, filter_24__6, filter_24__5, filter_24__4, 
                    filter_24__3, filter_24__2, filter_24__1, filter_24__0, 
                    filter_23__7, filter_23__6, filter_23__5, filter_23__4, 
                    filter_23__3, filter_23__2, filter_23__1, filter_23__0, 
                    filter_22__7, filter_22__6, filter_22__5, filter_22__4, 
                    filter_22__3, filter_22__2, filter_22__1, filter_22__0, 
                    filter_21__7, filter_21__6, filter_21__5, filter_21__4, 
                    filter_21__3, filter_21__2, filter_21__1, filter_21__0, 
                    filter_20__7, filter_20__6, filter_20__5, filter_20__4, 
                    filter_20__3, filter_20__2, filter_20__1, filter_20__0, 
                    filter_19__7, filter_19__6, filter_19__5, filter_19__4, 
                    filter_19__3, filter_19__2, filter_19__1, filter_19__0, 
                    filter_18__7, filter_18__6, filter_18__5, filter_18__4, 
                    filter_18__3, filter_18__2, filter_18__1, filter_18__0, 
                    filter_17__7, filter_17__6, filter_17__5, filter_17__4, 
                    filter_17__3, filter_17__2, filter_17__1, filter_17__0, 
                    filter_16__7, filter_16__6, filter_16__5, filter_16__4, 
                    filter_16__3, filter_16__2, filter_16__1, filter_16__0, 
                    filter_15__7, filter_15__6, filter_15__5, filter_15__4, 
                    filter_15__3, filter_15__2, filter_15__1, filter_15__0, 
                    filter_14__7, filter_14__6, filter_14__5, filter_14__4, 
                    filter_14__3, filter_14__2, filter_14__1, filter_14__0, 
                    filter_13__7, filter_13__6, filter_13__5, filter_13__4, 
                    filter_13__3, filter_13__2, filter_13__1, filter_13__0, 
                    filter_12__7, filter_12__6, filter_12__5, filter_12__4, 
                    filter_12__3, filter_12__2, filter_12__1, filter_12__0, 
                    filter_11__7, filter_11__6, filter_11__5, filter_11__4, 
                    filter_11__3, filter_11__2, filter_11__1, filter_11__0, 
                    filter_10__7, filter_10__6, filter_10__5, filter_10__4, 
                    filter_10__3, filter_10__2, filter_10__1, filter_10__0, 
                    filter_9__7, filter_9__6, filter_9__5, filter_9__4, 
                    filter_9__3, filter_9__2, filter_9__1, filter_9__0, 
                    filter_8__7, filter_8__6, filter_8__5, filter_8__4, 
                    filter_8__3, filter_8__2, filter_8__1, filter_8__0, 
                    filter_7__7, filter_7__6, filter_7__5, filter_7__4, 
                    filter_7__3, filter_7__2, filter_7__1, filter_7__0, 
                    filter_6__7, filter_6__6, filter_6__5, filter_6__4, 
                    filter_6__3, filter_6__2, filter_6__1, filter_6__0, 
                    filter_5__7, filter_5__6, filter_5__5, filter_5__4, 
                    filter_5__3, filter_5__2, filter_5__1, filter_5__0, 
                    filter_4__7, filter_4__6, filter_4__5, filter_4__4, 
                    filter_4__3, filter_4__2, filter_4__1, filter_4__0, 
                    filter_3__7, filter_3__6, filter_3__5, filter_3__4, 
                    filter_3__3, filter_3__2, filter_3__1, filter_3__0, 
                    filter_2__7, filter_2__6, filter_2__5, filter_2__4, 
                    filter_2__3, filter_2__2, filter_2__1, filter_2__0, 
                    filter_1__7, filter_1__6, filter_1__5, filter_1__4, 
                    filter_1__3, filter_1__2, filter_1__1, filter_1__0, 
                    filter_0__7, filter_0__6, filter_0__5, filter_0__4, 
                    filter_0__3, filter_0__2, filter_0__1, filter_0__0, 
                    window_24__15, window_24__14, window_24__13, window_24__12, 
                    window_24__11, window_24__10, window_24__9, window_24__8, 
                    window_24__7, window_24__6, window_24__5, window_24__4, 
                    window_24__3, window_24__2, window_24__1, window_24__0, 
                    window_23__15, window_23__14, window_23__13, window_23__12, 
                    window_23__11, window_23__10, window_23__9, window_23__8, 
                    window_23__7, window_23__6, window_23__5, window_23__4, 
                    window_23__3, window_23__2, window_23__1, window_23__0, 
                    window_22__15, window_22__14, window_22__13, window_22__12, 
                    window_22__11, window_22__10, window_22__9, window_22__8, 
                    window_22__7, window_22__6, window_22__5, window_22__4, 
                    window_22__3, window_22__2, window_22__1, window_22__0, 
                    window_21__15, window_21__14, window_21__13, window_21__12, 
                    window_21__11, window_21__10, window_21__9, window_21__8, 
                    window_21__7, window_21__6, window_21__5, window_21__4, 
                    window_21__3, window_21__2, window_21__1, window_21__0, 
                    window_20__15, window_20__14, window_20__13, window_20__12, 
                    window_20__11, window_20__10, window_20__9, window_20__8, 
                    window_20__7, window_20__6, window_20__5, window_20__4, 
                    window_20__3, window_20__2, window_20__1, window_20__0, 
                    window_19__15, window_19__14, window_19__13, window_19__12, 
                    window_19__11, window_19__10, window_19__9, window_19__8, 
                    window_19__7, window_19__6, window_19__5, window_19__4, 
                    window_19__3, window_19__2, window_19__1, window_19__0, 
                    window_18__15, window_18__14, window_18__13, window_18__12, 
                    window_18__11, window_18__10, window_18__9, window_18__8, 
                    window_18__7, window_18__6, window_18__5, window_18__4, 
                    window_18__3, window_18__2, window_18__1, window_18__0, 
                    window_17__15, window_17__14, window_17__13, window_17__12, 
                    window_17__11, window_17__10, window_17__9, window_17__8, 
                    window_17__7, window_17__6, window_17__5, window_17__4, 
                    window_17__3, window_17__2, window_17__1, window_17__0, 
                    window_16__15, window_16__14, window_16__13, window_16__12, 
                    window_16__11, window_16__10, window_16__9, window_16__8, 
                    window_16__7, window_16__6, window_16__5, window_16__4, 
                    window_16__3, window_16__2, window_16__1, window_16__0, 
                    window_15__15, window_15__14, window_15__13, window_15__12, 
                    window_15__11, window_15__10, window_15__9, window_15__8, 
                    window_15__7, window_15__6, window_15__5, window_15__4, 
                    window_15__3, window_15__2, window_15__1, window_15__0, 
                    window_14__15, window_14__14, window_14__13, window_14__12, 
                    window_14__11, window_14__10, window_14__9, window_14__8, 
                    window_14__7, window_14__6, window_14__5, window_14__4, 
                    window_14__3, window_14__2, window_14__1, window_14__0, 
                    window_13__15, window_13__14, window_13__13, window_13__12, 
                    window_13__11, window_13__10, window_13__9, window_13__8, 
                    window_13__7, window_13__6, window_13__5, window_13__4, 
                    window_13__3, window_13__2, window_13__1, window_13__0, 
                    window_12__15, window_12__14, window_12__13, window_12__12, 
                    window_12__11, window_12__10, window_12__9, window_12__8, 
                    window_12__7, window_12__6, window_12__5, window_12__4, 
                    window_12__3, window_12__2, window_12__1, window_12__0, 
                    window_11__15, window_11__14, window_11__13, window_11__12, 
                    window_11__11, window_11__10, window_11__9, window_11__8, 
                    window_11__7, window_11__6, window_11__5, window_11__4, 
                    window_11__3, window_11__2, window_11__1, window_11__0, 
                    window_10__15, window_10__14, window_10__13, window_10__12, 
                    window_10__11, window_10__10, window_10__9, window_10__8, 
                    window_10__7, window_10__6, window_10__5, window_10__4, 
                    window_10__3, window_10__2, window_10__1, window_10__0, 
                    window_9__15, window_9__14, window_9__13, window_9__12, 
                    window_9__11, window_9__10, window_9__9, window_9__8, 
                    window_9__7, window_9__6, window_9__5, window_9__4, 
                    window_9__3, window_9__2, window_9__1, window_9__0, 
                    window_8__15, window_8__14, window_8__13, window_8__12, 
                    window_8__11, window_8__10, window_8__9, window_8__8, 
                    window_8__7, window_8__6, window_8__5, window_8__4, 
                    window_8__3, window_8__2, window_8__1, window_8__0, 
                    window_7__15, window_7__14, window_7__13, window_7__12, 
                    window_7__11, window_7__10, window_7__9, window_7__8, 
                    window_7__7, window_7__6, window_7__5, window_7__4, 
                    window_7__3, window_7__2, window_7__1, window_7__0, 
                    window_6__15, window_6__14, window_6__13, window_6__12, 
                    window_6__11, window_6__10, window_6__9, window_6__8, 
                    window_6__7, window_6__6, window_6__5, window_6__4, 
                    window_6__3, window_6__2, window_6__1, window_6__0, 
                    window_5__15, window_5__14, window_5__13, window_5__12, 
                    window_5__11, window_5__10, window_5__9, window_5__8, 
                    window_5__7, window_5__6, window_5__5, window_5__4, 
                    window_5__3, window_5__2, window_5__1, window_5__0, 
                    window_4__15, window_4__14, window_4__13, window_4__12, 
                    window_4__11, window_4__10, window_4__9, window_4__8, 
                    window_4__7, window_4__6, window_4__5, window_4__4, 
                    window_4__3, window_4__2, window_4__1, window_4__0, 
                    window_3__15, window_3__14, window_3__13, window_3__12, 
                    window_3__11, window_3__10, window_3__9, window_3__8, 
                    window_3__7, window_3__6, window_3__5, window_3__4, 
                    window_3__3, window_3__2, window_3__1, window_3__0, 
                    window_2__15, window_2__14, window_2__13, window_2__12, 
                    window_2__11, window_2__10, window_2__9, window_2__8, 
                    window_2__7, window_2__6, window_2__5, window_2__4, 
                    window_2__3, window_2__2, window_2__1, window_2__0, 
                    window_1__15, window_1__14, window_1__13, window_1__12, 
                    window_1__11, window_1__10, window_1__9, window_1__8, 
                    window_1__7, window_1__6, window_1__5, window_1__4, 
                    window_1__3, window_1__2, window_1__1, window_1__0, 
                    window_0__15, window_0__14, window_0__13, window_0__12, 
                    window_0__11, window_0__10, window_0__9, window_0__8, 
                    window_0__7, window_0__6, window_0__5, window_0__4, 
                    window_0__3, window_0__2, window_0__1, window_0__0, 
                    outputs_24__15, outputs_24__14, outputs_24__13, 
                    outputs_24__12, outputs_24__11, outputs_24__10, 
                    outputs_24__9, outputs_24__8, outputs_24__7, outputs_24__6, 
                    outputs_24__5, outputs_24__4, outputs_24__3, outputs_24__2, 
                    outputs_24__1, outputs_24__0, outputs_23__15, outputs_23__14, 
                    outputs_23__13, outputs_23__12, outputs_23__11, 
                    outputs_23__10, outputs_23__9, outputs_23__8, outputs_23__7, 
                    outputs_23__6, outputs_23__5, outputs_23__4, outputs_23__3, 
                    outputs_23__2, outputs_23__1, outputs_23__0, outputs_22__15, 
                    outputs_22__14, outputs_22__13, outputs_22__12, 
                    outputs_22__11, outputs_22__10, outputs_22__9, outputs_22__8, 
                    outputs_22__7, outputs_22__6, outputs_22__5, outputs_22__4, 
                    outputs_22__3, outputs_22__2, outputs_22__1, outputs_22__0, 
                    outputs_21__15, outputs_21__14, outputs_21__13, 
                    outputs_21__12, outputs_21__11, outputs_21__10, 
                    outputs_21__9, outputs_21__8, outputs_21__7, outputs_21__6, 
                    outputs_21__5, outputs_21__4, outputs_21__3, outputs_21__2, 
                    outputs_21__1, outputs_21__0, outputs_20__15, outputs_20__14, 
                    outputs_20__13, outputs_20__12, outputs_20__11, 
                    outputs_20__10, outputs_20__9, outputs_20__8, outputs_20__7, 
                    outputs_20__6, outputs_20__5, outputs_20__4, outputs_20__3, 
                    outputs_20__2, outputs_20__1, outputs_20__0, outputs_19__15, 
                    outputs_19__14, outputs_19__13, outputs_19__12, 
                    outputs_19__11, outputs_19__10, outputs_19__9, outputs_19__8, 
                    outputs_19__7, outputs_19__6, outputs_19__5, outputs_19__4, 
                    outputs_19__3, outputs_19__2, outputs_19__1, outputs_19__0, 
                    outputs_18__15, outputs_18__14, outputs_18__13, 
                    outputs_18__12, outputs_18__11, outputs_18__10, 
                    outputs_18__9, outputs_18__8, outputs_18__7, outputs_18__6, 
                    outputs_18__5, outputs_18__4, outputs_18__3, outputs_18__2, 
                    outputs_18__1, outputs_18__0, outputs_17__15, outputs_17__14, 
                    outputs_17__13, outputs_17__12, outputs_17__11, 
                    outputs_17__10, outputs_17__9, outputs_17__8, outputs_17__7, 
                    outputs_17__6, outputs_17__5, outputs_17__4, outputs_17__3, 
                    outputs_17__2, outputs_17__1, outputs_17__0, outputs_16__15, 
                    outputs_16__14, outputs_16__13, outputs_16__12, 
                    outputs_16__11, outputs_16__10, outputs_16__9, outputs_16__8, 
                    outputs_16__7, outputs_16__6, outputs_16__5, outputs_16__4, 
                    outputs_16__3, outputs_16__2, outputs_16__1, outputs_16__0, 
                    outputs_15__15, outputs_15__14, outputs_15__13, 
                    outputs_15__12, outputs_15__11, outputs_15__10, 
                    outputs_15__9, outputs_15__8, outputs_15__7, outputs_15__6, 
                    outputs_15__5, outputs_15__4, outputs_15__3, outputs_15__2, 
                    outputs_15__1, outputs_15__0, outputs_14__15, outputs_14__14, 
                    outputs_14__13, outputs_14__12, outputs_14__11, 
                    outputs_14__10, outputs_14__9, outputs_14__8, outputs_14__7, 
                    outputs_14__6, outputs_14__5, outputs_14__4, outputs_14__3, 
                    outputs_14__2, outputs_14__1, outputs_14__0, outputs_13__15, 
                    outputs_13__14, outputs_13__13, outputs_13__12, 
                    outputs_13__11, outputs_13__10, outputs_13__9, outputs_13__8, 
                    outputs_13__7, outputs_13__6, outputs_13__5, outputs_13__4, 
                    outputs_13__3, outputs_13__2, outputs_13__1, outputs_13__0, 
                    outputs_12__15, outputs_12__14, outputs_12__13, 
                    outputs_12__12, outputs_12__11, outputs_12__10, 
                    outputs_12__9, outputs_12__8, outputs_12__7, outputs_12__6, 
                    outputs_12__5, outputs_12__4, outputs_12__3, outputs_12__2, 
                    outputs_12__1, outputs_12__0, outputs_11__15, outputs_11__14, 
                    outputs_11__13, outputs_11__12, outputs_11__11, 
                    outputs_11__10, outputs_11__9, outputs_11__8, outputs_11__7, 
                    outputs_11__6, outputs_11__5, outputs_11__4, outputs_11__3, 
                    outputs_11__2, outputs_11__1, outputs_11__0, outputs_10__15, 
                    outputs_10__14, outputs_10__13, outputs_10__12, 
                    outputs_10__11, outputs_10__10, outputs_10__9, outputs_10__8, 
                    outputs_10__7, outputs_10__6, outputs_10__5, outputs_10__4, 
                    outputs_10__3, outputs_10__2, outputs_10__1, outputs_10__0, 
                    outputs_9__15, outputs_9__14, outputs_9__13, outputs_9__12, 
                    outputs_9__11, outputs_9__10, outputs_9__9, outputs_9__8, 
                    outputs_9__7, outputs_9__6, outputs_9__5, outputs_9__4, 
                    outputs_9__3, outputs_9__2, outputs_9__1, outputs_9__0, 
                    outputs_8__15, outputs_8__14, outputs_8__13, outputs_8__12, 
                    outputs_8__11, outputs_8__10, outputs_8__9, outputs_8__8, 
                    outputs_8__7, outputs_8__6, outputs_8__5, outputs_8__4, 
                    outputs_8__3, outputs_8__2, outputs_8__1, outputs_8__0, 
                    outputs_7__15, outputs_7__14, outputs_7__13, outputs_7__12, 
                    outputs_7__11, outputs_7__10, outputs_7__9, outputs_7__8, 
                    outputs_7__7, outputs_7__6, outputs_7__5, outputs_7__4, 
                    outputs_7__3, outputs_7__2, outputs_7__1, outputs_7__0, 
                    outputs_6__15, outputs_6__14, outputs_6__13, outputs_6__12, 
                    outputs_6__11, outputs_6__10, outputs_6__9, outputs_6__8, 
                    outputs_6__7, outputs_6__6, outputs_6__5, outputs_6__4, 
                    outputs_6__3, outputs_6__2, outputs_6__1, outputs_6__0, 
                    outputs_5__15, outputs_5__14, outputs_5__13, outputs_5__12, 
                    outputs_5__11, outputs_5__10, outputs_5__9, outputs_5__8, 
                    outputs_5__7, outputs_5__6, outputs_5__5, outputs_5__4, 
                    outputs_5__3, outputs_5__2, outputs_5__1, outputs_5__0, 
                    outputs_4__15, outputs_4__14, outputs_4__13, outputs_4__12, 
                    outputs_4__11, outputs_4__10, outputs_4__9, outputs_4__8, 
                    outputs_4__7, outputs_4__6, outputs_4__5, outputs_4__4, 
                    outputs_4__3, outputs_4__2, outputs_4__1, outputs_4__0, 
                    outputs_3__15, outputs_3__14, outputs_3__13, outputs_3__12, 
                    outputs_3__11, outputs_3__10, outputs_3__9, outputs_3__8, 
                    outputs_3__7, outputs_3__6, outputs_3__5, outputs_3__4, 
                    outputs_3__3, outputs_3__2, outputs_3__1, outputs_3__0, 
                    outputs_2__15, outputs_2__14, outputs_2__13, outputs_2__12, 
                    outputs_2__11, outputs_2__10, outputs_2__9, outputs_2__8, 
                    outputs_2__7, outputs_2__6, outputs_2__5, outputs_2__4, 
                    outputs_2__3, outputs_2__2, outputs_2__1, outputs_2__0, 
                    outputs_1__15, outputs_1__14, outputs_1__13, outputs_1__12, 
                    outputs_1__11, outputs_1__10, outputs_1__9, outputs_1__8, 
                    outputs_1__7, outputs_1__6, outputs_1__5, outputs_1__4, 
                    outputs_1__3, outputs_1__2, outputs_1__1, outputs_1__0, 
                    outputs_0__15, outputs_0__14, outputs_0__13, outputs_0__12, 
                    outputs_0__11, outputs_0__10, outputs_0__9, outputs_0__8, 
                    outputs_0__7, outputs_0__6, outputs_0__5, outputs_0__4, 
                    outputs_0__3, outputs_0__2, outputs_0__1, outputs_0__0, clk, 
                    start, rst, done, working ) ;

    input filter_24__7 ;
    input filter_24__6 ;
    input filter_24__5 ;
    input filter_24__4 ;
    input filter_24__3 ;
    input filter_24__2 ;
    input filter_24__1 ;
    input filter_24__0 ;
    input filter_23__7 ;
    input filter_23__6 ;
    input filter_23__5 ;
    input filter_23__4 ;
    input filter_23__3 ;
    input filter_23__2 ;
    input filter_23__1 ;
    input filter_23__0 ;
    input filter_22__7 ;
    input filter_22__6 ;
    input filter_22__5 ;
    input filter_22__4 ;
    input filter_22__3 ;
    input filter_22__2 ;
    input filter_22__1 ;
    input filter_22__0 ;
    input filter_21__7 ;
    input filter_21__6 ;
    input filter_21__5 ;
    input filter_21__4 ;
    input filter_21__3 ;
    input filter_21__2 ;
    input filter_21__1 ;
    input filter_21__0 ;
    input filter_20__7 ;
    input filter_20__6 ;
    input filter_20__5 ;
    input filter_20__4 ;
    input filter_20__3 ;
    input filter_20__2 ;
    input filter_20__1 ;
    input filter_20__0 ;
    input filter_19__7 ;
    input filter_19__6 ;
    input filter_19__5 ;
    input filter_19__4 ;
    input filter_19__3 ;
    input filter_19__2 ;
    input filter_19__1 ;
    input filter_19__0 ;
    input filter_18__7 ;
    input filter_18__6 ;
    input filter_18__5 ;
    input filter_18__4 ;
    input filter_18__3 ;
    input filter_18__2 ;
    input filter_18__1 ;
    input filter_18__0 ;
    input filter_17__7 ;
    input filter_17__6 ;
    input filter_17__5 ;
    input filter_17__4 ;
    input filter_17__3 ;
    input filter_17__2 ;
    input filter_17__1 ;
    input filter_17__0 ;
    input filter_16__7 ;
    input filter_16__6 ;
    input filter_16__5 ;
    input filter_16__4 ;
    input filter_16__3 ;
    input filter_16__2 ;
    input filter_16__1 ;
    input filter_16__0 ;
    input filter_15__7 ;
    input filter_15__6 ;
    input filter_15__5 ;
    input filter_15__4 ;
    input filter_15__3 ;
    input filter_15__2 ;
    input filter_15__1 ;
    input filter_15__0 ;
    input filter_14__7 ;
    input filter_14__6 ;
    input filter_14__5 ;
    input filter_14__4 ;
    input filter_14__3 ;
    input filter_14__2 ;
    input filter_14__1 ;
    input filter_14__0 ;
    input filter_13__7 ;
    input filter_13__6 ;
    input filter_13__5 ;
    input filter_13__4 ;
    input filter_13__3 ;
    input filter_13__2 ;
    input filter_13__1 ;
    input filter_13__0 ;
    input filter_12__7 ;
    input filter_12__6 ;
    input filter_12__5 ;
    input filter_12__4 ;
    input filter_12__3 ;
    input filter_12__2 ;
    input filter_12__1 ;
    input filter_12__0 ;
    input filter_11__7 ;
    input filter_11__6 ;
    input filter_11__5 ;
    input filter_11__4 ;
    input filter_11__3 ;
    input filter_11__2 ;
    input filter_11__1 ;
    input filter_11__0 ;
    input filter_10__7 ;
    input filter_10__6 ;
    input filter_10__5 ;
    input filter_10__4 ;
    input filter_10__3 ;
    input filter_10__2 ;
    input filter_10__1 ;
    input filter_10__0 ;
    input filter_9__7 ;
    input filter_9__6 ;
    input filter_9__5 ;
    input filter_9__4 ;
    input filter_9__3 ;
    input filter_9__2 ;
    input filter_9__1 ;
    input filter_9__0 ;
    input filter_8__7 ;
    input filter_8__6 ;
    input filter_8__5 ;
    input filter_8__4 ;
    input filter_8__3 ;
    input filter_8__2 ;
    input filter_8__1 ;
    input filter_8__0 ;
    input filter_7__7 ;
    input filter_7__6 ;
    input filter_7__5 ;
    input filter_7__4 ;
    input filter_7__3 ;
    input filter_7__2 ;
    input filter_7__1 ;
    input filter_7__0 ;
    input filter_6__7 ;
    input filter_6__6 ;
    input filter_6__5 ;
    input filter_6__4 ;
    input filter_6__3 ;
    input filter_6__2 ;
    input filter_6__1 ;
    input filter_6__0 ;
    input filter_5__7 ;
    input filter_5__6 ;
    input filter_5__5 ;
    input filter_5__4 ;
    input filter_5__3 ;
    input filter_5__2 ;
    input filter_5__1 ;
    input filter_5__0 ;
    input filter_4__7 ;
    input filter_4__6 ;
    input filter_4__5 ;
    input filter_4__4 ;
    input filter_4__3 ;
    input filter_4__2 ;
    input filter_4__1 ;
    input filter_4__0 ;
    input filter_3__7 ;
    input filter_3__6 ;
    input filter_3__5 ;
    input filter_3__4 ;
    input filter_3__3 ;
    input filter_3__2 ;
    input filter_3__1 ;
    input filter_3__0 ;
    input filter_2__7 ;
    input filter_2__6 ;
    input filter_2__5 ;
    input filter_2__4 ;
    input filter_2__3 ;
    input filter_2__2 ;
    input filter_2__1 ;
    input filter_2__0 ;
    input filter_1__7 ;
    input filter_1__6 ;
    input filter_1__5 ;
    input filter_1__4 ;
    input filter_1__3 ;
    input filter_1__2 ;
    input filter_1__1 ;
    input filter_1__0 ;
    input filter_0__7 ;
    input filter_0__6 ;
    input filter_0__5 ;
    input filter_0__4 ;
    input filter_0__3 ;
    input filter_0__2 ;
    input filter_0__1 ;
    input filter_0__0 ;
    input window_24__15 ;
    input window_24__14 ;
    input window_24__13 ;
    input window_24__12 ;
    input window_24__11 ;
    input window_24__10 ;
    input window_24__9 ;
    input window_24__8 ;
    input window_24__7 ;
    input window_24__6 ;
    input window_24__5 ;
    input window_24__4 ;
    input window_24__3 ;
    input window_24__2 ;
    input window_24__1 ;
    input window_24__0 ;
    input window_23__15 ;
    input window_23__14 ;
    input window_23__13 ;
    input window_23__12 ;
    input window_23__11 ;
    input window_23__10 ;
    input window_23__9 ;
    input window_23__8 ;
    input window_23__7 ;
    input window_23__6 ;
    input window_23__5 ;
    input window_23__4 ;
    input window_23__3 ;
    input window_23__2 ;
    input window_23__1 ;
    input window_23__0 ;
    input window_22__15 ;
    input window_22__14 ;
    input window_22__13 ;
    input window_22__12 ;
    input window_22__11 ;
    input window_22__10 ;
    input window_22__9 ;
    input window_22__8 ;
    input window_22__7 ;
    input window_22__6 ;
    input window_22__5 ;
    input window_22__4 ;
    input window_22__3 ;
    input window_22__2 ;
    input window_22__1 ;
    input window_22__0 ;
    input window_21__15 ;
    input window_21__14 ;
    input window_21__13 ;
    input window_21__12 ;
    input window_21__11 ;
    input window_21__10 ;
    input window_21__9 ;
    input window_21__8 ;
    input window_21__7 ;
    input window_21__6 ;
    input window_21__5 ;
    input window_21__4 ;
    input window_21__3 ;
    input window_21__2 ;
    input window_21__1 ;
    input window_21__0 ;
    input window_20__15 ;
    input window_20__14 ;
    input window_20__13 ;
    input window_20__12 ;
    input window_20__11 ;
    input window_20__10 ;
    input window_20__9 ;
    input window_20__8 ;
    input window_20__7 ;
    input window_20__6 ;
    input window_20__5 ;
    input window_20__4 ;
    input window_20__3 ;
    input window_20__2 ;
    input window_20__1 ;
    input window_20__0 ;
    input window_19__15 ;
    input window_19__14 ;
    input window_19__13 ;
    input window_19__12 ;
    input window_19__11 ;
    input window_19__10 ;
    input window_19__9 ;
    input window_19__8 ;
    input window_19__7 ;
    input window_19__6 ;
    input window_19__5 ;
    input window_19__4 ;
    input window_19__3 ;
    input window_19__2 ;
    input window_19__1 ;
    input window_19__0 ;
    input window_18__15 ;
    input window_18__14 ;
    input window_18__13 ;
    input window_18__12 ;
    input window_18__11 ;
    input window_18__10 ;
    input window_18__9 ;
    input window_18__8 ;
    input window_18__7 ;
    input window_18__6 ;
    input window_18__5 ;
    input window_18__4 ;
    input window_18__3 ;
    input window_18__2 ;
    input window_18__1 ;
    input window_18__0 ;
    input window_17__15 ;
    input window_17__14 ;
    input window_17__13 ;
    input window_17__12 ;
    input window_17__11 ;
    input window_17__10 ;
    input window_17__9 ;
    input window_17__8 ;
    input window_17__7 ;
    input window_17__6 ;
    input window_17__5 ;
    input window_17__4 ;
    input window_17__3 ;
    input window_17__2 ;
    input window_17__1 ;
    input window_17__0 ;
    input window_16__15 ;
    input window_16__14 ;
    input window_16__13 ;
    input window_16__12 ;
    input window_16__11 ;
    input window_16__10 ;
    input window_16__9 ;
    input window_16__8 ;
    input window_16__7 ;
    input window_16__6 ;
    input window_16__5 ;
    input window_16__4 ;
    input window_16__3 ;
    input window_16__2 ;
    input window_16__1 ;
    input window_16__0 ;
    input window_15__15 ;
    input window_15__14 ;
    input window_15__13 ;
    input window_15__12 ;
    input window_15__11 ;
    input window_15__10 ;
    input window_15__9 ;
    input window_15__8 ;
    input window_15__7 ;
    input window_15__6 ;
    input window_15__5 ;
    input window_15__4 ;
    input window_15__3 ;
    input window_15__2 ;
    input window_15__1 ;
    input window_15__0 ;
    input window_14__15 ;
    input window_14__14 ;
    input window_14__13 ;
    input window_14__12 ;
    input window_14__11 ;
    input window_14__10 ;
    input window_14__9 ;
    input window_14__8 ;
    input window_14__7 ;
    input window_14__6 ;
    input window_14__5 ;
    input window_14__4 ;
    input window_14__3 ;
    input window_14__2 ;
    input window_14__1 ;
    input window_14__0 ;
    input window_13__15 ;
    input window_13__14 ;
    input window_13__13 ;
    input window_13__12 ;
    input window_13__11 ;
    input window_13__10 ;
    input window_13__9 ;
    input window_13__8 ;
    input window_13__7 ;
    input window_13__6 ;
    input window_13__5 ;
    input window_13__4 ;
    input window_13__3 ;
    input window_13__2 ;
    input window_13__1 ;
    input window_13__0 ;
    input window_12__15 ;
    input window_12__14 ;
    input window_12__13 ;
    input window_12__12 ;
    input window_12__11 ;
    input window_12__10 ;
    input window_12__9 ;
    input window_12__8 ;
    input window_12__7 ;
    input window_12__6 ;
    input window_12__5 ;
    input window_12__4 ;
    input window_12__3 ;
    input window_12__2 ;
    input window_12__1 ;
    input window_12__0 ;
    input window_11__15 ;
    input window_11__14 ;
    input window_11__13 ;
    input window_11__12 ;
    input window_11__11 ;
    input window_11__10 ;
    input window_11__9 ;
    input window_11__8 ;
    input window_11__7 ;
    input window_11__6 ;
    input window_11__5 ;
    input window_11__4 ;
    input window_11__3 ;
    input window_11__2 ;
    input window_11__1 ;
    input window_11__0 ;
    input window_10__15 ;
    input window_10__14 ;
    input window_10__13 ;
    input window_10__12 ;
    input window_10__11 ;
    input window_10__10 ;
    input window_10__9 ;
    input window_10__8 ;
    input window_10__7 ;
    input window_10__6 ;
    input window_10__5 ;
    input window_10__4 ;
    input window_10__3 ;
    input window_10__2 ;
    input window_10__1 ;
    input window_10__0 ;
    input window_9__15 ;
    input window_9__14 ;
    input window_9__13 ;
    input window_9__12 ;
    input window_9__11 ;
    input window_9__10 ;
    input window_9__9 ;
    input window_9__8 ;
    input window_9__7 ;
    input window_9__6 ;
    input window_9__5 ;
    input window_9__4 ;
    input window_9__3 ;
    input window_9__2 ;
    input window_9__1 ;
    input window_9__0 ;
    input window_8__15 ;
    input window_8__14 ;
    input window_8__13 ;
    input window_8__12 ;
    input window_8__11 ;
    input window_8__10 ;
    input window_8__9 ;
    input window_8__8 ;
    input window_8__7 ;
    input window_8__6 ;
    input window_8__5 ;
    input window_8__4 ;
    input window_8__3 ;
    input window_8__2 ;
    input window_8__1 ;
    input window_8__0 ;
    input window_7__15 ;
    input window_7__14 ;
    input window_7__13 ;
    input window_7__12 ;
    input window_7__11 ;
    input window_7__10 ;
    input window_7__9 ;
    input window_7__8 ;
    input window_7__7 ;
    input window_7__6 ;
    input window_7__5 ;
    input window_7__4 ;
    input window_7__3 ;
    input window_7__2 ;
    input window_7__1 ;
    input window_7__0 ;
    input window_6__15 ;
    input window_6__14 ;
    input window_6__13 ;
    input window_6__12 ;
    input window_6__11 ;
    input window_6__10 ;
    input window_6__9 ;
    input window_6__8 ;
    input window_6__7 ;
    input window_6__6 ;
    input window_6__5 ;
    input window_6__4 ;
    input window_6__3 ;
    input window_6__2 ;
    input window_6__1 ;
    input window_6__0 ;
    input window_5__15 ;
    input window_5__14 ;
    input window_5__13 ;
    input window_5__12 ;
    input window_5__11 ;
    input window_5__10 ;
    input window_5__9 ;
    input window_5__8 ;
    input window_5__7 ;
    input window_5__6 ;
    input window_5__5 ;
    input window_5__4 ;
    input window_5__3 ;
    input window_5__2 ;
    input window_5__1 ;
    input window_5__0 ;
    input window_4__15 ;
    input window_4__14 ;
    input window_4__13 ;
    input window_4__12 ;
    input window_4__11 ;
    input window_4__10 ;
    input window_4__9 ;
    input window_4__8 ;
    input window_4__7 ;
    input window_4__6 ;
    input window_4__5 ;
    input window_4__4 ;
    input window_4__3 ;
    input window_4__2 ;
    input window_4__1 ;
    input window_4__0 ;
    input window_3__15 ;
    input window_3__14 ;
    input window_3__13 ;
    input window_3__12 ;
    input window_3__11 ;
    input window_3__10 ;
    input window_3__9 ;
    input window_3__8 ;
    input window_3__7 ;
    input window_3__6 ;
    input window_3__5 ;
    input window_3__4 ;
    input window_3__3 ;
    input window_3__2 ;
    input window_3__1 ;
    input window_3__0 ;
    input window_2__15 ;
    input window_2__14 ;
    input window_2__13 ;
    input window_2__12 ;
    input window_2__11 ;
    input window_2__10 ;
    input window_2__9 ;
    input window_2__8 ;
    input window_2__7 ;
    input window_2__6 ;
    input window_2__5 ;
    input window_2__4 ;
    input window_2__3 ;
    input window_2__2 ;
    input window_2__1 ;
    input window_2__0 ;
    input window_1__15 ;
    input window_1__14 ;
    input window_1__13 ;
    input window_1__12 ;
    input window_1__11 ;
    input window_1__10 ;
    input window_1__9 ;
    input window_1__8 ;
    input window_1__7 ;
    input window_1__6 ;
    input window_1__5 ;
    input window_1__4 ;
    input window_1__3 ;
    input window_1__2 ;
    input window_1__1 ;
    input window_1__0 ;
    input window_0__15 ;
    input window_0__14 ;
    input window_0__13 ;
    input window_0__12 ;
    input window_0__11 ;
    input window_0__10 ;
    input window_0__9 ;
    input window_0__8 ;
    input window_0__7 ;
    input window_0__6 ;
    input window_0__5 ;
    input window_0__4 ;
    input window_0__3 ;
    input window_0__2 ;
    input window_0__1 ;
    input window_0__0 ;
    inout outputs_24__15 ;
    inout outputs_24__14 ;
    inout outputs_24__13 ;
    inout outputs_24__12 ;
    inout outputs_24__11 ;
    inout outputs_24__10 ;
    inout outputs_24__9 ;
    inout outputs_24__8 ;
    inout outputs_24__7 ;
    inout outputs_24__6 ;
    inout outputs_24__5 ;
    inout outputs_24__4 ;
    inout outputs_24__3 ;
    inout outputs_24__2 ;
    inout outputs_24__1 ;
    inout outputs_24__0 ;
    inout outputs_23__15 ;
    inout outputs_23__14 ;
    inout outputs_23__13 ;
    inout outputs_23__12 ;
    inout outputs_23__11 ;
    inout outputs_23__10 ;
    inout outputs_23__9 ;
    inout outputs_23__8 ;
    inout outputs_23__7 ;
    inout outputs_23__6 ;
    inout outputs_23__5 ;
    inout outputs_23__4 ;
    inout outputs_23__3 ;
    inout outputs_23__2 ;
    inout outputs_23__1 ;
    inout outputs_23__0 ;
    inout outputs_22__15 ;
    inout outputs_22__14 ;
    inout outputs_22__13 ;
    inout outputs_22__12 ;
    inout outputs_22__11 ;
    inout outputs_22__10 ;
    inout outputs_22__9 ;
    inout outputs_22__8 ;
    inout outputs_22__7 ;
    inout outputs_22__6 ;
    inout outputs_22__5 ;
    inout outputs_22__4 ;
    inout outputs_22__3 ;
    inout outputs_22__2 ;
    inout outputs_22__1 ;
    inout outputs_22__0 ;
    inout outputs_21__15 ;
    inout outputs_21__14 ;
    inout outputs_21__13 ;
    inout outputs_21__12 ;
    inout outputs_21__11 ;
    inout outputs_21__10 ;
    inout outputs_21__9 ;
    inout outputs_21__8 ;
    inout outputs_21__7 ;
    inout outputs_21__6 ;
    inout outputs_21__5 ;
    inout outputs_21__4 ;
    inout outputs_21__3 ;
    inout outputs_21__2 ;
    inout outputs_21__1 ;
    inout outputs_21__0 ;
    inout outputs_20__15 ;
    inout outputs_20__14 ;
    inout outputs_20__13 ;
    inout outputs_20__12 ;
    inout outputs_20__11 ;
    inout outputs_20__10 ;
    inout outputs_20__9 ;
    inout outputs_20__8 ;
    inout outputs_20__7 ;
    inout outputs_20__6 ;
    inout outputs_20__5 ;
    inout outputs_20__4 ;
    inout outputs_20__3 ;
    inout outputs_20__2 ;
    inout outputs_20__1 ;
    inout outputs_20__0 ;
    inout outputs_19__15 ;
    inout outputs_19__14 ;
    inout outputs_19__13 ;
    inout outputs_19__12 ;
    inout outputs_19__11 ;
    inout outputs_19__10 ;
    inout outputs_19__9 ;
    inout outputs_19__8 ;
    inout outputs_19__7 ;
    inout outputs_19__6 ;
    inout outputs_19__5 ;
    inout outputs_19__4 ;
    inout outputs_19__3 ;
    inout outputs_19__2 ;
    inout outputs_19__1 ;
    inout outputs_19__0 ;
    inout outputs_18__15 ;
    inout outputs_18__14 ;
    inout outputs_18__13 ;
    inout outputs_18__12 ;
    inout outputs_18__11 ;
    inout outputs_18__10 ;
    inout outputs_18__9 ;
    inout outputs_18__8 ;
    inout outputs_18__7 ;
    inout outputs_18__6 ;
    inout outputs_18__5 ;
    inout outputs_18__4 ;
    inout outputs_18__3 ;
    inout outputs_18__2 ;
    inout outputs_18__1 ;
    inout outputs_18__0 ;
    inout outputs_17__15 ;
    inout outputs_17__14 ;
    inout outputs_17__13 ;
    inout outputs_17__12 ;
    inout outputs_17__11 ;
    inout outputs_17__10 ;
    inout outputs_17__9 ;
    inout outputs_17__8 ;
    inout outputs_17__7 ;
    inout outputs_17__6 ;
    inout outputs_17__5 ;
    inout outputs_17__4 ;
    inout outputs_17__3 ;
    inout outputs_17__2 ;
    inout outputs_17__1 ;
    inout outputs_17__0 ;
    inout outputs_16__15 ;
    inout outputs_16__14 ;
    inout outputs_16__13 ;
    inout outputs_16__12 ;
    inout outputs_16__11 ;
    inout outputs_16__10 ;
    inout outputs_16__9 ;
    inout outputs_16__8 ;
    inout outputs_16__7 ;
    inout outputs_16__6 ;
    inout outputs_16__5 ;
    inout outputs_16__4 ;
    inout outputs_16__3 ;
    inout outputs_16__2 ;
    inout outputs_16__1 ;
    inout outputs_16__0 ;
    inout outputs_15__15 ;
    inout outputs_15__14 ;
    inout outputs_15__13 ;
    inout outputs_15__12 ;
    inout outputs_15__11 ;
    inout outputs_15__10 ;
    inout outputs_15__9 ;
    inout outputs_15__8 ;
    inout outputs_15__7 ;
    inout outputs_15__6 ;
    inout outputs_15__5 ;
    inout outputs_15__4 ;
    inout outputs_15__3 ;
    inout outputs_15__2 ;
    inout outputs_15__1 ;
    inout outputs_15__0 ;
    inout outputs_14__15 ;
    inout outputs_14__14 ;
    inout outputs_14__13 ;
    inout outputs_14__12 ;
    inout outputs_14__11 ;
    inout outputs_14__10 ;
    inout outputs_14__9 ;
    inout outputs_14__8 ;
    inout outputs_14__7 ;
    inout outputs_14__6 ;
    inout outputs_14__5 ;
    inout outputs_14__4 ;
    inout outputs_14__3 ;
    inout outputs_14__2 ;
    inout outputs_14__1 ;
    inout outputs_14__0 ;
    inout outputs_13__15 ;
    inout outputs_13__14 ;
    inout outputs_13__13 ;
    inout outputs_13__12 ;
    inout outputs_13__11 ;
    inout outputs_13__10 ;
    inout outputs_13__9 ;
    inout outputs_13__8 ;
    inout outputs_13__7 ;
    inout outputs_13__6 ;
    inout outputs_13__5 ;
    inout outputs_13__4 ;
    inout outputs_13__3 ;
    inout outputs_13__2 ;
    inout outputs_13__1 ;
    inout outputs_13__0 ;
    inout outputs_12__15 ;
    inout outputs_12__14 ;
    inout outputs_12__13 ;
    inout outputs_12__12 ;
    inout outputs_12__11 ;
    inout outputs_12__10 ;
    inout outputs_12__9 ;
    inout outputs_12__8 ;
    inout outputs_12__7 ;
    inout outputs_12__6 ;
    inout outputs_12__5 ;
    inout outputs_12__4 ;
    inout outputs_12__3 ;
    inout outputs_12__2 ;
    inout outputs_12__1 ;
    inout outputs_12__0 ;
    inout outputs_11__15 ;
    inout outputs_11__14 ;
    inout outputs_11__13 ;
    inout outputs_11__12 ;
    inout outputs_11__11 ;
    inout outputs_11__10 ;
    inout outputs_11__9 ;
    inout outputs_11__8 ;
    inout outputs_11__7 ;
    inout outputs_11__6 ;
    inout outputs_11__5 ;
    inout outputs_11__4 ;
    inout outputs_11__3 ;
    inout outputs_11__2 ;
    inout outputs_11__1 ;
    inout outputs_11__0 ;
    inout outputs_10__15 ;
    inout outputs_10__14 ;
    inout outputs_10__13 ;
    inout outputs_10__12 ;
    inout outputs_10__11 ;
    inout outputs_10__10 ;
    inout outputs_10__9 ;
    inout outputs_10__8 ;
    inout outputs_10__7 ;
    inout outputs_10__6 ;
    inout outputs_10__5 ;
    inout outputs_10__4 ;
    inout outputs_10__3 ;
    inout outputs_10__2 ;
    inout outputs_10__1 ;
    inout outputs_10__0 ;
    inout outputs_9__15 ;
    inout outputs_9__14 ;
    inout outputs_9__13 ;
    inout outputs_9__12 ;
    inout outputs_9__11 ;
    inout outputs_9__10 ;
    inout outputs_9__9 ;
    inout outputs_9__8 ;
    inout outputs_9__7 ;
    inout outputs_9__6 ;
    inout outputs_9__5 ;
    inout outputs_9__4 ;
    inout outputs_9__3 ;
    inout outputs_9__2 ;
    inout outputs_9__1 ;
    inout outputs_9__0 ;
    inout outputs_8__15 ;
    inout outputs_8__14 ;
    inout outputs_8__13 ;
    inout outputs_8__12 ;
    inout outputs_8__11 ;
    inout outputs_8__10 ;
    inout outputs_8__9 ;
    inout outputs_8__8 ;
    inout outputs_8__7 ;
    inout outputs_8__6 ;
    inout outputs_8__5 ;
    inout outputs_8__4 ;
    inout outputs_8__3 ;
    inout outputs_8__2 ;
    inout outputs_8__1 ;
    inout outputs_8__0 ;
    inout outputs_7__15 ;
    inout outputs_7__14 ;
    inout outputs_7__13 ;
    inout outputs_7__12 ;
    inout outputs_7__11 ;
    inout outputs_7__10 ;
    inout outputs_7__9 ;
    inout outputs_7__8 ;
    inout outputs_7__7 ;
    inout outputs_7__6 ;
    inout outputs_7__5 ;
    inout outputs_7__4 ;
    inout outputs_7__3 ;
    inout outputs_7__2 ;
    inout outputs_7__1 ;
    inout outputs_7__0 ;
    inout outputs_6__15 ;
    inout outputs_6__14 ;
    inout outputs_6__13 ;
    inout outputs_6__12 ;
    inout outputs_6__11 ;
    inout outputs_6__10 ;
    inout outputs_6__9 ;
    inout outputs_6__8 ;
    inout outputs_6__7 ;
    inout outputs_6__6 ;
    inout outputs_6__5 ;
    inout outputs_6__4 ;
    inout outputs_6__3 ;
    inout outputs_6__2 ;
    inout outputs_6__1 ;
    inout outputs_6__0 ;
    inout outputs_5__15 ;
    inout outputs_5__14 ;
    inout outputs_5__13 ;
    inout outputs_5__12 ;
    inout outputs_5__11 ;
    inout outputs_5__10 ;
    inout outputs_5__9 ;
    inout outputs_5__8 ;
    inout outputs_5__7 ;
    inout outputs_5__6 ;
    inout outputs_5__5 ;
    inout outputs_5__4 ;
    inout outputs_5__3 ;
    inout outputs_5__2 ;
    inout outputs_5__1 ;
    inout outputs_5__0 ;
    inout outputs_4__15 ;
    inout outputs_4__14 ;
    inout outputs_4__13 ;
    inout outputs_4__12 ;
    inout outputs_4__11 ;
    inout outputs_4__10 ;
    inout outputs_4__9 ;
    inout outputs_4__8 ;
    inout outputs_4__7 ;
    inout outputs_4__6 ;
    inout outputs_4__5 ;
    inout outputs_4__4 ;
    inout outputs_4__3 ;
    inout outputs_4__2 ;
    inout outputs_4__1 ;
    inout outputs_4__0 ;
    inout outputs_3__15 ;
    inout outputs_3__14 ;
    inout outputs_3__13 ;
    inout outputs_3__12 ;
    inout outputs_3__11 ;
    inout outputs_3__10 ;
    inout outputs_3__9 ;
    inout outputs_3__8 ;
    inout outputs_3__7 ;
    inout outputs_3__6 ;
    inout outputs_3__5 ;
    inout outputs_3__4 ;
    inout outputs_3__3 ;
    inout outputs_3__2 ;
    inout outputs_3__1 ;
    inout outputs_3__0 ;
    inout outputs_2__15 ;
    inout outputs_2__14 ;
    inout outputs_2__13 ;
    inout outputs_2__12 ;
    inout outputs_2__11 ;
    inout outputs_2__10 ;
    inout outputs_2__9 ;
    inout outputs_2__8 ;
    inout outputs_2__7 ;
    inout outputs_2__6 ;
    inout outputs_2__5 ;
    inout outputs_2__4 ;
    inout outputs_2__3 ;
    inout outputs_2__2 ;
    inout outputs_2__1 ;
    inout outputs_2__0 ;
    inout outputs_1__15 ;
    inout outputs_1__14 ;
    inout outputs_1__13 ;
    inout outputs_1__12 ;
    inout outputs_1__11 ;
    inout outputs_1__10 ;
    inout outputs_1__9 ;
    inout outputs_1__8 ;
    inout outputs_1__7 ;
    inout outputs_1__6 ;
    inout outputs_1__5 ;
    inout outputs_1__4 ;
    inout outputs_1__3 ;
    inout outputs_1__2 ;
    inout outputs_1__1 ;
    inout outputs_1__0 ;
    inout outputs_0__15 ;
    inout outputs_0__14 ;
    inout outputs_0__13 ;
    inout outputs_0__12 ;
    inout outputs_0__11 ;
    inout outputs_0__10 ;
    inout outputs_0__9 ;
    inout outputs_0__8 ;
    inout outputs_0__7 ;
    inout outputs_0__6 ;
    inout outputs_0__5 ;
    inout outputs_0__4 ;
    inout outputs_0__3 ;
    inout outputs_0__2 ;
    inout outputs_0__1 ;
    inout outputs_0__0 ;
    input clk ;
    input start ;
    input rst ;
    inout done ;
    inout working ;

    wire gen_24_cmp_pBs_30, gen_24_cmp_pBs_29, gen_24_cmp_pBs_28, 
         gen_24_cmp_pBs_27, gen_24_cmp_pBs_26, gen_24_cmp_pBs_25, 
         gen_24_cmp_pBs_24, gen_24_cmp_pBs_23, gen_24_cmp_pMux_30, 
         gen_24_cmp_pMux_29, gen_24_cmp_pMux_28, gen_24_cmp_pMux_27, 
         gen_24_cmp_pMux_26, gen_24_cmp_pMux_25, gen_24_cmp_pMux_24, 
         gen_24_cmp_pMux_23, gen_24_cmp_pMux_22, gen_24_cmp_pMux_21, 
         gen_24_cmp_pMux_20, gen_24_cmp_pMux_19, gen_24_cmp_pMux_18, 
         gen_24_cmp_pMux_17, gen_24_cmp_pMux_16, gen_24_cmp_pMux_15, 
         gen_24_cmp_pMux_14, gen_24_cmp_pMux_13, gen_24_cmp_pMux_12, 
         gen_24_cmp_pMux_11, gen_24_cmp_pMux_10, gen_24_cmp_pMux_9, 
         gen_24_cmp_pMux_8, gen_24_cmp_pMux_7, gen_24_cmp_pMux_6, 
         gen_24_cmp_pMux_5, gen_24_cmp_pMux_4, gen_24_cmp_pMux_3, 
         gen_24_cmp_pMux_2, gen_24_cmp_pMux_1, gen_24_cmp_pMux_0, 
         gen_24_cmp_pReg_30, gen_24_cmp_pReg_29, gen_24_cmp_pReg_28, 
         gen_24_cmp_pReg_27, gen_24_cmp_pReg_26, gen_24_cmp_pReg_25, 
         gen_24_cmp_pReg_24, gen_24_cmp_pReg_23, gen_24_cmp_pReg_22, 
         gen_24_cmp_pReg_21, gen_24_cmp_pReg_20, gen_24_cmp_pReg_19, 
         gen_24_cmp_pReg_18, gen_24_cmp_pReg_17, gen_24_cmp_pReg_16, 
         gen_24_cmp_pReg_15, gen_24_cmp_pReg_14, gen_24_cmp_pReg_13, 
         gen_24_cmp_pReg_12, gen_24_cmp_pReg_11, gen_24_cmp_pReg_10, 
         gen_24_cmp_pReg_9, gen_24_cmp_pReg_8, gen_24_cmp_pReg_7, 
         gen_24_cmp_pReg_6, gen_24_cmp_pReg_5, gen_24_cmp_pReg_4, 
         gen_24_cmp_pReg_3, gen_24_cmp_pReg_2, gen_24_cmp_pReg_1, 
         gen_24_cmp_pReg_0, gen_24_cmp_BSCmp_op2_0, gen_24_cmp_BSCmp_carryIn, 
         gen_23_cmp_pBs_30, gen_23_cmp_pBs_29, gen_23_cmp_pBs_28, 
         gen_23_cmp_pBs_27, gen_23_cmp_pBs_26, gen_23_cmp_pBs_25, 
         gen_23_cmp_pBs_24, gen_23_cmp_pBs_23, gen_23_cmp_pMux_30, 
         gen_23_cmp_pMux_29, gen_23_cmp_pMux_28, gen_23_cmp_pMux_27, 
         gen_23_cmp_pMux_26, gen_23_cmp_pMux_25, gen_23_cmp_pMux_24, 
         gen_23_cmp_pMux_23, gen_23_cmp_pMux_22, gen_23_cmp_pMux_21, 
         gen_23_cmp_pMux_20, gen_23_cmp_pMux_19, gen_23_cmp_pMux_18, 
         gen_23_cmp_pMux_17, gen_23_cmp_pMux_16, gen_23_cmp_pMux_15, 
         gen_23_cmp_pMux_14, gen_23_cmp_pMux_13, gen_23_cmp_pMux_12, 
         gen_23_cmp_pMux_11, gen_23_cmp_pMux_10, gen_23_cmp_pMux_9, 
         gen_23_cmp_pMux_8, gen_23_cmp_pMux_7, gen_23_cmp_pMux_6, 
         gen_23_cmp_pMux_5, gen_23_cmp_pMux_4, gen_23_cmp_pMux_3, 
         gen_23_cmp_pMux_2, gen_23_cmp_pMux_1, gen_23_cmp_pMux_0, 
         gen_23_cmp_pReg_30, gen_23_cmp_pReg_29, gen_23_cmp_pReg_28, 
         gen_23_cmp_pReg_27, gen_23_cmp_pReg_26, gen_23_cmp_pReg_25, 
         gen_23_cmp_pReg_24, gen_23_cmp_pReg_23, gen_23_cmp_pReg_22, 
         gen_23_cmp_pReg_21, gen_23_cmp_pReg_20, gen_23_cmp_pReg_19, 
         gen_23_cmp_pReg_18, gen_23_cmp_pReg_17, gen_23_cmp_pReg_16, 
         gen_23_cmp_pReg_15, gen_23_cmp_pReg_14, gen_23_cmp_pReg_13, 
         gen_23_cmp_pReg_12, gen_23_cmp_pReg_11, gen_23_cmp_pReg_10, 
         gen_23_cmp_pReg_9, gen_23_cmp_pReg_8, gen_23_cmp_pReg_7, 
         gen_23_cmp_pReg_6, gen_23_cmp_pReg_5, gen_23_cmp_pReg_4, 
         gen_23_cmp_pReg_3, gen_23_cmp_pReg_2, gen_23_cmp_pReg_1, 
         gen_23_cmp_pReg_0, gen_23_cmp_BSCmp_op2_0, gen_23_cmp_BSCmp_carryIn, 
         gen_22_cmp_pBs_30, gen_22_cmp_pBs_29, gen_22_cmp_pBs_28, 
         gen_22_cmp_pBs_27, gen_22_cmp_pBs_26, gen_22_cmp_pBs_25, 
         gen_22_cmp_pBs_24, gen_22_cmp_pBs_23, gen_22_cmp_pMux_30, 
         gen_22_cmp_pMux_29, gen_22_cmp_pMux_28, gen_22_cmp_pMux_27, 
         gen_22_cmp_pMux_26, gen_22_cmp_pMux_25, gen_22_cmp_pMux_24, 
         gen_22_cmp_pMux_23, gen_22_cmp_pMux_22, gen_22_cmp_pMux_21, 
         gen_22_cmp_pMux_20, gen_22_cmp_pMux_19, gen_22_cmp_pMux_18, 
         gen_22_cmp_pMux_17, gen_22_cmp_pMux_16, gen_22_cmp_pMux_15, 
         gen_22_cmp_pMux_14, gen_22_cmp_pMux_13, gen_22_cmp_pMux_12, 
         gen_22_cmp_pMux_11, gen_22_cmp_pMux_10, gen_22_cmp_pMux_9, 
         gen_22_cmp_pMux_8, gen_22_cmp_pMux_7, gen_22_cmp_pMux_6, 
         gen_22_cmp_pMux_5, gen_22_cmp_pMux_4, gen_22_cmp_pMux_3, 
         gen_22_cmp_pMux_2, gen_22_cmp_pMux_1, gen_22_cmp_pMux_0, 
         gen_22_cmp_pReg_30, gen_22_cmp_pReg_29, gen_22_cmp_pReg_28, 
         gen_22_cmp_pReg_27, gen_22_cmp_pReg_26, gen_22_cmp_pReg_25, 
         gen_22_cmp_pReg_24, gen_22_cmp_pReg_23, gen_22_cmp_pReg_22, 
         gen_22_cmp_pReg_21, gen_22_cmp_pReg_20, gen_22_cmp_pReg_19, 
         gen_22_cmp_pReg_18, gen_22_cmp_pReg_17, gen_22_cmp_pReg_16, 
         gen_22_cmp_pReg_15, gen_22_cmp_pReg_14, gen_22_cmp_pReg_13, 
         gen_22_cmp_pReg_12, gen_22_cmp_pReg_11, gen_22_cmp_pReg_10, 
         gen_22_cmp_pReg_9, gen_22_cmp_pReg_8, gen_22_cmp_pReg_7, 
         gen_22_cmp_pReg_6, gen_22_cmp_pReg_5, gen_22_cmp_pReg_4, 
         gen_22_cmp_pReg_3, gen_22_cmp_pReg_2, gen_22_cmp_pReg_1, 
         gen_22_cmp_pReg_0, gen_22_cmp_BSCmp_op2_0, gen_22_cmp_BSCmp_carryIn, 
         gen_21_cmp_pBs_30, gen_21_cmp_pBs_29, gen_21_cmp_pBs_28, 
         gen_21_cmp_pBs_27, gen_21_cmp_pBs_26, gen_21_cmp_pBs_25, 
         gen_21_cmp_pBs_24, gen_21_cmp_pBs_23, gen_21_cmp_pMux_30, 
         gen_21_cmp_pMux_29, gen_21_cmp_pMux_28, gen_21_cmp_pMux_27, 
         gen_21_cmp_pMux_26, gen_21_cmp_pMux_25, gen_21_cmp_pMux_24, 
         gen_21_cmp_pMux_23, gen_21_cmp_pMux_22, gen_21_cmp_pMux_21, 
         gen_21_cmp_pMux_20, gen_21_cmp_pMux_19, gen_21_cmp_pMux_18, 
         gen_21_cmp_pMux_17, gen_21_cmp_pMux_16, gen_21_cmp_pMux_15, 
         gen_21_cmp_pMux_14, gen_21_cmp_pMux_13, gen_21_cmp_pMux_12, 
         gen_21_cmp_pMux_11, gen_21_cmp_pMux_10, gen_21_cmp_pMux_9, 
         gen_21_cmp_pMux_8, gen_21_cmp_pMux_7, gen_21_cmp_pMux_6, 
         gen_21_cmp_pMux_5, gen_21_cmp_pMux_4, gen_21_cmp_pMux_3, 
         gen_21_cmp_pMux_2, gen_21_cmp_pMux_1, gen_21_cmp_pMux_0, 
         gen_21_cmp_pReg_30, gen_21_cmp_pReg_29, gen_21_cmp_pReg_28, 
         gen_21_cmp_pReg_27, gen_21_cmp_pReg_26, gen_21_cmp_pReg_25, 
         gen_21_cmp_pReg_24, gen_21_cmp_pReg_23, gen_21_cmp_pReg_22, 
         gen_21_cmp_pReg_21, gen_21_cmp_pReg_20, gen_21_cmp_pReg_19, 
         gen_21_cmp_pReg_18, gen_21_cmp_pReg_17, gen_21_cmp_pReg_16, 
         gen_21_cmp_pReg_15, gen_21_cmp_pReg_14, gen_21_cmp_pReg_13, 
         gen_21_cmp_pReg_12, gen_21_cmp_pReg_11, gen_21_cmp_pReg_10, 
         gen_21_cmp_pReg_9, gen_21_cmp_pReg_8, gen_21_cmp_pReg_7, 
         gen_21_cmp_pReg_6, gen_21_cmp_pReg_5, gen_21_cmp_pReg_4, 
         gen_21_cmp_pReg_3, gen_21_cmp_pReg_2, gen_21_cmp_pReg_1, 
         gen_21_cmp_pReg_0, gen_21_cmp_BSCmp_op2_0, gen_21_cmp_BSCmp_carryIn, 
         gen_20_cmp_pBs_30, gen_20_cmp_pBs_29, gen_20_cmp_pBs_28, 
         gen_20_cmp_pBs_27, gen_20_cmp_pBs_26, gen_20_cmp_pBs_25, 
         gen_20_cmp_pBs_24, gen_20_cmp_pBs_23, gen_20_cmp_pMux_30, 
         gen_20_cmp_pMux_29, gen_20_cmp_pMux_28, gen_20_cmp_pMux_27, 
         gen_20_cmp_pMux_26, gen_20_cmp_pMux_25, gen_20_cmp_pMux_24, 
         gen_20_cmp_pMux_23, gen_20_cmp_pMux_22, gen_20_cmp_pMux_21, 
         gen_20_cmp_pMux_20, gen_20_cmp_pMux_19, gen_20_cmp_pMux_18, 
         gen_20_cmp_pMux_17, gen_20_cmp_pMux_16, gen_20_cmp_pMux_15, 
         gen_20_cmp_pMux_14, gen_20_cmp_pMux_13, gen_20_cmp_pMux_12, 
         gen_20_cmp_pMux_11, gen_20_cmp_pMux_10, gen_20_cmp_pMux_9, 
         gen_20_cmp_pMux_8, gen_20_cmp_pMux_7, gen_20_cmp_pMux_6, 
         gen_20_cmp_pMux_5, gen_20_cmp_pMux_4, gen_20_cmp_pMux_3, 
         gen_20_cmp_pMux_2, gen_20_cmp_pMux_1, gen_20_cmp_pMux_0, 
         gen_20_cmp_pReg_30, gen_20_cmp_pReg_29, gen_20_cmp_pReg_28, 
         gen_20_cmp_pReg_27, gen_20_cmp_pReg_26, gen_20_cmp_pReg_25, 
         gen_20_cmp_pReg_24, gen_20_cmp_pReg_23, gen_20_cmp_pReg_22, 
         gen_20_cmp_pReg_21, gen_20_cmp_pReg_20, gen_20_cmp_pReg_19, 
         gen_20_cmp_pReg_18, gen_20_cmp_pReg_17, gen_20_cmp_pReg_16, 
         gen_20_cmp_pReg_15, gen_20_cmp_pReg_14, gen_20_cmp_pReg_13, 
         gen_20_cmp_pReg_12, gen_20_cmp_pReg_11, gen_20_cmp_pReg_10, 
         gen_20_cmp_pReg_9, gen_20_cmp_pReg_8, gen_20_cmp_pReg_7, 
         gen_20_cmp_pReg_6, gen_20_cmp_pReg_5, gen_20_cmp_pReg_4, 
         gen_20_cmp_pReg_3, gen_20_cmp_pReg_2, gen_20_cmp_pReg_1, 
         gen_20_cmp_pReg_0, gen_20_cmp_BSCmp_op2_0, gen_20_cmp_BSCmp_carryIn, 
         gen_19_cmp_pBs_30, gen_19_cmp_pBs_29, gen_19_cmp_pBs_28, 
         gen_19_cmp_pBs_27, gen_19_cmp_pBs_26, gen_19_cmp_pBs_25, 
         gen_19_cmp_pBs_24, gen_19_cmp_pBs_23, gen_19_cmp_pMux_30, 
         gen_19_cmp_pMux_29, gen_19_cmp_pMux_28, gen_19_cmp_pMux_27, 
         gen_19_cmp_pMux_26, gen_19_cmp_pMux_25, gen_19_cmp_pMux_24, 
         gen_19_cmp_pMux_23, gen_19_cmp_pMux_22, gen_19_cmp_pMux_21, 
         gen_19_cmp_pMux_20, gen_19_cmp_pMux_19, gen_19_cmp_pMux_18, 
         gen_19_cmp_pMux_17, gen_19_cmp_pMux_16, gen_19_cmp_pMux_15, 
         gen_19_cmp_pMux_14, gen_19_cmp_pMux_13, gen_19_cmp_pMux_12, 
         gen_19_cmp_pMux_11, gen_19_cmp_pMux_10, gen_19_cmp_pMux_9, 
         gen_19_cmp_pMux_8, gen_19_cmp_pMux_7, gen_19_cmp_pMux_6, 
         gen_19_cmp_pMux_5, gen_19_cmp_pMux_4, gen_19_cmp_pMux_3, 
         gen_19_cmp_pMux_2, gen_19_cmp_pMux_1, gen_19_cmp_pMux_0, 
         gen_19_cmp_pReg_30, gen_19_cmp_pReg_29, gen_19_cmp_pReg_28, 
         gen_19_cmp_pReg_27, gen_19_cmp_pReg_26, gen_19_cmp_pReg_25, 
         gen_19_cmp_pReg_24, gen_19_cmp_pReg_23, gen_19_cmp_pReg_22, 
         gen_19_cmp_pReg_21, gen_19_cmp_pReg_20, gen_19_cmp_pReg_19, 
         gen_19_cmp_pReg_18, gen_19_cmp_pReg_17, gen_19_cmp_pReg_16, 
         gen_19_cmp_pReg_15, gen_19_cmp_pReg_14, gen_19_cmp_pReg_13, 
         gen_19_cmp_pReg_12, gen_19_cmp_pReg_11, gen_19_cmp_pReg_10, 
         gen_19_cmp_pReg_9, gen_19_cmp_pReg_8, gen_19_cmp_pReg_7, 
         gen_19_cmp_pReg_6, gen_19_cmp_pReg_5, gen_19_cmp_pReg_4, 
         gen_19_cmp_pReg_3, gen_19_cmp_pReg_2, gen_19_cmp_pReg_1, 
         gen_19_cmp_pReg_0, gen_19_cmp_BSCmp_op2_0, gen_19_cmp_BSCmp_carryIn, 
         gen_18_cmp_pBs_30, gen_18_cmp_pBs_29, gen_18_cmp_pBs_28, 
         gen_18_cmp_pBs_27, gen_18_cmp_pBs_26, gen_18_cmp_pBs_25, 
         gen_18_cmp_pBs_24, gen_18_cmp_pBs_23, gen_18_cmp_pMux_30, 
         gen_18_cmp_pMux_29, gen_18_cmp_pMux_28, gen_18_cmp_pMux_27, 
         gen_18_cmp_pMux_26, gen_18_cmp_pMux_25, gen_18_cmp_pMux_24, 
         gen_18_cmp_pMux_23, gen_18_cmp_pMux_22, gen_18_cmp_pMux_21, 
         gen_18_cmp_pMux_20, gen_18_cmp_pMux_19, gen_18_cmp_pMux_18, 
         gen_18_cmp_pMux_17, gen_18_cmp_pMux_16, gen_18_cmp_pMux_15, 
         gen_18_cmp_pMux_14, gen_18_cmp_pMux_13, gen_18_cmp_pMux_12, 
         gen_18_cmp_pMux_11, gen_18_cmp_pMux_10, gen_18_cmp_pMux_9, 
         gen_18_cmp_pMux_8, gen_18_cmp_pMux_7, gen_18_cmp_pMux_6, 
         gen_18_cmp_pMux_5, gen_18_cmp_pMux_4, gen_18_cmp_pMux_3, 
         gen_18_cmp_pMux_2, gen_18_cmp_pMux_1, gen_18_cmp_pMux_0, 
         gen_18_cmp_pReg_30, gen_18_cmp_pReg_29, gen_18_cmp_pReg_28, 
         gen_18_cmp_pReg_27, gen_18_cmp_pReg_26, gen_18_cmp_pReg_25, 
         gen_18_cmp_pReg_24, gen_18_cmp_pReg_23, gen_18_cmp_pReg_22, 
         gen_18_cmp_pReg_21, gen_18_cmp_pReg_20, gen_18_cmp_pReg_19, 
         gen_18_cmp_pReg_18, gen_18_cmp_pReg_17, gen_18_cmp_pReg_16, 
         gen_18_cmp_pReg_15, gen_18_cmp_pReg_14, gen_18_cmp_pReg_13, 
         gen_18_cmp_pReg_12, gen_18_cmp_pReg_11, gen_18_cmp_pReg_10, 
         gen_18_cmp_pReg_9, gen_18_cmp_pReg_8, gen_18_cmp_pReg_7, 
         gen_18_cmp_pReg_6, gen_18_cmp_pReg_5, gen_18_cmp_pReg_4, 
         gen_18_cmp_pReg_3, gen_18_cmp_pReg_2, gen_18_cmp_pReg_1, 
         gen_18_cmp_pReg_0, gen_18_cmp_BSCmp_op2_0, gen_18_cmp_BSCmp_carryIn, 
         gen_17_cmp_pBs_30, gen_17_cmp_pBs_29, gen_17_cmp_pBs_28, 
         gen_17_cmp_pBs_27, gen_17_cmp_pBs_26, gen_17_cmp_pBs_25, 
         gen_17_cmp_pBs_24, gen_17_cmp_pBs_23, gen_17_cmp_pMux_30, 
         gen_17_cmp_pMux_29, gen_17_cmp_pMux_28, gen_17_cmp_pMux_27, 
         gen_17_cmp_pMux_26, gen_17_cmp_pMux_25, gen_17_cmp_pMux_24, 
         gen_17_cmp_pMux_23, gen_17_cmp_pMux_22, gen_17_cmp_pMux_21, 
         gen_17_cmp_pMux_20, gen_17_cmp_pMux_19, gen_17_cmp_pMux_18, 
         gen_17_cmp_pMux_17, gen_17_cmp_pMux_16, gen_17_cmp_pMux_15, 
         gen_17_cmp_pMux_14, gen_17_cmp_pMux_13, gen_17_cmp_pMux_12, 
         gen_17_cmp_pMux_11, gen_17_cmp_pMux_10, gen_17_cmp_pMux_9, 
         gen_17_cmp_pMux_8, gen_17_cmp_pMux_7, gen_17_cmp_pMux_6, 
         gen_17_cmp_pMux_5, gen_17_cmp_pMux_4, gen_17_cmp_pMux_3, 
         gen_17_cmp_pMux_2, gen_17_cmp_pMux_1, gen_17_cmp_pMux_0, 
         gen_17_cmp_pReg_30, gen_17_cmp_pReg_29, gen_17_cmp_pReg_28, 
         gen_17_cmp_pReg_27, gen_17_cmp_pReg_26, gen_17_cmp_pReg_25, 
         gen_17_cmp_pReg_24, gen_17_cmp_pReg_23, gen_17_cmp_pReg_22, 
         gen_17_cmp_pReg_21, gen_17_cmp_pReg_20, gen_17_cmp_pReg_19, 
         gen_17_cmp_pReg_18, gen_17_cmp_pReg_17, gen_17_cmp_pReg_16, 
         gen_17_cmp_pReg_15, gen_17_cmp_pReg_14, gen_17_cmp_pReg_13, 
         gen_17_cmp_pReg_12, gen_17_cmp_pReg_11, gen_17_cmp_pReg_10, 
         gen_17_cmp_pReg_9, gen_17_cmp_pReg_8, gen_17_cmp_pReg_7, 
         gen_17_cmp_pReg_6, gen_17_cmp_pReg_5, gen_17_cmp_pReg_4, 
         gen_17_cmp_pReg_3, gen_17_cmp_pReg_2, gen_17_cmp_pReg_1, 
         gen_17_cmp_pReg_0, gen_17_cmp_BSCmp_op2_0, gen_17_cmp_BSCmp_carryIn, 
         gen_16_cmp_pBs_30, gen_16_cmp_pBs_29, gen_16_cmp_pBs_28, 
         gen_16_cmp_pBs_27, gen_16_cmp_pBs_26, gen_16_cmp_pBs_25, 
         gen_16_cmp_pBs_24, gen_16_cmp_pBs_23, gen_16_cmp_pMux_30, 
         gen_16_cmp_pMux_29, gen_16_cmp_pMux_28, gen_16_cmp_pMux_27, 
         gen_16_cmp_pMux_26, gen_16_cmp_pMux_25, gen_16_cmp_pMux_24, 
         gen_16_cmp_pMux_23, gen_16_cmp_pMux_22, gen_16_cmp_pMux_21, 
         gen_16_cmp_pMux_20, gen_16_cmp_pMux_19, gen_16_cmp_pMux_18, 
         gen_16_cmp_pMux_17, gen_16_cmp_pMux_16, gen_16_cmp_pMux_15, 
         gen_16_cmp_pMux_14, gen_16_cmp_pMux_13, gen_16_cmp_pMux_12, 
         gen_16_cmp_pMux_11, gen_16_cmp_pMux_10, gen_16_cmp_pMux_9, 
         gen_16_cmp_pMux_8, gen_16_cmp_pMux_7, gen_16_cmp_pMux_6, 
         gen_16_cmp_pMux_5, gen_16_cmp_pMux_4, gen_16_cmp_pMux_3, 
         gen_16_cmp_pMux_2, gen_16_cmp_pMux_1, gen_16_cmp_pMux_0, 
         gen_16_cmp_pReg_30, gen_16_cmp_pReg_29, gen_16_cmp_pReg_28, 
         gen_16_cmp_pReg_27, gen_16_cmp_pReg_26, gen_16_cmp_pReg_25, 
         gen_16_cmp_pReg_24, gen_16_cmp_pReg_23, gen_16_cmp_pReg_22, 
         gen_16_cmp_pReg_21, gen_16_cmp_pReg_20, gen_16_cmp_pReg_19, 
         gen_16_cmp_pReg_18, gen_16_cmp_pReg_17, gen_16_cmp_pReg_16, 
         gen_16_cmp_pReg_15, gen_16_cmp_pReg_14, gen_16_cmp_pReg_13, 
         gen_16_cmp_pReg_12, gen_16_cmp_pReg_11, gen_16_cmp_pReg_10, 
         gen_16_cmp_pReg_9, gen_16_cmp_pReg_8, gen_16_cmp_pReg_7, 
         gen_16_cmp_pReg_6, gen_16_cmp_pReg_5, gen_16_cmp_pReg_4, 
         gen_16_cmp_pReg_3, gen_16_cmp_pReg_2, gen_16_cmp_pReg_1, 
         gen_16_cmp_pReg_0, gen_16_cmp_BSCmp_op2_0, gen_16_cmp_BSCmp_carryIn, 
         gen_15_cmp_pBs_30, gen_15_cmp_pBs_29, gen_15_cmp_pBs_28, 
         gen_15_cmp_pBs_27, gen_15_cmp_pBs_26, gen_15_cmp_pBs_25, 
         gen_15_cmp_pBs_24, gen_15_cmp_pBs_23, gen_15_cmp_pMux_30, 
         gen_15_cmp_pMux_29, gen_15_cmp_pMux_28, gen_15_cmp_pMux_27, 
         gen_15_cmp_pMux_26, gen_15_cmp_pMux_25, gen_15_cmp_pMux_24, 
         gen_15_cmp_pMux_23, gen_15_cmp_pMux_22, gen_15_cmp_pMux_21, 
         gen_15_cmp_pMux_20, gen_15_cmp_pMux_19, gen_15_cmp_pMux_18, 
         gen_15_cmp_pMux_17, gen_15_cmp_pMux_16, gen_15_cmp_pMux_15, 
         gen_15_cmp_pMux_14, gen_15_cmp_pMux_13, gen_15_cmp_pMux_12, 
         gen_15_cmp_pMux_11, gen_15_cmp_pMux_10, gen_15_cmp_pMux_9, 
         gen_15_cmp_pMux_8, gen_15_cmp_pMux_7, gen_15_cmp_pMux_6, 
         gen_15_cmp_pMux_5, gen_15_cmp_pMux_4, gen_15_cmp_pMux_3, 
         gen_15_cmp_pMux_2, gen_15_cmp_pMux_1, gen_15_cmp_pMux_0, 
         gen_15_cmp_pReg_30, gen_15_cmp_pReg_29, gen_15_cmp_pReg_28, 
         gen_15_cmp_pReg_27, gen_15_cmp_pReg_26, gen_15_cmp_pReg_25, 
         gen_15_cmp_pReg_24, gen_15_cmp_pReg_23, gen_15_cmp_pReg_22, 
         gen_15_cmp_pReg_21, gen_15_cmp_pReg_20, gen_15_cmp_pReg_19, 
         gen_15_cmp_pReg_18, gen_15_cmp_pReg_17, gen_15_cmp_pReg_16, 
         gen_15_cmp_pReg_15, gen_15_cmp_pReg_14, gen_15_cmp_pReg_13, 
         gen_15_cmp_pReg_12, gen_15_cmp_pReg_11, gen_15_cmp_pReg_10, 
         gen_15_cmp_pReg_9, gen_15_cmp_pReg_8, gen_15_cmp_pReg_7, 
         gen_15_cmp_pReg_6, gen_15_cmp_pReg_5, gen_15_cmp_pReg_4, 
         gen_15_cmp_pReg_3, gen_15_cmp_pReg_2, gen_15_cmp_pReg_1, 
         gen_15_cmp_pReg_0, gen_15_cmp_BSCmp_op2_0, gen_15_cmp_BSCmp_carryIn, 
         gen_14_cmp_pBs_30, gen_14_cmp_pBs_29, gen_14_cmp_pBs_28, 
         gen_14_cmp_pBs_27, gen_14_cmp_pBs_26, gen_14_cmp_pBs_25, 
         gen_14_cmp_pBs_24, gen_14_cmp_pBs_23, gen_14_cmp_pMux_30, 
         gen_14_cmp_pMux_29, gen_14_cmp_pMux_28, gen_14_cmp_pMux_27, 
         gen_14_cmp_pMux_26, gen_14_cmp_pMux_25, gen_14_cmp_pMux_24, 
         gen_14_cmp_pMux_23, gen_14_cmp_pMux_22, gen_14_cmp_pMux_21, 
         gen_14_cmp_pMux_20, gen_14_cmp_pMux_19, gen_14_cmp_pMux_18, 
         gen_14_cmp_pMux_17, gen_14_cmp_pMux_16, gen_14_cmp_pMux_15, 
         gen_14_cmp_pMux_14, gen_14_cmp_pMux_13, gen_14_cmp_pMux_12, 
         gen_14_cmp_pMux_11, gen_14_cmp_pMux_10, gen_14_cmp_pMux_9, 
         gen_14_cmp_pMux_8, gen_14_cmp_pMux_7, gen_14_cmp_pMux_6, 
         gen_14_cmp_pMux_5, gen_14_cmp_pMux_4, gen_14_cmp_pMux_3, 
         gen_14_cmp_pMux_2, gen_14_cmp_pMux_1, gen_14_cmp_pMux_0, 
         gen_14_cmp_pReg_30, gen_14_cmp_pReg_29, gen_14_cmp_pReg_28, 
         gen_14_cmp_pReg_27, gen_14_cmp_pReg_26, gen_14_cmp_pReg_25, 
         gen_14_cmp_pReg_24, gen_14_cmp_pReg_23, gen_14_cmp_pReg_22, 
         gen_14_cmp_pReg_21, gen_14_cmp_pReg_20, gen_14_cmp_pReg_19, 
         gen_14_cmp_pReg_18, gen_14_cmp_pReg_17, gen_14_cmp_pReg_16, 
         gen_14_cmp_pReg_15, gen_14_cmp_pReg_14, gen_14_cmp_pReg_13, 
         gen_14_cmp_pReg_12, gen_14_cmp_pReg_11, gen_14_cmp_pReg_10, 
         gen_14_cmp_pReg_9, gen_14_cmp_pReg_8, gen_14_cmp_pReg_7, 
         gen_14_cmp_pReg_6, gen_14_cmp_pReg_5, gen_14_cmp_pReg_4, 
         gen_14_cmp_pReg_3, gen_14_cmp_pReg_2, gen_14_cmp_pReg_1, 
         gen_14_cmp_pReg_0, gen_14_cmp_BSCmp_op2_0, gen_14_cmp_BSCmp_carryIn, 
         gen_13_cmp_pBs_30, gen_13_cmp_pBs_29, gen_13_cmp_pBs_28, 
         gen_13_cmp_pBs_27, gen_13_cmp_pBs_26, gen_13_cmp_pBs_25, 
         gen_13_cmp_pBs_24, gen_13_cmp_pBs_23, gen_13_cmp_pMux_30, 
         gen_13_cmp_pMux_29, gen_13_cmp_pMux_28, gen_13_cmp_pMux_27, 
         gen_13_cmp_pMux_26, gen_13_cmp_pMux_25, gen_13_cmp_pMux_24, 
         gen_13_cmp_pMux_23, gen_13_cmp_pMux_22, gen_13_cmp_pMux_21, 
         gen_13_cmp_pMux_20, gen_13_cmp_pMux_19, gen_13_cmp_pMux_18, 
         gen_13_cmp_pMux_17, gen_13_cmp_pMux_16, gen_13_cmp_pMux_15, 
         gen_13_cmp_pMux_14, gen_13_cmp_pMux_13, gen_13_cmp_pMux_12, 
         gen_13_cmp_pMux_11, gen_13_cmp_pMux_10, gen_13_cmp_pMux_9, 
         gen_13_cmp_pMux_8, gen_13_cmp_pMux_7, gen_13_cmp_pMux_6, 
         gen_13_cmp_pMux_5, gen_13_cmp_pMux_4, gen_13_cmp_pMux_3, 
         gen_13_cmp_pMux_2, gen_13_cmp_pMux_1, gen_13_cmp_pMux_0, 
         gen_13_cmp_pReg_30, gen_13_cmp_pReg_29, gen_13_cmp_pReg_28, 
         gen_13_cmp_pReg_27, gen_13_cmp_pReg_26, gen_13_cmp_pReg_25, 
         gen_13_cmp_pReg_24, gen_13_cmp_pReg_23, gen_13_cmp_pReg_22, 
         gen_13_cmp_pReg_21, gen_13_cmp_pReg_20, gen_13_cmp_pReg_19, 
         gen_13_cmp_pReg_18, gen_13_cmp_pReg_17, gen_13_cmp_pReg_16, 
         gen_13_cmp_pReg_15, gen_13_cmp_pReg_14, gen_13_cmp_pReg_13, 
         gen_13_cmp_pReg_12, gen_13_cmp_pReg_11, gen_13_cmp_pReg_10, 
         gen_13_cmp_pReg_9, gen_13_cmp_pReg_8, gen_13_cmp_pReg_7, 
         gen_13_cmp_pReg_6, gen_13_cmp_pReg_5, gen_13_cmp_pReg_4, 
         gen_13_cmp_pReg_3, gen_13_cmp_pReg_2, gen_13_cmp_pReg_1, 
         gen_13_cmp_pReg_0, gen_13_cmp_BSCmp_op2_0, gen_13_cmp_BSCmp_carryIn, 
         gen_12_cmp_pBs_30, gen_12_cmp_pBs_29, gen_12_cmp_pBs_28, 
         gen_12_cmp_pBs_27, gen_12_cmp_pBs_26, gen_12_cmp_pBs_25, 
         gen_12_cmp_pBs_24, gen_12_cmp_pBs_23, gen_12_cmp_pMux_30, 
         gen_12_cmp_pMux_29, gen_12_cmp_pMux_28, gen_12_cmp_pMux_27, 
         gen_12_cmp_pMux_26, gen_12_cmp_pMux_25, gen_12_cmp_pMux_24, 
         gen_12_cmp_pMux_23, gen_12_cmp_pMux_22, gen_12_cmp_pMux_21, 
         gen_12_cmp_pMux_20, gen_12_cmp_pMux_19, gen_12_cmp_pMux_18, 
         gen_12_cmp_pMux_17, gen_12_cmp_pMux_16, gen_12_cmp_pMux_15, 
         gen_12_cmp_pMux_14, gen_12_cmp_pMux_13, gen_12_cmp_pMux_12, 
         gen_12_cmp_pMux_11, gen_12_cmp_pMux_10, gen_12_cmp_pMux_9, 
         gen_12_cmp_pMux_8, gen_12_cmp_pMux_7, gen_12_cmp_pMux_6, 
         gen_12_cmp_pMux_5, gen_12_cmp_pMux_4, gen_12_cmp_pMux_3, 
         gen_12_cmp_pMux_2, gen_12_cmp_pMux_1, gen_12_cmp_pMux_0, 
         gen_12_cmp_pReg_30, gen_12_cmp_pReg_29, gen_12_cmp_pReg_28, 
         gen_12_cmp_pReg_27, gen_12_cmp_pReg_26, gen_12_cmp_pReg_25, 
         gen_12_cmp_pReg_24, gen_12_cmp_pReg_23, gen_12_cmp_pReg_22, 
         gen_12_cmp_pReg_21, gen_12_cmp_pReg_20, gen_12_cmp_pReg_19, 
         gen_12_cmp_pReg_18, gen_12_cmp_pReg_17, gen_12_cmp_pReg_16, 
         gen_12_cmp_pReg_15, gen_12_cmp_pReg_14, gen_12_cmp_pReg_13, 
         gen_12_cmp_pReg_12, gen_12_cmp_pReg_11, gen_12_cmp_pReg_10, 
         gen_12_cmp_pReg_9, gen_12_cmp_pReg_8, gen_12_cmp_pReg_7, 
         gen_12_cmp_pReg_6, gen_12_cmp_pReg_5, gen_12_cmp_pReg_4, 
         gen_12_cmp_pReg_3, gen_12_cmp_pReg_2, gen_12_cmp_pReg_1, 
         gen_12_cmp_pReg_0, gen_12_cmp_BSCmp_op2_0, gen_12_cmp_BSCmp_carryIn, 
         gen_11_cmp_pBs_30, gen_11_cmp_pBs_29, gen_11_cmp_pBs_28, 
         gen_11_cmp_pBs_27, gen_11_cmp_pBs_26, gen_11_cmp_pBs_25, 
         gen_11_cmp_pBs_24, gen_11_cmp_pBs_23, gen_11_cmp_pMux_30, 
         gen_11_cmp_pMux_29, gen_11_cmp_pMux_28, gen_11_cmp_pMux_27, 
         gen_11_cmp_pMux_26, gen_11_cmp_pMux_25, gen_11_cmp_pMux_24, 
         gen_11_cmp_pMux_23, gen_11_cmp_pMux_22, gen_11_cmp_pMux_21, 
         gen_11_cmp_pMux_20, gen_11_cmp_pMux_19, gen_11_cmp_pMux_18, 
         gen_11_cmp_pMux_17, gen_11_cmp_pMux_16, gen_11_cmp_pMux_15, 
         gen_11_cmp_pMux_14, gen_11_cmp_pMux_13, gen_11_cmp_pMux_12, 
         gen_11_cmp_pMux_11, gen_11_cmp_pMux_10, gen_11_cmp_pMux_9, 
         gen_11_cmp_pMux_8, gen_11_cmp_pMux_7, gen_11_cmp_pMux_6, 
         gen_11_cmp_pMux_5, gen_11_cmp_pMux_4, gen_11_cmp_pMux_3, 
         gen_11_cmp_pMux_2, gen_11_cmp_pMux_1, gen_11_cmp_pMux_0, 
         gen_11_cmp_pReg_30, gen_11_cmp_pReg_29, gen_11_cmp_pReg_28, 
         gen_11_cmp_pReg_27, gen_11_cmp_pReg_26, gen_11_cmp_pReg_25, 
         gen_11_cmp_pReg_24, gen_11_cmp_pReg_23, gen_11_cmp_pReg_22, 
         gen_11_cmp_pReg_21, gen_11_cmp_pReg_20, gen_11_cmp_pReg_19, 
         gen_11_cmp_pReg_18, gen_11_cmp_pReg_17, gen_11_cmp_pReg_16, 
         gen_11_cmp_pReg_15, gen_11_cmp_pReg_14, gen_11_cmp_pReg_13, 
         gen_11_cmp_pReg_12, gen_11_cmp_pReg_11, gen_11_cmp_pReg_10, 
         gen_11_cmp_pReg_9, gen_11_cmp_pReg_8, gen_11_cmp_pReg_7, 
         gen_11_cmp_pReg_6, gen_11_cmp_pReg_5, gen_11_cmp_pReg_4, 
         gen_11_cmp_pReg_3, gen_11_cmp_pReg_2, gen_11_cmp_pReg_1, 
         gen_11_cmp_pReg_0, gen_11_cmp_BSCmp_op2_0, gen_11_cmp_BSCmp_carryIn, 
         gen_10_cmp_pBs_30, gen_10_cmp_pBs_29, gen_10_cmp_pBs_28, 
         gen_10_cmp_pBs_27, gen_10_cmp_pBs_26, gen_10_cmp_pBs_25, 
         gen_10_cmp_pBs_24, gen_10_cmp_pBs_23, gen_10_cmp_pMux_30, 
         gen_10_cmp_pMux_29, gen_10_cmp_pMux_28, gen_10_cmp_pMux_27, 
         gen_10_cmp_pMux_26, gen_10_cmp_pMux_25, gen_10_cmp_pMux_24, 
         gen_10_cmp_pMux_23, gen_10_cmp_pMux_22, gen_10_cmp_pMux_21, 
         gen_10_cmp_pMux_20, gen_10_cmp_pMux_19, gen_10_cmp_pMux_18, 
         gen_10_cmp_pMux_17, gen_10_cmp_pMux_16, gen_10_cmp_pMux_15, 
         gen_10_cmp_pMux_14, gen_10_cmp_pMux_13, gen_10_cmp_pMux_12, 
         gen_10_cmp_pMux_11, gen_10_cmp_pMux_10, gen_10_cmp_pMux_9, 
         gen_10_cmp_pMux_8, gen_10_cmp_pMux_7, gen_10_cmp_pMux_6, 
         gen_10_cmp_pMux_5, gen_10_cmp_pMux_4, gen_10_cmp_pMux_3, 
         gen_10_cmp_pMux_2, gen_10_cmp_pMux_1, gen_10_cmp_pMux_0, 
         gen_10_cmp_pReg_30, gen_10_cmp_pReg_29, gen_10_cmp_pReg_28, 
         gen_10_cmp_pReg_27, gen_10_cmp_pReg_26, gen_10_cmp_pReg_25, 
         gen_10_cmp_pReg_24, gen_10_cmp_pReg_23, gen_10_cmp_pReg_22, 
         gen_10_cmp_pReg_21, gen_10_cmp_pReg_20, gen_10_cmp_pReg_19, 
         gen_10_cmp_pReg_18, gen_10_cmp_pReg_17, gen_10_cmp_pReg_16, 
         gen_10_cmp_pReg_15, gen_10_cmp_pReg_14, gen_10_cmp_pReg_13, 
         gen_10_cmp_pReg_12, gen_10_cmp_pReg_11, gen_10_cmp_pReg_10, 
         gen_10_cmp_pReg_9, gen_10_cmp_pReg_8, gen_10_cmp_pReg_7, 
         gen_10_cmp_pReg_6, gen_10_cmp_pReg_5, gen_10_cmp_pReg_4, 
         gen_10_cmp_pReg_3, gen_10_cmp_pReg_2, gen_10_cmp_pReg_1, 
         gen_10_cmp_pReg_0, gen_10_cmp_BSCmp_op2_0, gen_10_cmp_BSCmp_carryIn, 
         gen_9_cmp_pBs_30, gen_9_cmp_pBs_29, gen_9_cmp_pBs_28, gen_9_cmp_pBs_27, 
         gen_9_cmp_pBs_26, gen_9_cmp_pBs_25, gen_9_cmp_pBs_24, gen_9_cmp_pBs_23, 
         gen_9_cmp_pMux_30, gen_9_cmp_pMux_29, gen_9_cmp_pMux_28, 
         gen_9_cmp_pMux_27, gen_9_cmp_pMux_26, gen_9_cmp_pMux_25, 
         gen_9_cmp_pMux_24, gen_9_cmp_pMux_23, gen_9_cmp_pMux_22, 
         gen_9_cmp_pMux_21, gen_9_cmp_pMux_20, gen_9_cmp_pMux_19, 
         gen_9_cmp_pMux_18, gen_9_cmp_pMux_17, gen_9_cmp_pMux_16, 
         gen_9_cmp_pMux_15, gen_9_cmp_pMux_14, gen_9_cmp_pMux_13, 
         gen_9_cmp_pMux_12, gen_9_cmp_pMux_11, gen_9_cmp_pMux_10, 
         gen_9_cmp_pMux_9, gen_9_cmp_pMux_8, gen_9_cmp_pMux_7, gen_9_cmp_pMux_6, 
         gen_9_cmp_pMux_5, gen_9_cmp_pMux_4, gen_9_cmp_pMux_3, gen_9_cmp_pMux_2, 
         gen_9_cmp_pMux_1, gen_9_cmp_pMux_0, gen_9_cmp_pReg_30, 
         gen_9_cmp_pReg_29, gen_9_cmp_pReg_28, gen_9_cmp_pReg_27, 
         gen_9_cmp_pReg_26, gen_9_cmp_pReg_25, gen_9_cmp_pReg_24, 
         gen_9_cmp_pReg_23, gen_9_cmp_pReg_22, gen_9_cmp_pReg_21, 
         gen_9_cmp_pReg_20, gen_9_cmp_pReg_19, gen_9_cmp_pReg_18, 
         gen_9_cmp_pReg_17, gen_9_cmp_pReg_16, gen_9_cmp_pReg_15, 
         gen_9_cmp_pReg_14, gen_9_cmp_pReg_13, gen_9_cmp_pReg_12, 
         gen_9_cmp_pReg_11, gen_9_cmp_pReg_10, gen_9_cmp_pReg_9, 
         gen_9_cmp_pReg_8, gen_9_cmp_pReg_7, gen_9_cmp_pReg_6, gen_9_cmp_pReg_5, 
         gen_9_cmp_pReg_4, gen_9_cmp_pReg_3, gen_9_cmp_pReg_2, gen_9_cmp_pReg_1, 
         gen_9_cmp_pReg_0, gen_9_cmp_BSCmp_op2_0, gen_9_cmp_BSCmp_carryIn, 
         gen_8_cmp_pBs_30, gen_8_cmp_pBs_29, gen_8_cmp_pBs_28, gen_8_cmp_pBs_27, 
         gen_8_cmp_pBs_26, gen_8_cmp_pBs_25, gen_8_cmp_pBs_24, gen_8_cmp_pBs_23, 
         gen_8_cmp_pMux_30, gen_8_cmp_pMux_29, gen_8_cmp_pMux_28, 
         gen_8_cmp_pMux_27, gen_8_cmp_pMux_26, gen_8_cmp_pMux_25, 
         gen_8_cmp_pMux_24, gen_8_cmp_pMux_23, gen_8_cmp_pMux_22, 
         gen_8_cmp_pMux_21, gen_8_cmp_pMux_20, gen_8_cmp_pMux_19, 
         gen_8_cmp_pMux_18, gen_8_cmp_pMux_17, gen_8_cmp_pMux_16, 
         gen_8_cmp_pMux_15, gen_8_cmp_pMux_14, gen_8_cmp_pMux_13, 
         gen_8_cmp_pMux_12, gen_8_cmp_pMux_11, gen_8_cmp_pMux_10, 
         gen_8_cmp_pMux_9, gen_8_cmp_pMux_8, gen_8_cmp_pMux_7, gen_8_cmp_pMux_6, 
         gen_8_cmp_pMux_5, gen_8_cmp_pMux_4, gen_8_cmp_pMux_3, gen_8_cmp_pMux_2, 
         gen_8_cmp_pMux_1, gen_8_cmp_pMux_0, gen_8_cmp_pReg_30, 
         gen_8_cmp_pReg_29, gen_8_cmp_pReg_28, gen_8_cmp_pReg_27, 
         gen_8_cmp_pReg_26, gen_8_cmp_pReg_25, gen_8_cmp_pReg_24, 
         gen_8_cmp_pReg_23, gen_8_cmp_pReg_22, gen_8_cmp_pReg_21, 
         gen_8_cmp_pReg_20, gen_8_cmp_pReg_19, gen_8_cmp_pReg_18, 
         gen_8_cmp_pReg_17, gen_8_cmp_pReg_16, gen_8_cmp_pReg_15, 
         gen_8_cmp_pReg_14, gen_8_cmp_pReg_13, gen_8_cmp_pReg_12, 
         gen_8_cmp_pReg_11, gen_8_cmp_pReg_10, gen_8_cmp_pReg_9, 
         gen_8_cmp_pReg_8, gen_8_cmp_pReg_7, gen_8_cmp_pReg_6, gen_8_cmp_pReg_5, 
         gen_8_cmp_pReg_4, gen_8_cmp_pReg_3, gen_8_cmp_pReg_2, gen_8_cmp_pReg_1, 
         gen_8_cmp_pReg_0, gen_8_cmp_BSCmp_op2_0, gen_8_cmp_BSCmp_carryIn, 
         gen_7_cmp_pBs_30, gen_7_cmp_pBs_29, gen_7_cmp_pBs_28, gen_7_cmp_pBs_27, 
         gen_7_cmp_pBs_26, gen_7_cmp_pBs_25, gen_7_cmp_pBs_24, gen_7_cmp_pBs_23, 
         gen_7_cmp_pMux_30, gen_7_cmp_pMux_29, gen_7_cmp_pMux_28, 
         gen_7_cmp_pMux_27, gen_7_cmp_pMux_26, gen_7_cmp_pMux_25, 
         gen_7_cmp_pMux_24, gen_7_cmp_pMux_23, gen_7_cmp_pMux_22, 
         gen_7_cmp_pMux_21, gen_7_cmp_pMux_20, gen_7_cmp_pMux_19, 
         gen_7_cmp_pMux_18, gen_7_cmp_pMux_17, gen_7_cmp_pMux_16, 
         gen_7_cmp_pMux_15, gen_7_cmp_pMux_14, gen_7_cmp_pMux_13, 
         gen_7_cmp_pMux_12, gen_7_cmp_pMux_11, gen_7_cmp_pMux_10, 
         gen_7_cmp_pMux_9, gen_7_cmp_pMux_8, gen_7_cmp_pMux_7, gen_7_cmp_pMux_6, 
         gen_7_cmp_pMux_5, gen_7_cmp_pMux_4, gen_7_cmp_pMux_3, gen_7_cmp_pMux_2, 
         gen_7_cmp_pMux_1, gen_7_cmp_pMux_0, gen_7_cmp_pReg_30, 
         gen_7_cmp_pReg_29, gen_7_cmp_pReg_28, gen_7_cmp_pReg_27, 
         gen_7_cmp_pReg_26, gen_7_cmp_pReg_25, gen_7_cmp_pReg_24, 
         gen_7_cmp_pReg_23, gen_7_cmp_pReg_22, gen_7_cmp_pReg_21, 
         gen_7_cmp_pReg_20, gen_7_cmp_pReg_19, gen_7_cmp_pReg_18, 
         gen_7_cmp_pReg_17, gen_7_cmp_pReg_16, gen_7_cmp_pReg_15, 
         gen_7_cmp_pReg_14, gen_7_cmp_pReg_13, gen_7_cmp_pReg_12, 
         gen_7_cmp_pReg_11, gen_7_cmp_pReg_10, gen_7_cmp_pReg_9, 
         gen_7_cmp_pReg_8, gen_7_cmp_pReg_7, gen_7_cmp_pReg_6, gen_7_cmp_pReg_5, 
         gen_7_cmp_pReg_4, gen_7_cmp_pReg_3, gen_7_cmp_pReg_2, gen_7_cmp_pReg_1, 
         gen_7_cmp_pReg_0, gen_7_cmp_BSCmp_op2_0, gen_7_cmp_BSCmp_carryIn, 
         gen_6_cmp_pBs_30, gen_6_cmp_pBs_29, gen_6_cmp_pBs_28, gen_6_cmp_pBs_27, 
         gen_6_cmp_pBs_26, gen_6_cmp_pBs_25, gen_6_cmp_pBs_24, gen_6_cmp_pBs_23, 
         gen_6_cmp_pMux_30, gen_6_cmp_pMux_29, gen_6_cmp_pMux_28, 
         gen_6_cmp_pMux_27, gen_6_cmp_pMux_26, gen_6_cmp_pMux_25, 
         gen_6_cmp_pMux_24, gen_6_cmp_pMux_23, gen_6_cmp_pMux_22, 
         gen_6_cmp_pMux_21, gen_6_cmp_pMux_20, gen_6_cmp_pMux_19, 
         gen_6_cmp_pMux_18, gen_6_cmp_pMux_17, gen_6_cmp_pMux_16, 
         gen_6_cmp_pMux_15, gen_6_cmp_pMux_14, gen_6_cmp_pMux_13, 
         gen_6_cmp_pMux_12, gen_6_cmp_pMux_11, gen_6_cmp_pMux_10, 
         gen_6_cmp_pMux_9, gen_6_cmp_pMux_8, gen_6_cmp_pMux_7, gen_6_cmp_pMux_6, 
         gen_6_cmp_pMux_5, gen_6_cmp_pMux_4, gen_6_cmp_pMux_3, gen_6_cmp_pMux_2, 
         gen_6_cmp_pMux_1, gen_6_cmp_pMux_0, gen_6_cmp_pReg_30, 
         gen_6_cmp_pReg_29, gen_6_cmp_pReg_28, gen_6_cmp_pReg_27, 
         gen_6_cmp_pReg_26, gen_6_cmp_pReg_25, gen_6_cmp_pReg_24, 
         gen_6_cmp_pReg_23, gen_6_cmp_pReg_22, gen_6_cmp_pReg_21, 
         gen_6_cmp_pReg_20, gen_6_cmp_pReg_19, gen_6_cmp_pReg_18, 
         gen_6_cmp_pReg_17, gen_6_cmp_pReg_16, gen_6_cmp_pReg_15, 
         gen_6_cmp_pReg_14, gen_6_cmp_pReg_13, gen_6_cmp_pReg_12, 
         gen_6_cmp_pReg_11, gen_6_cmp_pReg_10, gen_6_cmp_pReg_9, 
         gen_6_cmp_pReg_8, gen_6_cmp_pReg_7, gen_6_cmp_pReg_6, gen_6_cmp_pReg_5, 
         gen_6_cmp_pReg_4, gen_6_cmp_pReg_3, gen_6_cmp_pReg_2, gen_6_cmp_pReg_1, 
         gen_6_cmp_pReg_0, gen_6_cmp_BSCmp_op2_0, gen_6_cmp_BSCmp_carryIn, 
         gen_5_cmp_pBs_30, gen_5_cmp_pBs_29, gen_5_cmp_pBs_28, gen_5_cmp_pBs_27, 
         gen_5_cmp_pBs_26, gen_5_cmp_pBs_25, gen_5_cmp_pBs_24, gen_5_cmp_pBs_23, 
         gen_5_cmp_pMux_30, gen_5_cmp_pMux_29, gen_5_cmp_pMux_28, 
         gen_5_cmp_pMux_27, gen_5_cmp_pMux_26, gen_5_cmp_pMux_25, 
         gen_5_cmp_pMux_24, gen_5_cmp_pMux_23, gen_5_cmp_pMux_22, 
         gen_5_cmp_pMux_21, gen_5_cmp_pMux_20, gen_5_cmp_pMux_19, 
         gen_5_cmp_pMux_18, gen_5_cmp_pMux_17, gen_5_cmp_pMux_16, 
         gen_5_cmp_pMux_15, gen_5_cmp_pMux_14, gen_5_cmp_pMux_13, 
         gen_5_cmp_pMux_12, gen_5_cmp_pMux_11, gen_5_cmp_pMux_10, 
         gen_5_cmp_pMux_9, gen_5_cmp_pMux_8, gen_5_cmp_pMux_7, gen_5_cmp_pMux_6, 
         gen_5_cmp_pMux_5, gen_5_cmp_pMux_4, gen_5_cmp_pMux_3, gen_5_cmp_pMux_2, 
         gen_5_cmp_pMux_1, gen_5_cmp_pMux_0, gen_5_cmp_pReg_30, 
         gen_5_cmp_pReg_29, gen_5_cmp_pReg_28, gen_5_cmp_pReg_27, 
         gen_5_cmp_pReg_26, gen_5_cmp_pReg_25, gen_5_cmp_pReg_24, 
         gen_5_cmp_pReg_23, gen_5_cmp_pReg_22, gen_5_cmp_pReg_21, 
         gen_5_cmp_pReg_20, gen_5_cmp_pReg_19, gen_5_cmp_pReg_18, 
         gen_5_cmp_pReg_17, gen_5_cmp_pReg_16, gen_5_cmp_pReg_15, 
         gen_5_cmp_pReg_14, gen_5_cmp_pReg_13, gen_5_cmp_pReg_12, 
         gen_5_cmp_pReg_11, gen_5_cmp_pReg_10, gen_5_cmp_pReg_9, 
         gen_5_cmp_pReg_8, gen_5_cmp_pReg_7, gen_5_cmp_pReg_6, gen_5_cmp_pReg_5, 
         gen_5_cmp_pReg_4, gen_5_cmp_pReg_3, gen_5_cmp_pReg_2, gen_5_cmp_pReg_1, 
         gen_5_cmp_pReg_0, gen_5_cmp_BSCmp_op2_0, gen_5_cmp_BSCmp_carryIn, 
         gen_4_cmp_pBs_30, gen_4_cmp_pBs_29, gen_4_cmp_pBs_28, gen_4_cmp_pBs_27, 
         gen_4_cmp_pBs_26, gen_4_cmp_pBs_25, gen_4_cmp_pBs_24, gen_4_cmp_pBs_23, 
         gen_4_cmp_pMux_30, gen_4_cmp_pMux_29, gen_4_cmp_pMux_28, 
         gen_4_cmp_pMux_27, gen_4_cmp_pMux_26, gen_4_cmp_pMux_25, 
         gen_4_cmp_pMux_24, gen_4_cmp_pMux_23, gen_4_cmp_pMux_22, 
         gen_4_cmp_pMux_21, gen_4_cmp_pMux_20, gen_4_cmp_pMux_19, 
         gen_4_cmp_pMux_18, gen_4_cmp_pMux_17, gen_4_cmp_pMux_16, 
         gen_4_cmp_pMux_15, gen_4_cmp_pMux_14, gen_4_cmp_pMux_13, 
         gen_4_cmp_pMux_12, gen_4_cmp_pMux_11, gen_4_cmp_pMux_10, 
         gen_4_cmp_pMux_9, gen_4_cmp_pMux_8, gen_4_cmp_pMux_7, gen_4_cmp_pMux_6, 
         gen_4_cmp_pMux_5, gen_4_cmp_pMux_4, gen_4_cmp_pMux_3, gen_4_cmp_pMux_2, 
         gen_4_cmp_pMux_1, gen_4_cmp_pMux_0, gen_4_cmp_pReg_30, 
         gen_4_cmp_pReg_29, gen_4_cmp_pReg_28, gen_4_cmp_pReg_27, 
         gen_4_cmp_pReg_26, gen_4_cmp_pReg_25, gen_4_cmp_pReg_24, 
         gen_4_cmp_pReg_23, gen_4_cmp_pReg_22, gen_4_cmp_pReg_21, 
         gen_4_cmp_pReg_20, gen_4_cmp_pReg_19, gen_4_cmp_pReg_18, 
         gen_4_cmp_pReg_17, gen_4_cmp_pReg_16, gen_4_cmp_pReg_15, 
         gen_4_cmp_pReg_14, gen_4_cmp_pReg_13, gen_4_cmp_pReg_12, 
         gen_4_cmp_pReg_11, gen_4_cmp_pReg_10, gen_4_cmp_pReg_9, 
         gen_4_cmp_pReg_8, gen_4_cmp_pReg_7, gen_4_cmp_pReg_6, gen_4_cmp_pReg_5, 
         gen_4_cmp_pReg_4, gen_4_cmp_pReg_3, gen_4_cmp_pReg_2, gen_4_cmp_pReg_1, 
         gen_4_cmp_pReg_0, gen_4_cmp_BSCmp_op2_0, gen_4_cmp_BSCmp_carryIn, 
         gen_3_cmp_pBs_30, gen_3_cmp_pBs_29, gen_3_cmp_pBs_28, gen_3_cmp_pBs_27, 
         gen_3_cmp_pBs_26, gen_3_cmp_pBs_25, gen_3_cmp_pBs_24, gen_3_cmp_pBs_23, 
         gen_3_cmp_pMux_30, gen_3_cmp_pMux_29, gen_3_cmp_pMux_28, 
         gen_3_cmp_pMux_27, gen_3_cmp_pMux_26, gen_3_cmp_pMux_25, 
         gen_3_cmp_pMux_24, gen_3_cmp_pMux_23, gen_3_cmp_pMux_22, 
         gen_3_cmp_pMux_21, gen_3_cmp_pMux_20, gen_3_cmp_pMux_19, 
         gen_3_cmp_pMux_18, gen_3_cmp_pMux_17, gen_3_cmp_pMux_16, 
         gen_3_cmp_pMux_15, gen_3_cmp_pMux_14, gen_3_cmp_pMux_13, 
         gen_3_cmp_pMux_12, gen_3_cmp_pMux_11, gen_3_cmp_pMux_10, 
         gen_3_cmp_pMux_9, gen_3_cmp_pMux_8, gen_3_cmp_pMux_7, gen_3_cmp_pMux_6, 
         gen_3_cmp_pMux_5, gen_3_cmp_pMux_4, gen_3_cmp_pMux_3, gen_3_cmp_pMux_2, 
         gen_3_cmp_pMux_1, gen_3_cmp_pMux_0, gen_3_cmp_pReg_30, 
         gen_3_cmp_pReg_29, gen_3_cmp_pReg_28, gen_3_cmp_pReg_27, 
         gen_3_cmp_pReg_26, gen_3_cmp_pReg_25, gen_3_cmp_pReg_24, 
         gen_3_cmp_pReg_23, gen_3_cmp_pReg_22, gen_3_cmp_pReg_21, 
         gen_3_cmp_pReg_20, gen_3_cmp_pReg_19, gen_3_cmp_pReg_18, 
         gen_3_cmp_pReg_17, gen_3_cmp_pReg_16, gen_3_cmp_pReg_15, 
         gen_3_cmp_pReg_14, gen_3_cmp_pReg_13, gen_3_cmp_pReg_12, 
         gen_3_cmp_pReg_11, gen_3_cmp_pReg_10, gen_3_cmp_pReg_9, 
         gen_3_cmp_pReg_8, gen_3_cmp_pReg_7, gen_3_cmp_pReg_6, gen_3_cmp_pReg_5, 
         gen_3_cmp_pReg_4, gen_3_cmp_pReg_3, gen_3_cmp_pReg_2, gen_3_cmp_pReg_1, 
         gen_3_cmp_pReg_0, gen_3_cmp_BSCmp_op2_0, gen_3_cmp_BSCmp_carryIn, 
         gen_2_cmp_pBs_30, gen_2_cmp_pBs_29, gen_2_cmp_pBs_28, gen_2_cmp_pBs_27, 
         gen_2_cmp_pBs_26, gen_2_cmp_pBs_25, gen_2_cmp_pBs_24, gen_2_cmp_pBs_23, 
         gen_2_cmp_pMux_30, gen_2_cmp_pMux_29, gen_2_cmp_pMux_28, 
         gen_2_cmp_pMux_27, gen_2_cmp_pMux_26, gen_2_cmp_pMux_25, 
         gen_2_cmp_pMux_24, gen_2_cmp_pMux_23, gen_2_cmp_pMux_22, 
         gen_2_cmp_pMux_21, gen_2_cmp_pMux_20, gen_2_cmp_pMux_19, 
         gen_2_cmp_pMux_18, gen_2_cmp_pMux_17, gen_2_cmp_pMux_16, 
         gen_2_cmp_pMux_15, gen_2_cmp_pMux_14, gen_2_cmp_pMux_13, 
         gen_2_cmp_pMux_12, gen_2_cmp_pMux_11, gen_2_cmp_pMux_10, 
         gen_2_cmp_pMux_9, gen_2_cmp_pMux_8, gen_2_cmp_pMux_7, gen_2_cmp_pMux_6, 
         gen_2_cmp_pMux_5, gen_2_cmp_pMux_4, gen_2_cmp_pMux_3, gen_2_cmp_pMux_2, 
         gen_2_cmp_pMux_1, gen_2_cmp_pMux_0, gen_2_cmp_pReg_30, 
         gen_2_cmp_pReg_29, gen_2_cmp_pReg_28, gen_2_cmp_pReg_27, 
         gen_2_cmp_pReg_26, gen_2_cmp_pReg_25, gen_2_cmp_pReg_24, 
         gen_2_cmp_pReg_23, gen_2_cmp_pReg_22, gen_2_cmp_pReg_21, 
         gen_2_cmp_pReg_20, gen_2_cmp_pReg_19, gen_2_cmp_pReg_18, 
         gen_2_cmp_pReg_17, gen_2_cmp_pReg_16, gen_2_cmp_pReg_15, 
         gen_2_cmp_pReg_14, gen_2_cmp_pReg_13, gen_2_cmp_pReg_12, 
         gen_2_cmp_pReg_11, gen_2_cmp_pReg_10, gen_2_cmp_pReg_9, 
         gen_2_cmp_pReg_8, gen_2_cmp_pReg_7, gen_2_cmp_pReg_6, gen_2_cmp_pReg_5, 
         gen_2_cmp_pReg_4, gen_2_cmp_pReg_3, gen_2_cmp_pReg_2, gen_2_cmp_pReg_1, 
         gen_2_cmp_pReg_0, gen_2_cmp_BSCmp_op2_0, gen_2_cmp_BSCmp_carryIn, 
         gen_1_cmp_pBs_30, gen_1_cmp_pBs_29, gen_1_cmp_pBs_28, gen_1_cmp_pBs_27, 
         gen_1_cmp_pBs_26, gen_1_cmp_pBs_25, gen_1_cmp_pBs_24, gen_1_cmp_pBs_23, 
         gen_1_cmp_pMux_30, gen_1_cmp_pMux_29, gen_1_cmp_pMux_28, 
         gen_1_cmp_pMux_27, gen_1_cmp_pMux_26, gen_1_cmp_pMux_25, 
         gen_1_cmp_pMux_24, gen_1_cmp_pMux_23, gen_1_cmp_pMux_22, 
         gen_1_cmp_pMux_21, gen_1_cmp_pMux_20, gen_1_cmp_pMux_19, 
         gen_1_cmp_pMux_18, gen_1_cmp_pMux_17, gen_1_cmp_pMux_16, 
         gen_1_cmp_pMux_15, gen_1_cmp_pMux_14, gen_1_cmp_pMux_13, 
         gen_1_cmp_pMux_12, gen_1_cmp_pMux_11, gen_1_cmp_pMux_10, 
         gen_1_cmp_pMux_9, gen_1_cmp_pMux_8, gen_1_cmp_pMux_7, gen_1_cmp_pMux_6, 
         gen_1_cmp_pMux_5, gen_1_cmp_pMux_4, gen_1_cmp_pMux_3, gen_1_cmp_pMux_2, 
         gen_1_cmp_pMux_1, gen_1_cmp_pMux_0, gen_1_cmp_pReg_30, 
         gen_1_cmp_pReg_29, gen_1_cmp_pReg_28, gen_1_cmp_pReg_27, 
         gen_1_cmp_pReg_26, gen_1_cmp_pReg_25, gen_1_cmp_pReg_24, 
         gen_1_cmp_pReg_23, gen_1_cmp_pReg_22, gen_1_cmp_pReg_21, 
         gen_1_cmp_pReg_20, gen_1_cmp_pReg_19, gen_1_cmp_pReg_18, 
         gen_1_cmp_pReg_17, gen_1_cmp_pReg_16, gen_1_cmp_pReg_15, 
         gen_1_cmp_pReg_14, gen_1_cmp_pReg_13, gen_1_cmp_pReg_12, 
         gen_1_cmp_pReg_11, gen_1_cmp_pReg_10, gen_1_cmp_pReg_9, 
         gen_1_cmp_pReg_8, gen_1_cmp_pReg_7, gen_1_cmp_pReg_6, gen_1_cmp_pReg_5, 
         gen_1_cmp_pReg_4, gen_1_cmp_pReg_3, gen_1_cmp_pReg_2, gen_1_cmp_pReg_1, 
         gen_1_cmp_pReg_0, gen_1_cmp_BSCmp_op2_0, gen_1_cmp_BSCmp_carryIn, 
         gen_0_cmp_pBs_30, gen_0_cmp_pBs_29, gen_0_cmp_pBs_28, gen_0_cmp_pBs_27, 
         gen_0_cmp_pBs_26, gen_0_cmp_pBs_25, gen_0_cmp_pBs_24, gen_0_cmp_pBs_23, 
         gen_0_cmp_pMux_30, gen_0_cmp_pMux_29, gen_0_cmp_pMux_28, 
         gen_0_cmp_pMux_27, gen_0_cmp_pMux_26, gen_0_cmp_pMux_25, 
         gen_0_cmp_pMux_24, gen_0_cmp_pMux_23, gen_0_cmp_pMux_22, 
         gen_0_cmp_pMux_21, gen_0_cmp_pMux_20, gen_0_cmp_pMux_19, 
         gen_0_cmp_pMux_18, gen_0_cmp_pMux_17, gen_0_cmp_pMux_16, 
         gen_0_cmp_pMux_15, gen_0_cmp_pMux_14, gen_0_cmp_pMux_13, 
         gen_0_cmp_pMux_12, gen_0_cmp_pMux_11, gen_0_cmp_pMux_10, 
         gen_0_cmp_pMux_9, gen_0_cmp_pMux_8, gen_0_cmp_pMux_7, gen_0_cmp_pMux_6, 
         gen_0_cmp_pMux_5, gen_0_cmp_pMux_4, gen_0_cmp_pMux_3, gen_0_cmp_pMux_2, 
         gen_0_cmp_pMux_1, gen_0_cmp_pMux_0, gen_0_cmp_pReg_30, 
         gen_0_cmp_pReg_29, gen_0_cmp_pReg_28, gen_0_cmp_pReg_27, 
         gen_0_cmp_pReg_26, gen_0_cmp_pReg_25, gen_0_cmp_pReg_24, 
         gen_0_cmp_pReg_23, gen_0_cmp_pReg_22, gen_0_cmp_pReg_21, 
         gen_0_cmp_pReg_20, gen_0_cmp_pReg_19, gen_0_cmp_pReg_18, 
         gen_0_cmp_pReg_17, gen_0_cmp_pReg_16, gen_0_cmp_pReg_15, 
         gen_0_cmp_pReg_14, gen_0_cmp_pReg_13, gen_0_cmp_pReg_12, 
         gen_0_cmp_pReg_11, gen_0_cmp_pReg_10, gen_0_cmp_pReg_9, 
         gen_0_cmp_pReg_8, gen_0_cmp_pReg_7, gen_0_cmp_pReg_6, gen_0_cmp_pReg_5, 
         gen_0_cmp_pReg_4, gen_0_cmp_pReg_3, gen_0_cmp_pReg_2, gen_0_cmp_pReg_1, 
         gen_0_cmp_pReg_0, gen_0_cmp_BSCmp_op2_0, gen_0_cmp_BSCmp_carryIn, 
         gen_24_cmp_BSCmp_op2_16, gen_24_cmp_BSCmp_op2_15, 
         gen_24_cmp_BSCmp_op2_14, gen_24_cmp_BSCmp_op2_13, 
         gen_24_cmp_BSCmp_op2_12, gen_24_cmp_BSCmp_op2_11, 
         gen_24_cmp_BSCmp_op2_10, gen_24_cmp_BSCmp_op2_9, gen_24_cmp_BSCmp_op2_8, 
         gen_24_cmp_BSCmp_op2_7, gen_24_cmp_BSCmp_op2_6, gen_24_cmp_BSCmp_op2_5, 
         gen_24_cmp_BSCmp_op2_4, gen_24_cmp_BSCmp_op2_3, gen_24_cmp_BSCmp_op2_2, 
         gen_24_cmp_BSCmp_op2_1, gen_23_cmp_BSCmp_op2_16, 
         gen_23_cmp_BSCmp_op2_15, gen_23_cmp_BSCmp_op2_14, 
         gen_23_cmp_BSCmp_op2_13, gen_23_cmp_BSCmp_op2_12, 
         gen_23_cmp_BSCmp_op2_11, gen_23_cmp_BSCmp_op2_10, 
         gen_23_cmp_BSCmp_op2_9, gen_23_cmp_BSCmp_op2_8, gen_23_cmp_BSCmp_op2_7, 
         gen_23_cmp_BSCmp_op2_6, gen_23_cmp_BSCmp_op2_5, gen_23_cmp_BSCmp_op2_4, 
         gen_23_cmp_BSCmp_op2_3, gen_23_cmp_BSCmp_op2_2, gen_23_cmp_BSCmp_op2_1, 
         gen_22_cmp_BSCmp_op2_16, gen_22_cmp_BSCmp_op2_15, 
         gen_22_cmp_BSCmp_op2_14, gen_22_cmp_BSCmp_op2_13, 
         gen_22_cmp_BSCmp_op2_12, gen_22_cmp_BSCmp_op2_11, 
         gen_22_cmp_BSCmp_op2_10, gen_22_cmp_BSCmp_op2_9, gen_22_cmp_BSCmp_op2_8, 
         gen_22_cmp_BSCmp_op2_7, gen_22_cmp_BSCmp_op2_6, gen_22_cmp_BSCmp_op2_5, 
         gen_22_cmp_BSCmp_op2_4, gen_22_cmp_BSCmp_op2_3, gen_22_cmp_BSCmp_op2_2, 
         gen_22_cmp_BSCmp_op2_1, gen_21_cmp_BSCmp_op2_16, 
         gen_21_cmp_BSCmp_op2_15, gen_21_cmp_BSCmp_op2_14, 
         gen_21_cmp_BSCmp_op2_13, gen_21_cmp_BSCmp_op2_12, 
         gen_21_cmp_BSCmp_op2_11, gen_21_cmp_BSCmp_op2_10, 
         gen_21_cmp_BSCmp_op2_9, gen_21_cmp_BSCmp_op2_8, gen_21_cmp_BSCmp_op2_7, 
         gen_21_cmp_BSCmp_op2_6, gen_21_cmp_BSCmp_op2_5, gen_21_cmp_BSCmp_op2_4, 
         gen_21_cmp_BSCmp_op2_3, gen_21_cmp_BSCmp_op2_2, gen_21_cmp_BSCmp_op2_1, 
         gen_20_cmp_BSCmp_op2_16, gen_20_cmp_BSCmp_op2_15, 
         gen_20_cmp_BSCmp_op2_14, gen_20_cmp_BSCmp_op2_13, 
         gen_20_cmp_BSCmp_op2_12, gen_20_cmp_BSCmp_op2_11, 
         gen_20_cmp_BSCmp_op2_10, gen_20_cmp_BSCmp_op2_9, gen_20_cmp_BSCmp_op2_8, 
         gen_20_cmp_BSCmp_op2_7, gen_20_cmp_BSCmp_op2_6, gen_20_cmp_BSCmp_op2_5, 
         gen_20_cmp_BSCmp_op2_4, gen_20_cmp_BSCmp_op2_3, gen_20_cmp_BSCmp_op2_2, 
         gen_20_cmp_BSCmp_op2_1, gen_19_cmp_BSCmp_op2_16, 
         gen_19_cmp_BSCmp_op2_15, gen_19_cmp_BSCmp_op2_14, 
         gen_19_cmp_BSCmp_op2_13, gen_19_cmp_BSCmp_op2_12, 
         gen_19_cmp_BSCmp_op2_11, gen_19_cmp_BSCmp_op2_10, 
         gen_19_cmp_BSCmp_op2_9, gen_19_cmp_BSCmp_op2_8, gen_19_cmp_BSCmp_op2_7, 
         gen_19_cmp_BSCmp_op2_6, gen_19_cmp_BSCmp_op2_5, gen_19_cmp_BSCmp_op2_4, 
         gen_19_cmp_BSCmp_op2_3, gen_19_cmp_BSCmp_op2_2, gen_19_cmp_BSCmp_op2_1, 
         gen_18_cmp_BSCmp_op2_16, gen_18_cmp_BSCmp_op2_15, 
         gen_18_cmp_BSCmp_op2_14, gen_18_cmp_BSCmp_op2_13, 
         gen_18_cmp_BSCmp_op2_12, gen_18_cmp_BSCmp_op2_11, 
         gen_18_cmp_BSCmp_op2_10, gen_18_cmp_BSCmp_op2_9, gen_18_cmp_BSCmp_op2_8, 
         gen_18_cmp_BSCmp_op2_7, gen_18_cmp_BSCmp_op2_6, gen_18_cmp_BSCmp_op2_5, 
         gen_18_cmp_BSCmp_op2_4, gen_18_cmp_BSCmp_op2_3, gen_18_cmp_BSCmp_op2_2, 
         gen_18_cmp_BSCmp_op2_1, gen_17_cmp_BSCmp_op2_16, 
         gen_17_cmp_BSCmp_op2_15, gen_17_cmp_BSCmp_op2_14, 
         gen_17_cmp_BSCmp_op2_13, gen_17_cmp_BSCmp_op2_12, 
         gen_17_cmp_BSCmp_op2_11, gen_17_cmp_BSCmp_op2_10, 
         gen_17_cmp_BSCmp_op2_9, gen_17_cmp_BSCmp_op2_8, gen_17_cmp_BSCmp_op2_7, 
         gen_17_cmp_BSCmp_op2_6, gen_17_cmp_BSCmp_op2_5, gen_17_cmp_BSCmp_op2_4, 
         gen_17_cmp_BSCmp_op2_3, gen_17_cmp_BSCmp_op2_2, gen_17_cmp_BSCmp_op2_1, 
         gen_16_cmp_BSCmp_op2_16, gen_16_cmp_BSCmp_op2_15, 
         gen_16_cmp_BSCmp_op2_14, gen_16_cmp_BSCmp_op2_13, 
         gen_16_cmp_BSCmp_op2_12, gen_16_cmp_BSCmp_op2_11, 
         gen_16_cmp_BSCmp_op2_10, gen_16_cmp_BSCmp_op2_9, gen_16_cmp_BSCmp_op2_8, 
         gen_16_cmp_BSCmp_op2_7, gen_16_cmp_BSCmp_op2_6, gen_16_cmp_BSCmp_op2_5, 
         gen_16_cmp_BSCmp_op2_4, gen_16_cmp_BSCmp_op2_3, gen_16_cmp_BSCmp_op2_2, 
         gen_16_cmp_BSCmp_op2_1, gen_15_cmp_BSCmp_op2_16, 
         gen_15_cmp_BSCmp_op2_15, gen_15_cmp_BSCmp_op2_14, 
         gen_15_cmp_BSCmp_op2_13, gen_15_cmp_BSCmp_op2_12, 
         gen_15_cmp_BSCmp_op2_11, gen_15_cmp_BSCmp_op2_10, 
         gen_15_cmp_BSCmp_op2_9, gen_15_cmp_BSCmp_op2_8, gen_15_cmp_BSCmp_op2_7, 
         gen_15_cmp_BSCmp_op2_6, gen_15_cmp_BSCmp_op2_5, gen_15_cmp_BSCmp_op2_4, 
         gen_15_cmp_BSCmp_op2_3, gen_15_cmp_BSCmp_op2_2, gen_15_cmp_BSCmp_op2_1, 
         gen_14_cmp_BSCmp_op2_16, gen_14_cmp_BSCmp_op2_15, 
         gen_14_cmp_BSCmp_op2_14, gen_14_cmp_BSCmp_op2_13, 
         gen_14_cmp_BSCmp_op2_12, gen_14_cmp_BSCmp_op2_11, 
         gen_14_cmp_BSCmp_op2_10, gen_14_cmp_BSCmp_op2_9, gen_14_cmp_BSCmp_op2_8, 
         gen_14_cmp_BSCmp_op2_7, gen_14_cmp_BSCmp_op2_6, gen_14_cmp_BSCmp_op2_5, 
         gen_14_cmp_BSCmp_op2_4, gen_14_cmp_BSCmp_op2_3, gen_14_cmp_BSCmp_op2_2, 
         gen_14_cmp_BSCmp_op2_1, gen_13_cmp_BSCmp_op2_16, 
         gen_13_cmp_BSCmp_op2_15, gen_13_cmp_BSCmp_op2_14, 
         gen_13_cmp_BSCmp_op2_13, gen_13_cmp_BSCmp_op2_12, 
         gen_13_cmp_BSCmp_op2_11, gen_13_cmp_BSCmp_op2_10, 
         gen_13_cmp_BSCmp_op2_9, gen_13_cmp_BSCmp_op2_8, gen_13_cmp_BSCmp_op2_7, 
         gen_13_cmp_BSCmp_op2_6, gen_13_cmp_BSCmp_op2_5, gen_13_cmp_BSCmp_op2_4, 
         gen_13_cmp_BSCmp_op2_3, gen_13_cmp_BSCmp_op2_2, gen_13_cmp_BSCmp_op2_1, 
         gen_12_cmp_BSCmp_op2_16, gen_12_cmp_BSCmp_op2_15, 
         gen_12_cmp_BSCmp_op2_14, gen_12_cmp_BSCmp_op2_13, 
         gen_12_cmp_BSCmp_op2_12, gen_12_cmp_BSCmp_op2_11, 
         gen_12_cmp_BSCmp_op2_10, gen_12_cmp_BSCmp_op2_9, gen_12_cmp_BSCmp_op2_8, 
         gen_12_cmp_BSCmp_op2_7, gen_12_cmp_BSCmp_op2_6, gen_12_cmp_BSCmp_op2_5, 
         gen_12_cmp_BSCmp_op2_4, gen_12_cmp_BSCmp_op2_3, gen_12_cmp_BSCmp_op2_2, 
         gen_12_cmp_BSCmp_op2_1, gen_11_cmp_BSCmp_op2_16, 
         gen_11_cmp_BSCmp_op2_15, gen_11_cmp_BSCmp_op2_14, 
         gen_11_cmp_BSCmp_op2_13, gen_11_cmp_BSCmp_op2_12, 
         gen_11_cmp_BSCmp_op2_11, gen_11_cmp_BSCmp_op2_10, 
         gen_11_cmp_BSCmp_op2_9, gen_11_cmp_BSCmp_op2_8, gen_11_cmp_BSCmp_op2_7, 
         gen_11_cmp_BSCmp_op2_6, gen_11_cmp_BSCmp_op2_5, gen_11_cmp_BSCmp_op2_4, 
         gen_11_cmp_BSCmp_op2_3, gen_11_cmp_BSCmp_op2_2, gen_11_cmp_BSCmp_op2_1, 
         gen_10_cmp_BSCmp_op2_16, gen_10_cmp_BSCmp_op2_15, 
         gen_10_cmp_BSCmp_op2_14, gen_10_cmp_BSCmp_op2_13, 
         gen_10_cmp_BSCmp_op2_12, gen_10_cmp_BSCmp_op2_11, 
         gen_10_cmp_BSCmp_op2_10, gen_10_cmp_BSCmp_op2_9, gen_10_cmp_BSCmp_op2_8, 
         gen_10_cmp_BSCmp_op2_7, gen_10_cmp_BSCmp_op2_6, gen_10_cmp_BSCmp_op2_5, 
         gen_10_cmp_BSCmp_op2_4, gen_10_cmp_BSCmp_op2_3, gen_10_cmp_BSCmp_op2_2, 
         gen_10_cmp_BSCmp_op2_1, gen_9_cmp_BSCmp_op2_16, gen_9_cmp_BSCmp_op2_15, 
         gen_9_cmp_BSCmp_op2_14, gen_9_cmp_BSCmp_op2_13, gen_9_cmp_BSCmp_op2_12, 
         gen_9_cmp_BSCmp_op2_11, gen_9_cmp_BSCmp_op2_10, gen_9_cmp_BSCmp_op2_9, 
         gen_9_cmp_BSCmp_op2_8, gen_9_cmp_BSCmp_op2_7, gen_9_cmp_BSCmp_op2_6, 
         gen_9_cmp_BSCmp_op2_5, gen_9_cmp_BSCmp_op2_4, gen_9_cmp_BSCmp_op2_3, 
         gen_9_cmp_BSCmp_op2_2, gen_9_cmp_BSCmp_op2_1, gen_8_cmp_BSCmp_op2_16, 
         gen_8_cmp_BSCmp_op2_15, gen_8_cmp_BSCmp_op2_14, gen_8_cmp_BSCmp_op2_13, 
         gen_8_cmp_BSCmp_op2_12, gen_8_cmp_BSCmp_op2_11, gen_8_cmp_BSCmp_op2_10, 
         gen_8_cmp_BSCmp_op2_9, gen_8_cmp_BSCmp_op2_8, gen_8_cmp_BSCmp_op2_7, 
         gen_8_cmp_BSCmp_op2_6, gen_8_cmp_BSCmp_op2_5, gen_8_cmp_BSCmp_op2_4, 
         gen_8_cmp_BSCmp_op2_3, gen_8_cmp_BSCmp_op2_2, gen_8_cmp_BSCmp_op2_1, 
         gen_7_cmp_BSCmp_op2_16, gen_7_cmp_BSCmp_op2_15, gen_7_cmp_BSCmp_op2_14, 
         gen_7_cmp_BSCmp_op2_13, gen_7_cmp_BSCmp_op2_12, gen_7_cmp_BSCmp_op2_11, 
         gen_7_cmp_BSCmp_op2_10, gen_7_cmp_BSCmp_op2_9, gen_7_cmp_BSCmp_op2_8, 
         gen_7_cmp_BSCmp_op2_7, gen_7_cmp_BSCmp_op2_6, gen_7_cmp_BSCmp_op2_5, 
         gen_7_cmp_BSCmp_op2_4, gen_7_cmp_BSCmp_op2_3, gen_7_cmp_BSCmp_op2_2, 
         gen_7_cmp_BSCmp_op2_1, gen_6_cmp_BSCmp_op2_16, gen_6_cmp_BSCmp_op2_15, 
         gen_6_cmp_BSCmp_op2_14, gen_6_cmp_BSCmp_op2_13, gen_6_cmp_BSCmp_op2_12, 
         gen_6_cmp_BSCmp_op2_11, gen_6_cmp_BSCmp_op2_10, gen_6_cmp_BSCmp_op2_9, 
         gen_6_cmp_BSCmp_op2_8, gen_6_cmp_BSCmp_op2_7, gen_6_cmp_BSCmp_op2_6, 
         gen_6_cmp_BSCmp_op2_5, gen_6_cmp_BSCmp_op2_4, gen_6_cmp_BSCmp_op2_3, 
         gen_6_cmp_BSCmp_op2_2, gen_6_cmp_BSCmp_op2_1, gen_5_cmp_BSCmp_op2_16, 
         gen_5_cmp_BSCmp_op2_15, gen_5_cmp_BSCmp_op2_14, gen_5_cmp_BSCmp_op2_13, 
         gen_5_cmp_BSCmp_op2_12, gen_5_cmp_BSCmp_op2_11, gen_5_cmp_BSCmp_op2_10, 
         gen_5_cmp_BSCmp_op2_9, gen_5_cmp_BSCmp_op2_8, gen_5_cmp_BSCmp_op2_7, 
         gen_5_cmp_BSCmp_op2_6, gen_5_cmp_BSCmp_op2_5, gen_5_cmp_BSCmp_op2_4, 
         gen_5_cmp_BSCmp_op2_3, gen_5_cmp_BSCmp_op2_2, gen_5_cmp_BSCmp_op2_1, 
         gen_4_cmp_BSCmp_op2_16, gen_4_cmp_BSCmp_op2_15, gen_4_cmp_BSCmp_op2_14, 
         gen_4_cmp_BSCmp_op2_13, gen_4_cmp_BSCmp_op2_12, gen_4_cmp_BSCmp_op2_11, 
         gen_4_cmp_BSCmp_op2_10, gen_4_cmp_BSCmp_op2_9, gen_4_cmp_BSCmp_op2_8, 
         gen_4_cmp_BSCmp_op2_7, gen_4_cmp_BSCmp_op2_6, gen_4_cmp_BSCmp_op2_5, 
         gen_4_cmp_BSCmp_op2_4, gen_4_cmp_BSCmp_op2_3, gen_4_cmp_BSCmp_op2_2, 
         gen_4_cmp_BSCmp_op2_1, gen_3_cmp_BSCmp_op2_16, gen_3_cmp_BSCmp_op2_15, 
         gen_3_cmp_BSCmp_op2_14, gen_3_cmp_BSCmp_op2_13, gen_3_cmp_BSCmp_op2_12, 
         gen_3_cmp_BSCmp_op2_11, gen_3_cmp_BSCmp_op2_10, gen_3_cmp_BSCmp_op2_9, 
         gen_3_cmp_BSCmp_op2_8, gen_3_cmp_BSCmp_op2_7, gen_3_cmp_BSCmp_op2_6, 
         gen_3_cmp_BSCmp_op2_5, gen_3_cmp_BSCmp_op2_4, gen_3_cmp_BSCmp_op2_3, 
         gen_3_cmp_BSCmp_op2_2, gen_3_cmp_BSCmp_op2_1, gen_2_cmp_BSCmp_op2_16, 
         gen_2_cmp_BSCmp_op2_15, gen_2_cmp_BSCmp_op2_14, gen_2_cmp_BSCmp_op2_13, 
         gen_2_cmp_BSCmp_op2_12, gen_2_cmp_BSCmp_op2_11, gen_2_cmp_BSCmp_op2_10, 
         gen_2_cmp_BSCmp_op2_9, gen_2_cmp_BSCmp_op2_8, gen_2_cmp_BSCmp_op2_7, 
         gen_2_cmp_BSCmp_op2_6, gen_2_cmp_BSCmp_op2_5, gen_2_cmp_BSCmp_op2_4, 
         gen_2_cmp_BSCmp_op2_3, gen_2_cmp_BSCmp_op2_2, gen_2_cmp_BSCmp_op2_1, 
         gen_1_cmp_BSCmp_op2_16, gen_1_cmp_BSCmp_op2_15, gen_1_cmp_BSCmp_op2_14, 
         gen_1_cmp_BSCmp_op2_13, gen_1_cmp_BSCmp_op2_12, gen_1_cmp_BSCmp_op2_11, 
         gen_1_cmp_BSCmp_op2_10, gen_1_cmp_BSCmp_op2_9, gen_1_cmp_BSCmp_op2_8, 
         gen_1_cmp_BSCmp_op2_7, gen_1_cmp_BSCmp_op2_6, gen_1_cmp_BSCmp_op2_5, 
         gen_1_cmp_BSCmp_op2_4, gen_1_cmp_BSCmp_op2_3, gen_1_cmp_BSCmp_op2_2, 
         gen_1_cmp_BSCmp_op2_1, gen_0_cmp_BSCmp_op2_16, gen_0_cmp_BSCmp_op2_15, 
         gen_0_cmp_BSCmp_op2_14, gen_0_cmp_BSCmp_op2_13, gen_0_cmp_BSCmp_op2_12, 
         gen_0_cmp_BSCmp_op2_11, gen_0_cmp_BSCmp_op2_10, gen_0_cmp_BSCmp_op2_9, 
         gen_0_cmp_BSCmp_op2_8, gen_0_cmp_BSCmp_op2_7, gen_0_cmp_BSCmp_op2_6, 
         gen_0_cmp_BSCmp_op2_5, gen_0_cmp_BSCmp_op2_4, gen_0_cmp_BSCmp_op2_3, 
         gen_0_cmp_BSCmp_op2_2, gen_0_cmp_BSCmp_op2_1, nx6, gen_0_cmp_mReg_0, 
         nx26, nx34, gen_0_cmp_mReg_1, nx46, nx48, nx58, nx62, gen_0_cmp_mReg_2, 
         nx74, nx76, nx80, nx84, gen_0_cmp_mReg_3, nx96, nx98, nx102, nx106, 
         gen_0_cmp_mReg_4, nx118, nx120, nx124, nx128, gen_0_cmp_mReg_5, nx140, 
         nx142, nx146, nx150, gen_0_cmp_mReg_6, nx162, nx164, nx168, nx172, 
         gen_0_cmp_mReg_7, nx184, nx186, nx190, nx194, gen_0_cmp_mReg_8, nx206, 
         nx208, nx212, nx216, gen_0_cmp_mReg_9, nx228, nx230, nx234, nx238, 
         gen_0_cmp_mReg_10, nx250, nx252, nx256, nx260, gen_0_cmp_mReg_11, nx272, 
         nx274, nx278, nx282, gen_0_cmp_mReg_12, nx294, nx296, nx300, nx304, 
         gen_0_cmp_mReg_13, nx316, nx318, nx322, nx326, gen_0_cmp_mReg_14, nx338, 
         nx340, nx344, nx348, gen_0_cmp_mReg_15, nx360, nx362, nx366, nx370, 
         nx376, nx380, nx392, gen_1_cmp_mReg_0, nx412, nx420, gen_1_cmp_mReg_1, 
         nx432, nx434, nx444, nx448, gen_1_cmp_mReg_2, nx460, nx462, nx466, 
         nx470, gen_1_cmp_mReg_3, nx482, nx484, nx488, nx492, gen_1_cmp_mReg_4, 
         nx504, nx506, nx510, nx514, gen_1_cmp_mReg_5, nx526, nx528, nx532, 
         nx536, gen_1_cmp_mReg_6, nx548, nx550, nx554, nx558, gen_1_cmp_mReg_7, 
         nx570, nx572, nx576, nx580, gen_1_cmp_mReg_8, nx592, nx594, nx598, 
         nx602, gen_1_cmp_mReg_9, nx614, nx616, nx620, nx624, gen_1_cmp_mReg_10, 
         nx636, nx638, nx642, nx646, gen_1_cmp_mReg_11, nx658, nx660, nx664, 
         nx668, gen_1_cmp_mReg_12, nx680, nx682, nx686, nx690, gen_1_cmp_mReg_13, 
         nx702, nx704, nx708, nx712, gen_1_cmp_mReg_14, nx724, nx726, nx730, 
         nx734, gen_1_cmp_mReg_15, nx746, nx748, nx752, nx756, nx762, nx766, 
         nx778, gen_2_cmp_mReg_0, nx798, nx806, gen_2_cmp_mReg_1, nx818, nx820, 
         nx830, nx834, gen_2_cmp_mReg_2, nx846, nx848, nx852, nx856, 
         gen_2_cmp_mReg_3, nx868, nx870, nx874, nx878, gen_2_cmp_mReg_4, nx890, 
         nx892, nx896, nx900, gen_2_cmp_mReg_5, nx912, nx914, nx918, nx922, 
         gen_2_cmp_mReg_6, nx934, nx936, nx940, nx944, gen_2_cmp_mReg_7, nx956, 
         nx958, nx962, nx966, gen_2_cmp_mReg_8, nx978, nx980, nx984, nx988, 
         gen_2_cmp_mReg_9, nx1000, nx1002, nx1006, nx1010, gen_2_cmp_mReg_10, 
         nx1022, nx1024, nx1028, nx1032, gen_2_cmp_mReg_11, nx1044, nx1046, 
         nx1050, nx1054, gen_2_cmp_mReg_12, nx1066, nx1068, nx1072, nx1076, 
         gen_2_cmp_mReg_13, nx1088, nx1090, nx1094, nx1098, gen_2_cmp_mReg_14, 
         nx1110, nx1112, nx1116, nx1120, gen_2_cmp_mReg_15, nx1132, nx1134, 
         nx1138, nx1142, nx1148, nx1152, nx1164, gen_3_cmp_mReg_0, nx1184, 
         nx1192, gen_3_cmp_mReg_1, nx1204, nx1206, nx1216, nx1220, 
         gen_3_cmp_mReg_2, nx1232, nx1234, nx1238, nx1242, gen_3_cmp_mReg_3, 
         nx1254, nx1256, nx1260, nx1264, gen_3_cmp_mReg_4, nx1276, nx1278, 
         nx1282, nx1286, gen_3_cmp_mReg_5, nx1298, nx1300, nx1304, nx1308, 
         gen_3_cmp_mReg_6, nx1320, nx1322, nx1326, nx1330, gen_3_cmp_mReg_7, 
         nx1342, nx1344, nx1348, nx1352, gen_3_cmp_mReg_8, nx1364, nx1366, 
         nx1370, nx1374, gen_3_cmp_mReg_9, nx1386, nx1388, nx1392, nx1396, 
         gen_3_cmp_mReg_10, nx1408, nx1410, nx1414, nx1418, gen_3_cmp_mReg_11, 
         nx1430, nx1432, nx1436, nx1440, gen_3_cmp_mReg_12, nx1452, nx1454, 
         nx1458, nx1462, gen_3_cmp_mReg_13, nx1474, nx1476, nx1480, nx1484, 
         gen_3_cmp_mReg_14, nx1496, nx1498, nx1502, nx1506, gen_3_cmp_mReg_15, 
         nx1518, nx1520, nx1524, nx1528, nx1534, nx1538, nx1550, 
         gen_4_cmp_mReg_0, nx1570, nx1578, gen_4_cmp_mReg_1, nx1590, nx1592, 
         nx1602, nx1606, gen_4_cmp_mReg_2, nx1618, nx1620, nx1624, nx1628, 
         gen_4_cmp_mReg_3, nx1640, nx1642, nx1646, nx1650, gen_4_cmp_mReg_4, 
         nx1662, nx1664, nx1668, nx1672, gen_4_cmp_mReg_5, nx1684, nx1686, 
         nx1690, nx1694, gen_4_cmp_mReg_6, nx1706, nx1708, nx1712, nx1716, 
         gen_4_cmp_mReg_7, nx1728, nx1730, nx1734, nx1738, gen_4_cmp_mReg_8, 
         nx1750, nx1752, nx1756, nx1760, gen_4_cmp_mReg_9, nx1772, nx1774, 
         nx1778, nx1782, gen_4_cmp_mReg_10, nx1794, nx1796, nx1800, nx1804, 
         gen_4_cmp_mReg_11, nx1816, nx1818, nx1822, nx1826, gen_4_cmp_mReg_12, 
         nx1838, nx1840, nx1844, nx1848, gen_4_cmp_mReg_13, nx1860, nx1862, 
         nx1866, nx1870, gen_4_cmp_mReg_14, nx1882, nx1884, nx1888, nx1892, 
         gen_4_cmp_mReg_15, nx1904, nx1906, nx1910, nx1914, nx1920, nx1924, 
         nx1936, gen_5_cmp_mReg_0, nx1956, nx1964, gen_5_cmp_mReg_1, nx1976, 
         nx1978, nx1988, nx1992, gen_5_cmp_mReg_2, nx2004, nx2006, nx2010, 
         nx2014, gen_5_cmp_mReg_3, nx2026, nx2028, nx2032, nx2036, 
         gen_5_cmp_mReg_4, nx2048, nx2050, nx2054, nx2058, gen_5_cmp_mReg_5, 
         nx2070, nx2072, nx2076, nx2080, gen_5_cmp_mReg_6, nx2092, nx2094, 
         nx2098, nx2102, gen_5_cmp_mReg_7, nx2114, nx2116, nx2120, nx2124, 
         gen_5_cmp_mReg_8, nx2136, nx2138, nx2142, nx2146, gen_5_cmp_mReg_9, 
         nx2158, nx2160, nx2164, nx2168, gen_5_cmp_mReg_10, nx2180, nx2182, 
         nx2186, nx2190, gen_5_cmp_mReg_11, nx2202, nx2204, nx2208, nx2212, 
         gen_5_cmp_mReg_12, nx2224, nx2226, nx2230, nx2234, gen_5_cmp_mReg_13, 
         nx2246, nx2248, nx2252, nx2256, gen_5_cmp_mReg_14, nx2268, nx2270, 
         nx2274, nx2278, gen_5_cmp_mReg_15, nx2290, nx2292, nx2296, nx2300, 
         nx2306, nx2310, nx2322, gen_6_cmp_mReg_0, nx2342, nx2350, 
         gen_6_cmp_mReg_1, nx2362, nx2364, nx2374, nx2378, gen_6_cmp_mReg_2, 
         nx2390, nx2392, nx2396, nx2400, gen_6_cmp_mReg_3, nx2412, nx2414, 
         nx2418, nx2422, gen_6_cmp_mReg_4, nx2434, nx2436, nx2440, nx2444, 
         gen_6_cmp_mReg_5, nx2456, nx2458, nx2462, nx2466, gen_6_cmp_mReg_6, 
         nx2478, nx2480, nx2484, nx2488, gen_6_cmp_mReg_7, nx2500, nx2502, 
         nx2506, nx2510, gen_6_cmp_mReg_8, nx2522, nx2524, nx2528, nx2532, 
         gen_6_cmp_mReg_9, nx2544, nx2546, nx2550, nx2554, gen_6_cmp_mReg_10, 
         nx2566, nx2568, nx2572, nx2576, gen_6_cmp_mReg_11, nx2588, nx2590, 
         nx2594, nx2598, gen_6_cmp_mReg_12, nx2610, nx2612, nx2616, nx2620, 
         gen_6_cmp_mReg_13, nx2632, nx2634, nx2638, nx2642, gen_6_cmp_mReg_14, 
         nx2654, nx2656, nx2660, nx2664, gen_6_cmp_mReg_15, nx2676, nx2678, 
         nx2682, nx2686, nx2692, nx2696, nx2708, gen_7_cmp_mReg_0, nx2728, 
         nx2736, gen_7_cmp_mReg_1, nx2748, nx2750, nx2760, nx2764, 
         gen_7_cmp_mReg_2, nx2776, nx2778, nx2782, nx2786, gen_7_cmp_mReg_3, 
         nx2798, nx2800, nx2804, nx2808, gen_7_cmp_mReg_4, nx2820, nx2822, 
         nx2826, nx2830, gen_7_cmp_mReg_5, nx2842, nx2844, nx2848, nx2852, 
         gen_7_cmp_mReg_6, nx2864, nx2866, nx2870, nx2874, gen_7_cmp_mReg_7, 
         nx2886, nx2888, nx2892, nx2896, gen_7_cmp_mReg_8, nx2908, nx2910, 
         nx2914, nx2918, gen_7_cmp_mReg_9, nx2930, nx2932, nx2936, nx2940, 
         gen_7_cmp_mReg_10, nx2952, nx2954, nx2958, nx2962, gen_7_cmp_mReg_11, 
         nx2974, nx2976, nx2980, nx2984, gen_7_cmp_mReg_12, nx2996, nx2998, 
         nx3002, nx3006, gen_7_cmp_mReg_13, nx3018, nx3020, nx3024, nx3028, 
         gen_7_cmp_mReg_14, nx3040, nx3042, nx3046, nx3050, gen_7_cmp_mReg_15, 
         nx3062, nx3064, nx3068, nx3072, nx3078, nx3082, nx3094, 
         gen_8_cmp_mReg_0, nx3114, nx3122, gen_8_cmp_mReg_1, nx3134, nx3136, 
         nx3146, nx3150, gen_8_cmp_mReg_2, nx3162, nx3164, nx3168, nx3172, 
         gen_8_cmp_mReg_3, nx3184, nx3186, nx3190, nx3194, gen_8_cmp_mReg_4, 
         nx3206, nx3208, nx3212, nx3216, gen_8_cmp_mReg_5, nx3228, nx3230, 
         nx3234, nx3238, gen_8_cmp_mReg_6, nx3250, nx3252, nx3256, nx3260, 
         gen_8_cmp_mReg_7, nx3272, nx3274, nx3278, nx3282, gen_8_cmp_mReg_8, 
         nx3294, nx3296, nx3300, nx3304, gen_8_cmp_mReg_9, nx3316, nx3318, 
         nx3322, nx3326, gen_8_cmp_mReg_10, nx3338, nx3340, nx3344, nx3348, 
         gen_8_cmp_mReg_11, nx3360, nx3362, nx3366, nx3370, gen_8_cmp_mReg_12, 
         nx3382, nx3384, nx3388, nx3392, gen_8_cmp_mReg_13, nx3404, nx3406, 
         nx3410, nx3414, gen_8_cmp_mReg_14, nx3426, nx3428, nx3432, nx3436, 
         gen_8_cmp_mReg_15, nx3448, nx3450, nx3454, nx3458, nx3464, nx3468, 
         nx3480, gen_9_cmp_mReg_0, nx3500, nx3508, gen_9_cmp_mReg_1, nx3520, 
         nx3522, nx3532, nx3536, gen_9_cmp_mReg_2, nx3548, nx3550, nx3554, 
         nx3558, gen_9_cmp_mReg_3, nx3570, nx3572, nx3576, nx3580, 
         gen_9_cmp_mReg_4, nx3592, nx3594, nx3598, nx3602, gen_9_cmp_mReg_5, 
         nx3614, nx3616, nx3620, nx3624, gen_9_cmp_mReg_6, nx3636, nx3638, 
         nx3642, nx3646, gen_9_cmp_mReg_7, nx3658, nx3660, nx3664, nx3668, 
         gen_9_cmp_mReg_8, nx3680, nx3682, nx3686, nx3690, gen_9_cmp_mReg_9, 
         nx3702, nx3704, nx3708, nx3712, gen_9_cmp_mReg_10, nx3724, nx3726, 
         nx3730, nx3734, gen_9_cmp_mReg_11, nx3746, nx3748, nx3752, nx3756, 
         gen_9_cmp_mReg_12, nx3768, nx3770, nx3774, nx3778, gen_9_cmp_mReg_13, 
         nx3790, nx3792, nx3796, nx3800, gen_9_cmp_mReg_14, nx3812, nx3814, 
         nx3818, nx3822, gen_9_cmp_mReg_15, nx3834, nx3836, nx3840, nx3844, 
         nx3850, nx3854, nx3866, gen_10_cmp_mReg_0, nx3886, nx3894, 
         gen_10_cmp_mReg_1, nx3906, nx3908, nx3918, nx3922, gen_10_cmp_mReg_2, 
         nx3934, nx3936, nx3940, nx3944, gen_10_cmp_mReg_3, nx3956, nx3958, 
         nx3962, nx3966, gen_10_cmp_mReg_4, nx3978, nx3980, nx3984, nx3988, 
         gen_10_cmp_mReg_5, nx4000, nx4002, nx4006, nx4010, gen_10_cmp_mReg_6, 
         nx4022, nx4024, nx4028, nx4032, gen_10_cmp_mReg_7, nx4044, nx4046, 
         nx4050, nx4054, gen_10_cmp_mReg_8, nx4066, nx4068, nx4072, nx4076, 
         gen_10_cmp_mReg_9, nx4088, nx4090, nx4094, nx4098, gen_10_cmp_mReg_10, 
         nx4110, nx4112, nx4116, nx4120, gen_10_cmp_mReg_11, nx4132, nx4134, 
         nx4138, nx4142, gen_10_cmp_mReg_12, nx4154, nx4156, nx4160, nx4164, 
         gen_10_cmp_mReg_13, nx4176, nx4178, nx4182, nx4186, gen_10_cmp_mReg_14, 
         nx4198, nx4200, nx4204, nx4208, gen_10_cmp_mReg_15, nx4220, nx4222, 
         nx4226, nx4230, nx4236, nx4240, nx4252, gen_11_cmp_mReg_0, nx4272, 
         nx4280, gen_11_cmp_mReg_1, nx4292, nx4294, nx4304, nx4308, 
         gen_11_cmp_mReg_2, nx4320, nx4322, nx4326, nx4330, gen_11_cmp_mReg_3, 
         nx4342, nx4344, nx4348, nx4352, gen_11_cmp_mReg_4, nx4364, nx4366, 
         nx4370, nx4374, gen_11_cmp_mReg_5, nx4386, nx4388, nx4392, nx4396, 
         gen_11_cmp_mReg_6, nx4408, nx4410, nx4414, nx4418, gen_11_cmp_mReg_7, 
         nx4430, nx4432, nx4436, nx4440, gen_11_cmp_mReg_8, nx4452, nx4454, 
         nx4458, nx4462, gen_11_cmp_mReg_9, nx4474, nx4476, nx4480, nx4484, 
         gen_11_cmp_mReg_10, nx4496, nx4498, nx4502, nx4506, gen_11_cmp_mReg_11, 
         nx4518, nx4520, nx4524, nx4528, gen_11_cmp_mReg_12, nx4540, nx4542, 
         nx4546, nx4550, gen_11_cmp_mReg_13, nx4562, nx4564, nx4568, nx4572, 
         gen_11_cmp_mReg_14, nx4584, nx4586, nx4590, nx4594, gen_11_cmp_mReg_15, 
         nx4606, nx4608, nx4612, nx4616, nx4622, nx4626, nx4638, 
         gen_12_cmp_mReg_0, nx4658, nx4666, gen_12_cmp_mReg_1, nx4678, nx4680, 
         nx4690, nx4694, gen_12_cmp_mReg_2, nx4706, nx4708, nx4712, nx4716, 
         gen_12_cmp_mReg_3, nx4728, nx4730, nx4734, nx4738, gen_12_cmp_mReg_4, 
         nx4750, nx4752, nx4756, nx4760, gen_12_cmp_mReg_5, nx4772, nx4774, 
         nx4778, nx4782, gen_12_cmp_mReg_6, nx4794, nx4796, nx4800, nx4804, 
         gen_12_cmp_mReg_7, nx4816, nx4818, nx4822, nx4826, gen_12_cmp_mReg_8, 
         nx4838, nx4840, nx4844, nx4848, gen_12_cmp_mReg_9, nx4860, nx4862, 
         nx4866, nx4870, gen_12_cmp_mReg_10, nx4882, nx4884, nx4888, nx4892, 
         gen_12_cmp_mReg_11, nx4904, nx4906, nx4910, nx4914, gen_12_cmp_mReg_12, 
         nx4926, nx4928, nx4932, nx4936, gen_12_cmp_mReg_13, nx4948, nx4950, 
         nx4954, nx4958, gen_12_cmp_mReg_14, nx4970, nx4972, nx4976, nx4980, 
         gen_12_cmp_mReg_15, nx4992, nx4994, nx4998, nx5002, nx5008, nx5012, 
         nx5024, gen_13_cmp_mReg_0, nx5044, nx5052, gen_13_cmp_mReg_1, nx5064, 
         nx5066, nx5076, nx5080, gen_13_cmp_mReg_2, nx5092, nx5094, nx5098, 
         nx5102, gen_13_cmp_mReg_3, nx5114, nx5116, nx5120, nx5124, 
         gen_13_cmp_mReg_4, nx5136, nx5138, nx5142, nx5146, gen_13_cmp_mReg_5, 
         nx5158, nx5160, nx5164, nx5168, gen_13_cmp_mReg_6, nx5180, nx5182, 
         nx5186, nx5190, gen_13_cmp_mReg_7, nx5202, nx5204, nx5208, nx5212, 
         gen_13_cmp_mReg_8, nx5224, nx5226, nx5230, nx5234, gen_13_cmp_mReg_9, 
         nx5246, nx5248, nx5252, nx5256, gen_13_cmp_mReg_10, nx5268, nx5270, 
         nx5274, nx5278, gen_13_cmp_mReg_11, nx5290, nx5292, nx5296, nx5300, 
         gen_13_cmp_mReg_12, nx5312, nx5314, nx5318, nx5322, gen_13_cmp_mReg_13, 
         nx5334, nx5336, nx5340, nx5344, gen_13_cmp_mReg_14, nx5356, nx5358, 
         nx5362, nx5366, gen_13_cmp_mReg_15, nx5378, nx5380, nx5384, nx5388, 
         nx5394, nx5398, nx5410, gen_14_cmp_mReg_0, nx5430, nx5438, 
         gen_14_cmp_mReg_1, nx5450, nx5452, nx5462, nx5466, gen_14_cmp_mReg_2, 
         nx5478, nx5480, nx5484, nx5488, gen_14_cmp_mReg_3, nx5500, nx5502, 
         nx5506, nx5510, gen_14_cmp_mReg_4, nx5522, nx5524, nx5528, nx5532, 
         gen_14_cmp_mReg_5, nx5544, nx5546, nx5550, nx5554, gen_14_cmp_mReg_6, 
         nx5566, nx5568, nx5572, nx5576, gen_14_cmp_mReg_7, nx5588, nx5590, 
         nx5594, nx5598, gen_14_cmp_mReg_8, nx5610, nx5612, nx5616, nx5620, 
         gen_14_cmp_mReg_9, nx5632, nx5634, nx5638, nx5642, gen_14_cmp_mReg_10, 
         nx5654, nx5656, nx5660, nx5664, gen_14_cmp_mReg_11, nx5676, nx5678, 
         nx5682, nx5686, gen_14_cmp_mReg_12, nx5698, nx5700, nx5704, nx5708, 
         gen_14_cmp_mReg_13, nx5720, nx5722, nx5726, nx5730, gen_14_cmp_mReg_14, 
         nx5742, nx5744, nx5748, nx5752, gen_14_cmp_mReg_15, nx5764, nx5766, 
         nx5770, nx5774, nx5780, nx5784, nx5796, gen_15_cmp_mReg_0, nx5816, 
         nx5824, gen_15_cmp_mReg_1, nx5836, nx5838, nx5848, nx5852, 
         gen_15_cmp_mReg_2, nx5864, nx5866, nx5870, nx5874, gen_15_cmp_mReg_3, 
         nx5886, nx5888, nx5892, nx5896, gen_15_cmp_mReg_4, nx5908, nx5910, 
         nx5914, nx5918, gen_15_cmp_mReg_5, nx5930, nx5932, nx5936, nx5940, 
         gen_15_cmp_mReg_6, nx5952, nx5954, nx5958, nx5962, gen_15_cmp_mReg_7, 
         nx5974, nx5976, nx5980, nx5984, gen_15_cmp_mReg_8, nx5996, nx5998, 
         nx6002, nx6006, gen_15_cmp_mReg_9, nx6018, nx6020, nx6024, nx6028, 
         gen_15_cmp_mReg_10, nx6040, nx6042, nx6046, nx6050, gen_15_cmp_mReg_11, 
         nx6062, nx6064, nx6068, nx6072, gen_15_cmp_mReg_12, nx6084, nx6086, 
         nx6090, nx6094, gen_15_cmp_mReg_13, nx6106, nx6108, nx6112, nx6116, 
         gen_15_cmp_mReg_14, nx6128, nx6130, nx6134, nx6138, gen_15_cmp_mReg_15, 
         nx6150, nx6152, nx6156, nx6160, nx6166, nx6170, nx6182, 
         gen_16_cmp_mReg_0, nx6202, nx6210, gen_16_cmp_mReg_1, nx6222, nx6224, 
         nx6234, nx6238, gen_16_cmp_mReg_2, nx6250, nx6252, nx6256, nx6260, 
         gen_16_cmp_mReg_3, nx6272, nx6274, nx6278, nx6282, gen_16_cmp_mReg_4, 
         nx6294, nx6296, nx6300, nx6304, gen_16_cmp_mReg_5, nx6316, nx6318, 
         nx6322, nx6326, gen_16_cmp_mReg_6, nx6338, nx6340, nx6344, nx6348, 
         gen_16_cmp_mReg_7, nx6360, nx6362, nx6366, nx6370, gen_16_cmp_mReg_8, 
         nx6382, nx6384, nx6388, nx6392, gen_16_cmp_mReg_9, nx6404, nx6406, 
         nx6410, nx6414, gen_16_cmp_mReg_10, nx6426, nx6428, nx6432, nx6436, 
         gen_16_cmp_mReg_11, nx6448, nx6450, nx6454, nx6458, gen_16_cmp_mReg_12, 
         nx6470, nx6472, nx6476, nx6480, gen_16_cmp_mReg_13, nx6492, nx6494, 
         nx6498, nx6502, gen_16_cmp_mReg_14, nx6514, nx6516, nx6520, nx6524, 
         gen_16_cmp_mReg_15, nx6536, nx6538, nx6542, nx6546, nx6552, nx6556, 
         nx6568, gen_17_cmp_mReg_0, nx6588, nx6596, gen_17_cmp_mReg_1, nx6608, 
         nx6610, nx6620, nx6624, gen_17_cmp_mReg_2, nx6636, nx6638, nx6642, 
         nx6646, gen_17_cmp_mReg_3, nx6658, nx6660, nx6664, nx6668, 
         gen_17_cmp_mReg_4, nx6680, nx6682, nx6686, nx6690, gen_17_cmp_mReg_5, 
         nx6702, nx6704, nx6708, nx6712, gen_17_cmp_mReg_6, nx6724, nx6726, 
         nx6730, nx6734, gen_17_cmp_mReg_7, nx6746, nx6748, nx6752, nx6756, 
         gen_17_cmp_mReg_8, nx6768, nx6770, nx6774, nx6778, gen_17_cmp_mReg_9, 
         nx6790, nx6792, nx6796, nx6800, gen_17_cmp_mReg_10, nx6812, nx6814, 
         nx6818, nx6822, gen_17_cmp_mReg_11, nx6834, nx6836, nx6840, nx6844, 
         gen_17_cmp_mReg_12, nx6856, nx6858, nx6862, nx6866, gen_17_cmp_mReg_13, 
         nx6878, nx6880, nx6884, nx6888, gen_17_cmp_mReg_14, nx6900, nx6902, 
         nx6906, nx6910, gen_17_cmp_mReg_15, nx6922, nx6924, nx6928, nx6932, 
         nx6938, nx6942, nx6954, gen_18_cmp_mReg_0, nx6974, nx6982, 
         gen_18_cmp_mReg_1, nx6994, nx6996, nx7006, nx7010, gen_18_cmp_mReg_2, 
         nx7022, nx7024, nx7028, nx7032, gen_18_cmp_mReg_3, nx7044, nx7046, 
         nx7050, nx7054, gen_18_cmp_mReg_4, nx7066, nx7068, nx7072, nx7076, 
         gen_18_cmp_mReg_5, nx7088, nx7090, nx7094, nx7098, gen_18_cmp_mReg_6, 
         nx7110, nx7112, nx7116, nx7120, gen_18_cmp_mReg_7, nx7132, nx7134, 
         nx7138, nx7142, gen_18_cmp_mReg_8, nx7154, nx7156, nx7160, nx7164, 
         gen_18_cmp_mReg_9, nx7176, nx7178, nx7182, nx7186, gen_18_cmp_mReg_10, 
         nx7198, nx7200, nx7204, nx7208, gen_18_cmp_mReg_11, nx7220, nx7222, 
         nx7226, nx7230, gen_18_cmp_mReg_12, nx7242, nx7244, nx7248, nx7252, 
         gen_18_cmp_mReg_13, nx7264, nx7266, nx7270, nx7274, gen_18_cmp_mReg_14, 
         nx7286, nx7288, nx7292, nx7296, gen_18_cmp_mReg_15, nx7308, nx7310, 
         nx7314, nx7318, nx7324, nx7328, nx7340, gen_19_cmp_mReg_0, nx7360, 
         nx7368, gen_19_cmp_mReg_1, nx7380, nx7382, nx7392, nx7396, 
         gen_19_cmp_mReg_2, nx7408, nx7410, nx7414, nx7418, gen_19_cmp_mReg_3, 
         nx7430, nx7432, nx7436, nx7440, gen_19_cmp_mReg_4, nx7452, nx7454, 
         nx7458, nx7462, gen_19_cmp_mReg_5, nx7474, nx7476, nx7480, nx7484, 
         gen_19_cmp_mReg_6, nx7496, nx7498, nx7502, nx7506, gen_19_cmp_mReg_7, 
         nx7518, nx7520, nx7524, nx7528, gen_19_cmp_mReg_8, nx7540, nx7542, 
         nx7546, nx7550, gen_19_cmp_mReg_9, nx7562, nx7564, nx7568, nx7572, 
         gen_19_cmp_mReg_10, nx7584, nx7586, nx7590, nx7594, gen_19_cmp_mReg_11, 
         nx7606, nx7608, nx7612, nx7616, gen_19_cmp_mReg_12, nx7628, nx7630, 
         nx7634, nx7638, gen_19_cmp_mReg_13, nx7650, nx7652, nx7656, nx7660, 
         gen_19_cmp_mReg_14, nx7672, nx7674, nx7678, nx7682, gen_19_cmp_mReg_15, 
         nx7694, nx7696, nx7700, nx7704, nx7710, nx7714, nx7726, 
         gen_20_cmp_mReg_0, nx7746, nx7754, gen_20_cmp_mReg_1, nx7766, nx7768, 
         nx7778, nx7782, gen_20_cmp_mReg_2, nx7794, nx7796, nx7800, nx7804, 
         gen_20_cmp_mReg_3, nx7816, nx7818, nx7822, nx7826, gen_20_cmp_mReg_4, 
         nx7838, nx7840, nx7844, nx7848, gen_20_cmp_mReg_5, nx7860, nx7862, 
         nx7866, nx7870, gen_20_cmp_mReg_6, nx7882, nx7884, nx7888, nx7892, 
         gen_20_cmp_mReg_7, nx7904, nx7906, nx7910, nx7914, gen_20_cmp_mReg_8, 
         nx7926, nx7928, nx7932, nx7936, gen_20_cmp_mReg_9, nx7948, nx7950, 
         nx7954, nx7958, gen_20_cmp_mReg_10, nx7970, nx7972, nx7976, nx7980, 
         gen_20_cmp_mReg_11, nx7992, nx7994, nx7998, nx8002, gen_20_cmp_mReg_12, 
         nx8014, nx8016, nx8020, nx8024, gen_20_cmp_mReg_13, nx8036, nx8038, 
         nx8042, nx8046, gen_20_cmp_mReg_14, nx8058, nx8060, nx8064, nx8068, 
         gen_20_cmp_mReg_15, nx8080, nx8082, nx8086, nx8090, nx8096, nx8100, 
         nx8112, gen_21_cmp_mReg_0, nx8132, nx8140, gen_21_cmp_mReg_1, nx8152, 
         nx8154, nx8164, nx8168, gen_21_cmp_mReg_2, nx8180, nx8182, nx8186, 
         nx8190, gen_21_cmp_mReg_3, nx8202, nx8204, nx8208, nx8212, 
         gen_21_cmp_mReg_4, nx8224, nx8226, nx8230, nx8234, gen_21_cmp_mReg_5, 
         nx8246, nx8248, nx8252, nx8256, gen_21_cmp_mReg_6, nx8268, nx8270, 
         nx8274, nx8278, gen_21_cmp_mReg_7, nx8290, nx8292, nx8296, nx8300, 
         gen_21_cmp_mReg_8, nx8312, nx8314, nx8318, nx8322, gen_21_cmp_mReg_9, 
         nx8334, nx8336, nx8340, nx8344, gen_21_cmp_mReg_10, nx8356, nx8358, 
         nx8362, nx8366, gen_21_cmp_mReg_11, nx8378, nx8380, nx8384, nx8388, 
         gen_21_cmp_mReg_12, nx8400, nx8402, nx8406, nx8410, gen_21_cmp_mReg_13, 
         nx8422, nx8424, nx8428, nx8432, gen_21_cmp_mReg_14, nx8444, nx8446, 
         nx8450, nx8454, gen_21_cmp_mReg_15, nx8466, nx8468, nx8472, nx8476, 
         nx8482, nx8486, nx8498, gen_22_cmp_mReg_0, nx8518, nx8526, 
         gen_22_cmp_mReg_1, nx8538, nx8540, nx8550, nx8554, gen_22_cmp_mReg_2, 
         nx8566, nx8568, nx8572, nx8576, gen_22_cmp_mReg_3, nx8588, nx8590, 
         nx8594, nx8598, gen_22_cmp_mReg_4, nx8610, nx8612, nx8616, nx8620, 
         gen_22_cmp_mReg_5, nx8632, nx8634, nx8638, nx8642, gen_22_cmp_mReg_6, 
         nx8654, nx8656, nx8660, nx8664, gen_22_cmp_mReg_7, nx8676, nx8678, 
         nx8682, nx8686, gen_22_cmp_mReg_8, nx8698, nx8700, nx8704, nx8708, 
         gen_22_cmp_mReg_9, nx8720, nx8722, nx8726, nx8730, gen_22_cmp_mReg_10, 
         nx8742, nx8744, nx8748, nx8752, gen_22_cmp_mReg_11, nx8764, nx8766, 
         nx8770, nx8774, gen_22_cmp_mReg_12, nx8786, nx8788, nx8792, nx8796, 
         gen_22_cmp_mReg_13, nx8808, nx8810, nx8814, nx8818, gen_22_cmp_mReg_14, 
         nx8830, nx8832, nx8836, nx8840, gen_22_cmp_mReg_15, nx8852, nx8854, 
         nx8858, nx8862, nx8868, nx8872, nx8884, gen_23_cmp_mReg_0, nx8904, 
         nx8912, gen_23_cmp_mReg_1, nx8924, nx8926, nx8936, nx8940, 
         gen_23_cmp_mReg_2, nx8952, nx8954, nx8958, nx8962, gen_23_cmp_mReg_3, 
         nx8974, nx8976, nx8980, nx8984, gen_23_cmp_mReg_4, nx8996, nx8998, 
         nx9002, nx9006, gen_23_cmp_mReg_5, nx9018, nx9020, nx9024, nx9028, 
         gen_23_cmp_mReg_6, nx9040, nx9042, nx9046, nx9050, gen_23_cmp_mReg_7, 
         nx9062, nx9064, nx9068, nx9072, gen_23_cmp_mReg_8, nx9084, nx9086, 
         nx9090, nx9094, gen_23_cmp_mReg_9, nx9106, nx9108, nx9112, nx9116, 
         gen_23_cmp_mReg_10, nx9128, nx9130, nx9134, nx9138, gen_23_cmp_mReg_11, 
         nx9150, nx9152, nx9156, nx9160, gen_23_cmp_mReg_12, nx9172, nx9174, 
         nx9178, nx9182, gen_23_cmp_mReg_13, nx9194, nx9196, nx9200, nx9204, 
         gen_23_cmp_mReg_14, nx9216, nx9218, nx9222, nx9226, gen_23_cmp_mReg_15, 
         nx9238, nx9240, nx9244, nx9248, nx9254, nx9258, nx9270, 
         gen_24_cmp_mReg_0, nx9290, nx9298, gen_24_cmp_mReg_1, nx9310, nx9312, 
         nx9322, nx9326, gen_24_cmp_mReg_2, nx9338, nx9340, nx9344, nx9348, 
         gen_24_cmp_mReg_3, nx9360, nx9362, nx9366, nx9370, gen_24_cmp_mReg_4, 
         nx9382, nx9384, nx9388, nx9392, gen_24_cmp_mReg_5, nx9404, nx9406, 
         nx9410, nx9414, gen_24_cmp_mReg_6, nx9426, nx9428, nx9432, nx9436, 
         gen_24_cmp_mReg_7, nx9448, nx9450, nx9454, nx9458, gen_24_cmp_mReg_8, 
         nx9470, nx9472, nx9476, nx9480, gen_24_cmp_mReg_9, nx9492, nx9494, 
         nx9498, nx9502, gen_24_cmp_mReg_10, nx9514, nx9516, nx9520, nx9524, 
         gen_24_cmp_mReg_11, nx9536, nx9538, nx9542, nx9546, gen_24_cmp_mReg_12, 
         nx9558, nx9560, nx9564, nx9568, gen_24_cmp_mReg_13, nx9580, nx9582, 
         nx9586, nx9590, gen_24_cmp_mReg_14, nx9602, nx9604, nx9608, nx9612, 
         gen_24_cmp_mReg_15, nx9624, nx9626, nx9630, nx9634, nx9640, nx9644, 
         nx9650, restartDetection, StartCaptuerCmp_d, nx9664, nx9670, nx2813, 
         nx2823, nx2833, nx2839, nx2853, nx2859, nx2862, nx2871, nx2873, nx2877, 
         nx2887, nx2893, nx2897, nx2903, nx2907, nx2911, nx2917, nx2923, nx2926, 
         nx2931, nx2937, nx2941, nx2947, nx2951, nx2955, nx2961, nx2967, nx2970, 
         nx2975, nx2981, nx2985, nx2991, nx2995, nx2999, nx3005, nx3011, nx3014, 
         nx3019, nx3025, nx3029, nx3035, nx3039, nx3043, nx3049, nx3055, nx3058, 
         nx3063, nx3069, nx3073, nx3079, nx3083, nx3087, nx3093, nx3099, nx3103, 
         nx3107, nx3115, nx3117, nx3121, nx3132, nx3139, nx3143, nx3149, nx3155, 
         nx3158, nx3163, nx3169, nx3173, nx3179, nx3183, nx3187, nx3193, nx3199, 
         nx3202, nx3207, nx3213, nx3217, nx3223, nx3227, nx3231, nx3237, nx3243, 
         nx3246, nx3251, nx3257, nx3261, nx3267, nx3271, nx3275, nx3281, nx3287, 
         nx3290, nx3295, nx3301, nx3305, nx3311, nx3315, nx3319, nx3325, nx3331, 
         nx3334, nx3339, nx3347, nx3353, nx3356, nx3363, nx3365, nx3369, nx3380, 
         nx3387, nx3391, nx3397, nx3401, nx3405, nx3411, nx3415, nx3419, nx3423, 
         nx3429, nx3433, nx3437, nx3443, nx3446, nx3453, nx3459, nx3463, nx3469, 
         nx3475, nx3479, nx3484, nx3488, nx3491, nx3497, nx3503, nx3507, nx3513, 
         nx3517, nx3521, nx3527, nx3533, nx3537, nx3543, nx3547, nx3551, nx3557, 
         nx3563, nx3566, nx3571, nx3577, nx3581, nx3587, nx3593, nx3599, nx3603, 
         nx3611, nx3613, nx3617, nx3629, nx3633, nx3637, nx3643, nx3647, nx3651, 
         nx3655, nx3661, nx3665, nx3669, nx3675, nx3678, nx3685, nx3691, nx3695, 
         nx3699, nx3705, nx3709, nx3713, nx3719, nx3722, nx3729, nx3735, nx3739, 
         nx3743, nx3749, nx3753, nx3757, nx3763, nx3766, nx3773, nx3779, nx3783, 
         nx3787, nx3793, nx3797, nx3801, nx3807, nx3810, nx3817, nx3823, nx3827, 
         nx3831, nx3839, nx3845, nx3849, nx3857, nx3859, nx3863, nx3873, nx3877, 
         nx3881, nx3887, nx3893, nx3897, nx3902, nx3907, nx3911, nx3915, nx3921, 
         nx3925, nx3930, nx3935, nx3939, nx3945, nx3951, nx3954, nx3961, nx3967, 
         nx3971, nx3975, nx3981, nx3985, nx3989, nx3995, nx3998, nx4005, nx4011, 
         nx4015, nx4019, nx4025, nx4029, nx4033, nx4039, nx4042, nx4049, nx4055, 
         nx4059, nx4063, nx4069, nx4073, nx4077, nx4084, nx4089, nx4093, nx4101, 
         nx4103, nx4106, nx4119, nx4125, nx4128, nx4133, nx4139, nx4143, nx4149, 
         nx4153, nx4157, nx4163, nx4169, nx4172, nx4177, nx4183, nx4187, nx4193, 
         nx4197, nx4201, nx4207, nx4213, nx4216, nx4221, nx4227, nx4231, nx4237, 
         nx4241, nx4245, nx4251, nx4256, nx4259, nx4263, nx4269, nx4273, nx4279, 
         nx4285, nx4288, nx4293, nx4299, nx4303, nx4309, nx4315, nx4318, nx4325, 
         nx4331, nx4337, nx4340, nx4349, nx4351, nx4355, nx4365, nx4371, nx4375, 
         nx4381, nx4385, nx4389, nx4395, nx4401, nx4404, nx4409, nx4415, nx4419, 
         nx4425, nx4429, nx4433, nx4439, nx4445, nx4448, nx4453, nx4459, nx4463, 
         nx4469, nx4473, nx4477, nx4483, nx4489, nx4492, nx4497, nx4503, nx4507, 
         nx4513, nx4517, nx4521, nx4527, nx4533, nx4536, nx4541, nx4547, nx4551, 
         nx4557, nx4561, nx4565, nx4571, nx4579, nx4583, nx4587, nx4595, nx4597, 
         nx4601, nx4613, nx4617, nx4621, nx4627, nx4633, nx4637, nx4642, nx4646, 
         nx4649, nx4655, nx4661, nx4665, nx4671, nx4675, nx4679, nx4685, nx4691, 
         nx4695, nx4701, nx4705, nx4709, nx4715, nx4721, nx4724, nx4729, nx4735, 
         nx4739, nx4745, nx4749, nx4753, nx4759, nx4765, nx4768, nx4773, nx4779, 
         nx4783, nx4789, nx4793, nx4797, nx4803, nx4809, nx4812, nx4817, nx4825, 
         nx4831, nx4834, nx4841, nx4843, nx4847, nx4858, nx4865, nx4869, nx4875, 
         nx4879, nx4883, nx4889, nx4893, nx4897, nx4901, nx4907, nx4911, nx4915, 
         nx4921, nx4924, nx4931, nx4937, nx4941, nx4945, nx4951, nx4955, nx4959, 
         nx4965, nx4968, nx4975, nx4981, nx4985, nx4989, nx4995, nx4999, nx5003, 
         nx5009, nx5013, nx5019, nx5025, nx5028, nx5032, nx5037, nx5041, nx5047, 
         nx5053, nx5057, nx5061, nx5069, nx5073, nx5077, nx5085, nx5087, nx5090, 
         nx5103, nx5109, nx5112, nx5119, nx5125, nx5129, nx5133, nx5139, nx5143, 
         nx5147, nx5153, nx5156, nx5163, nx5169, nx5173, nx5177, nx5183, nx5187, 
         nx5191, nx5197, nx5200, nx5207, nx5213, nx5217, nx5221, nx5227, nx5231, 
         nx5235, nx5241, nx5244, nx5251, nx5257, nx5261, nx5265, nx5271, nx5275, 
         nx5279, nx5285, nx5288, nx5295, nx5301, nx5305, nx5309, nx5317, nx5323, 
         nx5327, nx5335, nx5337, nx5341, nx5352, nx5357, nx5361, nx5367, nx5373, 
         nx5376, nx5383, nx5389, nx5393, nx5399, nx5405, nx5409, nx5414, nx5418, 
         nx5421, nx5427, nx5433, nx5437, nx5443, nx5447, nx5451, nx5457, nx5463, 
         nx5467, nx5473, nx5477, nx5481, nx5487, nx5493, nx5496, nx5501, nx5507, 
         nx5511, nx5517, nx5521, nx5525, nx5531, nx5537, nx5540, nx5545, nx5551, 
         nx5555, nx5561, nx5567, nx5573, nx5577, nx5585, nx5587, nx5591, nx5603, 
         nx5607, nx5611, nx5617, nx5621, nx5625, nx5629, nx5635, nx5639, nx5643, 
         nx5649, nx5652, nx5659, nx5665, nx5669, nx5673, nx5679, nx5683, nx5687, 
         nx5693, nx5696, nx5703, nx5709, nx5713, nx5717, nx5723, nx5727, nx5731, 
         nx5737, nx5740, nx5747, nx5753, nx5757, nx5761, nx5767, nx5771, nx5775, 
         nx5781, nx5785, nx5791, nx5797, nx5800, nx5804, nx5811, nx5817, nx5821, 
         nx5829, nx5831, nx5834, nx5847, nx5853, nx5857, nx5861, nx5867, nx5871, 
         nx5875, nx5881, nx5884, nx5891, nx5897, nx5901, nx5905, nx5911, nx5915, 
         nx5919, nx5925, nx5928, nx5935, nx5941, nx5945, nx5949, nx5955, nx5959, 
         nx5963, nx5969, nx5972, nx5979, nx5985, nx5989, nx5993, nx5999, nx6003, 
         nx6007, nx6013, nx6016, nx6023, nx6029, nx6033, nx6037, nx6043, nx6047, 
         nx6051, nx6058, nx6063, nx6067, nx6075, nx6077, nx6080, nx6093, nx6099, 
         nx6102, nx6107, nx6113, nx6117, nx6123, nx6127, nx6131, nx6137, nx6143, 
         nx6146, nx6151, nx6157, nx6161, nx6167, nx6171, nx6175, nx6181, nx6186, 
         nx6189, nx6193, nx6199, nx6203, nx6209, nx6215, nx6218, nx6223, nx6229, 
         nx6233, nx6239, nx6245, nx6248, nx6255, nx6261, nx6265, nx6269, nx6275, 
         nx6279, nx6283, nx6289, nx6292, nx6299, nx6305, nx6311, nx6314, nx6323, 
         nx6325, nx6329, nx6339, nx6345, nx6349, nx6355, nx6359, nx6363, nx6369, 
         nx6375, nx6378, nx6383, nx6389, nx6393, nx6399, nx6403, nx6407, nx6413, 
         nx6419, nx6422, nx6427, nx6433, nx6437, nx6443, nx6447, nx6451, nx6457, 
         nx6463, nx6466, nx6471, nx6477, nx6481, nx6487, nx6491, nx6495, nx6501, 
         nx6507, nx6510, nx6515, nx6521, nx6525, nx6531, nx6535, nx6539, nx6545, 
         nx6553, nx6557, nx6561, nx6569, nx6571, nx6574, nx6585, nx6591, nx6595, 
         nx6601, nx6605, nx6609, nx6615, nx6621, nx6625, nx6631, nx6635, nx6639, 
         nx6645, nx6651, nx6654, nx6659, nx6665, nx6669, nx6675, nx6679, nx6683, 
         nx6689, nx6695, nx6698, nx6703, nx6709, nx6713, nx6719, nx6723, nx6727, 
         nx6733, nx6739, nx6742, nx6747, nx6753, nx6757, nx6763, nx6767, nx6771, 
         nx6777, nx6783, nx6786, nx6791, nx6799, nx6805, nx6808, nx6815, nx6817, 
         nx6821, nx6832, nx6839, nx6843, nx6849, nx6853, nx6857, nx6863, nx6867, 
         nx6871, nx6875, nx6881, nx6885, nx6889, nx6895, nx6898, nx6905, nx6911, 
         nx6915, nx6919, nx6925, nx6929, nx6933, nx6939, nx6943, nx6949, nx6955, 
         nx6958, nx6962, nx6967, nx6971, nx6977, nx6983, nx6987, nx6991, nx6997, 
         nx7001, nx7007, nx7011, nx7015, nx7019, nx7025, nx7029, nx7033, nx7040, 
         nx7045, nx7049, nx7057, nx7059, nx7062, nx7075, nx7081, nx7084, nx7089, 
         nx7095, nx7099, nx7105, nx7109, nx7113, nx7119, nx7125, nx7128, nx7133, 
         nx7139, nx7143, nx7149, nx7153, nx7157, nx7163, nx7169, nx7172, nx7177, 
         nx7183, nx7187, nx7193, nx7197, nx7201, nx7207, nx7213, nx7216, nx7221, 
         nx7227, nx7231, nx7237, nx7241, nx7245, nx7251, nx7257, nx7260, nx7265, 
         nx7271, nx7275, nx7281, nx7287, nx7293, nx7297, nx7305, nx7307, nx7311, 
         nx7323, nx7329, nx7333, nx7339, nx7344, nx7347, nx7351, nx7357, nx7361, 
         nx7367, nx7373, nx7376, nx7381, nx7387, nx7391, nx7397, nx7403, nx7406, 
         nx7413, nx7419, nx7423, nx7427, nx7433, nx7437, nx7441, nx7447, nx7450, 
         nx7457, nx7463, nx7467, nx7471, nx7477, nx7481, nx7485, nx7491, nx7494, 
         nx7501, nx7507, nx7511, nx7515, nx7521, nx7525, nx7529, nx7536, nx7541, 
         nx7545, nx7553, nx7555, nx7558, nx7571, nx7577, nx7580, nx7585, nx7591, 
         nx7595, nx7601, nx7605, nx7609, nx7615, nx7621, nx7624, nx7629, nx7635, 
         nx7639, nx7645, nx7649, nx7653, nx7659, nx7665, nx7668, nx7673, nx7679, 
         nx7683, nx7689, nx7693, nx7697, nx7703, nx7709, nx7713, nx7719, nx7725, 
         nx7729, nx7733, nx7737, nx7741, nx7747, nx7753, nx7757, nx7762, nx7767, 
         nx7771, nx7775, nx7783, nx7789, nx7792, nx7801, nx7803, nx7807, nx7817, 
         nx7823, nx7827, nx7833, nx7837, nx7841, nx7847, nx7853, nx7856, nx7861, 
         nx7867, nx7871, nx7877, nx7881, nx7885, nx7891, nx7897, nx7900, nx7905, 
         nx7911, nx7915, nx7921, nx7925, nx7929, nx7935, nx7941, nx7944, nx7949, 
         nx7955, nx7959, nx7965, nx7969, nx7973, nx7979, nx7985, nx7988, nx7993, 
         nx7999, nx8003, nx8009, nx8013, nx8017, nx8023, nx8031, nx8035, nx8039, 
         nx8047, nx8049, nx8053, nx8065, nx8069, nx8073, nx8077, nx8083, nx8087, 
         nx8091, nx8097, nx8101, nx8107, nx8113, nx8116, nx8120, nx8125, nx8129, 
         nx8135, nx8141, nx8145, nx8149, nx8155, nx8159, nx8165, nx8169, nx8173, 
         nx8177, nx8183, nx8187, nx8191, nx8197, nx8200, nx8207, nx8213, nx8217, 
         nx8221, nx8227, nx8231, nx8235, nx8241, nx8244, nx8251, nx8257, nx8261, 
         nx8265, nx8273, nx8279, nx8283, nx8291, nx8293, nx8297, nx8308, nx8313, 
         nx8317, nx8323, nx8329, nx8332, nx8339, nx8345, nx8349, nx8353, nx8359, 
         nx8363, nx8367, nx8373, nx8376, nx8383, nx8389, nx8393, nx8397, nx8403, 
         nx8407, nx8411, nx8417, nx8420, nx8427, nx8433, nx8437, nx8441, nx8447, 
         nx8451, nx8455, nx8461, nx8464, nx8471, nx8477, nx8481, nx8487, nx8493, 
         nx8497, nx8502, nx8506, nx8509, nx8515, nx8523, nx8529, nx8533, nx8541, 
         nx8543, nx8547, nx8559, nx8563, nx8567, nx8573, nx8577, nx8581, nx8585, 
         nx8591, nx8595, nx8599, nx8605, nx8608, nx8615, nx8621, nx8625, nx8629, 
         nx8635, nx8639, nx8643, nx8649, nx8652, nx8659, nx8665, nx8669, nx8673, 
         nx8679, nx8683, nx8687, nx8693, nx8696, nx8703, nx8709, nx8713, nx8717, 
         nx8723, nx8727, nx8731, nx8737, nx8740, nx8747, nx8753, nx8757, nx8761, 
         nx8769, nx8775, nx8779, nx8787, nx8789, nx8793, nx8804, nx8809, nx8813, 
         nx8819, nx8825, nx8828, nx8835, nx8841, nx8845, nx8849, nx8855, nx8859, 
         nx8863, nx8869, nx8873, nx8879, nx8885, nx8888, nx8892, nx8897, nx8901, 
         nx8907, nx8913, nx8917, nx8921, nx8927, nx8931, nx8937, nx8941, nx8945, 
         nx8949, nx8955, nx8959, nx8963, nx8969, nx8972, nx8979, nx8985, nx8989, 
         nx8993, nx8999, nx9003, nx9007, nx9014, nx9017, nx9023, nx9027, nx9031, 
         nx9036, nx9039, nx9043, nx9049, nx9053, nx9057, nx9061, nx9065, nx9069, 
         nx9073, nx9077, nx9080, nx9085, nx9089, nx9093, nx9099, nx9102, nx9105, 
         nx9111, nx9115, nx9119, nx9124, nx9127, nx9131, nx9137, nx9141, nx9145, 
         nx9149, nx9153, nx9157, nx9161, nx9165, nx9168, nx9173, nx9177, nx9181, 
         nx9187, nx9190, nx9193, nx9199, nx9203, nx9207, nx9212, nx9215, nx9219, 
         nx9225, nx9229, nx9233, nx9237, nx9241, nx9245, nx9249, nx9253, nx9257, 
         nx9263, nx9267, nx9271, nx9275, nx9278, nx9281, nx9287, nx9291, nx9295, 
         nx9301, nx9305, nx9308, nx9315, nx9319, nx9323, nx9327, nx9333, nx9336, 
         nx9343, nx9353, nx9357, nx9361, nx9365, nx9373, nx9375, nx9377, nx9379, 
         nx9381, nx9389, nx9391, nx9393, nx9395, nx9397, nx9399, nx9401, nx9403, 
         nx9405, nx9407, nx9409, nx9411, nx9413, nx9415, nx9417, nx9419, nx9421, 
         nx9423, nx9425, nx9427, nx9429, nx9431, nx9433, nx9435, nx9437, nx9439, 
         nx9441, nx9443, nx9445, nx9447, nx9449, nx9451, nx9453, nx9455, nx9457, 
         nx9459, nx9461, nx9463, nx9465, nx9467, nx9469, nx9471, nx9473, nx9475, 
         nx9477, nx9479, nx9481, nx9483, nx9485, nx9487, nx9489, nx9491, nx9493, 
         nx9495, nx9497, nx9499, nx9501, nx9503, nx9505, nx9507, nx9509, nx9511, 
         nx9513, nx9515, nx9517, nx9519, nx9521, nx9523, nx9525, nx9527, nx9529, 
         nx9531, nx9533, nx9535, nx9537, nx9539, nx9541, nx9543, nx9545, nx9547, 
         nx9549, nx9551, nx9553, nx9555, nx9557, nx9559, nx9561, nx9563, nx9565, 
         nx9567, nx9569, nx9571, nx9573, nx9575, nx9577, nx9579, nx9581, nx9583, 
         nx9585, nx9587, nx9589, nx9591, nx9593, nx9595, nx9597, nx9599, nx9601, 
         nx9603, nx9605, nx9607, nx9609, nx9611, nx9613, nx9615, nx9617, nx9619, 
         nx9621, nx9623, nx9625, nx9627, nx9629, nx9631, nx9633, nx9635, nx9637, 
         nx9639, nx9641, nx9643, nx9645, nx9647, nx9649, nx9651, nx9653, nx9655, 
         nx9657, nx9659, nx9661, nx9663, nx9665, nx9667, nx9669, nx9671, nx9673, 
         nx9675, nx9677, nx9679, nx9681, nx9683, nx9685, nx9687, nx9689, nx9691, 
         nx9693, nx9695, nx9697, nx9699, nx9701, nx9703, nx9705, nx9707, nx9709, 
         nx9711, nx9713, nx9715, nx9717, nx9719, nx9721, nx9723, nx9725, nx9727, 
         nx9729, nx9731, nx9733, nx9735, nx9737, nx9739, nx9741, nx9743, nx9745, 
         nx9747, nx9749, nx9751, nx9753, nx9755, nx9757, nx9759, nx9761, nx9763, 
         nx9765, nx9767, nx9769, nx9771, nx9773, nx9775, nx9777, nx9779, nx9781, 
         nx9783, nx9785, nx9787, nx9789, nx9791, nx9793, nx9795, nx9797, nx9799, 
         nx9801, nx9803, nx9805, nx9807, nx9809, nx9811, nx9813, nx9815, nx9817, 
         nx9819, nx9821, nx9823, nx9825, nx9827, nx9829, nx9831, nx9833, nx9835, 
         nx9837, nx9839, nx9841, nx9843, nx9845, nx9847, nx9849, nx9851, nx9853, 
         nx9855, nx9857, nx9859, nx9861, nx9863, nx9865, nx9867, nx9869, nx9871, 
         nx9873, nx9875, nx9877, nx9879, nx9881, nx9883, nx9885, nx9887, nx9889, 
         nx9891, nx9893, nx9895, nx9897, nx9899, nx9901, nx9903, nx9905, nx9907, 
         nx9909, nx9911, nx9913, nx9915, nx9917, nx9919, nx9921, nx9923, nx9925, 
         nx9927, nx9929, nx9931, nx9933, nx9935, nx9937, nx9939, nx9941, nx9943, 
         nx9945, nx9947, nx9949, nx9951, nx9953, nx9955, nx9957, nx9959, nx9961, 
         nx9963, nx9965, nx9967, nx9969, nx9971, nx9973, nx9975, nx9977, nx9979, 
         nx9981, nx9983, nx9985, nx9987, nx9989, nx9991, nx9993, nx9995, nx9997, 
         nx9999, nx10001, nx10003, nx10005, nx10007, nx10009, nx10011, nx10013, 
         nx10015, nx10017, nx10019, nx10021, nx10023, nx10025, nx10027, nx10029, 
         nx10031, nx10033, nx10035, nx10037, nx10039, nx10041, nx10043, nx10045, 
         nx10047, nx10049, nx10051, nx10053, nx10055, nx10057, nx10059, nx10061, 
         nx10063, nx10065, nx10067, nx10069, nx10071, nx10073, nx10075, nx10077, 
         nx10079, nx10081, nx10083, nx10085, nx10087, nx10089, nx10091, nx10093, 
         nx10095, nx10097, nx10099, nx10101, nx10103, nx10105, nx10107, nx10109, 
         nx10111, nx10113, nx10115, nx10117, nx10119, nx10121, nx10123, nx10125, 
         nx10127, nx10129, nx10131, nx10133, nx10135, nx10137, nx10139, nx10141, 
         nx10143, nx10145, nx10147, nx10149, nx10151, nx10153, nx10155, nx10157, 
         nx10159, nx10161, nx10163, nx10165, nx10167, nx10169, nx10171, nx10173, 
         nx10175, nx10177, nx10179, nx10181, nx10183, nx10185, nx10187, nx10189, 
         nx10191, nx10193, nx10195, nx10197, nx10199, nx10201, nx10203, nx10205, 
         nx10207, nx10209, nx10211, nx10213, nx10215, nx10217, nx10219, nx10221, 
         nx10223, nx10225, nx10227, nx10229, nx10231, nx10233, nx10235, nx10237, 
         nx10239, nx10241, nx10243, nx10245, nx10247, nx10249, nx10251, nx10253, 
         nx10255, nx10257, nx10259, nx10261, nx10263, nx10265, nx10267, nx10269, 
         nx10271, nx10273, nx10275, nx10277, nx10279, nx10281, nx10283, nx10285, 
         nx10287, nx10289, nx10291, nx10293, nx10295, nx10297, nx10299, nx10301, 
         nx10303, nx10305, nx10307, nx10309, nx10311, nx10313, nx10315, nx10317, 
         nx10319, nx10321, nx10323, nx10325, nx10327, nx10329, nx10331, nx10333, 
         nx10335, nx10337, nx10339, nx10341, nx10343, nx10345, nx10347, nx10349, 
         nx10351, nx10353, nx10355, nx10357, nx10359, nx10361, nx10363, nx10365, 
         nx10367, nx10369, nx10371, nx10373, nx10375, nx10377, nx10379, nx10381, 
         nx10383, nx10385, nx10387, nx10389, nx10391, nx10393, nx10395, nx10397, 
         nx10399, nx10401, nx10403, nx10405, nx10407, nx10409, nx10411, nx10413, 
         nx10415, nx10417, nx10419, nx10421, nx10423, nx10425, nx10427, nx10429, 
         nx10431, nx10433, nx10435, nx10437, nx10439, nx10441, nx10443, nx10445, 
         nx10447, nx10449, nx10451, nx10453, nx10455, nx10457, nx10459, nx10461, 
         nx10463, nx10465, nx10467, nx10469, nx10471, nx10473, nx10475, nx10477, 
         nx10479, nx10481, nx10483, nx10485, nx10487, nx10489, nx10491, nx10493, 
         nx10495, nx10497, nx10499, nx10501, nx10503, nx10505, nx10507, nx10509, 
         nx10511, nx10513, nx10515, nx10517, nx10519, nx10521, nx10523, nx10525, 
         nx10527, nx10529, nx10531, nx10533, nx10535, nx10537, nx10539, nx10541, 
         nx10543, nx10545, nx10547, nx10549, nx10551, nx10553, nx10555, nx10557, 
         nx10559, nx10561, nx10563, nx10565, nx10567, nx10569, nx10571, nx10573, 
         nx10575, nx10577, nx10579, nx10581, nx10583, nx10585, nx10587, nx10589, 
         nx10591, nx10593, nx10595, nx10597, nx10599, nx10601, nx10603, nx10605, 
         nx10607, nx10609, nx10611, nx10613, nx10615, nx10617, nx10619, nx10621, 
         nx10623, nx10625, nx10627, nx10629, nx10631, nx10633, nx10635, nx10637, 
         nx10639, nx10641, nx10643, nx10645, nx10647, nx10649, nx10651, nx10653, 
         nx10655, nx10657, nx10659, nx10661, nx10663, nx10665, nx10667, nx10669, 
         nx10671, nx10673, nx10675, nx10677, nx10679, nx10681, nx10683, nx10685, 
         nx10687, nx10689, nx10691, nx10693, nx10695, nx10697, nx10699, nx10701, 
         nx10703, nx10705, nx10707, nx10709, nx10711, nx10713, nx10715, nx10717, 
         nx10719, nx10721, nx10723, nx10725, nx10727, nx10729, nx10731, nx10733, 
         nx10735, nx10737, nx10739, nx10741, nx10743, nx10745, nx10747, nx10749, 
         nx10751, nx10753, nx10755, nx10757, nx10759, nx10761, nx10763, nx10765, 
         nx10767, nx10769, nx10771, nx10773, nx10775, nx10777, nx10779, nx10781, 
         nx10783, nx10785, nx10787, nx10789, nx10791, nx10793, nx10795, nx10797, 
         nx10799, nx10801, nx10803, nx10805, nx10807, nx10809, nx10811, nx10813, 
         nx10815, nx10817, nx10819, nx10821, nx10823, nx10825, nx10827, nx10829, 
         nx10831, nx10833, nx10835, nx10837, nx10839, nx10841, nx10843, nx10845, 
         nx10847, nx10849, nx10851, nx10853, nx10855, nx10857, nx10859, nx10861, 
         nx10863, nx10865, nx10867, nx10869, nx10871, nx10873, nx10875, nx10877, 
         nx10879, nx10881, nx10883, nx10885, nx10887, nx10889, nx10891, nx10893, 
         nx10895, nx10897, nx10899, nx10901, nx10903, nx10905, nx10907, nx10909, 
         nx10911, nx10913, nx10915, nx10917, nx10919, nx10921, nx10923, nx10925, 
         nx10927, nx10929, nx10931, nx10933, nx10935, nx10937, nx10939, nx10941, 
         nx10943, nx10945, nx10947, nx10949, nx10951, nx10953, nx10955, nx10957, 
         nx10959, nx10961, nx10963, nx10965, nx10967, nx10969, nx10971, nx10973, 
         nx10975, nx10977, nx10979, nx10981, nx10983, nx10985, nx10987, nx10989, 
         nx10991, nx10993, nx10995, nx10997, nx10999, nx11001, nx11003, nx11005, 
         nx11007, nx11009, nx11011, nx11013, nx11015, nx11017, nx11019, nx11021, 
         nx11023, nx11025, nx11027, nx11029, nx11031, nx11033, nx11035, nx11037, 
         nx11039, nx11041, nx11043, nx11045, nx11047, nx11049, nx11051, nx11053, 
         nx11055, nx11057, nx11059, nx11061, nx11063, nx11065, nx11067, nx11069, 
         nx11071, nx11073, nx11075, nx11077, nx11079, nx11081, nx11083, nx11085, 
         nx11087, nx11089, nx11091, nx11093, nx11095, nx11097, nx11099, nx11101, 
         nx11103, nx11105, nx11107, nx11109, nx11111, nx11113, nx11115, nx11117, 
         nx11119, nx11121, nx11123, nx11125, nx11127, nx11129, nx11131, nx11133, 
         nx11135, nx11137, nx11139, nx11141, nx11143, nx11145, nx11147, nx11157, 
         nx11159, nx11161, nx11163, nx11165, nx11167, nx11169, nx11171, nx11173, 
         nx11175, nx11177, nx11179, nx11181, nx11183, nx11185, nx11187, nx11189, 
         nx11191, nx11197, nx11199, nx11201, nx11203;
    wire [130:0] \$dummy ;




    Reg_33 gen_24_cmp_pRegCmp (.D ({working,working,gen_24_cmp_pBs_30,
           gen_24_cmp_pBs_29,gen_24_cmp_pBs_28,gen_24_cmp_pBs_27,
           gen_24_cmp_pBs_26,gen_24_cmp_pBs_25,gen_24_cmp_pBs_24,
           gen_24_cmp_pBs_23,outputs_24__15,outputs_24__14,outputs_24__13,
           outputs_24__12,outputs_24__11,outputs_24__10,outputs_24__9,
           outputs_24__8,outputs_24__7,outputs_24__6,outputs_24__5,outputs_24__4
           ,outputs_24__3,outputs_24__2,outputs_24__1,outputs_24__0,
           gen_24_cmp_pMux_8,gen_24_cmp_pMux_7,gen_24_cmp_pMux_6,
           gen_24_cmp_pMux_5,gen_24_cmp_pMux_4,gen_24_cmp_pMux_3,nx9399}), .en (
           nx11159), .clk (nx9391), .rst (rst), .Q ({\$dummy [0],\$dummy [1],
           gen_24_cmp_pReg_30,gen_24_cmp_pReg_29,gen_24_cmp_pReg_28,
           gen_24_cmp_pReg_27,gen_24_cmp_pReg_26,gen_24_cmp_pReg_25,
           gen_24_cmp_pReg_24,gen_24_cmp_pReg_23,gen_24_cmp_pReg_22,
           gen_24_cmp_pReg_21,gen_24_cmp_pReg_20,gen_24_cmp_pReg_19,
           gen_24_cmp_pReg_18,gen_24_cmp_pReg_17,gen_24_cmp_pReg_16,
           gen_24_cmp_pReg_15,gen_24_cmp_pReg_14,gen_24_cmp_pReg_13,
           gen_24_cmp_pReg_12,gen_24_cmp_pReg_11,gen_24_cmp_pReg_10,
           gen_24_cmp_pReg_9,gen_24_cmp_pReg_8,gen_24_cmp_pReg_7,
           gen_24_cmp_pReg_6,gen_24_cmp_pReg_5,gen_24_cmp_pReg_4,
           gen_24_cmp_pReg_3,gen_24_cmp_pReg_2,gen_24_cmp_pReg_1,
           gen_24_cmp_pReg_0})) ;
    BinaryMux_33 gen_24_cmp_MuxCmp (.a ({working,working,gen_24_cmp_pReg_30,
                 gen_24_cmp_pReg_29,gen_24_cmp_pReg_28,gen_24_cmp_pReg_27,
                 gen_24_cmp_pReg_26,gen_24_cmp_pReg_25,gen_24_cmp_pReg_24,
                 gen_24_cmp_pReg_23,gen_24_cmp_pReg_22,gen_24_cmp_pReg_21,
                 gen_24_cmp_pReg_20,gen_24_cmp_pReg_19,gen_24_cmp_pReg_18,
                 gen_24_cmp_pReg_17,gen_24_cmp_pReg_16,gen_24_cmp_pReg_15,
                 gen_24_cmp_pReg_14,gen_24_cmp_pReg_13,gen_24_cmp_pReg_12,
                 gen_24_cmp_pReg_11,gen_24_cmp_pReg_10,gen_24_cmp_pReg_9,
                 gen_24_cmp_pReg_8,gen_24_cmp_pReg_7,gen_24_cmp_pReg_6,
                 gen_24_cmp_pReg_5,gen_24_cmp_pReg_4,gen_24_cmp_pReg_3,
                 gen_24_cmp_pReg_2,gen_24_cmp_pReg_1,gen_24_cmp_pReg_0}), .b ({
                 working,working,working,working,working,working,working,working
                 ,working,working,working,working,working,working,working,
                 working,working,working,working,working,working,working,working
                 ,working,filter_24__7,filter_24__6,filter_24__5,filter_24__4,
                 filter_24__3,filter_24__2,filter_24__1,filter_24__0,working}), 
                 .sel (nx11173), .f ({\$dummy [2],\$dummy [3],gen_24_cmp_pMux_30
                 ,gen_24_cmp_pMux_29,gen_24_cmp_pMux_28,gen_24_cmp_pMux_27,
                 gen_24_cmp_pMux_26,gen_24_cmp_pMux_25,gen_24_cmp_pMux_24,
                 gen_24_cmp_pMux_23,gen_24_cmp_pMux_22,gen_24_cmp_pMux_21,
                 gen_24_cmp_pMux_20,gen_24_cmp_pMux_19,gen_24_cmp_pMux_18,
                 gen_24_cmp_pMux_17,gen_24_cmp_pMux_16,gen_24_cmp_pMux_15,
                 gen_24_cmp_pMux_14,gen_24_cmp_pMux_13,gen_24_cmp_pMux_12,
                 gen_24_cmp_pMux_11,gen_24_cmp_pMux_10,gen_24_cmp_pMux_9,
                 gen_24_cmp_pMux_8,gen_24_cmp_pMux_7,gen_24_cmp_pMux_6,
                 gen_24_cmp_pMux_5,gen_24_cmp_pMux_4,gen_24_cmp_pMux_3,
                 gen_24_cmp_pMux_2,gen_24_cmp_pMux_1,gen_24_cmp_pMux_0})) ;
    NBitAdder_24 gen_24_cmp_BSCmp_AdderCmp (.a ({working,working,
                 gen_24_cmp_pMux_30,gen_24_cmp_pMux_29,gen_24_cmp_pMux_28,
                 gen_24_cmp_pMux_27,gen_24_cmp_pMux_26,gen_24_cmp_pMux_25,
                 gen_24_cmp_pMux_24,gen_24_cmp_pMux_23,gen_24_cmp_pMux_22,
                 gen_24_cmp_pMux_21,gen_24_cmp_pMux_20,gen_24_cmp_pMux_19,
                 gen_24_cmp_pMux_18,gen_24_cmp_pMux_17,gen_24_cmp_pMux_16,
                 gen_24_cmp_pMux_15,gen_24_cmp_pMux_14,gen_24_cmp_pMux_13,
                 gen_24_cmp_pMux_12,gen_24_cmp_pMux_11,gen_24_cmp_pMux_10,
                 gen_24_cmp_pMux_9}), .b ({nx9703,nx9703,nx9701,nx9709,nx9707,
                 nx9705,nx9703,nx9701,gen_24_cmp_BSCmp_op2_15,
                 gen_24_cmp_BSCmp_op2_14,gen_24_cmp_BSCmp_op2_13,
                 gen_24_cmp_BSCmp_op2_12,gen_24_cmp_BSCmp_op2_11,
                 gen_24_cmp_BSCmp_op2_10,gen_24_cmp_BSCmp_op2_9,
                 gen_24_cmp_BSCmp_op2_8,gen_24_cmp_BSCmp_op2_7,
                 gen_24_cmp_BSCmp_op2_6,gen_24_cmp_BSCmp_op2_5,
                 gen_24_cmp_BSCmp_op2_4,gen_24_cmp_BSCmp_op2_3,
                 gen_24_cmp_BSCmp_op2_2,gen_24_cmp_BSCmp_op2_1,
                 gen_24_cmp_BSCmp_op2_0}), .carryIn (gen_24_cmp_BSCmp_carryIn), 
                 .sum ({gen_24_cmp_pBs_30,gen_24_cmp_pBs_29,gen_24_cmp_pBs_28,
                 gen_24_cmp_pBs_27,gen_24_cmp_pBs_26,gen_24_cmp_pBs_25,
                 gen_24_cmp_pBs_24,gen_24_cmp_pBs_23,outputs_24__15,
                 outputs_24__14,outputs_24__13,outputs_24__12,outputs_24__11,
                 outputs_24__10,outputs_24__9,outputs_24__8,outputs_24__7,
                 outputs_24__6,outputs_24__5,outputs_24__4,outputs_24__3,
                 outputs_24__2,outputs_24__1,outputs_24__0}), .carryOut (
                 \$dummy [4])) ;
    Reg_33 gen_23_cmp_pRegCmp (.D ({working,working,gen_23_cmp_pBs_30,
           gen_23_cmp_pBs_29,gen_23_cmp_pBs_28,gen_23_cmp_pBs_27,
           gen_23_cmp_pBs_26,gen_23_cmp_pBs_25,gen_23_cmp_pBs_24,
           gen_23_cmp_pBs_23,outputs_23__15,outputs_23__14,outputs_23__13,
           outputs_23__12,outputs_23__11,outputs_23__10,outputs_23__9,
           outputs_23__8,outputs_23__7,outputs_23__6,outputs_23__5,outputs_23__4
           ,outputs_23__3,outputs_23__2,outputs_23__1,outputs_23__0,
           gen_23_cmp_pMux_8,gen_23_cmp_pMux_7,gen_23_cmp_pMux_6,
           gen_23_cmp_pMux_5,gen_23_cmp_pMux_4,gen_23_cmp_pMux_3,nx9411}), .en (
           nx11159), .clk (nx9391), .rst (rst), .Q ({\$dummy [5],\$dummy [6],
           gen_23_cmp_pReg_30,gen_23_cmp_pReg_29,gen_23_cmp_pReg_28,
           gen_23_cmp_pReg_27,gen_23_cmp_pReg_26,gen_23_cmp_pReg_25,
           gen_23_cmp_pReg_24,gen_23_cmp_pReg_23,gen_23_cmp_pReg_22,
           gen_23_cmp_pReg_21,gen_23_cmp_pReg_20,gen_23_cmp_pReg_19,
           gen_23_cmp_pReg_18,gen_23_cmp_pReg_17,gen_23_cmp_pReg_16,
           gen_23_cmp_pReg_15,gen_23_cmp_pReg_14,gen_23_cmp_pReg_13,
           gen_23_cmp_pReg_12,gen_23_cmp_pReg_11,gen_23_cmp_pReg_10,
           gen_23_cmp_pReg_9,gen_23_cmp_pReg_8,gen_23_cmp_pReg_7,
           gen_23_cmp_pReg_6,gen_23_cmp_pReg_5,gen_23_cmp_pReg_4,
           gen_23_cmp_pReg_3,gen_23_cmp_pReg_2,gen_23_cmp_pReg_1,
           gen_23_cmp_pReg_0})) ;
    BinaryMux_33 gen_23_cmp_MuxCmp (.a ({working,working,gen_23_cmp_pReg_30,
                 gen_23_cmp_pReg_29,gen_23_cmp_pReg_28,gen_23_cmp_pReg_27,
                 gen_23_cmp_pReg_26,gen_23_cmp_pReg_25,gen_23_cmp_pReg_24,
                 gen_23_cmp_pReg_23,gen_23_cmp_pReg_22,gen_23_cmp_pReg_21,
                 gen_23_cmp_pReg_20,gen_23_cmp_pReg_19,gen_23_cmp_pReg_18,
                 gen_23_cmp_pReg_17,gen_23_cmp_pReg_16,gen_23_cmp_pReg_15,
                 gen_23_cmp_pReg_14,gen_23_cmp_pReg_13,gen_23_cmp_pReg_12,
                 gen_23_cmp_pReg_11,gen_23_cmp_pReg_10,gen_23_cmp_pReg_9,
                 gen_23_cmp_pReg_8,gen_23_cmp_pReg_7,gen_23_cmp_pReg_6,
                 gen_23_cmp_pReg_5,gen_23_cmp_pReg_4,gen_23_cmp_pReg_3,
                 gen_23_cmp_pReg_2,gen_23_cmp_pReg_1,gen_23_cmp_pReg_0}), .b ({
                 working,working,working,working,working,working,working,working
                 ,working,working,working,working,working,working,working,
                 working,working,working,working,working,working,working,working
                 ,working,filter_23__7,filter_23__6,filter_23__5,filter_23__4,
                 filter_23__3,filter_23__2,filter_23__1,filter_23__0,working}), 
                 .sel (nx11173), .f ({\$dummy [7],\$dummy [8],gen_23_cmp_pMux_30
                 ,gen_23_cmp_pMux_29,gen_23_cmp_pMux_28,gen_23_cmp_pMux_27,
                 gen_23_cmp_pMux_26,gen_23_cmp_pMux_25,gen_23_cmp_pMux_24,
                 gen_23_cmp_pMux_23,gen_23_cmp_pMux_22,gen_23_cmp_pMux_21,
                 gen_23_cmp_pMux_20,gen_23_cmp_pMux_19,gen_23_cmp_pMux_18,
                 gen_23_cmp_pMux_17,gen_23_cmp_pMux_16,gen_23_cmp_pMux_15,
                 gen_23_cmp_pMux_14,gen_23_cmp_pMux_13,gen_23_cmp_pMux_12,
                 gen_23_cmp_pMux_11,gen_23_cmp_pMux_10,gen_23_cmp_pMux_9,
                 gen_23_cmp_pMux_8,gen_23_cmp_pMux_7,gen_23_cmp_pMux_6,
                 gen_23_cmp_pMux_5,gen_23_cmp_pMux_4,gen_23_cmp_pMux_3,
                 gen_23_cmp_pMux_2,gen_23_cmp_pMux_1,gen_23_cmp_pMux_0})) ;
    NBitAdder_24 gen_23_cmp_BSCmp_AdderCmp (.a ({working,working,
                 gen_23_cmp_pMux_30,gen_23_cmp_pMux_29,gen_23_cmp_pMux_28,
                 gen_23_cmp_pMux_27,gen_23_cmp_pMux_26,gen_23_cmp_pMux_25,
                 gen_23_cmp_pMux_24,gen_23_cmp_pMux_23,gen_23_cmp_pMux_22,
                 gen_23_cmp_pMux_21,gen_23_cmp_pMux_20,gen_23_cmp_pMux_19,
                 gen_23_cmp_pMux_18,gen_23_cmp_pMux_17,gen_23_cmp_pMux_16,
                 gen_23_cmp_pMux_15,gen_23_cmp_pMux_14,gen_23_cmp_pMux_13,
                 gen_23_cmp_pMux_12,gen_23_cmp_pMux_11,gen_23_cmp_pMux_10,
                 gen_23_cmp_pMux_9}), .b ({nx9715,nx9715,nx9713,nx9721,nx9719,
                 nx9717,nx9715,nx9713,gen_23_cmp_BSCmp_op2_15,
                 gen_23_cmp_BSCmp_op2_14,gen_23_cmp_BSCmp_op2_13,
                 gen_23_cmp_BSCmp_op2_12,gen_23_cmp_BSCmp_op2_11,
                 gen_23_cmp_BSCmp_op2_10,gen_23_cmp_BSCmp_op2_9,
                 gen_23_cmp_BSCmp_op2_8,gen_23_cmp_BSCmp_op2_7,
                 gen_23_cmp_BSCmp_op2_6,gen_23_cmp_BSCmp_op2_5,
                 gen_23_cmp_BSCmp_op2_4,gen_23_cmp_BSCmp_op2_3,
                 gen_23_cmp_BSCmp_op2_2,gen_23_cmp_BSCmp_op2_1,
                 gen_23_cmp_BSCmp_op2_0}), .carryIn (gen_23_cmp_BSCmp_carryIn), 
                 .sum ({gen_23_cmp_pBs_30,gen_23_cmp_pBs_29,gen_23_cmp_pBs_28,
                 gen_23_cmp_pBs_27,gen_23_cmp_pBs_26,gen_23_cmp_pBs_25,
                 gen_23_cmp_pBs_24,gen_23_cmp_pBs_23,outputs_23__15,
                 outputs_23__14,outputs_23__13,outputs_23__12,outputs_23__11,
                 outputs_23__10,outputs_23__9,outputs_23__8,outputs_23__7,
                 outputs_23__6,outputs_23__5,outputs_23__4,outputs_23__3,
                 outputs_23__2,outputs_23__1,outputs_23__0}), .carryOut (
                 \$dummy [9])) ;
    Reg_33 gen_22_cmp_pRegCmp (.D ({working,working,gen_22_cmp_pBs_30,
           gen_22_cmp_pBs_29,gen_22_cmp_pBs_28,gen_22_cmp_pBs_27,
           gen_22_cmp_pBs_26,gen_22_cmp_pBs_25,gen_22_cmp_pBs_24,
           gen_22_cmp_pBs_23,outputs_22__15,outputs_22__14,outputs_22__13,
           outputs_22__12,outputs_22__11,outputs_22__10,outputs_22__9,
           outputs_22__8,outputs_22__7,outputs_22__6,outputs_22__5,outputs_22__4
           ,outputs_22__3,outputs_22__2,outputs_22__1,outputs_22__0,
           gen_22_cmp_pMux_8,gen_22_cmp_pMux_7,gen_22_cmp_pMux_6,
           gen_22_cmp_pMux_5,gen_22_cmp_pMux_4,gen_22_cmp_pMux_3,nx9423}), .en (
           nx11159), .clk (nx9391), .rst (rst), .Q ({\$dummy [10],\$dummy [11],
           gen_22_cmp_pReg_30,gen_22_cmp_pReg_29,gen_22_cmp_pReg_28,
           gen_22_cmp_pReg_27,gen_22_cmp_pReg_26,gen_22_cmp_pReg_25,
           gen_22_cmp_pReg_24,gen_22_cmp_pReg_23,gen_22_cmp_pReg_22,
           gen_22_cmp_pReg_21,gen_22_cmp_pReg_20,gen_22_cmp_pReg_19,
           gen_22_cmp_pReg_18,gen_22_cmp_pReg_17,gen_22_cmp_pReg_16,
           gen_22_cmp_pReg_15,gen_22_cmp_pReg_14,gen_22_cmp_pReg_13,
           gen_22_cmp_pReg_12,gen_22_cmp_pReg_11,gen_22_cmp_pReg_10,
           gen_22_cmp_pReg_9,gen_22_cmp_pReg_8,gen_22_cmp_pReg_7,
           gen_22_cmp_pReg_6,gen_22_cmp_pReg_5,gen_22_cmp_pReg_4,
           gen_22_cmp_pReg_3,gen_22_cmp_pReg_2,gen_22_cmp_pReg_1,
           gen_22_cmp_pReg_0})) ;
    BinaryMux_33 gen_22_cmp_MuxCmp (.a ({working,working,gen_22_cmp_pReg_30,
                 gen_22_cmp_pReg_29,gen_22_cmp_pReg_28,gen_22_cmp_pReg_27,
                 gen_22_cmp_pReg_26,gen_22_cmp_pReg_25,gen_22_cmp_pReg_24,
                 gen_22_cmp_pReg_23,gen_22_cmp_pReg_22,gen_22_cmp_pReg_21,
                 gen_22_cmp_pReg_20,gen_22_cmp_pReg_19,gen_22_cmp_pReg_18,
                 gen_22_cmp_pReg_17,gen_22_cmp_pReg_16,gen_22_cmp_pReg_15,
                 gen_22_cmp_pReg_14,gen_22_cmp_pReg_13,gen_22_cmp_pReg_12,
                 gen_22_cmp_pReg_11,gen_22_cmp_pReg_10,gen_22_cmp_pReg_9,
                 gen_22_cmp_pReg_8,gen_22_cmp_pReg_7,gen_22_cmp_pReg_6,
                 gen_22_cmp_pReg_5,gen_22_cmp_pReg_4,gen_22_cmp_pReg_3,
                 gen_22_cmp_pReg_2,gen_22_cmp_pReg_1,gen_22_cmp_pReg_0}), .b ({
                 working,working,working,working,working,working,working,working
                 ,working,working,working,working,working,working,working,
                 working,working,working,working,working,working,working,working
                 ,working,filter_22__7,filter_22__6,filter_22__5,filter_22__4,
                 filter_22__3,filter_22__2,filter_22__1,filter_22__0,working}), 
                 .sel (nx11173), .f ({\$dummy [12],\$dummy [13],
                 gen_22_cmp_pMux_30,gen_22_cmp_pMux_29,gen_22_cmp_pMux_28,
                 gen_22_cmp_pMux_27,gen_22_cmp_pMux_26,gen_22_cmp_pMux_25,
                 gen_22_cmp_pMux_24,gen_22_cmp_pMux_23,gen_22_cmp_pMux_22,
                 gen_22_cmp_pMux_21,gen_22_cmp_pMux_20,gen_22_cmp_pMux_19,
                 gen_22_cmp_pMux_18,gen_22_cmp_pMux_17,gen_22_cmp_pMux_16,
                 gen_22_cmp_pMux_15,gen_22_cmp_pMux_14,gen_22_cmp_pMux_13,
                 gen_22_cmp_pMux_12,gen_22_cmp_pMux_11,gen_22_cmp_pMux_10,
                 gen_22_cmp_pMux_9,gen_22_cmp_pMux_8,gen_22_cmp_pMux_7,
                 gen_22_cmp_pMux_6,gen_22_cmp_pMux_5,gen_22_cmp_pMux_4,
                 gen_22_cmp_pMux_3,gen_22_cmp_pMux_2,gen_22_cmp_pMux_1,
                 gen_22_cmp_pMux_0})) ;
    NBitAdder_24 gen_22_cmp_BSCmp_AdderCmp (.a ({working,working,
                 gen_22_cmp_pMux_30,gen_22_cmp_pMux_29,gen_22_cmp_pMux_28,
                 gen_22_cmp_pMux_27,gen_22_cmp_pMux_26,gen_22_cmp_pMux_25,
                 gen_22_cmp_pMux_24,gen_22_cmp_pMux_23,gen_22_cmp_pMux_22,
                 gen_22_cmp_pMux_21,gen_22_cmp_pMux_20,gen_22_cmp_pMux_19,
                 gen_22_cmp_pMux_18,gen_22_cmp_pMux_17,gen_22_cmp_pMux_16,
                 gen_22_cmp_pMux_15,gen_22_cmp_pMux_14,gen_22_cmp_pMux_13,
                 gen_22_cmp_pMux_12,gen_22_cmp_pMux_11,gen_22_cmp_pMux_10,
                 gen_22_cmp_pMux_9}), .b ({nx9727,nx9727,nx9725,nx9733,nx9731,
                 nx9729,nx9727,nx9725,gen_22_cmp_BSCmp_op2_15,
                 gen_22_cmp_BSCmp_op2_14,gen_22_cmp_BSCmp_op2_13,
                 gen_22_cmp_BSCmp_op2_12,gen_22_cmp_BSCmp_op2_11,
                 gen_22_cmp_BSCmp_op2_10,gen_22_cmp_BSCmp_op2_9,
                 gen_22_cmp_BSCmp_op2_8,gen_22_cmp_BSCmp_op2_7,
                 gen_22_cmp_BSCmp_op2_6,gen_22_cmp_BSCmp_op2_5,
                 gen_22_cmp_BSCmp_op2_4,gen_22_cmp_BSCmp_op2_3,
                 gen_22_cmp_BSCmp_op2_2,gen_22_cmp_BSCmp_op2_1,
                 gen_22_cmp_BSCmp_op2_0}), .carryIn (gen_22_cmp_BSCmp_carryIn), 
                 .sum ({gen_22_cmp_pBs_30,gen_22_cmp_pBs_29,gen_22_cmp_pBs_28,
                 gen_22_cmp_pBs_27,gen_22_cmp_pBs_26,gen_22_cmp_pBs_25,
                 gen_22_cmp_pBs_24,gen_22_cmp_pBs_23,outputs_22__15,
                 outputs_22__14,outputs_22__13,outputs_22__12,outputs_22__11,
                 outputs_22__10,outputs_22__9,outputs_22__8,outputs_22__7,
                 outputs_22__6,outputs_22__5,outputs_22__4,outputs_22__3,
                 outputs_22__2,outputs_22__1,outputs_22__0}), .carryOut (
                 \$dummy [14])) ;
    Reg_33 gen_21_cmp_pRegCmp (.D ({working,working,gen_21_cmp_pBs_30,
           gen_21_cmp_pBs_29,gen_21_cmp_pBs_28,gen_21_cmp_pBs_27,
           gen_21_cmp_pBs_26,gen_21_cmp_pBs_25,gen_21_cmp_pBs_24,
           gen_21_cmp_pBs_23,outputs_21__15,outputs_21__14,outputs_21__13,
           outputs_21__12,outputs_21__11,outputs_21__10,outputs_21__9,
           outputs_21__8,outputs_21__7,outputs_21__6,outputs_21__5,outputs_21__4
           ,outputs_21__3,outputs_21__2,outputs_21__1,outputs_21__0,
           gen_21_cmp_pMux_8,gen_21_cmp_pMux_7,gen_21_cmp_pMux_6,
           gen_21_cmp_pMux_5,gen_21_cmp_pMux_4,gen_21_cmp_pMux_3,nx9435}), .en (
           nx11161), .clk (nx9391), .rst (rst), .Q ({\$dummy [15],\$dummy [16],
           gen_21_cmp_pReg_30,gen_21_cmp_pReg_29,gen_21_cmp_pReg_28,
           gen_21_cmp_pReg_27,gen_21_cmp_pReg_26,gen_21_cmp_pReg_25,
           gen_21_cmp_pReg_24,gen_21_cmp_pReg_23,gen_21_cmp_pReg_22,
           gen_21_cmp_pReg_21,gen_21_cmp_pReg_20,gen_21_cmp_pReg_19,
           gen_21_cmp_pReg_18,gen_21_cmp_pReg_17,gen_21_cmp_pReg_16,
           gen_21_cmp_pReg_15,gen_21_cmp_pReg_14,gen_21_cmp_pReg_13,
           gen_21_cmp_pReg_12,gen_21_cmp_pReg_11,gen_21_cmp_pReg_10,
           gen_21_cmp_pReg_9,gen_21_cmp_pReg_8,gen_21_cmp_pReg_7,
           gen_21_cmp_pReg_6,gen_21_cmp_pReg_5,gen_21_cmp_pReg_4,
           gen_21_cmp_pReg_3,gen_21_cmp_pReg_2,gen_21_cmp_pReg_1,
           gen_21_cmp_pReg_0})) ;
    BinaryMux_33 gen_21_cmp_MuxCmp (.a ({working,working,gen_21_cmp_pReg_30,
                 gen_21_cmp_pReg_29,gen_21_cmp_pReg_28,gen_21_cmp_pReg_27,
                 gen_21_cmp_pReg_26,gen_21_cmp_pReg_25,gen_21_cmp_pReg_24,
                 gen_21_cmp_pReg_23,gen_21_cmp_pReg_22,gen_21_cmp_pReg_21,
                 gen_21_cmp_pReg_20,gen_21_cmp_pReg_19,gen_21_cmp_pReg_18,
                 gen_21_cmp_pReg_17,gen_21_cmp_pReg_16,gen_21_cmp_pReg_15,
                 gen_21_cmp_pReg_14,gen_21_cmp_pReg_13,gen_21_cmp_pReg_12,
                 gen_21_cmp_pReg_11,gen_21_cmp_pReg_10,gen_21_cmp_pReg_9,
                 gen_21_cmp_pReg_8,gen_21_cmp_pReg_7,gen_21_cmp_pReg_6,
                 gen_21_cmp_pReg_5,gen_21_cmp_pReg_4,gen_21_cmp_pReg_3,
                 gen_21_cmp_pReg_2,gen_21_cmp_pReg_1,gen_21_cmp_pReg_0}), .b ({
                 working,working,working,working,working,working,working,working
                 ,working,working,working,working,working,working,working,
                 working,working,working,working,working,working,working,working
                 ,working,filter_21__7,filter_21__6,filter_21__5,filter_21__4,
                 filter_21__3,filter_21__2,filter_21__1,filter_21__0,working}), 
                 .sel (nx11175), .f ({\$dummy [17],\$dummy [18],
                 gen_21_cmp_pMux_30,gen_21_cmp_pMux_29,gen_21_cmp_pMux_28,
                 gen_21_cmp_pMux_27,gen_21_cmp_pMux_26,gen_21_cmp_pMux_25,
                 gen_21_cmp_pMux_24,gen_21_cmp_pMux_23,gen_21_cmp_pMux_22,
                 gen_21_cmp_pMux_21,gen_21_cmp_pMux_20,gen_21_cmp_pMux_19,
                 gen_21_cmp_pMux_18,gen_21_cmp_pMux_17,gen_21_cmp_pMux_16,
                 gen_21_cmp_pMux_15,gen_21_cmp_pMux_14,gen_21_cmp_pMux_13,
                 gen_21_cmp_pMux_12,gen_21_cmp_pMux_11,gen_21_cmp_pMux_10,
                 gen_21_cmp_pMux_9,gen_21_cmp_pMux_8,gen_21_cmp_pMux_7,
                 gen_21_cmp_pMux_6,gen_21_cmp_pMux_5,gen_21_cmp_pMux_4,
                 gen_21_cmp_pMux_3,gen_21_cmp_pMux_2,gen_21_cmp_pMux_1,
                 gen_21_cmp_pMux_0})) ;
    NBitAdder_24 gen_21_cmp_BSCmp_AdderCmp (.a ({working,working,
                 gen_21_cmp_pMux_30,gen_21_cmp_pMux_29,gen_21_cmp_pMux_28,
                 gen_21_cmp_pMux_27,gen_21_cmp_pMux_26,gen_21_cmp_pMux_25,
                 gen_21_cmp_pMux_24,gen_21_cmp_pMux_23,gen_21_cmp_pMux_22,
                 gen_21_cmp_pMux_21,gen_21_cmp_pMux_20,gen_21_cmp_pMux_19,
                 gen_21_cmp_pMux_18,gen_21_cmp_pMux_17,gen_21_cmp_pMux_16,
                 gen_21_cmp_pMux_15,gen_21_cmp_pMux_14,gen_21_cmp_pMux_13,
                 gen_21_cmp_pMux_12,gen_21_cmp_pMux_11,gen_21_cmp_pMux_10,
                 gen_21_cmp_pMux_9}), .b ({nx9739,nx9739,nx9737,nx9745,nx9743,
                 nx9741,nx9739,nx9737,gen_21_cmp_BSCmp_op2_15,
                 gen_21_cmp_BSCmp_op2_14,gen_21_cmp_BSCmp_op2_13,
                 gen_21_cmp_BSCmp_op2_12,gen_21_cmp_BSCmp_op2_11,
                 gen_21_cmp_BSCmp_op2_10,gen_21_cmp_BSCmp_op2_9,
                 gen_21_cmp_BSCmp_op2_8,gen_21_cmp_BSCmp_op2_7,
                 gen_21_cmp_BSCmp_op2_6,gen_21_cmp_BSCmp_op2_5,
                 gen_21_cmp_BSCmp_op2_4,gen_21_cmp_BSCmp_op2_3,
                 gen_21_cmp_BSCmp_op2_2,gen_21_cmp_BSCmp_op2_1,
                 gen_21_cmp_BSCmp_op2_0}), .carryIn (gen_21_cmp_BSCmp_carryIn), 
                 .sum ({gen_21_cmp_pBs_30,gen_21_cmp_pBs_29,gen_21_cmp_pBs_28,
                 gen_21_cmp_pBs_27,gen_21_cmp_pBs_26,gen_21_cmp_pBs_25,
                 gen_21_cmp_pBs_24,gen_21_cmp_pBs_23,outputs_21__15,
                 outputs_21__14,outputs_21__13,outputs_21__12,outputs_21__11,
                 outputs_21__10,outputs_21__9,outputs_21__8,outputs_21__7,
                 outputs_21__6,outputs_21__5,outputs_21__4,outputs_21__3,
                 outputs_21__2,outputs_21__1,outputs_21__0}), .carryOut (
                 \$dummy [19])) ;
    Reg_33 gen_20_cmp_pRegCmp (.D ({working,working,gen_20_cmp_pBs_30,
           gen_20_cmp_pBs_29,gen_20_cmp_pBs_28,gen_20_cmp_pBs_27,
           gen_20_cmp_pBs_26,gen_20_cmp_pBs_25,gen_20_cmp_pBs_24,
           gen_20_cmp_pBs_23,outputs_20__15,outputs_20__14,outputs_20__13,
           outputs_20__12,outputs_20__11,outputs_20__10,outputs_20__9,
           outputs_20__8,outputs_20__7,outputs_20__6,outputs_20__5,outputs_20__4
           ,outputs_20__3,outputs_20__2,outputs_20__1,outputs_20__0,
           gen_20_cmp_pMux_8,gen_20_cmp_pMux_7,gen_20_cmp_pMux_6,
           gen_20_cmp_pMux_5,gen_20_cmp_pMux_4,gen_20_cmp_pMux_3,nx9447}), .en (
           nx11161), .clk (nx9391), .rst (rst), .Q ({\$dummy [20],\$dummy [21],
           gen_20_cmp_pReg_30,gen_20_cmp_pReg_29,gen_20_cmp_pReg_28,
           gen_20_cmp_pReg_27,gen_20_cmp_pReg_26,gen_20_cmp_pReg_25,
           gen_20_cmp_pReg_24,gen_20_cmp_pReg_23,gen_20_cmp_pReg_22,
           gen_20_cmp_pReg_21,gen_20_cmp_pReg_20,gen_20_cmp_pReg_19,
           gen_20_cmp_pReg_18,gen_20_cmp_pReg_17,gen_20_cmp_pReg_16,
           gen_20_cmp_pReg_15,gen_20_cmp_pReg_14,gen_20_cmp_pReg_13,
           gen_20_cmp_pReg_12,gen_20_cmp_pReg_11,gen_20_cmp_pReg_10,
           gen_20_cmp_pReg_9,gen_20_cmp_pReg_8,gen_20_cmp_pReg_7,
           gen_20_cmp_pReg_6,gen_20_cmp_pReg_5,gen_20_cmp_pReg_4,
           gen_20_cmp_pReg_3,gen_20_cmp_pReg_2,gen_20_cmp_pReg_1,
           gen_20_cmp_pReg_0})) ;
    BinaryMux_33 gen_20_cmp_MuxCmp (.a ({working,working,gen_20_cmp_pReg_30,
                 gen_20_cmp_pReg_29,gen_20_cmp_pReg_28,gen_20_cmp_pReg_27,
                 gen_20_cmp_pReg_26,gen_20_cmp_pReg_25,gen_20_cmp_pReg_24,
                 gen_20_cmp_pReg_23,gen_20_cmp_pReg_22,gen_20_cmp_pReg_21,
                 gen_20_cmp_pReg_20,gen_20_cmp_pReg_19,gen_20_cmp_pReg_18,
                 gen_20_cmp_pReg_17,gen_20_cmp_pReg_16,gen_20_cmp_pReg_15,
                 gen_20_cmp_pReg_14,gen_20_cmp_pReg_13,gen_20_cmp_pReg_12,
                 gen_20_cmp_pReg_11,gen_20_cmp_pReg_10,gen_20_cmp_pReg_9,
                 gen_20_cmp_pReg_8,gen_20_cmp_pReg_7,gen_20_cmp_pReg_6,
                 gen_20_cmp_pReg_5,gen_20_cmp_pReg_4,gen_20_cmp_pReg_3,
                 gen_20_cmp_pReg_2,gen_20_cmp_pReg_1,gen_20_cmp_pReg_0}), .b ({
                 working,working,working,working,working,working,working,working
                 ,working,working,working,working,working,working,working,
                 working,working,working,working,working,working,working,working
                 ,working,filter_20__7,filter_20__6,filter_20__5,filter_20__4,
                 filter_20__3,filter_20__2,filter_20__1,filter_20__0,working}), 
                 .sel (nx11175), .f ({\$dummy [22],\$dummy [23],
                 gen_20_cmp_pMux_30,gen_20_cmp_pMux_29,gen_20_cmp_pMux_28,
                 gen_20_cmp_pMux_27,gen_20_cmp_pMux_26,gen_20_cmp_pMux_25,
                 gen_20_cmp_pMux_24,gen_20_cmp_pMux_23,gen_20_cmp_pMux_22,
                 gen_20_cmp_pMux_21,gen_20_cmp_pMux_20,gen_20_cmp_pMux_19,
                 gen_20_cmp_pMux_18,gen_20_cmp_pMux_17,gen_20_cmp_pMux_16,
                 gen_20_cmp_pMux_15,gen_20_cmp_pMux_14,gen_20_cmp_pMux_13,
                 gen_20_cmp_pMux_12,gen_20_cmp_pMux_11,gen_20_cmp_pMux_10,
                 gen_20_cmp_pMux_9,gen_20_cmp_pMux_8,gen_20_cmp_pMux_7,
                 gen_20_cmp_pMux_6,gen_20_cmp_pMux_5,gen_20_cmp_pMux_4,
                 gen_20_cmp_pMux_3,gen_20_cmp_pMux_2,gen_20_cmp_pMux_1,
                 gen_20_cmp_pMux_0})) ;
    NBitAdder_24 gen_20_cmp_BSCmp_AdderCmp (.a ({working,working,
                 gen_20_cmp_pMux_30,gen_20_cmp_pMux_29,gen_20_cmp_pMux_28,
                 gen_20_cmp_pMux_27,gen_20_cmp_pMux_26,gen_20_cmp_pMux_25,
                 gen_20_cmp_pMux_24,gen_20_cmp_pMux_23,gen_20_cmp_pMux_22,
                 gen_20_cmp_pMux_21,gen_20_cmp_pMux_20,gen_20_cmp_pMux_19,
                 gen_20_cmp_pMux_18,gen_20_cmp_pMux_17,gen_20_cmp_pMux_16,
                 gen_20_cmp_pMux_15,gen_20_cmp_pMux_14,gen_20_cmp_pMux_13,
                 gen_20_cmp_pMux_12,gen_20_cmp_pMux_11,gen_20_cmp_pMux_10,
                 gen_20_cmp_pMux_9}), .b ({nx9751,nx9751,nx9749,nx9757,nx9755,
                 nx9753,nx9751,nx9749,gen_20_cmp_BSCmp_op2_15,
                 gen_20_cmp_BSCmp_op2_14,gen_20_cmp_BSCmp_op2_13,
                 gen_20_cmp_BSCmp_op2_12,gen_20_cmp_BSCmp_op2_11,
                 gen_20_cmp_BSCmp_op2_10,gen_20_cmp_BSCmp_op2_9,
                 gen_20_cmp_BSCmp_op2_8,gen_20_cmp_BSCmp_op2_7,
                 gen_20_cmp_BSCmp_op2_6,gen_20_cmp_BSCmp_op2_5,
                 gen_20_cmp_BSCmp_op2_4,gen_20_cmp_BSCmp_op2_3,
                 gen_20_cmp_BSCmp_op2_2,gen_20_cmp_BSCmp_op2_1,
                 gen_20_cmp_BSCmp_op2_0}), .carryIn (gen_20_cmp_BSCmp_carryIn), 
                 .sum ({gen_20_cmp_pBs_30,gen_20_cmp_pBs_29,gen_20_cmp_pBs_28,
                 gen_20_cmp_pBs_27,gen_20_cmp_pBs_26,gen_20_cmp_pBs_25,
                 gen_20_cmp_pBs_24,gen_20_cmp_pBs_23,outputs_20__15,
                 outputs_20__14,outputs_20__13,outputs_20__12,outputs_20__11,
                 outputs_20__10,outputs_20__9,outputs_20__8,outputs_20__7,
                 outputs_20__6,outputs_20__5,outputs_20__4,outputs_20__3,
                 outputs_20__2,outputs_20__1,outputs_20__0}), .carryOut (
                 \$dummy [24])) ;
    Reg_33 gen_19_cmp_pRegCmp (.D ({working,working,gen_19_cmp_pBs_30,
           gen_19_cmp_pBs_29,gen_19_cmp_pBs_28,gen_19_cmp_pBs_27,
           gen_19_cmp_pBs_26,gen_19_cmp_pBs_25,gen_19_cmp_pBs_24,
           gen_19_cmp_pBs_23,outputs_19__15,outputs_19__14,outputs_19__13,
           outputs_19__12,outputs_19__11,outputs_19__10,outputs_19__9,
           outputs_19__8,outputs_19__7,outputs_19__6,outputs_19__5,outputs_19__4
           ,outputs_19__3,outputs_19__2,outputs_19__1,outputs_19__0,
           gen_19_cmp_pMux_8,gen_19_cmp_pMux_7,gen_19_cmp_pMux_6,
           gen_19_cmp_pMux_5,gen_19_cmp_pMux_4,gen_19_cmp_pMux_3,nx9459}), .en (
           nx11161), .clk (nx9391), .rst (rst), .Q ({\$dummy [25],\$dummy [26],
           gen_19_cmp_pReg_30,gen_19_cmp_pReg_29,gen_19_cmp_pReg_28,
           gen_19_cmp_pReg_27,gen_19_cmp_pReg_26,gen_19_cmp_pReg_25,
           gen_19_cmp_pReg_24,gen_19_cmp_pReg_23,gen_19_cmp_pReg_22,
           gen_19_cmp_pReg_21,gen_19_cmp_pReg_20,gen_19_cmp_pReg_19,
           gen_19_cmp_pReg_18,gen_19_cmp_pReg_17,gen_19_cmp_pReg_16,
           gen_19_cmp_pReg_15,gen_19_cmp_pReg_14,gen_19_cmp_pReg_13,
           gen_19_cmp_pReg_12,gen_19_cmp_pReg_11,gen_19_cmp_pReg_10,
           gen_19_cmp_pReg_9,gen_19_cmp_pReg_8,gen_19_cmp_pReg_7,
           gen_19_cmp_pReg_6,gen_19_cmp_pReg_5,gen_19_cmp_pReg_4,
           gen_19_cmp_pReg_3,gen_19_cmp_pReg_2,gen_19_cmp_pReg_1,
           gen_19_cmp_pReg_0})) ;
    BinaryMux_33 gen_19_cmp_MuxCmp (.a ({working,working,gen_19_cmp_pReg_30,
                 gen_19_cmp_pReg_29,gen_19_cmp_pReg_28,gen_19_cmp_pReg_27,
                 gen_19_cmp_pReg_26,gen_19_cmp_pReg_25,gen_19_cmp_pReg_24,
                 gen_19_cmp_pReg_23,gen_19_cmp_pReg_22,gen_19_cmp_pReg_21,
                 gen_19_cmp_pReg_20,gen_19_cmp_pReg_19,gen_19_cmp_pReg_18,
                 gen_19_cmp_pReg_17,gen_19_cmp_pReg_16,gen_19_cmp_pReg_15,
                 gen_19_cmp_pReg_14,gen_19_cmp_pReg_13,gen_19_cmp_pReg_12,
                 gen_19_cmp_pReg_11,gen_19_cmp_pReg_10,gen_19_cmp_pReg_9,
                 gen_19_cmp_pReg_8,gen_19_cmp_pReg_7,gen_19_cmp_pReg_6,
                 gen_19_cmp_pReg_5,gen_19_cmp_pReg_4,gen_19_cmp_pReg_3,
                 gen_19_cmp_pReg_2,gen_19_cmp_pReg_1,gen_19_cmp_pReg_0}), .b ({
                 working,working,working,working,working,working,working,working
                 ,working,working,working,working,working,working,working,
                 working,working,working,working,working,working,working,working
                 ,working,filter_19__7,filter_19__6,filter_19__5,filter_19__4,
                 filter_19__3,filter_19__2,filter_19__1,filter_19__0,working}), 
                 .sel (nx11175), .f ({\$dummy [27],\$dummy [28],
                 gen_19_cmp_pMux_30,gen_19_cmp_pMux_29,gen_19_cmp_pMux_28,
                 gen_19_cmp_pMux_27,gen_19_cmp_pMux_26,gen_19_cmp_pMux_25,
                 gen_19_cmp_pMux_24,gen_19_cmp_pMux_23,gen_19_cmp_pMux_22,
                 gen_19_cmp_pMux_21,gen_19_cmp_pMux_20,gen_19_cmp_pMux_19,
                 gen_19_cmp_pMux_18,gen_19_cmp_pMux_17,gen_19_cmp_pMux_16,
                 gen_19_cmp_pMux_15,gen_19_cmp_pMux_14,gen_19_cmp_pMux_13,
                 gen_19_cmp_pMux_12,gen_19_cmp_pMux_11,gen_19_cmp_pMux_10,
                 gen_19_cmp_pMux_9,gen_19_cmp_pMux_8,gen_19_cmp_pMux_7,
                 gen_19_cmp_pMux_6,gen_19_cmp_pMux_5,gen_19_cmp_pMux_4,
                 gen_19_cmp_pMux_3,gen_19_cmp_pMux_2,gen_19_cmp_pMux_1,
                 gen_19_cmp_pMux_0})) ;
    NBitAdder_24 gen_19_cmp_BSCmp_AdderCmp (.a ({working,working,
                 gen_19_cmp_pMux_30,gen_19_cmp_pMux_29,gen_19_cmp_pMux_28,
                 gen_19_cmp_pMux_27,gen_19_cmp_pMux_26,gen_19_cmp_pMux_25,
                 gen_19_cmp_pMux_24,gen_19_cmp_pMux_23,gen_19_cmp_pMux_22,
                 gen_19_cmp_pMux_21,gen_19_cmp_pMux_20,gen_19_cmp_pMux_19,
                 gen_19_cmp_pMux_18,gen_19_cmp_pMux_17,gen_19_cmp_pMux_16,
                 gen_19_cmp_pMux_15,gen_19_cmp_pMux_14,gen_19_cmp_pMux_13,
                 gen_19_cmp_pMux_12,gen_19_cmp_pMux_11,gen_19_cmp_pMux_10,
                 gen_19_cmp_pMux_9}), .b ({nx9763,nx9763,nx9761,nx9769,nx9767,
                 nx9765,nx9763,nx9761,gen_19_cmp_BSCmp_op2_15,
                 gen_19_cmp_BSCmp_op2_14,gen_19_cmp_BSCmp_op2_13,
                 gen_19_cmp_BSCmp_op2_12,gen_19_cmp_BSCmp_op2_11,
                 gen_19_cmp_BSCmp_op2_10,gen_19_cmp_BSCmp_op2_9,
                 gen_19_cmp_BSCmp_op2_8,gen_19_cmp_BSCmp_op2_7,
                 gen_19_cmp_BSCmp_op2_6,gen_19_cmp_BSCmp_op2_5,
                 gen_19_cmp_BSCmp_op2_4,gen_19_cmp_BSCmp_op2_3,
                 gen_19_cmp_BSCmp_op2_2,gen_19_cmp_BSCmp_op2_1,
                 gen_19_cmp_BSCmp_op2_0}), .carryIn (gen_19_cmp_BSCmp_carryIn), 
                 .sum ({gen_19_cmp_pBs_30,gen_19_cmp_pBs_29,gen_19_cmp_pBs_28,
                 gen_19_cmp_pBs_27,gen_19_cmp_pBs_26,gen_19_cmp_pBs_25,
                 gen_19_cmp_pBs_24,gen_19_cmp_pBs_23,outputs_19__15,
                 outputs_19__14,outputs_19__13,outputs_19__12,outputs_19__11,
                 outputs_19__10,outputs_19__9,outputs_19__8,outputs_19__7,
                 outputs_19__6,outputs_19__5,outputs_19__4,outputs_19__3,
                 outputs_19__2,outputs_19__1,outputs_19__0}), .carryOut (
                 \$dummy [29])) ;
    Reg_33 gen_18_cmp_pRegCmp (.D ({working,working,gen_18_cmp_pBs_30,
           gen_18_cmp_pBs_29,gen_18_cmp_pBs_28,gen_18_cmp_pBs_27,
           gen_18_cmp_pBs_26,gen_18_cmp_pBs_25,gen_18_cmp_pBs_24,
           gen_18_cmp_pBs_23,outputs_18__15,outputs_18__14,outputs_18__13,
           outputs_18__12,outputs_18__11,outputs_18__10,outputs_18__9,
           outputs_18__8,outputs_18__7,outputs_18__6,outputs_18__5,outputs_18__4
           ,outputs_18__3,outputs_18__2,outputs_18__1,outputs_18__0,
           gen_18_cmp_pMux_8,gen_18_cmp_pMux_7,gen_18_cmp_pMux_6,
           gen_18_cmp_pMux_5,gen_18_cmp_pMux_4,gen_18_cmp_pMux_3,nx9471}), .en (
           nx9375), .clk (nx9391), .rst (rst), .Q ({\$dummy [30],\$dummy [31],
           gen_18_cmp_pReg_30,gen_18_cmp_pReg_29,gen_18_cmp_pReg_28,
           gen_18_cmp_pReg_27,gen_18_cmp_pReg_26,gen_18_cmp_pReg_25,
           gen_18_cmp_pReg_24,gen_18_cmp_pReg_23,gen_18_cmp_pReg_22,
           gen_18_cmp_pReg_21,gen_18_cmp_pReg_20,gen_18_cmp_pReg_19,
           gen_18_cmp_pReg_18,gen_18_cmp_pReg_17,gen_18_cmp_pReg_16,
           gen_18_cmp_pReg_15,gen_18_cmp_pReg_14,gen_18_cmp_pReg_13,
           gen_18_cmp_pReg_12,gen_18_cmp_pReg_11,gen_18_cmp_pReg_10,
           gen_18_cmp_pReg_9,gen_18_cmp_pReg_8,gen_18_cmp_pReg_7,
           gen_18_cmp_pReg_6,gen_18_cmp_pReg_5,gen_18_cmp_pReg_4,
           gen_18_cmp_pReg_3,gen_18_cmp_pReg_2,gen_18_cmp_pReg_1,
           gen_18_cmp_pReg_0})) ;
    BinaryMux_33 gen_18_cmp_MuxCmp (.a ({working,working,gen_18_cmp_pReg_30,
                 gen_18_cmp_pReg_29,gen_18_cmp_pReg_28,gen_18_cmp_pReg_27,
                 gen_18_cmp_pReg_26,gen_18_cmp_pReg_25,gen_18_cmp_pReg_24,
                 gen_18_cmp_pReg_23,gen_18_cmp_pReg_22,gen_18_cmp_pReg_21,
                 gen_18_cmp_pReg_20,gen_18_cmp_pReg_19,gen_18_cmp_pReg_18,
                 gen_18_cmp_pReg_17,gen_18_cmp_pReg_16,gen_18_cmp_pReg_15,
                 gen_18_cmp_pReg_14,gen_18_cmp_pReg_13,gen_18_cmp_pReg_12,
                 gen_18_cmp_pReg_11,gen_18_cmp_pReg_10,gen_18_cmp_pReg_9,
                 gen_18_cmp_pReg_8,gen_18_cmp_pReg_7,gen_18_cmp_pReg_6,
                 gen_18_cmp_pReg_5,gen_18_cmp_pReg_4,gen_18_cmp_pReg_3,
                 gen_18_cmp_pReg_2,gen_18_cmp_pReg_1,gen_18_cmp_pReg_0}), .b ({
                 working,working,working,working,working,working,working,working
                 ,working,working,working,working,working,working,working,
                 working,working,working,working,working,working,working,working
                 ,working,filter_18__7,filter_18__6,filter_18__5,filter_18__4,
                 filter_18__3,filter_18__2,filter_18__1,filter_18__0,working}), 
                 .sel (nx11177), .f ({\$dummy [32],\$dummy [33],
                 gen_18_cmp_pMux_30,gen_18_cmp_pMux_29,gen_18_cmp_pMux_28,
                 gen_18_cmp_pMux_27,gen_18_cmp_pMux_26,gen_18_cmp_pMux_25,
                 gen_18_cmp_pMux_24,gen_18_cmp_pMux_23,gen_18_cmp_pMux_22,
                 gen_18_cmp_pMux_21,gen_18_cmp_pMux_20,gen_18_cmp_pMux_19,
                 gen_18_cmp_pMux_18,gen_18_cmp_pMux_17,gen_18_cmp_pMux_16,
                 gen_18_cmp_pMux_15,gen_18_cmp_pMux_14,gen_18_cmp_pMux_13,
                 gen_18_cmp_pMux_12,gen_18_cmp_pMux_11,gen_18_cmp_pMux_10,
                 gen_18_cmp_pMux_9,gen_18_cmp_pMux_8,gen_18_cmp_pMux_7,
                 gen_18_cmp_pMux_6,gen_18_cmp_pMux_5,gen_18_cmp_pMux_4,
                 gen_18_cmp_pMux_3,gen_18_cmp_pMux_2,gen_18_cmp_pMux_1,
                 gen_18_cmp_pMux_0})) ;
    NBitAdder_24 gen_18_cmp_BSCmp_AdderCmp (.a ({working,working,
                 gen_18_cmp_pMux_30,gen_18_cmp_pMux_29,gen_18_cmp_pMux_28,
                 gen_18_cmp_pMux_27,gen_18_cmp_pMux_26,gen_18_cmp_pMux_25,
                 gen_18_cmp_pMux_24,gen_18_cmp_pMux_23,gen_18_cmp_pMux_22,
                 gen_18_cmp_pMux_21,gen_18_cmp_pMux_20,gen_18_cmp_pMux_19,
                 gen_18_cmp_pMux_18,gen_18_cmp_pMux_17,gen_18_cmp_pMux_16,
                 gen_18_cmp_pMux_15,gen_18_cmp_pMux_14,gen_18_cmp_pMux_13,
                 gen_18_cmp_pMux_12,gen_18_cmp_pMux_11,gen_18_cmp_pMux_10,
                 gen_18_cmp_pMux_9}), .b ({nx9775,nx9775,nx9773,nx9781,nx9779,
                 nx9777,nx9775,nx9773,gen_18_cmp_BSCmp_op2_15,
                 gen_18_cmp_BSCmp_op2_14,gen_18_cmp_BSCmp_op2_13,
                 gen_18_cmp_BSCmp_op2_12,gen_18_cmp_BSCmp_op2_11,
                 gen_18_cmp_BSCmp_op2_10,gen_18_cmp_BSCmp_op2_9,
                 gen_18_cmp_BSCmp_op2_8,gen_18_cmp_BSCmp_op2_7,
                 gen_18_cmp_BSCmp_op2_6,gen_18_cmp_BSCmp_op2_5,
                 gen_18_cmp_BSCmp_op2_4,gen_18_cmp_BSCmp_op2_3,
                 gen_18_cmp_BSCmp_op2_2,gen_18_cmp_BSCmp_op2_1,
                 gen_18_cmp_BSCmp_op2_0}), .carryIn (gen_18_cmp_BSCmp_carryIn), 
                 .sum ({gen_18_cmp_pBs_30,gen_18_cmp_pBs_29,gen_18_cmp_pBs_28,
                 gen_18_cmp_pBs_27,gen_18_cmp_pBs_26,gen_18_cmp_pBs_25,
                 gen_18_cmp_pBs_24,gen_18_cmp_pBs_23,outputs_18__15,
                 outputs_18__14,outputs_18__13,outputs_18__12,outputs_18__11,
                 outputs_18__10,outputs_18__9,outputs_18__8,outputs_18__7,
                 outputs_18__6,outputs_18__5,outputs_18__4,outputs_18__3,
                 outputs_18__2,outputs_18__1,outputs_18__0}), .carryOut (
                 \$dummy [34])) ;
    Reg_33 gen_17_cmp_pRegCmp (.D ({working,working,gen_17_cmp_pBs_30,
           gen_17_cmp_pBs_29,gen_17_cmp_pBs_28,gen_17_cmp_pBs_27,
           gen_17_cmp_pBs_26,gen_17_cmp_pBs_25,gen_17_cmp_pBs_24,
           gen_17_cmp_pBs_23,outputs_17__15,outputs_17__14,outputs_17__13,
           outputs_17__12,outputs_17__11,outputs_17__10,outputs_17__9,
           outputs_17__8,outputs_17__7,outputs_17__6,outputs_17__5,outputs_17__4
           ,outputs_17__3,outputs_17__2,outputs_17__1,outputs_17__0,
           gen_17_cmp_pMux_8,gen_17_cmp_pMux_7,gen_17_cmp_pMux_6,
           gen_17_cmp_pMux_5,gen_17_cmp_pMux_4,gen_17_cmp_pMux_3,nx9483}), .en (
           nx11163), .clk (nx9393), .rst (rst), .Q ({\$dummy [35],\$dummy [36],
           gen_17_cmp_pReg_30,gen_17_cmp_pReg_29,gen_17_cmp_pReg_28,
           gen_17_cmp_pReg_27,gen_17_cmp_pReg_26,gen_17_cmp_pReg_25,
           gen_17_cmp_pReg_24,gen_17_cmp_pReg_23,gen_17_cmp_pReg_22,
           gen_17_cmp_pReg_21,gen_17_cmp_pReg_20,gen_17_cmp_pReg_19,
           gen_17_cmp_pReg_18,gen_17_cmp_pReg_17,gen_17_cmp_pReg_16,
           gen_17_cmp_pReg_15,gen_17_cmp_pReg_14,gen_17_cmp_pReg_13,
           gen_17_cmp_pReg_12,gen_17_cmp_pReg_11,gen_17_cmp_pReg_10,
           gen_17_cmp_pReg_9,gen_17_cmp_pReg_8,gen_17_cmp_pReg_7,
           gen_17_cmp_pReg_6,gen_17_cmp_pReg_5,gen_17_cmp_pReg_4,
           gen_17_cmp_pReg_3,gen_17_cmp_pReg_2,gen_17_cmp_pReg_1,
           gen_17_cmp_pReg_0})) ;
    BinaryMux_33 gen_17_cmp_MuxCmp (.a ({working,working,gen_17_cmp_pReg_30,
                 gen_17_cmp_pReg_29,gen_17_cmp_pReg_28,gen_17_cmp_pReg_27,
                 gen_17_cmp_pReg_26,gen_17_cmp_pReg_25,gen_17_cmp_pReg_24,
                 gen_17_cmp_pReg_23,gen_17_cmp_pReg_22,gen_17_cmp_pReg_21,
                 gen_17_cmp_pReg_20,gen_17_cmp_pReg_19,gen_17_cmp_pReg_18,
                 gen_17_cmp_pReg_17,gen_17_cmp_pReg_16,gen_17_cmp_pReg_15,
                 gen_17_cmp_pReg_14,gen_17_cmp_pReg_13,gen_17_cmp_pReg_12,
                 gen_17_cmp_pReg_11,gen_17_cmp_pReg_10,gen_17_cmp_pReg_9,
                 gen_17_cmp_pReg_8,gen_17_cmp_pReg_7,gen_17_cmp_pReg_6,
                 gen_17_cmp_pReg_5,gen_17_cmp_pReg_4,gen_17_cmp_pReg_3,
                 gen_17_cmp_pReg_2,gen_17_cmp_pReg_1,gen_17_cmp_pReg_0}), .b ({
                 working,working,working,working,working,working,working,working
                 ,working,working,working,working,working,working,working,
                 working,working,working,working,working,working,working,working
                 ,working,filter_17__7,filter_17__6,filter_17__5,filter_17__4,
                 filter_17__3,filter_17__2,filter_17__1,filter_17__0,working}), 
                 .sel (nx11179), .f ({\$dummy [37],\$dummy [38],
                 gen_17_cmp_pMux_30,gen_17_cmp_pMux_29,gen_17_cmp_pMux_28,
                 gen_17_cmp_pMux_27,gen_17_cmp_pMux_26,gen_17_cmp_pMux_25,
                 gen_17_cmp_pMux_24,gen_17_cmp_pMux_23,gen_17_cmp_pMux_22,
                 gen_17_cmp_pMux_21,gen_17_cmp_pMux_20,gen_17_cmp_pMux_19,
                 gen_17_cmp_pMux_18,gen_17_cmp_pMux_17,gen_17_cmp_pMux_16,
                 gen_17_cmp_pMux_15,gen_17_cmp_pMux_14,gen_17_cmp_pMux_13,
                 gen_17_cmp_pMux_12,gen_17_cmp_pMux_11,gen_17_cmp_pMux_10,
                 gen_17_cmp_pMux_9,gen_17_cmp_pMux_8,gen_17_cmp_pMux_7,
                 gen_17_cmp_pMux_6,gen_17_cmp_pMux_5,gen_17_cmp_pMux_4,
                 gen_17_cmp_pMux_3,gen_17_cmp_pMux_2,gen_17_cmp_pMux_1,
                 gen_17_cmp_pMux_0})) ;
    NBitAdder_24 gen_17_cmp_BSCmp_AdderCmp (.a ({working,working,
                 gen_17_cmp_pMux_30,gen_17_cmp_pMux_29,gen_17_cmp_pMux_28,
                 gen_17_cmp_pMux_27,gen_17_cmp_pMux_26,gen_17_cmp_pMux_25,
                 gen_17_cmp_pMux_24,gen_17_cmp_pMux_23,gen_17_cmp_pMux_22,
                 gen_17_cmp_pMux_21,gen_17_cmp_pMux_20,gen_17_cmp_pMux_19,
                 gen_17_cmp_pMux_18,gen_17_cmp_pMux_17,gen_17_cmp_pMux_16,
                 gen_17_cmp_pMux_15,gen_17_cmp_pMux_14,gen_17_cmp_pMux_13,
                 gen_17_cmp_pMux_12,gen_17_cmp_pMux_11,gen_17_cmp_pMux_10,
                 gen_17_cmp_pMux_9}), .b ({nx9787,nx9787,nx9785,nx9793,nx9791,
                 nx9789,nx9787,nx9785,gen_17_cmp_BSCmp_op2_15,
                 gen_17_cmp_BSCmp_op2_14,gen_17_cmp_BSCmp_op2_13,
                 gen_17_cmp_BSCmp_op2_12,gen_17_cmp_BSCmp_op2_11,
                 gen_17_cmp_BSCmp_op2_10,gen_17_cmp_BSCmp_op2_9,
                 gen_17_cmp_BSCmp_op2_8,gen_17_cmp_BSCmp_op2_7,
                 gen_17_cmp_BSCmp_op2_6,gen_17_cmp_BSCmp_op2_5,
                 gen_17_cmp_BSCmp_op2_4,gen_17_cmp_BSCmp_op2_3,
                 gen_17_cmp_BSCmp_op2_2,gen_17_cmp_BSCmp_op2_1,
                 gen_17_cmp_BSCmp_op2_0}), .carryIn (gen_17_cmp_BSCmp_carryIn), 
                 .sum ({gen_17_cmp_pBs_30,gen_17_cmp_pBs_29,gen_17_cmp_pBs_28,
                 gen_17_cmp_pBs_27,gen_17_cmp_pBs_26,gen_17_cmp_pBs_25,
                 gen_17_cmp_pBs_24,gen_17_cmp_pBs_23,outputs_17__15,
                 outputs_17__14,outputs_17__13,outputs_17__12,outputs_17__11,
                 outputs_17__10,outputs_17__9,outputs_17__8,outputs_17__7,
                 outputs_17__6,outputs_17__5,outputs_17__4,outputs_17__3,
                 outputs_17__2,outputs_17__1,outputs_17__0}), .carryOut (
                 \$dummy [39])) ;
    Reg_33 gen_16_cmp_pRegCmp (.D ({working,working,gen_16_cmp_pBs_30,
           gen_16_cmp_pBs_29,gen_16_cmp_pBs_28,gen_16_cmp_pBs_27,
           gen_16_cmp_pBs_26,gen_16_cmp_pBs_25,gen_16_cmp_pBs_24,
           gen_16_cmp_pBs_23,outputs_16__15,outputs_16__14,outputs_16__13,
           outputs_16__12,outputs_16__11,outputs_16__10,outputs_16__9,
           outputs_16__8,outputs_16__7,outputs_16__6,outputs_16__5,outputs_16__4
           ,outputs_16__3,outputs_16__2,outputs_16__1,outputs_16__0,
           gen_16_cmp_pMux_8,gen_16_cmp_pMux_7,gen_16_cmp_pMux_6,
           gen_16_cmp_pMux_5,gen_16_cmp_pMux_4,gen_16_cmp_pMux_3,nx9495}), .en (
           nx11163), .clk (nx9393), .rst (rst), .Q ({\$dummy [40],\$dummy [41],
           gen_16_cmp_pReg_30,gen_16_cmp_pReg_29,gen_16_cmp_pReg_28,
           gen_16_cmp_pReg_27,gen_16_cmp_pReg_26,gen_16_cmp_pReg_25,
           gen_16_cmp_pReg_24,gen_16_cmp_pReg_23,gen_16_cmp_pReg_22,
           gen_16_cmp_pReg_21,gen_16_cmp_pReg_20,gen_16_cmp_pReg_19,
           gen_16_cmp_pReg_18,gen_16_cmp_pReg_17,gen_16_cmp_pReg_16,
           gen_16_cmp_pReg_15,gen_16_cmp_pReg_14,gen_16_cmp_pReg_13,
           gen_16_cmp_pReg_12,gen_16_cmp_pReg_11,gen_16_cmp_pReg_10,
           gen_16_cmp_pReg_9,gen_16_cmp_pReg_8,gen_16_cmp_pReg_7,
           gen_16_cmp_pReg_6,gen_16_cmp_pReg_5,gen_16_cmp_pReg_4,
           gen_16_cmp_pReg_3,gen_16_cmp_pReg_2,gen_16_cmp_pReg_1,
           gen_16_cmp_pReg_0})) ;
    BinaryMux_33 gen_16_cmp_MuxCmp (.a ({working,working,gen_16_cmp_pReg_30,
                 gen_16_cmp_pReg_29,gen_16_cmp_pReg_28,gen_16_cmp_pReg_27,
                 gen_16_cmp_pReg_26,gen_16_cmp_pReg_25,gen_16_cmp_pReg_24,
                 gen_16_cmp_pReg_23,gen_16_cmp_pReg_22,gen_16_cmp_pReg_21,
                 gen_16_cmp_pReg_20,gen_16_cmp_pReg_19,gen_16_cmp_pReg_18,
                 gen_16_cmp_pReg_17,gen_16_cmp_pReg_16,gen_16_cmp_pReg_15,
                 gen_16_cmp_pReg_14,gen_16_cmp_pReg_13,gen_16_cmp_pReg_12,
                 gen_16_cmp_pReg_11,gen_16_cmp_pReg_10,gen_16_cmp_pReg_9,
                 gen_16_cmp_pReg_8,gen_16_cmp_pReg_7,gen_16_cmp_pReg_6,
                 gen_16_cmp_pReg_5,gen_16_cmp_pReg_4,gen_16_cmp_pReg_3,
                 gen_16_cmp_pReg_2,gen_16_cmp_pReg_1,gen_16_cmp_pReg_0}), .b ({
                 working,working,working,working,working,working,working,working
                 ,working,working,working,working,working,working,working,
                 working,working,working,working,working,working,working,working
                 ,working,filter_16__7,filter_16__6,filter_16__5,filter_16__4,
                 filter_16__3,filter_16__2,filter_16__1,filter_16__0,working}), 
                 .sel (nx11179), .f ({\$dummy [42],\$dummy [43],
                 gen_16_cmp_pMux_30,gen_16_cmp_pMux_29,gen_16_cmp_pMux_28,
                 gen_16_cmp_pMux_27,gen_16_cmp_pMux_26,gen_16_cmp_pMux_25,
                 gen_16_cmp_pMux_24,gen_16_cmp_pMux_23,gen_16_cmp_pMux_22,
                 gen_16_cmp_pMux_21,gen_16_cmp_pMux_20,gen_16_cmp_pMux_19,
                 gen_16_cmp_pMux_18,gen_16_cmp_pMux_17,gen_16_cmp_pMux_16,
                 gen_16_cmp_pMux_15,gen_16_cmp_pMux_14,gen_16_cmp_pMux_13,
                 gen_16_cmp_pMux_12,gen_16_cmp_pMux_11,gen_16_cmp_pMux_10,
                 gen_16_cmp_pMux_9,gen_16_cmp_pMux_8,gen_16_cmp_pMux_7,
                 gen_16_cmp_pMux_6,gen_16_cmp_pMux_5,gen_16_cmp_pMux_4,
                 gen_16_cmp_pMux_3,gen_16_cmp_pMux_2,gen_16_cmp_pMux_1,
                 gen_16_cmp_pMux_0})) ;
    NBitAdder_24 gen_16_cmp_BSCmp_AdderCmp (.a ({working,working,
                 gen_16_cmp_pMux_30,gen_16_cmp_pMux_29,gen_16_cmp_pMux_28,
                 gen_16_cmp_pMux_27,gen_16_cmp_pMux_26,gen_16_cmp_pMux_25,
                 gen_16_cmp_pMux_24,gen_16_cmp_pMux_23,gen_16_cmp_pMux_22,
                 gen_16_cmp_pMux_21,gen_16_cmp_pMux_20,gen_16_cmp_pMux_19,
                 gen_16_cmp_pMux_18,gen_16_cmp_pMux_17,gen_16_cmp_pMux_16,
                 gen_16_cmp_pMux_15,gen_16_cmp_pMux_14,gen_16_cmp_pMux_13,
                 gen_16_cmp_pMux_12,gen_16_cmp_pMux_11,gen_16_cmp_pMux_10,
                 gen_16_cmp_pMux_9}), .b ({nx9799,nx9799,nx9797,nx9805,nx9803,
                 nx9801,nx9799,nx9797,gen_16_cmp_BSCmp_op2_15,
                 gen_16_cmp_BSCmp_op2_14,gen_16_cmp_BSCmp_op2_13,
                 gen_16_cmp_BSCmp_op2_12,gen_16_cmp_BSCmp_op2_11,
                 gen_16_cmp_BSCmp_op2_10,gen_16_cmp_BSCmp_op2_9,
                 gen_16_cmp_BSCmp_op2_8,gen_16_cmp_BSCmp_op2_7,
                 gen_16_cmp_BSCmp_op2_6,gen_16_cmp_BSCmp_op2_5,
                 gen_16_cmp_BSCmp_op2_4,gen_16_cmp_BSCmp_op2_3,
                 gen_16_cmp_BSCmp_op2_2,gen_16_cmp_BSCmp_op2_1,
                 gen_16_cmp_BSCmp_op2_0}), .carryIn (gen_16_cmp_BSCmp_carryIn), 
                 .sum ({gen_16_cmp_pBs_30,gen_16_cmp_pBs_29,gen_16_cmp_pBs_28,
                 gen_16_cmp_pBs_27,gen_16_cmp_pBs_26,gen_16_cmp_pBs_25,
                 gen_16_cmp_pBs_24,gen_16_cmp_pBs_23,outputs_16__15,
                 outputs_16__14,outputs_16__13,outputs_16__12,outputs_16__11,
                 outputs_16__10,outputs_16__9,outputs_16__8,outputs_16__7,
                 outputs_16__6,outputs_16__5,outputs_16__4,outputs_16__3,
                 outputs_16__2,outputs_16__1,outputs_16__0}), .carryOut (
                 \$dummy [44])) ;
    Reg_33 gen_15_cmp_pRegCmp (.D ({working,working,gen_15_cmp_pBs_30,
           gen_15_cmp_pBs_29,gen_15_cmp_pBs_28,gen_15_cmp_pBs_27,
           gen_15_cmp_pBs_26,gen_15_cmp_pBs_25,gen_15_cmp_pBs_24,
           gen_15_cmp_pBs_23,outputs_15__15,outputs_15__14,outputs_15__13,
           outputs_15__12,outputs_15__11,outputs_15__10,outputs_15__9,
           outputs_15__8,outputs_15__7,outputs_15__6,outputs_15__5,outputs_15__4
           ,outputs_15__3,outputs_15__2,outputs_15__1,outputs_15__0,
           gen_15_cmp_pMux_8,gen_15_cmp_pMux_7,gen_15_cmp_pMux_6,
           gen_15_cmp_pMux_5,gen_15_cmp_pMux_4,gen_15_cmp_pMux_3,nx9507}), .en (
           nx11163), .clk (nx9393), .rst (rst), .Q ({\$dummy [45],\$dummy [46],
           gen_15_cmp_pReg_30,gen_15_cmp_pReg_29,gen_15_cmp_pReg_28,
           gen_15_cmp_pReg_27,gen_15_cmp_pReg_26,gen_15_cmp_pReg_25,
           gen_15_cmp_pReg_24,gen_15_cmp_pReg_23,gen_15_cmp_pReg_22,
           gen_15_cmp_pReg_21,gen_15_cmp_pReg_20,gen_15_cmp_pReg_19,
           gen_15_cmp_pReg_18,gen_15_cmp_pReg_17,gen_15_cmp_pReg_16,
           gen_15_cmp_pReg_15,gen_15_cmp_pReg_14,gen_15_cmp_pReg_13,
           gen_15_cmp_pReg_12,gen_15_cmp_pReg_11,gen_15_cmp_pReg_10,
           gen_15_cmp_pReg_9,gen_15_cmp_pReg_8,gen_15_cmp_pReg_7,
           gen_15_cmp_pReg_6,gen_15_cmp_pReg_5,gen_15_cmp_pReg_4,
           gen_15_cmp_pReg_3,gen_15_cmp_pReg_2,gen_15_cmp_pReg_1,
           gen_15_cmp_pReg_0})) ;
    BinaryMux_33 gen_15_cmp_MuxCmp (.a ({working,working,gen_15_cmp_pReg_30,
                 gen_15_cmp_pReg_29,gen_15_cmp_pReg_28,gen_15_cmp_pReg_27,
                 gen_15_cmp_pReg_26,gen_15_cmp_pReg_25,gen_15_cmp_pReg_24,
                 gen_15_cmp_pReg_23,gen_15_cmp_pReg_22,gen_15_cmp_pReg_21,
                 gen_15_cmp_pReg_20,gen_15_cmp_pReg_19,gen_15_cmp_pReg_18,
                 gen_15_cmp_pReg_17,gen_15_cmp_pReg_16,gen_15_cmp_pReg_15,
                 gen_15_cmp_pReg_14,gen_15_cmp_pReg_13,gen_15_cmp_pReg_12,
                 gen_15_cmp_pReg_11,gen_15_cmp_pReg_10,gen_15_cmp_pReg_9,
                 gen_15_cmp_pReg_8,gen_15_cmp_pReg_7,gen_15_cmp_pReg_6,
                 gen_15_cmp_pReg_5,gen_15_cmp_pReg_4,gen_15_cmp_pReg_3,
                 gen_15_cmp_pReg_2,gen_15_cmp_pReg_1,gen_15_cmp_pReg_0}), .b ({
                 working,working,working,working,working,working,working,working
                 ,working,working,working,working,working,working,working,
                 working,working,working,working,working,working,working,working
                 ,working,filter_15__7,filter_15__6,filter_15__5,filter_15__4,
                 filter_15__3,filter_15__2,filter_15__1,filter_15__0,working}), 
                 .sel (nx11179), .f ({\$dummy [47],\$dummy [48],
                 gen_15_cmp_pMux_30,gen_15_cmp_pMux_29,gen_15_cmp_pMux_28,
                 gen_15_cmp_pMux_27,gen_15_cmp_pMux_26,gen_15_cmp_pMux_25,
                 gen_15_cmp_pMux_24,gen_15_cmp_pMux_23,gen_15_cmp_pMux_22,
                 gen_15_cmp_pMux_21,gen_15_cmp_pMux_20,gen_15_cmp_pMux_19,
                 gen_15_cmp_pMux_18,gen_15_cmp_pMux_17,gen_15_cmp_pMux_16,
                 gen_15_cmp_pMux_15,gen_15_cmp_pMux_14,gen_15_cmp_pMux_13,
                 gen_15_cmp_pMux_12,gen_15_cmp_pMux_11,gen_15_cmp_pMux_10,
                 gen_15_cmp_pMux_9,gen_15_cmp_pMux_8,gen_15_cmp_pMux_7,
                 gen_15_cmp_pMux_6,gen_15_cmp_pMux_5,gen_15_cmp_pMux_4,
                 gen_15_cmp_pMux_3,gen_15_cmp_pMux_2,gen_15_cmp_pMux_1,
                 gen_15_cmp_pMux_0})) ;
    NBitAdder_24 gen_15_cmp_BSCmp_AdderCmp (.a ({working,working,
                 gen_15_cmp_pMux_30,gen_15_cmp_pMux_29,gen_15_cmp_pMux_28,
                 gen_15_cmp_pMux_27,gen_15_cmp_pMux_26,gen_15_cmp_pMux_25,
                 gen_15_cmp_pMux_24,gen_15_cmp_pMux_23,gen_15_cmp_pMux_22,
                 gen_15_cmp_pMux_21,gen_15_cmp_pMux_20,gen_15_cmp_pMux_19,
                 gen_15_cmp_pMux_18,gen_15_cmp_pMux_17,gen_15_cmp_pMux_16,
                 gen_15_cmp_pMux_15,gen_15_cmp_pMux_14,gen_15_cmp_pMux_13,
                 gen_15_cmp_pMux_12,gen_15_cmp_pMux_11,gen_15_cmp_pMux_10,
                 gen_15_cmp_pMux_9}), .b ({nx9811,nx9811,nx9809,nx9817,nx9815,
                 nx9813,nx9811,nx9809,gen_15_cmp_BSCmp_op2_15,
                 gen_15_cmp_BSCmp_op2_14,gen_15_cmp_BSCmp_op2_13,
                 gen_15_cmp_BSCmp_op2_12,gen_15_cmp_BSCmp_op2_11,
                 gen_15_cmp_BSCmp_op2_10,gen_15_cmp_BSCmp_op2_9,
                 gen_15_cmp_BSCmp_op2_8,gen_15_cmp_BSCmp_op2_7,
                 gen_15_cmp_BSCmp_op2_6,gen_15_cmp_BSCmp_op2_5,
                 gen_15_cmp_BSCmp_op2_4,gen_15_cmp_BSCmp_op2_3,
                 gen_15_cmp_BSCmp_op2_2,gen_15_cmp_BSCmp_op2_1,
                 gen_15_cmp_BSCmp_op2_0}), .carryIn (gen_15_cmp_BSCmp_carryIn), 
                 .sum ({gen_15_cmp_pBs_30,gen_15_cmp_pBs_29,gen_15_cmp_pBs_28,
                 gen_15_cmp_pBs_27,gen_15_cmp_pBs_26,gen_15_cmp_pBs_25,
                 gen_15_cmp_pBs_24,gen_15_cmp_pBs_23,outputs_15__15,
                 outputs_15__14,outputs_15__13,outputs_15__12,outputs_15__11,
                 outputs_15__10,outputs_15__9,outputs_15__8,outputs_15__7,
                 outputs_15__6,outputs_15__5,outputs_15__4,outputs_15__3,
                 outputs_15__2,outputs_15__1,outputs_15__0}), .carryOut (
                 \$dummy [49])) ;
    Reg_33 gen_14_cmp_pRegCmp (.D ({working,working,gen_14_cmp_pBs_30,
           gen_14_cmp_pBs_29,gen_14_cmp_pBs_28,gen_14_cmp_pBs_27,
           gen_14_cmp_pBs_26,gen_14_cmp_pBs_25,gen_14_cmp_pBs_24,
           gen_14_cmp_pBs_23,outputs_14__15,outputs_14__14,outputs_14__13,
           outputs_14__12,outputs_14__11,outputs_14__10,outputs_14__9,
           outputs_14__8,outputs_14__7,outputs_14__6,outputs_14__5,outputs_14__4
           ,outputs_14__3,outputs_14__2,outputs_14__1,outputs_14__0,
           gen_14_cmp_pMux_8,gen_14_cmp_pMux_7,gen_14_cmp_pMux_6,
           gen_14_cmp_pMux_5,gen_14_cmp_pMux_4,gen_14_cmp_pMux_3,nx9519}), .en (
           nx11165), .clk (nx9393), .rst (rst), .Q ({\$dummy [50],\$dummy [51],
           gen_14_cmp_pReg_30,gen_14_cmp_pReg_29,gen_14_cmp_pReg_28,
           gen_14_cmp_pReg_27,gen_14_cmp_pReg_26,gen_14_cmp_pReg_25,
           gen_14_cmp_pReg_24,gen_14_cmp_pReg_23,gen_14_cmp_pReg_22,
           gen_14_cmp_pReg_21,gen_14_cmp_pReg_20,gen_14_cmp_pReg_19,
           gen_14_cmp_pReg_18,gen_14_cmp_pReg_17,gen_14_cmp_pReg_16,
           gen_14_cmp_pReg_15,gen_14_cmp_pReg_14,gen_14_cmp_pReg_13,
           gen_14_cmp_pReg_12,gen_14_cmp_pReg_11,gen_14_cmp_pReg_10,
           gen_14_cmp_pReg_9,gen_14_cmp_pReg_8,gen_14_cmp_pReg_7,
           gen_14_cmp_pReg_6,gen_14_cmp_pReg_5,gen_14_cmp_pReg_4,
           gen_14_cmp_pReg_3,gen_14_cmp_pReg_2,gen_14_cmp_pReg_1,
           gen_14_cmp_pReg_0})) ;
    BinaryMux_33 gen_14_cmp_MuxCmp (.a ({working,working,gen_14_cmp_pReg_30,
                 gen_14_cmp_pReg_29,gen_14_cmp_pReg_28,gen_14_cmp_pReg_27,
                 gen_14_cmp_pReg_26,gen_14_cmp_pReg_25,gen_14_cmp_pReg_24,
                 gen_14_cmp_pReg_23,gen_14_cmp_pReg_22,gen_14_cmp_pReg_21,
                 gen_14_cmp_pReg_20,gen_14_cmp_pReg_19,gen_14_cmp_pReg_18,
                 gen_14_cmp_pReg_17,gen_14_cmp_pReg_16,gen_14_cmp_pReg_15,
                 gen_14_cmp_pReg_14,gen_14_cmp_pReg_13,gen_14_cmp_pReg_12,
                 gen_14_cmp_pReg_11,gen_14_cmp_pReg_10,gen_14_cmp_pReg_9,
                 gen_14_cmp_pReg_8,gen_14_cmp_pReg_7,gen_14_cmp_pReg_6,
                 gen_14_cmp_pReg_5,gen_14_cmp_pReg_4,gen_14_cmp_pReg_3,
                 gen_14_cmp_pReg_2,gen_14_cmp_pReg_1,gen_14_cmp_pReg_0}), .b ({
                 working,working,working,working,working,working,working,working
                 ,working,working,working,working,working,working,working,
                 working,working,working,working,working,working,working,working
                 ,working,filter_14__7,filter_14__6,filter_14__5,filter_14__4,
                 filter_14__3,filter_14__2,filter_14__1,filter_14__0,working}), 
                 .sel (nx11181), .f ({\$dummy [52],\$dummy [53],
                 gen_14_cmp_pMux_30,gen_14_cmp_pMux_29,gen_14_cmp_pMux_28,
                 gen_14_cmp_pMux_27,gen_14_cmp_pMux_26,gen_14_cmp_pMux_25,
                 gen_14_cmp_pMux_24,gen_14_cmp_pMux_23,gen_14_cmp_pMux_22,
                 gen_14_cmp_pMux_21,gen_14_cmp_pMux_20,gen_14_cmp_pMux_19,
                 gen_14_cmp_pMux_18,gen_14_cmp_pMux_17,gen_14_cmp_pMux_16,
                 gen_14_cmp_pMux_15,gen_14_cmp_pMux_14,gen_14_cmp_pMux_13,
                 gen_14_cmp_pMux_12,gen_14_cmp_pMux_11,gen_14_cmp_pMux_10,
                 gen_14_cmp_pMux_9,gen_14_cmp_pMux_8,gen_14_cmp_pMux_7,
                 gen_14_cmp_pMux_6,gen_14_cmp_pMux_5,gen_14_cmp_pMux_4,
                 gen_14_cmp_pMux_3,gen_14_cmp_pMux_2,gen_14_cmp_pMux_1,
                 gen_14_cmp_pMux_0})) ;
    NBitAdder_24 gen_14_cmp_BSCmp_AdderCmp (.a ({working,working,
                 gen_14_cmp_pMux_30,gen_14_cmp_pMux_29,gen_14_cmp_pMux_28,
                 gen_14_cmp_pMux_27,gen_14_cmp_pMux_26,gen_14_cmp_pMux_25,
                 gen_14_cmp_pMux_24,gen_14_cmp_pMux_23,gen_14_cmp_pMux_22,
                 gen_14_cmp_pMux_21,gen_14_cmp_pMux_20,gen_14_cmp_pMux_19,
                 gen_14_cmp_pMux_18,gen_14_cmp_pMux_17,gen_14_cmp_pMux_16,
                 gen_14_cmp_pMux_15,gen_14_cmp_pMux_14,gen_14_cmp_pMux_13,
                 gen_14_cmp_pMux_12,gen_14_cmp_pMux_11,gen_14_cmp_pMux_10,
                 gen_14_cmp_pMux_9}), .b ({nx9823,nx9823,nx9821,nx9829,nx9827,
                 nx9825,nx9823,nx9821,gen_14_cmp_BSCmp_op2_15,
                 gen_14_cmp_BSCmp_op2_14,gen_14_cmp_BSCmp_op2_13,
                 gen_14_cmp_BSCmp_op2_12,gen_14_cmp_BSCmp_op2_11,
                 gen_14_cmp_BSCmp_op2_10,gen_14_cmp_BSCmp_op2_9,
                 gen_14_cmp_BSCmp_op2_8,gen_14_cmp_BSCmp_op2_7,
                 gen_14_cmp_BSCmp_op2_6,gen_14_cmp_BSCmp_op2_5,
                 gen_14_cmp_BSCmp_op2_4,gen_14_cmp_BSCmp_op2_3,
                 gen_14_cmp_BSCmp_op2_2,gen_14_cmp_BSCmp_op2_1,
                 gen_14_cmp_BSCmp_op2_0}), .carryIn (gen_14_cmp_BSCmp_carryIn), 
                 .sum ({gen_14_cmp_pBs_30,gen_14_cmp_pBs_29,gen_14_cmp_pBs_28,
                 gen_14_cmp_pBs_27,gen_14_cmp_pBs_26,gen_14_cmp_pBs_25,
                 gen_14_cmp_pBs_24,gen_14_cmp_pBs_23,outputs_14__15,
                 outputs_14__14,outputs_14__13,outputs_14__12,outputs_14__11,
                 outputs_14__10,outputs_14__9,outputs_14__8,outputs_14__7,
                 outputs_14__6,outputs_14__5,outputs_14__4,outputs_14__3,
                 outputs_14__2,outputs_14__1,outputs_14__0}), .carryOut (
                 \$dummy [54])) ;
    Reg_33 gen_13_cmp_pRegCmp (.D ({working,working,gen_13_cmp_pBs_30,
           gen_13_cmp_pBs_29,gen_13_cmp_pBs_28,gen_13_cmp_pBs_27,
           gen_13_cmp_pBs_26,gen_13_cmp_pBs_25,gen_13_cmp_pBs_24,
           gen_13_cmp_pBs_23,outputs_13__15,outputs_13__14,outputs_13__13,
           outputs_13__12,outputs_13__11,outputs_13__10,outputs_13__9,
           outputs_13__8,outputs_13__7,outputs_13__6,outputs_13__5,outputs_13__4
           ,outputs_13__3,outputs_13__2,outputs_13__1,outputs_13__0,
           gen_13_cmp_pMux_8,gen_13_cmp_pMux_7,gen_13_cmp_pMux_6,
           gen_13_cmp_pMux_5,gen_13_cmp_pMux_4,gen_13_cmp_pMux_3,nx9531}), .en (
           nx11165), .clk (nx9393), .rst (rst), .Q ({\$dummy [55],\$dummy [56],
           gen_13_cmp_pReg_30,gen_13_cmp_pReg_29,gen_13_cmp_pReg_28,
           gen_13_cmp_pReg_27,gen_13_cmp_pReg_26,gen_13_cmp_pReg_25,
           gen_13_cmp_pReg_24,gen_13_cmp_pReg_23,gen_13_cmp_pReg_22,
           gen_13_cmp_pReg_21,gen_13_cmp_pReg_20,gen_13_cmp_pReg_19,
           gen_13_cmp_pReg_18,gen_13_cmp_pReg_17,gen_13_cmp_pReg_16,
           gen_13_cmp_pReg_15,gen_13_cmp_pReg_14,gen_13_cmp_pReg_13,
           gen_13_cmp_pReg_12,gen_13_cmp_pReg_11,gen_13_cmp_pReg_10,
           gen_13_cmp_pReg_9,gen_13_cmp_pReg_8,gen_13_cmp_pReg_7,
           gen_13_cmp_pReg_6,gen_13_cmp_pReg_5,gen_13_cmp_pReg_4,
           gen_13_cmp_pReg_3,gen_13_cmp_pReg_2,gen_13_cmp_pReg_1,
           gen_13_cmp_pReg_0})) ;
    BinaryMux_33 gen_13_cmp_MuxCmp (.a ({working,working,gen_13_cmp_pReg_30,
                 gen_13_cmp_pReg_29,gen_13_cmp_pReg_28,gen_13_cmp_pReg_27,
                 gen_13_cmp_pReg_26,gen_13_cmp_pReg_25,gen_13_cmp_pReg_24,
                 gen_13_cmp_pReg_23,gen_13_cmp_pReg_22,gen_13_cmp_pReg_21,
                 gen_13_cmp_pReg_20,gen_13_cmp_pReg_19,gen_13_cmp_pReg_18,
                 gen_13_cmp_pReg_17,gen_13_cmp_pReg_16,gen_13_cmp_pReg_15,
                 gen_13_cmp_pReg_14,gen_13_cmp_pReg_13,gen_13_cmp_pReg_12,
                 gen_13_cmp_pReg_11,gen_13_cmp_pReg_10,gen_13_cmp_pReg_9,
                 gen_13_cmp_pReg_8,gen_13_cmp_pReg_7,gen_13_cmp_pReg_6,
                 gen_13_cmp_pReg_5,gen_13_cmp_pReg_4,gen_13_cmp_pReg_3,
                 gen_13_cmp_pReg_2,gen_13_cmp_pReg_1,gen_13_cmp_pReg_0}), .b ({
                 working,working,working,working,working,working,working,working
                 ,working,working,working,working,working,working,working,
                 working,working,working,working,working,working,working,working
                 ,working,filter_13__7,filter_13__6,filter_13__5,filter_13__4,
                 filter_13__3,filter_13__2,filter_13__1,filter_13__0,working}), 
                 .sel (nx11181), .f ({\$dummy [57],\$dummy [58],
                 gen_13_cmp_pMux_30,gen_13_cmp_pMux_29,gen_13_cmp_pMux_28,
                 gen_13_cmp_pMux_27,gen_13_cmp_pMux_26,gen_13_cmp_pMux_25,
                 gen_13_cmp_pMux_24,gen_13_cmp_pMux_23,gen_13_cmp_pMux_22,
                 gen_13_cmp_pMux_21,gen_13_cmp_pMux_20,gen_13_cmp_pMux_19,
                 gen_13_cmp_pMux_18,gen_13_cmp_pMux_17,gen_13_cmp_pMux_16,
                 gen_13_cmp_pMux_15,gen_13_cmp_pMux_14,gen_13_cmp_pMux_13,
                 gen_13_cmp_pMux_12,gen_13_cmp_pMux_11,gen_13_cmp_pMux_10,
                 gen_13_cmp_pMux_9,gen_13_cmp_pMux_8,gen_13_cmp_pMux_7,
                 gen_13_cmp_pMux_6,gen_13_cmp_pMux_5,gen_13_cmp_pMux_4,
                 gen_13_cmp_pMux_3,gen_13_cmp_pMux_2,gen_13_cmp_pMux_1,
                 gen_13_cmp_pMux_0})) ;
    NBitAdder_24 gen_13_cmp_BSCmp_AdderCmp (.a ({working,working,
                 gen_13_cmp_pMux_30,gen_13_cmp_pMux_29,gen_13_cmp_pMux_28,
                 gen_13_cmp_pMux_27,gen_13_cmp_pMux_26,gen_13_cmp_pMux_25,
                 gen_13_cmp_pMux_24,gen_13_cmp_pMux_23,gen_13_cmp_pMux_22,
                 gen_13_cmp_pMux_21,gen_13_cmp_pMux_20,gen_13_cmp_pMux_19,
                 gen_13_cmp_pMux_18,gen_13_cmp_pMux_17,gen_13_cmp_pMux_16,
                 gen_13_cmp_pMux_15,gen_13_cmp_pMux_14,gen_13_cmp_pMux_13,
                 gen_13_cmp_pMux_12,gen_13_cmp_pMux_11,gen_13_cmp_pMux_10,
                 gen_13_cmp_pMux_9}), .b ({nx9835,nx9835,nx9833,nx9841,nx9839,
                 nx9837,nx9835,nx9833,gen_13_cmp_BSCmp_op2_15,
                 gen_13_cmp_BSCmp_op2_14,gen_13_cmp_BSCmp_op2_13,
                 gen_13_cmp_BSCmp_op2_12,gen_13_cmp_BSCmp_op2_11,
                 gen_13_cmp_BSCmp_op2_10,gen_13_cmp_BSCmp_op2_9,
                 gen_13_cmp_BSCmp_op2_8,gen_13_cmp_BSCmp_op2_7,
                 gen_13_cmp_BSCmp_op2_6,gen_13_cmp_BSCmp_op2_5,
                 gen_13_cmp_BSCmp_op2_4,gen_13_cmp_BSCmp_op2_3,
                 gen_13_cmp_BSCmp_op2_2,gen_13_cmp_BSCmp_op2_1,
                 gen_13_cmp_BSCmp_op2_0}), .carryIn (gen_13_cmp_BSCmp_carryIn), 
                 .sum ({gen_13_cmp_pBs_30,gen_13_cmp_pBs_29,gen_13_cmp_pBs_28,
                 gen_13_cmp_pBs_27,gen_13_cmp_pBs_26,gen_13_cmp_pBs_25,
                 gen_13_cmp_pBs_24,gen_13_cmp_pBs_23,outputs_13__15,
                 outputs_13__14,outputs_13__13,outputs_13__12,outputs_13__11,
                 outputs_13__10,outputs_13__9,outputs_13__8,outputs_13__7,
                 outputs_13__6,outputs_13__5,outputs_13__4,outputs_13__3,
                 outputs_13__2,outputs_13__1,outputs_13__0}), .carryOut (
                 \$dummy [59])) ;
    Reg_33 gen_12_cmp_pRegCmp (.D ({working,working,gen_12_cmp_pBs_30,
           gen_12_cmp_pBs_29,gen_12_cmp_pBs_28,gen_12_cmp_pBs_27,
           gen_12_cmp_pBs_26,gen_12_cmp_pBs_25,gen_12_cmp_pBs_24,
           gen_12_cmp_pBs_23,outputs_12__15,outputs_12__14,outputs_12__13,
           outputs_12__12,outputs_12__11,outputs_12__10,outputs_12__9,
           outputs_12__8,outputs_12__7,outputs_12__6,outputs_12__5,outputs_12__4
           ,outputs_12__3,outputs_12__2,outputs_12__1,outputs_12__0,
           gen_12_cmp_pMux_8,gen_12_cmp_pMux_7,gen_12_cmp_pMux_6,
           gen_12_cmp_pMux_5,gen_12_cmp_pMux_4,gen_12_cmp_pMux_3,nx9543}), .en (
           nx11165), .clk (nx9393), .rst (rst), .Q ({\$dummy [60],\$dummy [61],
           gen_12_cmp_pReg_30,gen_12_cmp_pReg_29,gen_12_cmp_pReg_28,
           gen_12_cmp_pReg_27,gen_12_cmp_pReg_26,gen_12_cmp_pReg_25,
           gen_12_cmp_pReg_24,gen_12_cmp_pReg_23,gen_12_cmp_pReg_22,
           gen_12_cmp_pReg_21,gen_12_cmp_pReg_20,gen_12_cmp_pReg_19,
           gen_12_cmp_pReg_18,gen_12_cmp_pReg_17,gen_12_cmp_pReg_16,
           gen_12_cmp_pReg_15,gen_12_cmp_pReg_14,gen_12_cmp_pReg_13,
           gen_12_cmp_pReg_12,gen_12_cmp_pReg_11,gen_12_cmp_pReg_10,
           gen_12_cmp_pReg_9,gen_12_cmp_pReg_8,gen_12_cmp_pReg_7,
           gen_12_cmp_pReg_6,gen_12_cmp_pReg_5,gen_12_cmp_pReg_4,
           gen_12_cmp_pReg_3,gen_12_cmp_pReg_2,gen_12_cmp_pReg_1,
           gen_12_cmp_pReg_0})) ;
    BinaryMux_33 gen_12_cmp_MuxCmp (.a ({working,working,gen_12_cmp_pReg_30,
                 gen_12_cmp_pReg_29,gen_12_cmp_pReg_28,gen_12_cmp_pReg_27,
                 gen_12_cmp_pReg_26,gen_12_cmp_pReg_25,gen_12_cmp_pReg_24,
                 gen_12_cmp_pReg_23,gen_12_cmp_pReg_22,gen_12_cmp_pReg_21,
                 gen_12_cmp_pReg_20,gen_12_cmp_pReg_19,gen_12_cmp_pReg_18,
                 gen_12_cmp_pReg_17,gen_12_cmp_pReg_16,gen_12_cmp_pReg_15,
                 gen_12_cmp_pReg_14,gen_12_cmp_pReg_13,gen_12_cmp_pReg_12,
                 gen_12_cmp_pReg_11,gen_12_cmp_pReg_10,gen_12_cmp_pReg_9,
                 gen_12_cmp_pReg_8,gen_12_cmp_pReg_7,gen_12_cmp_pReg_6,
                 gen_12_cmp_pReg_5,gen_12_cmp_pReg_4,gen_12_cmp_pReg_3,
                 gen_12_cmp_pReg_2,gen_12_cmp_pReg_1,gen_12_cmp_pReg_0}), .b ({
                 working,working,working,working,working,working,working,working
                 ,working,working,working,working,working,working,working,
                 working,working,working,working,working,working,working,working
                 ,working,filter_12__7,filter_12__6,filter_12__5,filter_12__4,
                 filter_12__3,filter_12__2,filter_12__1,filter_12__0,working}), 
                 .sel (nx11181), .f ({\$dummy [62],\$dummy [63],
                 gen_12_cmp_pMux_30,gen_12_cmp_pMux_29,gen_12_cmp_pMux_28,
                 gen_12_cmp_pMux_27,gen_12_cmp_pMux_26,gen_12_cmp_pMux_25,
                 gen_12_cmp_pMux_24,gen_12_cmp_pMux_23,gen_12_cmp_pMux_22,
                 gen_12_cmp_pMux_21,gen_12_cmp_pMux_20,gen_12_cmp_pMux_19,
                 gen_12_cmp_pMux_18,gen_12_cmp_pMux_17,gen_12_cmp_pMux_16,
                 gen_12_cmp_pMux_15,gen_12_cmp_pMux_14,gen_12_cmp_pMux_13,
                 gen_12_cmp_pMux_12,gen_12_cmp_pMux_11,gen_12_cmp_pMux_10,
                 gen_12_cmp_pMux_9,gen_12_cmp_pMux_8,gen_12_cmp_pMux_7,
                 gen_12_cmp_pMux_6,gen_12_cmp_pMux_5,gen_12_cmp_pMux_4,
                 gen_12_cmp_pMux_3,gen_12_cmp_pMux_2,gen_12_cmp_pMux_1,
                 gen_12_cmp_pMux_0})) ;
    NBitAdder_24 gen_12_cmp_BSCmp_AdderCmp (.a ({working,working,
                 gen_12_cmp_pMux_30,gen_12_cmp_pMux_29,gen_12_cmp_pMux_28,
                 gen_12_cmp_pMux_27,gen_12_cmp_pMux_26,gen_12_cmp_pMux_25,
                 gen_12_cmp_pMux_24,gen_12_cmp_pMux_23,gen_12_cmp_pMux_22,
                 gen_12_cmp_pMux_21,gen_12_cmp_pMux_20,gen_12_cmp_pMux_19,
                 gen_12_cmp_pMux_18,gen_12_cmp_pMux_17,gen_12_cmp_pMux_16,
                 gen_12_cmp_pMux_15,gen_12_cmp_pMux_14,gen_12_cmp_pMux_13,
                 gen_12_cmp_pMux_12,gen_12_cmp_pMux_11,gen_12_cmp_pMux_10,
                 gen_12_cmp_pMux_9}), .b ({nx9847,nx9847,nx9845,nx9853,nx9851,
                 nx9849,nx9847,nx9845,gen_12_cmp_BSCmp_op2_15,
                 gen_12_cmp_BSCmp_op2_14,gen_12_cmp_BSCmp_op2_13,
                 gen_12_cmp_BSCmp_op2_12,gen_12_cmp_BSCmp_op2_11,
                 gen_12_cmp_BSCmp_op2_10,gen_12_cmp_BSCmp_op2_9,
                 gen_12_cmp_BSCmp_op2_8,gen_12_cmp_BSCmp_op2_7,
                 gen_12_cmp_BSCmp_op2_6,gen_12_cmp_BSCmp_op2_5,
                 gen_12_cmp_BSCmp_op2_4,gen_12_cmp_BSCmp_op2_3,
                 gen_12_cmp_BSCmp_op2_2,gen_12_cmp_BSCmp_op2_1,
                 gen_12_cmp_BSCmp_op2_0}), .carryIn (gen_12_cmp_BSCmp_carryIn), 
                 .sum ({gen_12_cmp_pBs_30,gen_12_cmp_pBs_29,gen_12_cmp_pBs_28,
                 gen_12_cmp_pBs_27,gen_12_cmp_pBs_26,gen_12_cmp_pBs_25,
                 gen_12_cmp_pBs_24,gen_12_cmp_pBs_23,outputs_12__15,
                 outputs_12__14,outputs_12__13,outputs_12__12,outputs_12__11,
                 outputs_12__10,outputs_12__9,outputs_12__8,outputs_12__7,
                 outputs_12__6,outputs_12__5,outputs_12__4,outputs_12__3,
                 outputs_12__2,outputs_12__1,outputs_12__0}), .carryOut (
                 \$dummy [64])) ;
    Reg_33 gen_11_cmp_pRegCmp (.D ({working,working,gen_11_cmp_pBs_30,
           gen_11_cmp_pBs_29,gen_11_cmp_pBs_28,gen_11_cmp_pBs_27,
           gen_11_cmp_pBs_26,gen_11_cmp_pBs_25,gen_11_cmp_pBs_24,
           gen_11_cmp_pBs_23,outputs_11__15,outputs_11__14,outputs_11__13,
           outputs_11__12,outputs_11__11,outputs_11__10,outputs_11__9,
           outputs_11__8,outputs_11__7,outputs_11__6,outputs_11__5,outputs_11__4
           ,outputs_11__3,outputs_11__2,outputs_11__1,outputs_11__0,
           gen_11_cmp_pMux_8,gen_11_cmp_pMux_7,gen_11_cmp_pMux_6,
           gen_11_cmp_pMux_5,gen_11_cmp_pMux_4,gen_11_cmp_pMux_3,nx9555}), .en (
           nx9377), .clk (nx9393), .rst (rst), .Q ({\$dummy [65],\$dummy [66],
           gen_11_cmp_pReg_30,gen_11_cmp_pReg_29,gen_11_cmp_pReg_28,
           gen_11_cmp_pReg_27,gen_11_cmp_pReg_26,gen_11_cmp_pReg_25,
           gen_11_cmp_pReg_24,gen_11_cmp_pReg_23,gen_11_cmp_pReg_22,
           gen_11_cmp_pReg_21,gen_11_cmp_pReg_20,gen_11_cmp_pReg_19,
           gen_11_cmp_pReg_18,gen_11_cmp_pReg_17,gen_11_cmp_pReg_16,
           gen_11_cmp_pReg_15,gen_11_cmp_pReg_14,gen_11_cmp_pReg_13,
           gen_11_cmp_pReg_12,gen_11_cmp_pReg_11,gen_11_cmp_pReg_10,
           gen_11_cmp_pReg_9,gen_11_cmp_pReg_8,gen_11_cmp_pReg_7,
           gen_11_cmp_pReg_6,gen_11_cmp_pReg_5,gen_11_cmp_pReg_4,
           gen_11_cmp_pReg_3,gen_11_cmp_pReg_2,gen_11_cmp_pReg_1,
           gen_11_cmp_pReg_0})) ;
    BinaryMux_33 gen_11_cmp_MuxCmp (.a ({working,working,gen_11_cmp_pReg_30,
                 gen_11_cmp_pReg_29,gen_11_cmp_pReg_28,gen_11_cmp_pReg_27,
                 gen_11_cmp_pReg_26,gen_11_cmp_pReg_25,gen_11_cmp_pReg_24,
                 gen_11_cmp_pReg_23,gen_11_cmp_pReg_22,gen_11_cmp_pReg_21,
                 gen_11_cmp_pReg_20,gen_11_cmp_pReg_19,gen_11_cmp_pReg_18,
                 gen_11_cmp_pReg_17,gen_11_cmp_pReg_16,gen_11_cmp_pReg_15,
                 gen_11_cmp_pReg_14,gen_11_cmp_pReg_13,gen_11_cmp_pReg_12,
                 gen_11_cmp_pReg_11,gen_11_cmp_pReg_10,gen_11_cmp_pReg_9,
                 gen_11_cmp_pReg_8,gen_11_cmp_pReg_7,gen_11_cmp_pReg_6,
                 gen_11_cmp_pReg_5,gen_11_cmp_pReg_4,gen_11_cmp_pReg_3,
                 gen_11_cmp_pReg_2,gen_11_cmp_pReg_1,gen_11_cmp_pReg_0}), .b ({
                 working,working,working,working,working,working,working,working
                 ,working,working,working,working,working,working,working,
                 working,working,working,working,working,working,working,working
                 ,working,filter_11__7,filter_11__6,filter_11__5,filter_11__4,
                 filter_11__3,filter_11__2,filter_11__1,filter_11__0,working}), 
                 .sel (nx11183), .f ({\$dummy [67],\$dummy [68],
                 gen_11_cmp_pMux_30,gen_11_cmp_pMux_29,gen_11_cmp_pMux_28,
                 gen_11_cmp_pMux_27,gen_11_cmp_pMux_26,gen_11_cmp_pMux_25,
                 gen_11_cmp_pMux_24,gen_11_cmp_pMux_23,gen_11_cmp_pMux_22,
                 gen_11_cmp_pMux_21,gen_11_cmp_pMux_20,gen_11_cmp_pMux_19,
                 gen_11_cmp_pMux_18,gen_11_cmp_pMux_17,gen_11_cmp_pMux_16,
                 gen_11_cmp_pMux_15,gen_11_cmp_pMux_14,gen_11_cmp_pMux_13,
                 gen_11_cmp_pMux_12,gen_11_cmp_pMux_11,gen_11_cmp_pMux_10,
                 gen_11_cmp_pMux_9,gen_11_cmp_pMux_8,gen_11_cmp_pMux_7,
                 gen_11_cmp_pMux_6,gen_11_cmp_pMux_5,gen_11_cmp_pMux_4,
                 gen_11_cmp_pMux_3,gen_11_cmp_pMux_2,gen_11_cmp_pMux_1,
                 gen_11_cmp_pMux_0})) ;
    NBitAdder_24 gen_11_cmp_BSCmp_AdderCmp (.a ({working,working,
                 gen_11_cmp_pMux_30,gen_11_cmp_pMux_29,gen_11_cmp_pMux_28,
                 gen_11_cmp_pMux_27,gen_11_cmp_pMux_26,gen_11_cmp_pMux_25,
                 gen_11_cmp_pMux_24,gen_11_cmp_pMux_23,gen_11_cmp_pMux_22,
                 gen_11_cmp_pMux_21,gen_11_cmp_pMux_20,gen_11_cmp_pMux_19,
                 gen_11_cmp_pMux_18,gen_11_cmp_pMux_17,gen_11_cmp_pMux_16,
                 gen_11_cmp_pMux_15,gen_11_cmp_pMux_14,gen_11_cmp_pMux_13,
                 gen_11_cmp_pMux_12,gen_11_cmp_pMux_11,gen_11_cmp_pMux_10,
                 gen_11_cmp_pMux_9}), .b ({nx9859,nx9859,nx9857,nx9865,nx9863,
                 nx9861,nx9859,nx9857,gen_11_cmp_BSCmp_op2_15,
                 gen_11_cmp_BSCmp_op2_14,gen_11_cmp_BSCmp_op2_13,
                 gen_11_cmp_BSCmp_op2_12,gen_11_cmp_BSCmp_op2_11,
                 gen_11_cmp_BSCmp_op2_10,gen_11_cmp_BSCmp_op2_9,
                 gen_11_cmp_BSCmp_op2_8,gen_11_cmp_BSCmp_op2_7,
                 gen_11_cmp_BSCmp_op2_6,gen_11_cmp_BSCmp_op2_5,
                 gen_11_cmp_BSCmp_op2_4,gen_11_cmp_BSCmp_op2_3,
                 gen_11_cmp_BSCmp_op2_2,gen_11_cmp_BSCmp_op2_1,
                 gen_11_cmp_BSCmp_op2_0}), .carryIn (gen_11_cmp_BSCmp_carryIn), 
                 .sum ({gen_11_cmp_pBs_30,gen_11_cmp_pBs_29,gen_11_cmp_pBs_28,
                 gen_11_cmp_pBs_27,gen_11_cmp_pBs_26,gen_11_cmp_pBs_25,
                 gen_11_cmp_pBs_24,gen_11_cmp_pBs_23,outputs_11__15,
                 outputs_11__14,outputs_11__13,outputs_11__12,outputs_11__11,
                 outputs_11__10,outputs_11__9,outputs_11__8,outputs_11__7,
                 outputs_11__6,outputs_11__5,outputs_11__4,outputs_11__3,
                 outputs_11__2,outputs_11__1,outputs_11__0}), .carryOut (
                 \$dummy [69])) ;
    Reg_33 gen_10_cmp_pRegCmp (.D ({working,working,gen_10_cmp_pBs_30,
           gen_10_cmp_pBs_29,gen_10_cmp_pBs_28,gen_10_cmp_pBs_27,
           gen_10_cmp_pBs_26,gen_10_cmp_pBs_25,gen_10_cmp_pBs_24,
           gen_10_cmp_pBs_23,outputs_10__15,outputs_10__14,outputs_10__13,
           outputs_10__12,outputs_10__11,outputs_10__10,outputs_10__9,
           outputs_10__8,outputs_10__7,outputs_10__6,outputs_10__5,outputs_10__4
           ,outputs_10__3,outputs_10__2,outputs_10__1,outputs_10__0,
           gen_10_cmp_pMux_8,gen_10_cmp_pMux_7,gen_10_cmp_pMux_6,
           gen_10_cmp_pMux_5,gen_10_cmp_pMux_4,gen_10_cmp_pMux_3,nx9567}), .en (
           nx11167), .clk (nx9395), .rst (rst), .Q ({\$dummy [70],\$dummy [71],
           gen_10_cmp_pReg_30,gen_10_cmp_pReg_29,gen_10_cmp_pReg_28,
           gen_10_cmp_pReg_27,gen_10_cmp_pReg_26,gen_10_cmp_pReg_25,
           gen_10_cmp_pReg_24,gen_10_cmp_pReg_23,gen_10_cmp_pReg_22,
           gen_10_cmp_pReg_21,gen_10_cmp_pReg_20,gen_10_cmp_pReg_19,
           gen_10_cmp_pReg_18,gen_10_cmp_pReg_17,gen_10_cmp_pReg_16,
           gen_10_cmp_pReg_15,gen_10_cmp_pReg_14,gen_10_cmp_pReg_13,
           gen_10_cmp_pReg_12,gen_10_cmp_pReg_11,gen_10_cmp_pReg_10,
           gen_10_cmp_pReg_9,gen_10_cmp_pReg_8,gen_10_cmp_pReg_7,
           gen_10_cmp_pReg_6,gen_10_cmp_pReg_5,gen_10_cmp_pReg_4,
           gen_10_cmp_pReg_3,gen_10_cmp_pReg_2,gen_10_cmp_pReg_1,
           gen_10_cmp_pReg_0})) ;
    BinaryMux_33 gen_10_cmp_MuxCmp (.a ({working,working,gen_10_cmp_pReg_30,
                 gen_10_cmp_pReg_29,gen_10_cmp_pReg_28,gen_10_cmp_pReg_27,
                 gen_10_cmp_pReg_26,gen_10_cmp_pReg_25,gen_10_cmp_pReg_24,
                 gen_10_cmp_pReg_23,gen_10_cmp_pReg_22,gen_10_cmp_pReg_21,
                 gen_10_cmp_pReg_20,gen_10_cmp_pReg_19,gen_10_cmp_pReg_18,
                 gen_10_cmp_pReg_17,gen_10_cmp_pReg_16,gen_10_cmp_pReg_15,
                 gen_10_cmp_pReg_14,gen_10_cmp_pReg_13,gen_10_cmp_pReg_12,
                 gen_10_cmp_pReg_11,gen_10_cmp_pReg_10,gen_10_cmp_pReg_9,
                 gen_10_cmp_pReg_8,gen_10_cmp_pReg_7,gen_10_cmp_pReg_6,
                 gen_10_cmp_pReg_5,gen_10_cmp_pReg_4,gen_10_cmp_pReg_3,
                 gen_10_cmp_pReg_2,gen_10_cmp_pReg_1,gen_10_cmp_pReg_0}), .b ({
                 working,working,working,working,working,working,working,working
                 ,working,working,working,working,working,working,working,
                 working,working,working,working,working,working,working,working
                 ,working,filter_10__7,filter_10__6,filter_10__5,filter_10__4,
                 filter_10__3,filter_10__2,filter_10__1,filter_10__0,working}), 
                 .sel (nx11185), .f ({\$dummy [72],\$dummy [73],
                 gen_10_cmp_pMux_30,gen_10_cmp_pMux_29,gen_10_cmp_pMux_28,
                 gen_10_cmp_pMux_27,gen_10_cmp_pMux_26,gen_10_cmp_pMux_25,
                 gen_10_cmp_pMux_24,gen_10_cmp_pMux_23,gen_10_cmp_pMux_22,
                 gen_10_cmp_pMux_21,gen_10_cmp_pMux_20,gen_10_cmp_pMux_19,
                 gen_10_cmp_pMux_18,gen_10_cmp_pMux_17,gen_10_cmp_pMux_16,
                 gen_10_cmp_pMux_15,gen_10_cmp_pMux_14,gen_10_cmp_pMux_13,
                 gen_10_cmp_pMux_12,gen_10_cmp_pMux_11,gen_10_cmp_pMux_10,
                 gen_10_cmp_pMux_9,gen_10_cmp_pMux_8,gen_10_cmp_pMux_7,
                 gen_10_cmp_pMux_6,gen_10_cmp_pMux_5,gen_10_cmp_pMux_4,
                 gen_10_cmp_pMux_3,gen_10_cmp_pMux_2,gen_10_cmp_pMux_1,
                 gen_10_cmp_pMux_0})) ;
    NBitAdder_24 gen_10_cmp_BSCmp_AdderCmp (.a ({working,working,
                 gen_10_cmp_pMux_30,gen_10_cmp_pMux_29,gen_10_cmp_pMux_28,
                 gen_10_cmp_pMux_27,gen_10_cmp_pMux_26,gen_10_cmp_pMux_25,
                 gen_10_cmp_pMux_24,gen_10_cmp_pMux_23,gen_10_cmp_pMux_22,
                 gen_10_cmp_pMux_21,gen_10_cmp_pMux_20,gen_10_cmp_pMux_19,
                 gen_10_cmp_pMux_18,gen_10_cmp_pMux_17,gen_10_cmp_pMux_16,
                 gen_10_cmp_pMux_15,gen_10_cmp_pMux_14,gen_10_cmp_pMux_13,
                 gen_10_cmp_pMux_12,gen_10_cmp_pMux_11,gen_10_cmp_pMux_10,
                 gen_10_cmp_pMux_9}), .b ({nx9871,nx9871,nx9869,nx9877,nx9875,
                 nx9873,nx9871,nx9869,gen_10_cmp_BSCmp_op2_15,
                 gen_10_cmp_BSCmp_op2_14,gen_10_cmp_BSCmp_op2_13,
                 gen_10_cmp_BSCmp_op2_12,gen_10_cmp_BSCmp_op2_11,
                 gen_10_cmp_BSCmp_op2_10,gen_10_cmp_BSCmp_op2_9,
                 gen_10_cmp_BSCmp_op2_8,gen_10_cmp_BSCmp_op2_7,
                 gen_10_cmp_BSCmp_op2_6,gen_10_cmp_BSCmp_op2_5,
                 gen_10_cmp_BSCmp_op2_4,gen_10_cmp_BSCmp_op2_3,
                 gen_10_cmp_BSCmp_op2_2,gen_10_cmp_BSCmp_op2_1,
                 gen_10_cmp_BSCmp_op2_0}), .carryIn (gen_10_cmp_BSCmp_carryIn), 
                 .sum ({gen_10_cmp_pBs_30,gen_10_cmp_pBs_29,gen_10_cmp_pBs_28,
                 gen_10_cmp_pBs_27,gen_10_cmp_pBs_26,gen_10_cmp_pBs_25,
                 gen_10_cmp_pBs_24,gen_10_cmp_pBs_23,outputs_10__15,
                 outputs_10__14,outputs_10__13,outputs_10__12,outputs_10__11,
                 outputs_10__10,outputs_10__9,outputs_10__8,outputs_10__7,
                 outputs_10__6,outputs_10__5,outputs_10__4,outputs_10__3,
                 outputs_10__2,outputs_10__1,outputs_10__0}), .carryOut (
                 \$dummy [74])) ;
    Reg_33 gen_9_cmp_pRegCmp (.D ({working,working,gen_9_cmp_pBs_30,
           gen_9_cmp_pBs_29,gen_9_cmp_pBs_28,gen_9_cmp_pBs_27,gen_9_cmp_pBs_26,
           gen_9_cmp_pBs_25,gen_9_cmp_pBs_24,gen_9_cmp_pBs_23,outputs_9__15,
           outputs_9__14,outputs_9__13,outputs_9__12,outputs_9__11,outputs_9__10
           ,outputs_9__9,outputs_9__8,outputs_9__7,outputs_9__6,outputs_9__5,
           outputs_9__4,outputs_9__3,outputs_9__2,outputs_9__1,outputs_9__0,
           gen_9_cmp_pMux_8,gen_9_cmp_pMux_7,gen_9_cmp_pMux_6,gen_9_cmp_pMux_5,
           gen_9_cmp_pMux_4,gen_9_cmp_pMux_3,nx9579}), .en (nx11167), .clk (
           nx9395), .rst (rst), .Q ({\$dummy [75],\$dummy [76],gen_9_cmp_pReg_30
           ,gen_9_cmp_pReg_29,gen_9_cmp_pReg_28,gen_9_cmp_pReg_27,
           gen_9_cmp_pReg_26,gen_9_cmp_pReg_25,gen_9_cmp_pReg_24,
           gen_9_cmp_pReg_23,gen_9_cmp_pReg_22,gen_9_cmp_pReg_21,
           gen_9_cmp_pReg_20,gen_9_cmp_pReg_19,gen_9_cmp_pReg_18,
           gen_9_cmp_pReg_17,gen_9_cmp_pReg_16,gen_9_cmp_pReg_15,
           gen_9_cmp_pReg_14,gen_9_cmp_pReg_13,gen_9_cmp_pReg_12,
           gen_9_cmp_pReg_11,gen_9_cmp_pReg_10,gen_9_cmp_pReg_9,gen_9_cmp_pReg_8
           ,gen_9_cmp_pReg_7,gen_9_cmp_pReg_6,gen_9_cmp_pReg_5,gen_9_cmp_pReg_4,
           gen_9_cmp_pReg_3,gen_9_cmp_pReg_2,gen_9_cmp_pReg_1,gen_9_cmp_pReg_0})
           ) ;
    BinaryMux_33 gen_9_cmp_MuxCmp (.a ({working,working,gen_9_cmp_pReg_30,
                 gen_9_cmp_pReg_29,gen_9_cmp_pReg_28,gen_9_cmp_pReg_27,
                 gen_9_cmp_pReg_26,gen_9_cmp_pReg_25,gen_9_cmp_pReg_24,
                 gen_9_cmp_pReg_23,gen_9_cmp_pReg_22,gen_9_cmp_pReg_21,
                 gen_9_cmp_pReg_20,gen_9_cmp_pReg_19,gen_9_cmp_pReg_18,
                 gen_9_cmp_pReg_17,gen_9_cmp_pReg_16,gen_9_cmp_pReg_15,
                 gen_9_cmp_pReg_14,gen_9_cmp_pReg_13,gen_9_cmp_pReg_12,
                 gen_9_cmp_pReg_11,gen_9_cmp_pReg_10,gen_9_cmp_pReg_9,
                 gen_9_cmp_pReg_8,gen_9_cmp_pReg_7,gen_9_cmp_pReg_6,
                 gen_9_cmp_pReg_5,gen_9_cmp_pReg_4,gen_9_cmp_pReg_3,
                 gen_9_cmp_pReg_2,gen_9_cmp_pReg_1,gen_9_cmp_pReg_0}), .b ({
                 working,working,working,working,working,working,working,working
                 ,working,working,working,working,working,working,working,
                 working,working,working,working,working,working,working,working
                 ,working,filter_9__7,filter_9__6,filter_9__5,filter_9__4,
                 filter_9__3,filter_9__2,filter_9__1,filter_9__0,working}), .sel (
                 nx11185), .f ({\$dummy [77],\$dummy [78],gen_9_cmp_pMux_30,
                 gen_9_cmp_pMux_29,gen_9_cmp_pMux_28,gen_9_cmp_pMux_27,
                 gen_9_cmp_pMux_26,gen_9_cmp_pMux_25,gen_9_cmp_pMux_24,
                 gen_9_cmp_pMux_23,gen_9_cmp_pMux_22,gen_9_cmp_pMux_21,
                 gen_9_cmp_pMux_20,gen_9_cmp_pMux_19,gen_9_cmp_pMux_18,
                 gen_9_cmp_pMux_17,gen_9_cmp_pMux_16,gen_9_cmp_pMux_15,
                 gen_9_cmp_pMux_14,gen_9_cmp_pMux_13,gen_9_cmp_pMux_12,
                 gen_9_cmp_pMux_11,gen_9_cmp_pMux_10,gen_9_cmp_pMux_9,
                 gen_9_cmp_pMux_8,gen_9_cmp_pMux_7,gen_9_cmp_pMux_6,
                 gen_9_cmp_pMux_5,gen_9_cmp_pMux_4,gen_9_cmp_pMux_3,
                 gen_9_cmp_pMux_2,gen_9_cmp_pMux_1,gen_9_cmp_pMux_0})) ;
    NBitAdder_24 gen_9_cmp_BSCmp_AdderCmp (.a ({working,working,
                 gen_9_cmp_pMux_30,gen_9_cmp_pMux_29,gen_9_cmp_pMux_28,
                 gen_9_cmp_pMux_27,gen_9_cmp_pMux_26,gen_9_cmp_pMux_25,
                 gen_9_cmp_pMux_24,gen_9_cmp_pMux_23,gen_9_cmp_pMux_22,
                 gen_9_cmp_pMux_21,gen_9_cmp_pMux_20,gen_9_cmp_pMux_19,
                 gen_9_cmp_pMux_18,gen_9_cmp_pMux_17,gen_9_cmp_pMux_16,
                 gen_9_cmp_pMux_15,gen_9_cmp_pMux_14,gen_9_cmp_pMux_13,
                 gen_9_cmp_pMux_12,gen_9_cmp_pMux_11,gen_9_cmp_pMux_10,
                 gen_9_cmp_pMux_9}), .b ({nx9883,nx9883,nx9881,nx9889,nx9887,
                 nx9885,nx9883,nx9881,gen_9_cmp_BSCmp_op2_15,
                 gen_9_cmp_BSCmp_op2_14,gen_9_cmp_BSCmp_op2_13,
                 gen_9_cmp_BSCmp_op2_12,gen_9_cmp_BSCmp_op2_11,
                 gen_9_cmp_BSCmp_op2_10,gen_9_cmp_BSCmp_op2_9,
                 gen_9_cmp_BSCmp_op2_8,gen_9_cmp_BSCmp_op2_7,
                 gen_9_cmp_BSCmp_op2_6,gen_9_cmp_BSCmp_op2_5,
                 gen_9_cmp_BSCmp_op2_4,gen_9_cmp_BSCmp_op2_3,
                 gen_9_cmp_BSCmp_op2_2,gen_9_cmp_BSCmp_op2_1,
                 gen_9_cmp_BSCmp_op2_0}), .carryIn (gen_9_cmp_BSCmp_carryIn), .sum (
                 {gen_9_cmp_pBs_30,gen_9_cmp_pBs_29,gen_9_cmp_pBs_28,
                 gen_9_cmp_pBs_27,gen_9_cmp_pBs_26,gen_9_cmp_pBs_25,
                 gen_9_cmp_pBs_24,gen_9_cmp_pBs_23,outputs_9__15,outputs_9__14,
                 outputs_9__13,outputs_9__12,outputs_9__11,outputs_9__10,
                 outputs_9__9,outputs_9__8,outputs_9__7,outputs_9__6,
                 outputs_9__5,outputs_9__4,outputs_9__3,outputs_9__2,
                 outputs_9__1,outputs_9__0}), .carryOut (\$dummy [79])) ;
    Reg_33 gen_8_cmp_pRegCmp (.D ({working,working,gen_8_cmp_pBs_30,
           gen_8_cmp_pBs_29,gen_8_cmp_pBs_28,gen_8_cmp_pBs_27,gen_8_cmp_pBs_26,
           gen_8_cmp_pBs_25,gen_8_cmp_pBs_24,gen_8_cmp_pBs_23,outputs_8__15,
           outputs_8__14,outputs_8__13,outputs_8__12,outputs_8__11,outputs_8__10
           ,outputs_8__9,outputs_8__8,outputs_8__7,outputs_8__6,outputs_8__5,
           outputs_8__4,outputs_8__3,outputs_8__2,outputs_8__1,outputs_8__0,
           gen_8_cmp_pMux_8,gen_8_cmp_pMux_7,gen_8_cmp_pMux_6,gen_8_cmp_pMux_5,
           gen_8_cmp_pMux_4,gen_8_cmp_pMux_3,nx9591}), .en (nx11167), .clk (
           nx9395), .rst (rst), .Q ({\$dummy [80],\$dummy [81],gen_8_cmp_pReg_30
           ,gen_8_cmp_pReg_29,gen_8_cmp_pReg_28,gen_8_cmp_pReg_27,
           gen_8_cmp_pReg_26,gen_8_cmp_pReg_25,gen_8_cmp_pReg_24,
           gen_8_cmp_pReg_23,gen_8_cmp_pReg_22,gen_8_cmp_pReg_21,
           gen_8_cmp_pReg_20,gen_8_cmp_pReg_19,gen_8_cmp_pReg_18,
           gen_8_cmp_pReg_17,gen_8_cmp_pReg_16,gen_8_cmp_pReg_15,
           gen_8_cmp_pReg_14,gen_8_cmp_pReg_13,gen_8_cmp_pReg_12,
           gen_8_cmp_pReg_11,gen_8_cmp_pReg_10,gen_8_cmp_pReg_9,gen_8_cmp_pReg_8
           ,gen_8_cmp_pReg_7,gen_8_cmp_pReg_6,gen_8_cmp_pReg_5,gen_8_cmp_pReg_4,
           gen_8_cmp_pReg_3,gen_8_cmp_pReg_2,gen_8_cmp_pReg_1,gen_8_cmp_pReg_0})
           ) ;
    BinaryMux_33 gen_8_cmp_MuxCmp (.a ({working,working,gen_8_cmp_pReg_30,
                 gen_8_cmp_pReg_29,gen_8_cmp_pReg_28,gen_8_cmp_pReg_27,
                 gen_8_cmp_pReg_26,gen_8_cmp_pReg_25,gen_8_cmp_pReg_24,
                 gen_8_cmp_pReg_23,gen_8_cmp_pReg_22,gen_8_cmp_pReg_21,
                 gen_8_cmp_pReg_20,gen_8_cmp_pReg_19,gen_8_cmp_pReg_18,
                 gen_8_cmp_pReg_17,gen_8_cmp_pReg_16,gen_8_cmp_pReg_15,
                 gen_8_cmp_pReg_14,gen_8_cmp_pReg_13,gen_8_cmp_pReg_12,
                 gen_8_cmp_pReg_11,gen_8_cmp_pReg_10,gen_8_cmp_pReg_9,
                 gen_8_cmp_pReg_8,gen_8_cmp_pReg_7,gen_8_cmp_pReg_6,
                 gen_8_cmp_pReg_5,gen_8_cmp_pReg_4,gen_8_cmp_pReg_3,
                 gen_8_cmp_pReg_2,gen_8_cmp_pReg_1,gen_8_cmp_pReg_0}), .b ({
                 working,working,working,working,working,working,working,working
                 ,working,working,working,working,working,working,working,
                 working,working,working,working,working,working,working,working
                 ,working,filter_8__7,filter_8__6,filter_8__5,filter_8__4,
                 filter_8__3,filter_8__2,filter_8__1,filter_8__0,working}), .sel (
                 nx11185), .f ({\$dummy [82],\$dummy [83],gen_8_cmp_pMux_30,
                 gen_8_cmp_pMux_29,gen_8_cmp_pMux_28,gen_8_cmp_pMux_27,
                 gen_8_cmp_pMux_26,gen_8_cmp_pMux_25,gen_8_cmp_pMux_24,
                 gen_8_cmp_pMux_23,gen_8_cmp_pMux_22,gen_8_cmp_pMux_21,
                 gen_8_cmp_pMux_20,gen_8_cmp_pMux_19,gen_8_cmp_pMux_18,
                 gen_8_cmp_pMux_17,gen_8_cmp_pMux_16,gen_8_cmp_pMux_15,
                 gen_8_cmp_pMux_14,gen_8_cmp_pMux_13,gen_8_cmp_pMux_12,
                 gen_8_cmp_pMux_11,gen_8_cmp_pMux_10,gen_8_cmp_pMux_9,
                 gen_8_cmp_pMux_8,gen_8_cmp_pMux_7,gen_8_cmp_pMux_6,
                 gen_8_cmp_pMux_5,gen_8_cmp_pMux_4,gen_8_cmp_pMux_3,
                 gen_8_cmp_pMux_2,gen_8_cmp_pMux_1,gen_8_cmp_pMux_0})) ;
    NBitAdder_24 gen_8_cmp_BSCmp_AdderCmp (.a ({working,working,
                 gen_8_cmp_pMux_30,gen_8_cmp_pMux_29,gen_8_cmp_pMux_28,
                 gen_8_cmp_pMux_27,gen_8_cmp_pMux_26,gen_8_cmp_pMux_25,
                 gen_8_cmp_pMux_24,gen_8_cmp_pMux_23,gen_8_cmp_pMux_22,
                 gen_8_cmp_pMux_21,gen_8_cmp_pMux_20,gen_8_cmp_pMux_19,
                 gen_8_cmp_pMux_18,gen_8_cmp_pMux_17,gen_8_cmp_pMux_16,
                 gen_8_cmp_pMux_15,gen_8_cmp_pMux_14,gen_8_cmp_pMux_13,
                 gen_8_cmp_pMux_12,gen_8_cmp_pMux_11,gen_8_cmp_pMux_10,
                 gen_8_cmp_pMux_9}), .b ({nx9895,nx9895,nx9893,nx9901,nx9899,
                 nx9897,nx9895,nx9893,gen_8_cmp_BSCmp_op2_15,
                 gen_8_cmp_BSCmp_op2_14,gen_8_cmp_BSCmp_op2_13,
                 gen_8_cmp_BSCmp_op2_12,gen_8_cmp_BSCmp_op2_11,
                 gen_8_cmp_BSCmp_op2_10,gen_8_cmp_BSCmp_op2_9,
                 gen_8_cmp_BSCmp_op2_8,gen_8_cmp_BSCmp_op2_7,
                 gen_8_cmp_BSCmp_op2_6,gen_8_cmp_BSCmp_op2_5,
                 gen_8_cmp_BSCmp_op2_4,gen_8_cmp_BSCmp_op2_3,
                 gen_8_cmp_BSCmp_op2_2,gen_8_cmp_BSCmp_op2_1,
                 gen_8_cmp_BSCmp_op2_0}), .carryIn (gen_8_cmp_BSCmp_carryIn), .sum (
                 {gen_8_cmp_pBs_30,gen_8_cmp_pBs_29,gen_8_cmp_pBs_28,
                 gen_8_cmp_pBs_27,gen_8_cmp_pBs_26,gen_8_cmp_pBs_25,
                 gen_8_cmp_pBs_24,gen_8_cmp_pBs_23,outputs_8__15,outputs_8__14,
                 outputs_8__13,outputs_8__12,outputs_8__11,outputs_8__10,
                 outputs_8__9,outputs_8__8,outputs_8__7,outputs_8__6,
                 outputs_8__5,outputs_8__4,outputs_8__3,outputs_8__2,
                 outputs_8__1,outputs_8__0}), .carryOut (\$dummy [84])) ;
    Reg_33 gen_7_cmp_pRegCmp (.D ({working,working,gen_7_cmp_pBs_30,
           gen_7_cmp_pBs_29,gen_7_cmp_pBs_28,gen_7_cmp_pBs_27,gen_7_cmp_pBs_26,
           gen_7_cmp_pBs_25,gen_7_cmp_pBs_24,gen_7_cmp_pBs_23,outputs_7__15,
           outputs_7__14,outputs_7__13,outputs_7__12,outputs_7__11,outputs_7__10
           ,outputs_7__9,outputs_7__8,outputs_7__7,outputs_7__6,outputs_7__5,
           outputs_7__4,outputs_7__3,outputs_7__2,outputs_7__1,outputs_7__0,
           gen_7_cmp_pMux_8,gen_7_cmp_pMux_7,gen_7_cmp_pMux_6,gen_7_cmp_pMux_5,
           gen_7_cmp_pMux_4,gen_7_cmp_pMux_3,nx9603}), .en (nx11169), .clk (
           nx9395), .rst (rst), .Q ({\$dummy [85],\$dummy [86],gen_7_cmp_pReg_30
           ,gen_7_cmp_pReg_29,gen_7_cmp_pReg_28,gen_7_cmp_pReg_27,
           gen_7_cmp_pReg_26,gen_7_cmp_pReg_25,gen_7_cmp_pReg_24,
           gen_7_cmp_pReg_23,gen_7_cmp_pReg_22,gen_7_cmp_pReg_21,
           gen_7_cmp_pReg_20,gen_7_cmp_pReg_19,gen_7_cmp_pReg_18,
           gen_7_cmp_pReg_17,gen_7_cmp_pReg_16,gen_7_cmp_pReg_15,
           gen_7_cmp_pReg_14,gen_7_cmp_pReg_13,gen_7_cmp_pReg_12,
           gen_7_cmp_pReg_11,gen_7_cmp_pReg_10,gen_7_cmp_pReg_9,gen_7_cmp_pReg_8
           ,gen_7_cmp_pReg_7,gen_7_cmp_pReg_6,gen_7_cmp_pReg_5,gen_7_cmp_pReg_4,
           gen_7_cmp_pReg_3,gen_7_cmp_pReg_2,gen_7_cmp_pReg_1,gen_7_cmp_pReg_0})
           ) ;
    BinaryMux_33 gen_7_cmp_MuxCmp (.a ({working,working,gen_7_cmp_pReg_30,
                 gen_7_cmp_pReg_29,gen_7_cmp_pReg_28,gen_7_cmp_pReg_27,
                 gen_7_cmp_pReg_26,gen_7_cmp_pReg_25,gen_7_cmp_pReg_24,
                 gen_7_cmp_pReg_23,gen_7_cmp_pReg_22,gen_7_cmp_pReg_21,
                 gen_7_cmp_pReg_20,gen_7_cmp_pReg_19,gen_7_cmp_pReg_18,
                 gen_7_cmp_pReg_17,gen_7_cmp_pReg_16,gen_7_cmp_pReg_15,
                 gen_7_cmp_pReg_14,gen_7_cmp_pReg_13,gen_7_cmp_pReg_12,
                 gen_7_cmp_pReg_11,gen_7_cmp_pReg_10,gen_7_cmp_pReg_9,
                 gen_7_cmp_pReg_8,gen_7_cmp_pReg_7,gen_7_cmp_pReg_6,
                 gen_7_cmp_pReg_5,gen_7_cmp_pReg_4,gen_7_cmp_pReg_3,
                 gen_7_cmp_pReg_2,gen_7_cmp_pReg_1,gen_7_cmp_pReg_0}), .b ({
                 working,working,working,working,working,working,working,working
                 ,working,working,working,working,working,working,working,
                 working,working,working,working,working,working,working,working
                 ,working,filter_7__7,filter_7__6,filter_7__5,filter_7__4,
                 filter_7__3,filter_7__2,filter_7__1,filter_7__0,working}), .sel (
                 nx11187), .f ({\$dummy [87],\$dummy [88],gen_7_cmp_pMux_30,
                 gen_7_cmp_pMux_29,gen_7_cmp_pMux_28,gen_7_cmp_pMux_27,
                 gen_7_cmp_pMux_26,gen_7_cmp_pMux_25,gen_7_cmp_pMux_24,
                 gen_7_cmp_pMux_23,gen_7_cmp_pMux_22,gen_7_cmp_pMux_21,
                 gen_7_cmp_pMux_20,gen_7_cmp_pMux_19,gen_7_cmp_pMux_18,
                 gen_7_cmp_pMux_17,gen_7_cmp_pMux_16,gen_7_cmp_pMux_15,
                 gen_7_cmp_pMux_14,gen_7_cmp_pMux_13,gen_7_cmp_pMux_12,
                 gen_7_cmp_pMux_11,gen_7_cmp_pMux_10,gen_7_cmp_pMux_9,
                 gen_7_cmp_pMux_8,gen_7_cmp_pMux_7,gen_7_cmp_pMux_6,
                 gen_7_cmp_pMux_5,gen_7_cmp_pMux_4,gen_7_cmp_pMux_3,
                 gen_7_cmp_pMux_2,gen_7_cmp_pMux_1,gen_7_cmp_pMux_0})) ;
    NBitAdder_24 gen_7_cmp_BSCmp_AdderCmp (.a ({working,working,
                 gen_7_cmp_pMux_30,gen_7_cmp_pMux_29,gen_7_cmp_pMux_28,
                 gen_7_cmp_pMux_27,gen_7_cmp_pMux_26,gen_7_cmp_pMux_25,
                 gen_7_cmp_pMux_24,gen_7_cmp_pMux_23,gen_7_cmp_pMux_22,
                 gen_7_cmp_pMux_21,gen_7_cmp_pMux_20,gen_7_cmp_pMux_19,
                 gen_7_cmp_pMux_18,gen_7_cmp_pMux_17,gen_7_cmp_pMux_16,
                 gen_7_cmp_pMux_15,gen_7_cmp_pMux_14,gen_7_cmp_pMux_13,
                 gen_7_cmp_pMux_12,gen_7_cmp_pMux_11,gen_7_cmp_pMux_10,
                 gen_7_cmp_pMux_9}), .b ({nx9907,nx9907,nx9905,nx9913,nx9911,
                 nx9909,nx9907,nx9905,gen_7_cmp_BSCmp_op2_15,
                 gen_7_cmp_BSCmp_op2_14,gen_7_cmp_BSCmp_op2_13,
                 gen_7_cmp_BSCmp_op2_12,gen_7_cmp_BSCmp_op2_11,
                 gen_7_cmp_BSCmp_op2_10,gen_7_cmp_BSCmp_op2_9,
                 gen_7_cmp_BSCmp_op2_8,gen_7_cmp_BSCmp_op2_7,
                 gen_7_cmp_BSCmp_op2_6,gen_7_cmp_BSCmp_op2_5,
                 gen_7_cmp_BSCmp_op2_4,gen_7_cmp_BSCmp_op2_3,
                 gen_7_cmp_BSCmp_op2_2,gen_7_cmp_BSCmp_op2_1,
                 gen_7_cmp_BSCmp_op2_0}), .carryIn (gen_7_cmp_BSCmp_carryIn), .sum (
                 {gen_7_cmp_pBs_30,gen_7_cmp_pBs_29,gen_7_cmp_pBs_28,
                 gen_7_cmp_pBs_27,gen_7_cmp_pBs_26,gen_7_cmp_pBs_25,
                 gen_7_cmp_pBs_24,gen_7_cmp_pBs_23,outputs_7__15,outputs_7__14,
                 outputs_7__13,outputs_7__12,outputs_7__11,outputs_7__10,
                 outputs_7__9,outputs_7__8,outputs_7__7,outputs_7__6,
                 outputs_7__5,outputs_7__4,outputs_7__3,outputs_7__2,
                 outputs_7__1,outputs_7__0}), .carryOut (\$dummy [89])) ;
    Reg_33 gen_6_cmp_pRegCmp (.D ({working,working,gen_6_cmp_pBs_30,
           gen_6_cmp_pBs_29,gen_6_cmp_pBs_28,gen_6_cmp_pBs_27,gen_6_cmp_pBs_26,
           gen_6_cmp_pBs_25,gen_6_cmp_pBs_24,gen_6_cmp_pBs_23,outputs_6__15,
           outputs_6__14,outputs_6__13,outputs_6__12,outputs_6__11,outputs_6__10
           ,outputs_6__9,outputs_6__8,outputs_6__7,outputs_6__6,outputs_6__5,
           outputs_6__4,outputs_6__3,outputs_6__2,outputs_6__1,outputs_6__0,
           gen_6_cmp_pMux_8,gen_6_cmp_pMux_7,gen_6_cmp_pMux_6,gen_6_cmp_pMux_5,
           gen_6_cmp_pMux_4,gen_6_cmp_pMux_3,nx9615}), .en (nx11169), .clk (
           nx9395), .rst (rst), .Q ({\$dummy [90],\$dummy [91],gen_6_cmp_pReg_30
           ,gen_6_cmp_pReg_29,gen_6_cmp_pReg_28,gen_6_cmp_pReg_27,
           gen_6_cmp_pReg_26,gen_6_cmp_pReg_25,gen_6_cmp_pReg_24,
           gen_6_cmp_pReg_23,gen_6_cmp_pReg_22,gen_6_cmp_pReg_21,
           gen_6_cmp_pReg_20,gen_6_cmp_pReg_19,gen_6_cmp_pReg_18,
           gen_6_cmp_pReg_17,gen_6_cmp_pReg_16,gen_6_cmp_pReg_15,
           gen_6_cmp_pReg_14,gen_6_cmp_pReg_13,gen_6_cmp_pReg_12,
           gen_6_cmp_pReg_11,gen_6_cmp_pReg_10,gen_6_cmp_pReg_9,gen_6_cmp_pReg_8
           ,gen_6_cmp_pReg_7,gen_6_cmp_pReg_6,gen_6_cmp_pReg_5,gen_6_cmp_pReg_4,
           gen_6_cmp_pReg_3,gen_6_cmp_pReg_2,gen_6_cmp_pReg_1,gen_6_cmp_pReg_0})
           ) ;
    BinaryMux_33 gen_6_cmp_MuxCmp (.a ({working,working,gen_6_cmp_pReg_30,
                 gen_6_cmp_pReg_29,gen_6_cmp_pReg_28,gen_6_cmp_pReg_27,
                 gen_6_cmp_pReg_26,gen_6_cmp_pReg_25,gen_6_cmp_pReg_24,
                 gen_6_cmp_pReg_23,gen_6_cmp_pReg_22,gen_6_cmp_pReg_21,
                 gen_6_cmp_pReg_20,gen_6_cmp_pReg_19,gen_6_cmp_pReg_18,
                 gen_6_cmp_pReg_17,gen_6_cmp_pReg_16,gen_6_cmp_pReg_15,
                 gen_6_cmp_pReg_14,gen_6_cmp_pReg_13,gen_6_cmp_pReg_12,
                 gen_6_cmp_pReg_11,gen_6_cmp_pReg_10,gen_6_cmp_pReg_9,
                 gen_6_cmp_pReg_8,gen_6_cmp_pReg_7,gen_6_cmp_pReg_6,
                 gen_6_cmp_pReg_5,gen_6_cmp_pReg_4,gen_6_cmp_pReg_3,
                 gen_6_cmp_pReg_2,gen_6_cmp_pReg_1,gen_6_cmp_pReg_0}), .b ({
                 working,working,working,working,working,working,working,working
                 ,working,working,working,working,working,working,working,
                 working,working,working,working,working,working,working,working
                 ,working,filter_6__7,filter_6__6,filter_6__5,filter_6__4,
                 filter_6__3,filter_6__2,filter_6__1,filter_6__0,working}), .sel (
                 nx11187), .f ({\$dummy [92],\$dummy [93],gen_6_cmp_pMux_30,
                 gen_6_cmp_pMux_29,gen_6_cmp_pMux_28,gen_6_cmp_pMux_27,
                 gen_6_cmp_pMux_26,gen_6_cmp_pMux_25,gen_6_cmp_pMux_24,
                 gen_6_cmp_pMux_23,gen_6_cmp_pMux_22,gen_6_cmp_pMux_21,
                 gen_6_cmp_pMux_20,gen_6_cmp_pMux_19,gen_6_cmp_pMux_18,
                 gen_6_cmp_pMux_17,gen_6_cmp_pMux_16,gen_6_cmp_pMux_15,
                 gen_6_cmp_pMux_14,gen_6_cmp_pMux_13,gen_6_cmp_pMux_12,
                 gen_6_cmp_pMux_11,gen_6_cmp_pMux_10,gen_6_cmp_pMux_9,
                 gen_6_cmp_pMux_8,gen_6_cmp_pMux_7,gen_6_cmp_pMux_6,
                 gen_6_cmp_pMux_5,gen_6_cmp_pMux_4,gen_6_cmp_pMux_3,
                 gen_6_cmp_pMux_2,gen_6_cmp_pMux_1,gen_6_cmp_pMux_0})) ;
    NBitAdder_24 gen_6_cmp_BSCmp_AdderCmp (.a ({working,working,
                 gen_6_cmp_pMux_30,gen_6_cmp_pMux_29,gen_6_cmp_pMux_28,
                 gen_6_cmp_pMux_27,gen_6_cmp_pMux_26,gen_6_cmp_pMux_25,
                 gen_6_cmp_pMux_24,gen_6_cmp_pMux_23,gen_6_cmp_pMux_22,
                 gen_6_cmp_pMux_21,gen_6_cmp_pMux_20,gen_6_cmp_pMux_19,
                 gen_6_cmp_pMux_18,gen_6_cmp_pMux_17,gen_6_cmp_pMux_16,
                 gen_6_cmp_pMux_15,gen_6_cmp_pMux_14,gen_6_cmp_pMux_13,
                 gen_6_cmp_pMux_12,gen_6_cmp_pMux_11,gen_6_cmp_pMux_10,
                 gen_6_cmp_pMux_9}), .b ({nx9919,nx9919,nx9917,nx9925,nx9923,
                 nx9921,nx9919,nx9917,gen_6_cmp_BSCmp_op2_15,
                 gen_6_cmp_BSCmp_op2_14,gen_6_cmp_BSCmp_op2_13,
                 gen_6_cmp_BSCmp_op2_12,gen_6_cmp_BSCmp_op2_11,
                 gen_6_cmp_BSCmp_op2_10,gen_6_cmp_BSCmp_op2_9,
                 gen_6_cmp_BSCmp_op2_8,gen_6_cmp_BSCmp_op2_7,
                 gen_6_cmp_BSCmp_op2_6,gen_6_cmp_BSCmp_op2_5,
                 gen_6_cmp_BSCmp_op2_4,gen_6_cmp_BSCmp_op2_3,
                 gen_6_cmp_BSCmp_op2_2,gen_6_cmp_BSCmp_op2_1,
                 gen_6_cmp_BSCmp_op2_0}), .carryIn (gen_6_cmp_BSCmp_carryIn), .sum (
                 {gen_6_cmp_pBs_30,gen_6_cmp_pBs_29,gen_6_cmp_pBs_28,
                 gen_6_cmp_pBs_27,gen_6_cmp_pBs_26,gen_6_cmp_pBs_25,
                 gen_6_cmp_pBs_24,gen_6_cmp_pBs_23,outputs_6__15,outputs_6__14,
                 outputs_6__13,outputs_6__12,outputs_6__11,outputs_6__10,
                 outputs_6__9,outputs_6__8,outputs_6__7,outputs_6__6,
                 outputs_6__5,outputs_6__4,outputs_6__3,outputs_6__2,
                 outputs_6__1,outputs_6__0}), .carryOut (\$dummy [94])) ;
    Reg_33 gen_5_cmp_pRegCmp (.D ({working,working,gen_5_cmp_pBs_30,
           gen_5_cmp_pBs_29,gen_5_cmp_pBs_28,gen_5_cmp_pBs_27,gen_5_cmp_pBs_26,
           gen_5_cmp_pBs_25,gen_5_cmp_pBs_24,gen_5_cmp_pBs_23,outputs_5__15,
           outputs_5__14,outputs_5__13,outputs_5__12,outputs_5__11,outputs_5__10
           ,outputs_5__9,outputs_5__8,outputs_5__7,outputs_5__6,outputs_5__5,
           outputs_5__4,outputs_5__3,outputs_5__2,outputs_5__1,outputs_5__0,
           gen_5_cmp_pMux_8,gen_5_cmp_pMux_7,gen_5_cmp_pMux_6,gen_5_cmp_pMux_5,
           gen_5_cmp_pMux_4,gen_5_cmp_pMux_3,nx9627}), .en (nx11169), .clk (
           nx9395), .rst (rst), .Q ({\$dummy [95],\$dummy [96],gen_5_cmp_pReg_30
           ,gen_5_cmp_pReg_29,gen_5_cmp_pReg_28,gen_5_cmp_pReg_27,
           gen_5_cmp_pReg_26,gen_5_cmp_pReg_25,gen_5_cmp_pReg_24,
           gen_5_cmp_pReg_23,gen_5_cmp_pReg_22,gen_5_cmp_pReg_21,
           gen_5_cmp_pReg_20,gen_5_cmp_pReg_19,gen_5_cmp_pReg_18,
           gen_5_cmp_pReg_17,gen_5_cmp_pReg_16,gen_5_cmp_pReg_15,
           gen_5_cmp_pReg_14,gen_5_cmp_pReg_13,gen_5_cmp_pReg_12,
           gen_5_cmp_pReg_11,gen_5_cmp_pReg_10,gen_5_cmp_pReg_9,gen_5_cmp_pReg_8
           ,gen_5_cmp_pReg_7,gen_5_cmp_pReg_6,gen_5_cmp_pReg_5,gen_5_cmp_pReg_4,
           gen_5_cmp_pReg_3,gen_5_cmp_pReg_2,gen_5_cmp_pReg_1,gen_5_cmp_pReg_0})
           ) ;
    BinaryMux_33 gen_5_cmp_MuxCmp (.a ({working,working,gen_5_cmp_pReg_30,
                 gen_5_cmp_pReg_29,gen_5_cmp_pReg_28,gen_5_cmp_pReg_27,
                 gen_5_cmp_pReg_26,gen_5_cmp_pReg_25,gen_5_cmp_pReg_24,
                 gen_5_cmp_pReg_23,gen_5_cmp_pReg_22,gen_5_cmp_pReg_21,
                 gen_5_cmp_pReg_20,gen_5_cmp_pReg_19,gen_5_cmp_pReg_18,
                 gen_5_cmp_pReg_17,gen_5_cmp_pReg_16,gen_5_cmp_pReg_15,
                 gen_5_cmp_pReg_14,gen_5_cmp_pReg_13,gen_5_cmp_pReg_12,
                 gen_5_cmp_pReg_11,gen_5_cmp_pReg_10,gen_5_cmp_pReg_9,
                 gen_5_cmp_pReg_8,gen_5_cmp_pReg_7,gen_5_cmp_pReg_6,
                 gen_5_cmp_pReg_5,gen_5_cmp_pReg_4,gen_5_cmp_pReg_3,
                 gen_5_cmp_pReg_2,gen_5_cmp_pReg_1,gen_5_cmp_pReg_0}), .b ({
                 working,working,working,working,working,working,working,working
                 ,working,working,working,working,working,working,working,
                 working,working,working,working,working,working,working,working
                 ,working,filter_5__7,filter_5__6,filter_5__5,filter_5__4,
                 filter_5__3,filter_5__2,filter_5__1,filter_5__0,working}), .sel (
                 nx11187), .f ({\$dummy [97],\$dummy [98],gen_5_cmp_pMux_30,
                 gen_5_cmp_pMux_29,gen_5_cmp_pMux_28,gen_5_cmp_pMux_27,
                 gen_5_cmp_pMux_26,gen_5_cmp_pMux_25,gen_5_cmp_pMux_24,
                 gen_5_cmp_pMux_23,gen_5_cmp_pMux_22,gen_5_cmp_pMux_21,
                 gen_5_cmp_pMux_20,gen_5_cmp_pMux_19,gen_5_cmp_pMux_18,
                 gen_5_cmp_pMux_17,gen_5_cmp_pMux_16,gen_5_cmp_pMux_15,
                 gen_5_cmp_pMux_14,gen_5_cmp_pMux_13,gen_5_cmp_pMux_12,
                 gen_5_cmp_pMux_11,gen_5_cmp_pMux_10,gen_5_cmp_pMux_9,
                 gen_5_cmp_pMux_8,gen_5_cmp_pMux_7,gen_5_cmp_pMux_6,
                 gen_5_cmp_pMux_5,gen_5_cmp_pMux_4,gen_5_cmp_pMux_3,
                 gen_5_cmp_pMux_2,gen_5_cmp_pMux_1,gen_5_cmp_pMux_0})) ;
    NBitAdder_24 gen_5_cmp_BSCmp_AdderCmp (.a ({working,working,
                 gen_5_cmp_pMux_30,gen_5_cmp_pMux_29,gen_5_cmp_pMux_28,
                 gen_5_cmp_pMux_27,gen_5_cmp_pMux_26,gen_5_cmp_pMux_25,
                 gen_5_cmp_pMux_24,gen_5_cmp_pMux_23,gen_5_cmp_pMux_22,
                 gen_5_cmp_pMux_21,gen_5_cmp_pMux_20,gen_5_cmp_pMux_19,
                 gen_5_cmp_pMux_18,gen_5_cmp_pMux_17,gen_5_cmp_pMux_16,
                 gen_5_cmp_pMux_15,gen_5_cmp_pMux_14,gen_5_cmp_pMux_13,
                 gen_5_cmp_pMux_12,gen_5_cmp_pMux_11,gen_5_cmp_pMux_10,
                 gen_5_cmp_pMux_9}), .b ({nx9931,nx9931,nx9929,nx9937,nx9935,
                 nx9933,nx9931,nx9929,gen_5_cmp_BSCmp_op2_15,
                 gen_5_cmp_BSCmp_op2_14,gen_5_cmp_BSCmp_op2_13,
                 gen_5_cmp_BSCmp_op2_12,gen_5_cmp_BSCmp_op2_11,
                 gen_5_cmp_BSCmp_op2_10,gen_5_cmp_BSCmp_op2_9,
                 gen_5_cmp_BSCmp_op2_8,gen_5_cmp_BSCmp_op2_7,
                 gen_5_cmp_BSCmp_op2_6,gen_5_cmp_BSCmp_op2_5,
                 gen_5_cmp_BSCmp_op2_4,gen_5_cmp_BSCmp_op2_3,
                 gen_5_cmp_BSCmp_op2_2,gen_5_cmp_BSCmp_op2_1,
                 gen_5_cmp_BSCmp_op2_0}), .carryIn (gen_5_cmp_BSCmp_carryIn), .sum (
                 {gen_5_cmp_pBs_30,gen_5_cmp_pBs_29,gen_5_cmp_pBs_28,
                 gen_5_cmp_pBs_27,gen_5_cmp_pBs_26,gen_5_cmp_pBs_25,
                 gen_5_cmp_pBs_24,gen_5_cmp_pBs_23,outputs_5__15,outputs_5__14,
                 outputs_5__13,outputs_5__12,outputs_5__11,outputs_5__10,
                 outputs_5__9,outputs_5__8,outputs_5__7,outputs_5__6,
                 outputs_5__5,outputs_5__4,outputs_5__3,outputs_5__2,
                 outputs_5__1,outputs_5__0}), .carryOut (\$dummy [99])) ;
    Reg_33 gen_4_cmp_pRegCmp (.D ({working,working,gen_4_cmp_pBs_30,
           gen_4_cmp_pBs_29,gen_4_cmp_pBs_28,gen_4_cmp_pBs_27,gen_4_cmp_pBs_26,
           gen_4_cmp_pBs_25,gen_4_cmp_pBs_24,gen_4_cmp_pBs_23,outputs_4__15,
           outputs_4__14,outputs_4__13,outputs_4__12,outputs_4__11,outputs_4__10
           ,outputs_4__9,outputs_4__8,outputs_4__7,outputs_4__6,outputs_4__5,
           outputs_4__4,outputs_4__3,outputs_4__2,outputs_4__1,outputs_4__0,
           gen_4_cmp_pMux_8,gen_4_cmp_pMux_7,gen_4_cmp_pMux_6,gen_4_cmp_pMux_5,
           gen_4_cmp_pMux_4,gen_4_cmp_pMux_3,nx9639}), .en (nx9379), .clk (
           nx9395), .rst (rst), .Q ({\$dummy [100],\$dummy [101],
           gen_4_cmp_pReg_30,gen_4_cmp_pReg_29,gen_4_cmp_pReg_28,
           gen_4_cmp_pReg_27,gen_4_cmp_pReg_26,gen_4_cmp_pReg_25,
           gen_4_cmp_pReg_24,gen_4_cmp_pReg_23,gen_4_cmp_pReg_22,
           gen_4_cmp_pReg_21,gen_4_cmp_pReg_20,gen_4_cmp_pReg_19,
           gen_4_cmp_pReg_18,gen_4_cmp_pReg_17,gen_4_cmp_pReg_16,
           gen_4_cmp_pReg_15,gen_4_cmp_pReg_14,gen_4_cmp_pReg_13,
           gen_4_cmp_pReg_12,gen_4_cmp_pReg_11,gen_4_cmp_pReg_10,
           gen_4_cmp_pReg_9,gen_4_cmp_pReg_8,gen_4_cmp_pReg_7,gen_4_cmp_pReg_6,
           gen_4_cmp_pReg_5,gen_4_cmp_pReg_4,gen_4_cmp_pReg_3,gen_4_cmp_pReg_2,
           gen_4_cmp_pReg_1,gen_4_cmp_pReg_0})) ;
    BinaryMux_33 gen_4_cmp_MuxCmp (.a ({working,working,gen_4_cmp_pReg_30,
                 gen_4_cmp_pReg_29,gen_4_cmp_pReg_28,gen_4_cmp_pReg_27,
                 gen_4_cmp_pReg_26,gen_4_cmp_pReg_25,gen_4_cmp_pReg_24,
                 gen_4_cmp_pReg_23,gen_4_cmp_pReg_22,gen_4_cmp_pReg_21,
                 gen_4_cmp_pReg_20,gen_4_cmp_pReg_19,gen_4_cmp_pReg_18,
                 gen_4_cmp_pReg_17,gen_4_cmp_pReg_16,gen_4_cmp_pReg_15,
                 gen_4_cmp_pReg_14,gen_4_cmp_pReg_13,gen_4_cmp_pReg_12,
                 gen_4_cmp_pReg_11,gen_4_cmp_pReg_10,gen_4_cmp_pReg_9,
                 gen_4_cmp_pReg_8,gen_4_cmp_pReg_7,gen_4_cmp_pReg_6,
                 gen_4_cmp_pReg_5,gen_4_cmp_pReg_4,gen_4_cmp_pReg_3,
                 gen_4_cmp_pReg_2,gen_4_cmp_pReg_1,gen_4_cmp_pReg_0}), .b ({
                 working,working,working,working,working,working,working,working
                 ,working,working,working,working,working,working,working,
                 working,working,working,working,working,working,working,working
                 ,working,filter_4__7,filter_4__6,filter_4__5,filter_4__4,
                 filter_4__3,filter_4__2,filter_4__1,filter_4__0,working}), .sel (
                 nx11189), .f ({\$dummy [102],\$dummy [103],gen_4_cmp_pMux_30,
                 gen_4_cmp_pMux_29,gen_4_cmp_pMux_28,gen_4_cmp_pMux_27,
                 gen_4_cmp_pMux_26,gen_4_cmp_pMux_25,gen_4_cmp_pMux_24,
                 gen_4_cmp_pMux_23,gen_4_cmp_pMux_22,gen_4_cmp_pMux_21,
                 gen_4_cmp_pMux_20,gen_4_cmp_pMux_19,gen_4_cmp_pMux_18,
                 gen_4_cmp_pMux_17,gen_4_cmp_pMux_16,gen_4_cmp_pMux_15,
                 gen_4_cmp_pMux_14,gen_4_cmp_pMux_13,gen_4_cmp_pMux_12,
                 gen_4_cmp_pMux_11,gen_4_cmp_pMux_10,gen_4_cmp_pMux_9,
                 gen_4_cmp_pMux_8,gen_4_cmp_pMux_7,gen_4_cmp_pMux_6,
                 gen_4_cmp_pMux_5,gen_4_cmp_pMux_4,gen_4_cmp_pMux_3,
                 gen_4_cmp_pMux_2,gen_4_cmp_pMux_1,gen_4_cmp_pMux_0})) ;
    NBitAdder_24 gen_4_cmp_BSCmp_AdderCmp (.a ({working,working,
                 gen_4_cmp_pMux_30,gen_4_cmp_pMux_29,gen_4_cmp_pMux_28,
                 gen_4_cmp_pMux_27,gen_4_cmp_pMux_26,gen_4_cmp_pMux_25,
                 gen_4_cmp_pMux_24,gen_4_cmp_pMux_23,gen_4_cmp_pMux_22,
                 gen_4_cmp_pMux_21,gen_4_cmp_pMux_20,gen_4_cmp_pMux_19,
                 gen_4_cmp_pMux_18,gen_4_cmp_pMux_17,gen_4_cmp_pMux_16,
                 gen_4_cmp_pMux_15,gen_4_cmp_pMux_14,gen_4_cmp_pMux_13,
                 gen_4_cmp_pMux_12,gen_4_cmp_pMux_11,gen_4_cmp_pMux_10,
                 gen_4_cmp_pMux_9}), .b ({nx9943,nx9943,nx9941,nx9949,nx9947,
                 nx9945,nx9943,nx9941,gen_4_cmp_BSCmp_op2_15,
                 gen_4_cmp_BSCmp_op2_14,gen_4_cmp_BSCmp_op2_13,
                 gen_4_cmp_BSCmp_op2_12,gen_4_cmp_BSCmp_op2_11,
                 gen_4_cmp_BSCmp_op2_10,gen_4_cmp_BSCmp_op2_9,
                 gen_4_cmp_BSCmp_op2_8,gen_4_cmp_BSCmp_op2_7,
                 gen_4_cmp_BSCmp_op2_6,gen_4_cmp_BSCmp_op2_5,
                 gen_4_cmp_BSCmp_op2_4,gen_4_cmp_BSCmp_op2_3,
                 gen_4_cmp_BSCmp_op2_2,gen_4_cmp_BSCmp_op2_1,
                 gen_4_cmp_BSCmp_op2_0}), .carryIn (gen_4_cmp_BSCmp_carryIn), .sum (
                 {gen_4_cmp_pBs_30,gen_4_cmp_pBs_29,gen_4_cmp_pBs_28,
                 gen_4_cmp_pBs_27,gen_4_cmp_pBs_26,gen_4_cmp_pBs_25,
                 gen_4_cmp_pBs_24,gen_4_cmp_pBs_23,outputs_4__15,outputs_4__14,
                 outputs_4__13,outputs_4__12,outputs_4__11,outputs_4__10,
                 outputs_4__9,outputs_4__8,outputs_4__7,outputs_4__6,
                 outputs_4__5,outputs_4__4,outputs_4__3,outputs_4__2,
                 outputs_4__1,outputs_4__0}), .carryOut (\$dummy [104])) ;
    Reg_33 gen_3_cmp_pRegCmp (.D ({working,working,gen_3_cmp_pBs_30,
           gen_3_cmp_pBs_29,gen_3_cmp_pBs_28,gen_3_cmp_pBs_27,gen_3_cmp_pBs_26,
           gen_3_cmp_pBs_25,gen_3_cmp_pBs_24,gen_3_cmp_pBs_23,outputs_3__15,
           outputs_3__14,outputs_3__13,outputs_3__12,outputs_3__11,outputs_3__10
           ,outputs_3__9,outputs_3__8,outputs_3__7,outputs_3__6,outputs_3__5,
           outputs_3__4,outputs_3__3,outputs_3__2,outputs_3__1,outputs_3__0,
           gen_3_cmp_pMux_8,gen_3_cmp_pMux_7,gen_3_cmp_pMux_6,gen_3_cmp_pMux_5,
           gen_3_cmp_pMux_4,gen_3_cmp_pMux_3,nx9651}), .en (nx11171), .clk (
           nx9397), .rst (rst), .Q ({\$dummy [105],\$dummy [106],
           gen_3_cmp_pReg_30,gen_3_cmp_pReg_29,gen_3_cmp_pReg_28,
           gen_3_cmp_pReg_27,gen_3_cmp_pReg_26,gen_3_cmp_pReg_25,
           gen_3_cmp_pReg_24,gen_3_cmp_pReg_23,gen_3_cmp_pReg_22,
           gen_3_cmp_pReg_21,gen_3_cmp_pReg_20,gen_3_cmp_pReg_19,
           gen_3_cmp_pReg_18,gen_3_cmp_pReg_17,gen_3_cmp_pReg_16,
           gen_3_cmp_pReg_15,gen_3_cmp_pReg_14,gen_3_cmp_pReg_13,
           gen_3_cmp_pReg_12,gen_3_cmp_pReg_11,gen_3_cmp_pReg_10,
           gen_3_cmp_pReg_9,gen_3_cmp_pReg_8,gen_3_cmp_pReg_7,gen_3_cmp_pReg_6,
           gen_3_cmp_pReg_5,gen_3_cmp_pReg_4,gen_3_cmp_pReg_3,gen_3_cmp_pReg_2,
           gen_3_cmp_pReg_1,gen_3_cmp_pReg_0})) ;
    BinaryMux_33 gen_3_cmp_MuxCmp (.a ({working,working,gen_3_cmp_pReg_30,
                 gen_3_cmp_pReg_29,gen_3_cmp_pReg_28,gen_3_cmp_pReg_27,
                 gen_3_cmp_pReg_26,gen_3_cmp_pReg_25,gen_3_cmp_pReg_24,
                 gen_3_cmp_pReg_23,gen_3_cmp_pReg_22,gen_3_cmp_pReg_21,
                 gen_3_cmp_pReg_20,gen_3_cmp_pReg_19,gen_3_cmp_pReg_18,
                 gen_3_cmp_pReg_17,gen_3_cmp_pReg_16,gen_3_cmp_pReg_15,
                 gen_3_cmp_pReg_14,gen_3_cmp_pReg_13,gen_3_cmp_pReg_12,
                 gen_3_cmp_pReg_11,gen_3_cmp_pReg_10,gen_3_cmp_pReg_9,
                 gen_3_cmp_pReg_8,gen_3_cmp_pReg_7,gen_3_cmp_pReg_6,
                 gen_3_cmp_pReg_5,gen_3_cmp_pReg_4,gen_3_cmp_pReg_3,
                 gen_3_cmp_pReg_2,gen_3_cmp_pReg_1,gen_3_cmp_pReg_0}), .b ({
                 working,working,working,working,working,working,working,working
                 ,working,working,working,working,working,working,working,
                 working,working,working,working,working,working,working,working
                 ,working,filter_3__7,filter_3__6,filter_3__5,filter_3__4,
                 filter_3__3,filter_3__2,filter_3__1,filter_3__0,working}), .sel (
                 nx11191), .f ({\$dummy [107],\$dummy [108],gen_3_cmp_pMux_30,
                 gen_3_cmp_pMux_29,gen_3_cmp_pMux_28,gen_3_cmp_pMux_27,
                 gen_3_cmp_pMux_26,gen_3_cmp_pMux_25,gen_3_cmp_pMux_24,
                 gen_3_cmp_pMux_23,gen_3_cmp_pMux_22,gen_3_cmp_pMux_21,
                 gen_3_cmp_pMux_20,gen_3_cmp_pMux_19,gen_3_cmp_pMux_18,
                 gen_3_cmp_pMux_17,gen_3_cmp_pMux_16,gen_3_cmp_pMux_15,
                 gen_3_cmp_pMux_14,gen_3_cmp_pMux_13,gen_3_cmp_pMux_12,
                 gen_3_cmp_pMux_11,gen_3_cmp_pMux_10,gen_3_cmp_pMux_9,
                 gen_3_cmp_pMux_8,gen_3_cmp_pMux_7,gen_3_cmp_pMux_6,
                 gen_3_cmp_pMux_5,gen_3_cmp_pMux_4,gen_3_cmp_pMux_3,
                 gen_3_cmp_pMux_2,gen_3_cmp_pMux_1,gen_3_cmp_pMux_0})) ;
    NBitAdder_24 gen_3_cmp_BSCmp_AdderCmp (.a ({working,working,
                 gen_3_cmp_pMux_30,gen_3_cmp_pMux_29,gen_3_cmp_pMux_28,
                 gen_3_cmp_pMux_27,gen_3_cmp_pMux_26,gen_3_cmp_pMux_25,
                 gen_3_cmp_pMux_24,gen_3_cmp_pMux_23,gen_3_cmp_pMux_22,
                 gen_3_cmp_pMux_21,gen_3_cmp_pMux_20,gen_3_cmp_pMux_19,
                 gen_3_cmp_pMux_18,gen_3_cmp_pMux_17,gen_3_cmp_pMux_16,
                 gen_3_cmp_pMux_15,gen_3_cmp_pMux_14,gen_3_cmp_pMux_13,
                 gen_3_cmp_pMux_12,gen_3_cmp_pMux_11,gen_3_cmp_pMux_10,
                 gen_3_cmp_pMux_9}), .b ({nx9955,nx9955,nx9953,nx9961,nx9959,
                 nx9957,nx9955,nx9953,gen_3_cmp_BSCmp_op2_15,
                 gen_3_cmp_BSCmp_op2_14,gen_3_cmp_BSCmp_op2_13,
                 gen_3_cmp_BSCmp_op2_12,gen_3_cmp_BSCmp_op2_11,
                 gen_3_cmp_BSCmp_op2_10,gen_3_cmp_BSCmp_op2_9,
                 gen_3_cmp_BSCmp_op2_8,gen_3_cmp_BSCmp_op2_7,
                 gen_3_cmp_BSCmp_op2_6,gen_3_cmp_BSCmp_op2_5,
                 gen_3_cmp_BSCmp_op2_4,gen_3_cmp_BSCmp_op2_3,
                 gen_3_cmp_BSCmp_op2_2,gen_3_cmp_BSCmp_op2_1,
                 gen_3_cmp_BSCmp_op2_0}), .carryIn (gen_3_cmp_BSCmp_carryIn), .sum (
                 {gen_3_cmp_pBs_30,gen_3_cmp_pBs_29,gen_3_cmp_pBs_28,
                 gen_3_cmp_pBs_27,gen_3_cmp_pBs_26,gen_3_cmp_pBs_25,
                 gen_3_cmp_pBs_24,gen_3_cmp_pBs_23,outputs_3__15,outputs_3__14,
                 outputs_3__13,outputs_3__12,outputs_3__11,outputs_3__10,
                 outputs_3__9,outputs_3__8,outputs_3__7,outputs_3__6,
                 outputs_3__5,outputs_3__4,outputs_3__3,outputs_3__2,
                 outputs_3__1,outputs_3__0}), .carryOut (\$dummy [109])) ;
    Reg_33 gen_2_cmp_pRegCmp (.D ({working,working,gen_2_cmp_pBs_30,
           gen_2_cmp_pBs_29,gen_2_cmp_pBs_28,gen_2_cmp_pBs_27,gen_2_cmp_pBs_26,
           gen_2_cmp_pBs_25,gen_2_cmp_pBs_24,gen_2_cmp_pBs_23,outputs_2__15,
           outputs_2__14,outputs_2__13,outputs_2__12,outputs_2__11,outputs_2__10
           ,outputs_2__9,outputs_2__8,outputs_2__7,outputs_2__6,outputs_2__5,
           outputs_2__4,outputs_2__3,outputs_2__2,outputs_2__1,outputs_2__0,
           gen_2_cmp_pMux_8,gen_2_cmp_pMux_7,gen_2_cmp_pMux_6,gen_2_cmp_pMux_5,
           gen_2_cmp_pMux_4,gen_2_cmp_pMux_3,nx9663}), .en (nx11171), .clk (
           nx9397), .rst (rst), .Q ({\$dummy [110],\$dummy [111],
           gen_2_cmp_pReg_30,gen_2_cmp_pReg_29,gen_2_cmp_pReg_28,
           gen_2_cmp_pReg_27,gen_2_cmp_pReg_26,gen_2_cmp_pReg_25,
           gen_2_cmp_pReg_24,gen_2_cmp_pReg_23,gen_2_cmp_pReg_22,
           gen_2_cmp_pReg_21,gen_2_cmp_pReg_20,gen_2_cmp_pReg_19,
           gen_2_cmp_pReg_18,gen_2_cmp_pReg_17,gen_2_cmp_pReg_16,
           gen_2_cmp_pReg_15,gen_2_cmp_pReg_14,gen_2_cmp_pReg_13,
           gen_2_cmp_pReg_12,gen_2_cmp_pReg_11,gen_2_cmp_pReg_10,
           gen_2_cmp_pReg_9,gen_2_cmp_pReg_8,gen_2_cmp_pReg_7,gen_2_cmp_pReg_6,
           gen_2_cmp_pReg_5,gen_2_cmp_pReg_4,gen_2_cmp_pReg_3,gen_2_cmp_pReg_2,
           gen_2_cmp_pReg_1,gen_2_cmp_pReg_0})) ;
    BinaryMux_33 gen_2_cmp_MuxCmp (.a ({working,working,gen_2_cmp_pReg_30,
                 gen_2_cmp_pReg_29,gen_2_cmp_pReg_28,gen_2_cmp_pReg_27,
                 gen_2_cmp_pReg_26,gen_2_cmp_pReg_25,gen_2_cmp_pReg_24,
                 gen_2_cmp_pReg_23,gen_2_cmp_pReg_22,gen_2_cmp_pReg_21,
                 gen_2_cmp_pReg_20,gen_2_cmp_pReg_19,gen_2_cmp_pReg_18,
                 gen_2_cmp_pReg_17,gen_2_cmp_pReg_16,gen_2_cmp_pReg_15,
                 gen_2_cmp_pReg_14,gen_2_cmp_pReg_13,gen_2_cmp_pReg_12,
                 gen_2_cmp_pReg_11,gen_2_cmp_pReg_10,gen_2_cmp_pReg_9,
                 gen_2_cmp_pReg_8,gen_2_cmp_pReg_7,gen_2_cmp_pReg_6,
                 gen_2_cmp_pReg_5,gen_2_cmp_pReg_4,gen_2_cmp_pReg_3,
                 gen_2_cmp_pReg_2,gen_2_cmp_pReg_1,gen_2_cmp_pReg_0}), .b ({
                 working,working,working,working,working,working,working,working
                 ,working,working,working,working,working,working,working,
                 working,working,working,working,working,working,working,working
                 ,working,filter_2__7,filter_2__6,filter_2__5,filter_2__4,
                 filter_2__3,filter_2__2,filter_2__1,filter_2__0,working}), .sel (
                 nx11191), .f ({\$dummy [112],\$dummy [113],gen_2_cmp_pMux_30,
                 gen_2_cmp_pMux_29,gen_2_cmp_pMux_28,gen_2_cmp_pMux_27,
                 gen_2_cmp_pMux_26,gen_2_cmp_pMux_25,gen_2_cmp_pMux_24,
                 gen_2_cmp_pMux_23,gen_2_cmp_pMux_22,gen_2_cmp_pMux_21,
                 gen_2_cmp_pMux_20,gen_2_cmp_pMux_19,gen_2_cmp_pMux_18,
                 gen_2_cmp_pMux_17,gen_2_cmp_pMux_16,gen_2_cmp_pMux_15,
                 gen_2_cmp_pMux_14,gen_2_cmp_pMux_13,gen_2_cmp_pMux_12,
                 gen_2_cmp_pMux_11,gen_2_cmp_pMux_10,gen_2_cmp_pMux_9,
                 gen_2_cmp_pMux_8,gen_2_cmp_pMux_7,gen_2_cmp_pMux_6,
                 gen_2_cmp_pMux_5,gen_2_cmp_pMux_4,gen_2_cmp_pMux_3,
                 gen_2_cmp_pMux_2,gen_2_cmp_pMux_1,gen_2_cmp_pMux_0})) ;
    NBitAdder_24 gen_2_cmp_BSCmp_AdderCmp (.a ({working,working,
                 gen_2_cmp_pMux_30,gen_2_cmp_pMux_29,gen_2_cmp_pMux_28,
                 gen_2_cmp_pMux_27,gen_2_cmp_pMux_26,gen_2_cmp_pMux_25,
                 gen_2_cmp_pMux_24,gen_2_cmp_pMux_23,gen_2_cmp_pMux_22,
                 gen_2_cmp_pMux_21,gen_2_cmp_pMux_20,gen_2_cmp_pMux_19,
                 gen_2_cmp_pMux_18,gen_2_cmp_pMux_17,gen_2_cmp_pMux_16,
                 gen_2_cmp_pMux_15,gen_2_cmp_pMux_14,gen_2_cmp_pMux_13,
                 gen_2_cmp_pMux_12,gen_2_cmp_pMux_11,gen_2_cmp_pMux_10,
                 gen_2_cmp_pMux_9}), .b ({nx9967,nx9967,nx9965,nx9973,nx9971,
                 nx9969,nx9967,nx9965,gen_2_cmp_BSCmp_op2_15,
                 gen_2_cmp_BSCmp_op2_14,gen_2_cmp_BSCmp_op2_13,
                 gen_2_cmp_BSCmp_op2_12,gen_2_cmp_BSCmp_op2_11,
                 gen_2_cmp_BSCmp_op2_10,gen_2_cmp_BSCmp_op2_9,
                 gen_2_cmp_BSCmp_op2_8,gen_2_cmp_BSCmp_op2_7,
                 gen_2_cmp_BSCmp_op2_6,gen_2_cmp_BSCmp_op2_5,
                 gen_2_cmp_BSCmp_op2_4,gen_2_cmp_BSCmp_op2_3,
                 gen_2_cmp_BSCmp_op2_2,gen_2_cmp_BSCmp_op2_1,
                 gen_2_cmp_BSCmp_op2_0}), .carryIn (gen_2_cmp_BSCmp_carryIn), .sum (
                 {gen_2_cmp_pBs_30,gen_2_cmp_pBs_29,gen_2_cmp_pBs_28,
                 gen_2_cmp_pBs_27,gen_2_cmp_pBs_26,gen_2_cmp_pBs_25,
                 gen_2_cmp_pBs_24,gen_2_cmp_pBs_23,outputs_2__15,outputs_2__14,
                 outputs_2__13,outputs_2__12,outputs_2__11,outputs_2__10,
                 outputs_2__9,outputs_2__8,outputs_2__7,outputs_2__6,
                 outputs_2__5,outputs_2__4,outputs_2__3,outputs_2__2,
                 outputs_2__1,outputs_2__0}), .carryOut (\$dummy [114])) ;
    Reg_33 gen_1_cmp_pRegCmp (.D ({working,working,gen_1_cmp_pBs_30,
           gen_1_cmp_pBs_29,gen_1_cmp_pBs_28,gen_1_cmp_pBs_27,gen_1_cmp_pBs_26,
           gen_1_cmp_pBs_25,gen_1_cmp_pBs_24,gen_1_cmp_pBs_23,outputs_1__15,
           outputs_1__14,outputs_1__13,outputs_1__12,outputs_1__11,outputs_1__10
           ,outputs_1__9,outputs_1__8,outputs_1__7,outputs_1__6,outputs_1__5,
           outputs_1__4,outputs_1__3,outputs_1__2,outputs_1__1,outputs_1__0,
           gen_1_cmp_pMux_8,gen_1_cmp_pMux_7,gen_1_cmp_pMux_6,gen_1_cmp_pMux_5,
           gen_1_cmp_pMux_4,gen_1_cmp_pMux_3,nx9675}), .en (nx11171), .clk (
           nx9397), .rst (rst), .Q ({\$dummy [115],\$dummy [116],
           gen_1_cmp_pReg_30,gen_1_cmp_pReg_29,gen_1_cmp_pReg_28,
           gen_1_cmp_pReg_27,gen_1_cmp_pReg_26,gen_1_cmp_pReg_25,
           gen_1_cmp_pReg_24,gen_1_cmp_pReg_23,gen_1_cmp_pReg_22,
           gen_1_cmp_pReg_21,gen_1_cmp_pReg_20,gen_1_cmp_pReg_19,
           gen_1_cmp_pReg_18,gen_1_cmp_pReg_17,gen_1_cmp_pReg_16,
           gen_1_cmp_pReg_15,gen_1_cmp_pReg_14,gen_1_cmp_pReg_13,
           gen_1_cmp_pReg_12,gen_1_cmp_pReg_11,gen_1_cmp_pReg_10,
           gen_1_cmp_pReg_9,gen_1_cmp_pReg_8,gen_1_cmp_pReg_7,gen_1_cmp_pReg_6,
           gen_1_cmp_pReg_5,gen_1_cmp_pReg_4,gen_1_cmp_pReg_3,gen_1_cmp_pReg_2,
           gen_1_cmp_pReg_1,gen_1_cmp_pReg_0})) ;
    BinaryMux_33 gen_1_cmp_MuxCmp (.a ({working,working,gen_1_cmp_pReg_30,
                 gen_1_cmp_pReg_29,gen_1_cmp_pReg_28,gen_1_cmp_pReg_27,
                 gen_1_cmp_pReg_26,gen_1_cmp_pReg_25,gen_1_cmp_pReg_24,
                 gen_1_cmp_pReg_23,gen_1_cmp_pReg_22,gen_1_cmp_pReg_21,
                 gen_1_cmp_pReg_20,gen_1_cmp_pReg_19,gen_1_cmp_pReg_18,
                 gen_1_cmp_pReg_17,gen_1_cmp_pReg_16,gen_1_cmp_pReg_15,
                 gen_1_cmp_pReg_14,gen_1_cmp_pReg_13,gen_1_cmp_pReg_12,
                 gen_1_cmp_pReg_11,gen_1_cmp_pReg_10,gen_1_cmp_pReg_9,
                 gen_1_cmp_pReg_8,gen_1_cmp_pReg_7,gen_1_cmp_pReg_6,
                 gen_1_cmp_pReg_5,gen_1_cmp_pReg_4,gen_1_cmp_pReg_3,
                 gen_1_cmp_pReg_2,gen_1_cmp_pReg_1,gen_1_cmp_pReg_0}), .b ({
                 working,working,working,working,working,working,working,working
                 ,working,working,working,working,working,working,working,
                 working,working,working,working,working,working,working,working
                 ,working,filter_1__7,filter_1__6,filter_1__5,filter_1__4,
                 filter_1__3,filter_1__2,filter_1__1,filter_1__0,working}), .sel (
                 nx9389), .f ({\$dummy [117],\$dummy [118],gen_1_cmp_pMux_30,
                 gen_1_cmp_pMux_29,gen_1_cmp_pMux_28,gen_1_cmp_pMux_27,
                 gen_1_cmp_pMux_26,gen_1_cmp_pMux_25,gen_1_cmp_pMux_24,
                 gen_1_cmp_pMux_23,gen_1_cmp_pMux_22,gen_1_cmp_pMux_21,
                 gen_1_cmp_pMux_20,gen_1_cmp_pMux_19,gen_1_cmp_pMux_18,
                 gen_1_cmp_pMux_17,gen_1_cmp_pMux_16,gen_1_cmp_pMux_15,
                 gen_1_cmp_pMux_14,gen_1_cmp_pMux_13,gen_1_cmp_pMux_12,
                 gen_1_cmp_pMux_11,gen_1_cmp_pMux_10,gen_1_cmp_pMux_9,
                 gen_1_cmp_pMux_8,gen_1_cmp_pMux_7,gen_1_cmp_pMux_6,
                 gen_1_cmp_pMux_5,gen_1_cmp_pMux_4,gen_1_cmp_pMux_3,
                 gen_1_cmp_pMux_2,gen_1_cmp_pMux_1,gen_1_cmp_pMux_0})) ;
    NBitAdder_24 gen_1_cmp_BSCmp_AdderCmp (.a ({working,working,
                 gen_1_cmp_pMux_30,gen_1_cmp_pMux_29,gen_1_cmp_pMux_28,
                 gen_1_cmp_pMux_27,gen_1_cmp_pMux_26,gen_1_cmp_pMux_25,
                 gen_1_cmp_pMux_24,gen_1_cmp_pMux_23,gen_1_cmp_pMux_22,
                 gen_1_cmp_pMux_21,gen_1_cmp_pMux_20,gen_1_cmp_pMux_19,
                 gen_1_cmp_pMux_18,gen_1_cmp_pMux_17,gen_1_cmp_pMux_16,
                 gen_1_cmp_pMux_15,gen_1_cmp_pMux_14,gen_1_cmp_pMux_13,
                 gen_1_cmp_pMux_12,gen_1_cmp_pMux_11,gen_1_cmp_pMux_10,
                 gen_1_cmp_pMux_9}), .b ({nx9979,nx9979,nx9977,nx9985,nx9983,
                 nx9981,nx9979,nx9977,gen_1_cmp_BSCmp_op2_15,
                 gen_1_cmp_BSCmp_op2_14,gen_1_cmp_BSCmp_op2_13,
                 gen_1_cmp_BSCmp_op2_12,gen_1_cmp_BSCmp_op2_11,
                 gen_1_cmp_BSCmp_op2_10,gen_1_cmp_BSCmp_op2_9,
                 gen_1_cmp_BSCmp_op2_8,gen_1_cmp_BSCmp_op2_7,
                 gen_1_cmp_BSCmp_op2_6,gen_1_cmp_BSCmp_op2_5,
                 gen_1_cmp_BSCmp_op2_4,gen_1_cmp_BSCmp_op2_3,
                 gen_1_cmp_BSCmp_op2_2,gen_1_cmp_BSCmp_op2_1,
                 gen_1_cmp_BSCmp_op2_0}), .carryIn (gen_1_cmp_BSCmp_carryIn), .sum (
                 {gen_1_cmp_pBs_30,gen_1_cmp_pBs_29,gen_1_cmp_pBs_28,
                 gen_1_cmp_pBs_27,gen_1_cmp_pBs_26,gen_1_cmp_pBs_25,
                 gen_1_cmp_pBs_24,gen_1_cmp_pBs_23,outputs_1__15,outputs_1__14,
                 outputs_1__13,outputs_1__12,outputs_1__11,outputs_1__10,
                 outputs_1__9,outputs_1__8,outputs_1__7,outputs_1__6,
                 outputs_1__5,outputs_1__4,outputs_1__3,outputs_1__2,
                 outputs_1__1,outputs_1__0}), .carryOut (\$dummy [119])) ;
    Reg_33 gen_0_cmp_pRegCmp (.D ({working,working,gen_0_cmp_pBs_30,
           gen_0_cmp_pBs_29,gen_0_cmp_pBs_28,gen_0_cmp_pBs_27,gen_0_cmp_pBs_26,
           gen_0_cmp_pBs_25,gen_0_cmp_pBs_24,gen_0_cmp_pBs_23,outputs_0__15,
           outputs_0__14,outputs_0__13,outputs_0__12,outputs_0__11,outputs_0__10
           ,outputs_0__9,outputs_0__8,outputs_0__7,outputs_0__6,outputs_0__5,
           outputs_0__4,outputs_0__3,outputs_0__2,outputs_0__1,outputs_0__0,
           gen_0_cmp_pMux_8,gen_0_cmp_pMux_7,gen_0_cmp_pMux_6,gen_0_cmp_pMux_5,
           gen_0_cmp_pMux_4,gen_0_cmp_pMux_3,nx9687}), .en (nx9381), .clk (
           nx9397), .rst (rst), .Q ({\$dummy [120],\$dummy [121],
           gen_0_cmp_pReg_30,gen_0_cmp_pReg_29,gen_0_cmp_pReg_28,
           gen_0_cmp_pReg_27,gen_0_cmp_pReg_26,gen_0_cmp_pReg_25,
           gen_0_cmp_pReg_24,gen_0_cmp_pReg_23,gen_0_cmp_pReg_22,
           gen_0_cmp_pReg_21,gen_0_cmp_pReg_20,gen_0_cmp_pReg_19,
           gen_0_cmp_pReg_18,gen_0_cmp_pReg_17,gen_0_cmp_pReg_16,
           gen_0_cmp_pReg_15,gen_0_cmp_pReg_14,gen_0_cmp_pReg_13,
           gen_0_cmp_pReg_12,gen_0_cmp_pReg_11,gen_0_cmp_pReg_10,
           gen_0_cmp_pReg_9,gen_0_cmp_pReg_8,gen_0_cmp_pReg_7,gen_0_cmp_pReg_6,
           gen_0_cmp_pReg_5,gen_0_cmp_pReg_4,gen_0_cmp_pReg_3,gen_0_cmp_pReg_2,
           gen_0_cmp_pReg_1,gen_0_cmp_pReg_0})) ;
    BinaryMux_33 gen_0_cmp_MuxCmp (.a ({working,working,gen_0_cmp_pReg_30,
                 gen_0_cmp_pReg_29,gen_0_cmp_pReg_28,gen_0_cmp_pReg_27,
                 gen_0_cmp_pReg_26,gen_0_cmp_pReg_25,gen_0_cmp_pReg_24,
                 gen_0_cmp_pReg_23,gen_0_cmp_pReg_22,gen_0_cmp_pReg_21,
                 gen_0_cmp_pReg_20,gen_0_cmp_pReg_19,gen_0_cmp_pReg_18,
                 gen_0_cmp_pReg_17,gen_0_cmp_pReg_16,gen_0_cmp_pReg_15,
                 gen_0_cmp_pReg_14,gen_0_cmp_pReg_13,gen_0_cmp_pReg_12,
                 gen_0_cmp_pReg_11,gen_0_cmp_pReg_10,gen_0_cmp_pReg_9,
                 gen_0_cmp_pReg_8,gen_0_cmp_pReg_7,gen_0_cmp_pReg_6,
                 gen_0_cmp_pReg_5,gen_0_cmp_pReg_4,gen_0_cmp_pReg_3,
                 gen_0_cmp_pReg_2,gen_0_cmp_pReg_1,gen_0_cmp_pReg_0}), .b ({
                 working,working,working,working,working,working,working,working
                 ,working,working,working,working,working,working,working,
                 working,working,working,working,working,working,working,working
                 ,working,filter_0__7,filter_0__6,filter_0__5,filter_0__4,
                 filter_0__3,filter_0__2,filter_0__1,filter_0__0,working}), .sel (
                 nx9389), .f ({\$dummy [122],\$dummy [123],gen_0_cmp_pMux_30,
                 gen_0_cmp_pMux_29,gen_0_cmp_pMux_28,gen_0_cmp_pMux_27,
                 gen_0_cmp_pMux_26,gen_0_cmp_pMux_25,gen_0_cmp_pMux_24,
                 gen_0_cmp_pMux_23,gen_0_cmp_pMux_22,gen_0_cmp_pMux_21,
                 gen_0_cmp_pMux_20,gen_0_cmp_pMux_19,gen_0_cmp_pMux_18,
                 gen_0_cmp_pMux_17,gen_0_cmp_pMux_16,gen_0_cmp_pMux_15,
                 gen_0_cmp_pMux_14,gen_0_cmp_pMux_13,gen_0_cmp_pMux_12,
                 gen_0_cmp_pMux_11,gen_0_cmp_pMux_10,gen_0_cmp_pMux_9,
                 gen_0_cmp_pMux_8,gen_0_cmp_pMux_7,gen_0_cmp_pMux_6,
                 gen_0_cmp_pMux_5,gen_0_cmp_pMux_4,gen_0_cmp_pMux_3,
                 gen_0_cmp_pMux_2,gen_0_cmp_pMux_1,gen_0_cmp_pMux_0})) ;
    NBitAdder_24 gen_0_cmp_BSCmp_AdderCmp (.a ({working,working,
                 gen_0_cmp_pMux_30,gen_0_cmp_pMux_29,gen_0_cmp_pMux_28,
                 gen_0_cmp_pMux_27,gen_0_cmp_pMux_26,gen_0_cmp_pMux_25,
                 gen_0_cmp_pMux_24,gen_0_cmp_pMux_23,gen_0_cmp_pMux_22,
                 gen_0_cmp_pMux_21,gen_0_cmp_pMux_20,gen_0_cmp_pMux_19,
                 gen_0_cmp_pMux_18,gen_0_cmp_pMux_17,gen_0_cmp_pMux_16,
                 gen_0_cmp_pMux_15,gen_0_cmp_pMux_14,gen_0_cmp_pMux_13,
                 gen_0_cmp_pMux_12,gen_0_cmp_pMux_11,gen_0_cmp_pMux_10,
                 gen_0_cmp_pMux_9}), .b ({nx9991,nx9991,nx9989,nx9997,nx9995,
                 nx9993,nx9991,nx9989,gen_0_cmp_BSCmp_op2_15,
                 gen_0_cmp_BSCmp_op2_14,gen_0_cmp_BSCmp_op2_13,
                 gen_0_cmp_BSCmp_op2_12,gen_0_cmp_BSCmp_op2_11,
                 gen_0_cmp_BSCmp_op2_10,gen_0_cmp_BSCmp_op2_9,
                 gen_0_cmp_BSCmp_op2_8,gen_0_cmp_BSCmp_op2_7,
                 gen_0_cmp_BSCmp_op2_6,gen_0_cmp_BSCmp_op2_5,
                 gen_0_cmp_BSCmp_op2_4,gen_0_cmp_BSCmp_op2_3,
                 gen_0_cmp_BSCmp_op2_2,gen_0_cmp_BSCmp_op2_1,
                 gen_0_cmp_BSCmp_op2_0}), .carryIn (gen_0_cmp_BSCmp_carryIn), .sum (
                 {gen_0_cmp_pBs_30,gen_0_cmp_pBs_29,gen_0_cmp_pBs_28,
                 gen_0_cmp_pBs_27,gen_0_cmp_pBs_26,gen_0_cmp_pBs_25,
                 gen_0_cmp_pBs_24,gen_0_cmp_pBs_23,outputs_0__15,outputs_0__14,
                 outputs_0__13,outputs_0__12,outputs_0__11,outputs_0__10,
                 outputs_0__9,outputs_0__8,outputs_0__7,outputs_0__6,
                 outputs_0__5,outputs_0__4,outputs_0__3,outputs_0__2,
                 outputs_0__1,outputs_0__0}), .carryOut (\$dummy [124])) ;
    fake_vcc ix9651 (.Y (nx9650)) ;
    fake_gnd ix2325 (.Y (working)) ;
    nand02 ix67 (.Y (gen_0_cmp_BSCmp_op2_1), .A0 (nx2853), .A1 (nx2873)) ;
    nor02_2x ix2854 (.Y (nx2853), .A0 (nx62), .A1 (nx58)) ;
    nor03_2x ix63 (.Y (nx62), .A0 (gen_0_cmp_mReg_0), .A1 (nx9693), .A2 (nx10151
             )) ;
    dffr gen_0_cmp_mRegCmp_reg_Q_0 (.Q (gen_0_cmp_mReg_0), .QB (nx2859), .D (
         window_0__0), .CLK (start), .R (rst)) ;
    inv01 ix2864 (.Y (nx2862), .A (gen_0_cmp_pMux_0)) ;
    nor03_2x ix59 (.Y (nx58), .A0 (nx2859), .A1 (nx10157), .A2 (nx10167)) ;
    inv02 ix2872 (.Y (nx2871), .A (gen_0_cmp_pMux_2)) ;
    nor02_2x ix2874 (.Y (nx2873), .A0 (nx48), .A1 (nx46)) ;
    nor03_2x ix49 (.Y (nx48), .A0 (nx2877), .A1 (nx9687), .A2 (nx10175)) ;
    dffr gen_0_cmp_mRegCmp_reg_Q_1 (.Q (gen_0_cmp_mReg_1), .QB (nx2877), .D (
         window_0__1), .CLK (start), .R (rst)) ;
    nor03_2x ix47 (.Y (nx46), .A0 (gen_0_cmp_mReg_1), .A1 (nx9999), .A2 (nx10183
             )) ;
    nor03_2x ix7 (.Y (nx6), .A0 (nx9693), .A1 (nx2871), .A2 (gen_0_cmp_pMux_0)
             ) ;
    nand02 ix89 (.Y (gen_0_cmp_BSCmp_op2_2), .A0 (nx2887), .A1 (nx2893)) ;
    nor02_2x ix2888 (.Y (nx2887), .A0 (nx84), .A1 (nx80)) ;
    nor03_2x ix85 (.Y (nx84), .A0 (gen_0_cmp_mReg_1), .A1 (nx9693), .A2 (nx10151
             )) ;
    nor03_2x ix81 (.Y (nx80), .A0 (nx2877), .A1 (nx10157), .A2 (nx10167)) ;
    nor02_2x ix2894 (.Y (nx2893), .A0 (nx76), .A1 (nx74)) ;
    nor03_2x ix77 (.Y (nx76), .A0 (nx2897), .A1 (nx9687), .A2 (nx10175)) ;
    dffr gen_0_cmp_mRegCmp_reg_Q_2 (.Q (gen_0_cmp_mReg_2), .QB (nx2897), .D (
         window_0__2), .CLK (start), .R (rst)) ;
    nor03_2x ix75 (.Y (nx74), .A0 (gen_0_cmp_mReg_2), .A1 (nx9999), .A2 (nx10183
             )) ;
    nand02 ix111 (.Y (gen_0_cmp_BSCmp_op2_3), .A0 (nx2903), .A1 (nx2907)) ;
    nor02_2x ix2904 (.Y (nx2903), .A0 (nx106), .A1 (nx102)) ;
    nor03_2x ix107 (.Y (nx106), .A0 (gen_0_cmp_mReg_2), .A1 (nx9693), .A2 (
             nx10151)) ;
    nor03_2x ix103 (.Y (nx102), .A0 (nx2897), .A1 (nx10157), .A2 (nx10167)) ;
    nor02_2x ix2908 (.Y (nx2907), .A0 (nx98), .A1 (nx96)) ;
    nor03_2x ix99 (.Y (nx98), .A0 (nx2911), .A1 (nx9687), .A2 (nx10175)) ;
    dffr gen_0_cmp_mRegCmp_reg_Q_3 (.Q (gen_0_cmp_mReg_3), .QB (nx2911), .D (
         window_0__3), .CLK (start), .R (rst)) ;
    nor03_2x ix97 (.Y (nx96), .A0 (gen_0_cmp_mReg_3), .A1 (nx9999), .A2 (nx10183
             )) ;
    nand02 ix133 (.Y (gen_0_cmp_BSCmp_op2_4), .A0 (nx2917), .A1 (nx2923)) ;
    nor02_2x ix2918 (.Y (nx2917), .A0 (nx128), .A1 (nx124)) ;
    nor03_2x ix129 (.Y (nx128), .A0 (gen_0_cmp_mReg_3), .A1 (nx9693), .A2 (
             nx10151)) ;
    nor03_2x ix125 (.Y (nx124), .A0 (nx2911), .A1 (nx10157), .A2 (nx10167)) ;
    nor02_2x ix2924 (.Y (nx2923), .A0 (nx120), .A1 (nx118)) ;
    nor03_2x ix121 (.Y (nx120), .A0 (nx2926), .A1 (nx9687), .A2 (nx10175)) ;
    dffr gen_0_cmp_mRegCmp_reg_Q_4 (.Q (gen_0_cmp_mReg_4), .QB (nx2926), .D (
         window_0__4), .CLK (start), .R (rst)) ;
    nor03_2x ix119 (.Y (nx118), .A0 (gen_0_cmp_mReg_4), .A1 (nx9999), .A2 (
             nx10183)) ;
    nand02 ix155 (.Y (gen_0_cmp_BSCmp_op2_5), .A0 (nx2931), .A1 (nx2937)) ;
    nor02_2x ix2932 (.Y (nx2931), .A0 (nx150), .A1 (nx146)) ;
    nor03_2x ix151 (.Y (nx150), .A0 (gen_0_cmp_mReg_4), .A1 (nx9693), .A2 (
             nx10151)) ;
    nor03_2x ix147 (.Y (nx146), .A0 (nx2926), .A1 (nx10157), .A2 (nx10167)) ;
    nor02_2x ix2938 (.Y (nx2937), .A0 (nx142), .A1 (nx140)) ;
    nor03_2x ix143 (.Y (nx142), .A0 (nx2941), .A1 (nx9689), .A2 (nx10175)) ;
    dffr gen_0_cmp_mRegCmp_reg_Q_5 (.Q (gen_0_cmp_mReg_5), .QB (nx2941), .D (
         window_0__5), .CLK (start), .R (rst)) ;
    nor03_2x ix141 (.Y (nx140), .A0 (gen_0_cmp_mReg_5), .A1 (nx9999), .A2 (
             nx10183)) ;
    nand02 ix177 (.Y (gen_0_cmp_BSCmp_op2_6), .A0 (nx2947), .A1 (nx2951)) ;
    nor02_2x ix2948 (.Y (nx2947), .A0 (nx172), .A1 (nx168)) ;
    nor03_2x ix173 (.Y (nx172), .A0 (gen_0_cmp_mReg_5), .A1 (nx9695), .A2 (
             nx10151)) ;
    nor03_2x ix169 (.Y (nx168), .A0 (nx2941), .A1 (nx10157), .A2 (nx10167)) ;
    nor02_2x ix2952 (.Y (nx2951), .A0 (nx164), .A1 (nx162)) ;
    nor03_2x ix165 (.Y (nx164), .A0 (nx2955), .A1 (nx9689), .A2 (nx10175)) ;
    dffr gen_0_cmp_mRegCmp_reg_Q_6 (.Q (gen_0_cmp_mReg_6), .QB (nx2955), .D (
         window_0__6), .CLK (start), .R (rst)) ;
    nor03_2x ix163 (.Y (nx162), .A0 (gen_0_cmp_mReg_6), .A1 (nx9999), .A2 (
             nx10183)) ;
    nand02 ix199 (.Y (gen_0_cmp_BSCmp_op2_7), .A0 (nx2961), .A1 (nx2967)) ;
    nor02_2x ix2962 (.Y (nx2961), .A0 (nx194), .A1 (nx190)) ;
    nor03_2x ix195 (.Y (nx194), .A0 (gen_0_cmp_mReg_6), .A1 (nx9695), .A2 (
             nx10153)) ;
    nor03_2x ix191 (.Y (nx190), .A0 (nx2955), .A1 (nx10159), .A2 (nx10169)) ;
    nor02_2x ix2968 (.Y (nx2967), .A0 (nx186), .A1 (nx184)) ;
    nor03_2x ix187 (.Y (nx186), .A0 (nx2970), .A1 (nx9689), .A2 (nx10177)) ;
    dffr gen_0_cmp_mRegCmp_reg_Q_7 (.Q (gen_0_cmp_mReg_7), .QB (nx2970), .D (
         window_0__7), .CLK (start), .R (rst)) ;
    nor03_2x ix185 (.Y (nx184), .A0 (gen_0_cmp_mReg_7), .A1 (nx9999), .A2 (
             nx10185)) ;
    nand02 ix221 (.Y (gen_0_cmp_BSCmp_op2_8), .A0 (nx2975), .A1 (nx2981)) ;
    nor02_2x ix2976 (.Y (nx2975), .A0 (nx216), .A1 (nx212)) ;
    nor03_2x ix217 (.Y (nx216), .A0 (gen_0_cmp_mReg_7), .A1 (nx9695), .A2 (
             nx10153)) ;
    nor03_2x ix213 (.Y (nx212), .A0 (nx2970), .A1 (nx10159), .A2 (nx10169)) ;
    nor02_2x ix2982 (.Y (nx2981), .A0 (nx208), .A1 (nx206)) ;
    nor03_2x ix209 (.Y (nx208), .A0 (nx2985), .A1 (nx9689), .A2 (nx10177)) ;
    dffr gen_0_cmp_mRegCmp_reg_Q_8 (.Q (gen_0_cmp_mReg_8), .QB (nx2985), .D (
         window_0__8), .CLK (start), .R (rst)) ;
    nor03_2x ix207 (.Y (nx206), .A0 (gen_0_cmp_mReg_8), .A1 (nx10001), .A2 (
             nx10185)) ;
    nand02 ix243 (.Y (gen_0_cmp_BSCmp_op2_9), .A0 (nx2991), .A1 (nx2995)) ;
    nor02_2x ix2992 (.Y (nx2991), .A0 (nx238), .A1 (nx234)) ;
    nor03_2x ix239 (.Y (nx238), .A0 (gen_0_cmp_mReg_8), .A1 (nx9695), .A2 (
             nx10153)) ;
    nor03_2x ix235 (.Y (nx234), .A0 (nx2985), .A1 (nx10159), .A2 (nx10169)) ;
    nor02_2x ix2996 (.Y (nx2995), .A0 (nx230), .A1 (nx228)) ;
    nor03_2x ix231 (.Y (nx230), .A0 (nx2999), .A1 (nx9689), .A2 (nx10177)) ;
    dffr gen_0_cmp_mRegCmp_reg_Q_9 (.Q (gen_0_cmp_mReg_9), .QB (nx2999), .D (
         window_0__9), .CLK (start), .R (rst)) ;
    nor03_2x ix229 (.Y (nx228), .A0 (gen_0_cmp_mReg_9), .A1 (nx10001), .A2 (
             nx10185)) ;
    nand02 ix265 (.Y (gen_0_cmp_BSCmp_op2_10), .A0 (nx3005), .A1 (nx3011)) ;
    nor02_2x ix3006 (.Y (nx3005), .A0 (nx260), .A1 (nx256)) ;
    nor03_2x ix261 (.Y (nx260), .A0 (gen_0_cmp_mReg_9), .A1 (nx9695), .A2 (
             nx10153)) ;
    nor03_2x ix257 (.Y (nx256), .A0 (nx2999), .A1 (nx10159), .A2 (nx10169)) ;
    nor02_2x ix3012 (.Y (nx3011), .A0 (nx252), .A1 (nx250)) ;
    nor03_2x ix253 (.Y (nx252), .A0 (nx3014), .A1 (nx9689), .A2 (nx10177)) ;
    dffr gen_0_cmp_mRegCmp_reg_Q_10 (.Q (gen_0_cmp_mReg_10), .QB (nx3014), .D (
         window_0__10), .CLK (start), .R (rst)) ;
    nor03_2x ix251 (.Y (nx250), .A0 (gen_0_cmp_mReg_10), .A1 (nx10001), .A2 (
             nx10185)) ;
    nand02 ix287 (.Y (gen_0_cmp_BSCmp_op2_11), .A0 (nx3019), .A1 (nx3025)) ;
    nor02_2x ix3020 (.Y (nx3019), .A0 (nx282), .A1 (nx278)) ;
    nor03_2x ix283 (.Y (nx282), .A0 (gen_0_cmp_mReg_10), .A1 (nx9695), .A2 (
             nx10153)) ;
    nor03_2x ix279 (.Y (nx278), .A0 (nx3014), .A1 (nx10159), .A2 (nx10169)) ;
    nor02_2x ix3026 (.Y (nx3025), .A0 (nx274), .A1 (nx272)) ;
    nor03_2x ix275 (.Y (nx274), .A0 (nx3029), .A1 (nx9689), .A2 (nx10177)) ;
    dffr gen_0_cmp_mRegCmp_reg_Q_11 (.Q (gen_0_cmp_mReg_11), .QB (nx3029), .D (
         window_0__11), .CLK (start), .R (rst)) ;
    nor03_2x ix273 (.Y (nx272), .A0 (gen_0_cmp_mReg_11), .A1 (nx10001), .A2 (
             nx10185)) ;
    nand02 ix309 (.Y (gen_0_cmp_BSCmp_op2_12), .A0 (nx3035), .A1 (nx3039)) ;
    nor02_2x ix3036 (.Y (nx3035), .A0 (nx304), .A1 (nx300)) ;
    nor03_2x ix305 (.Y (nx304), .A0 (gen_0_cmp_mReg_11), .A1 (nx9695), .A2 (
             nx10153)) ;
    nor03_2x ix301 (.Y (nx300), .A0 (nx3029), .A1 (nx10159), .A2 (nx10169)) ;
    nor02_2x ix3040 (.Y (nx3039), .A0 (nx296), .A1 (nx294)) ;
    nor03_2x ix297 (.Y (nx296), .A0 (nx3043), .A1 (nx9691), .A2 (nx10177)) ;
    dffr gen_0_cmp_mRegCmp_reg_Q_12 (.Q (gen_0_cmp_mReg_12), .QB (nx3043), .D (
         window_0__12), .CLK (start), .R (rst)) ;
    nor03_2x ix295 (.Y (nx294), .A0 (gen_0_cmp_mReg_12), .A1 (nx10001), .A2 (
             nx10185)) ;
    nand02 ix331 (.Y (gen_0_cmp_BSCmp_op2_13), .A0 (nx3049), .A1 (nx3055)) ;
    nor02_2x ix3050 (.Y (nx3049), .A0 (nx326), .A1 (nx322)) ;
    nor03_2x ix327 (.Y (nx326), .A0 (gen_0_cmp_mReg_12), .A1 (nx9697), .A2 (
             nx10155)) ;
    nor03_2x ix323 (.Y (nx322), .A0 (nx3043), .A1 (nx10159), .A2 (nx10171)) ;
    nor02_2x ix3056 (.Y (nx3055), .A0 (nx318), .A1 (nx316)) ;
    nor03_2x ix319 (.Y (nx318), .A0 (nx3058), .A1 (nx9691), .A2 (nx10179)) ;
    dffr gen_0_cmp_mRegCmp_reg_Q_13 (.Q (gen_0_cmp_mReg_13), .QB (nx3058), .D (
         window_0__13), .CLK (start), .R (rst)) ;
    nor03_2x ix317 (.Y (nx316), .A0 (gen_0_cmp_mReg_13), .A1 (nx10001), .A2 (
             nx10187)) ;
    nand02 ix353 (.Y (gen_0_cmp_BSCmp_op2_14), .A0 (nx3063), .A1 (nx3069)) ;
    nor02_2x ix3064 (.Y (nx3063), .A0 (nx348), .A1 (nx344)) ;
    nor03_2x ix349 (.Y (nx348), .A0 (gen_0_cmp_mReg_13), .A1 (nx9697), .A2 (
             nx10155)) ;
    nor03_2x ix345 (.Y (nx344), .A0 (nx3058), .A1 (nx10161), .A2 (nx10171)) ;
    nor02_2x ix3070 (.Y (nx3069), .A0 (nx340), .A1 (nx338)) ;
    nor03_2x ix341 (.Y (nx340), .A0 (nx3073), .A1 (nx9691), .A2 (nx10179)) ;
    dffr gen_0_cmp_mRegCmp_reg_Q_14 (.Q (gen_0_cmp_mReg_14), .QB (nx3073), .D (
         window_0__14), .CLK (start), .R (rst)) ;
    nor03_2x ix339 (.Y (nx338), .A0 (gen_0_cmp_mReg_14), .A1 (nx10001), .A2 (
             nx10187)) ;
    nand02 ix375 (.Y (gen_0_cmp_BSCmp_op2_15), .A0 (nx3079), .A1 (nx3083)) ;
    nor02_2x ix3080 (.Y (nx3079), .A0 (nx370), .A1 (nx366)) ;
    nor03_2x ix371 (.Y (nx370), .A0 (gen_0_cmp_mReg_14), .A1 (nx9697), .A2 (
             nx10155)) ;
    nor03_2x ix367 (.Y (nx366), .A0 (nx3073), .A1 (nx10161), .A2 (nx10171)) ;
    nor02_2x ix3084 (.Y (nx3083), .A0 (nx362), .A1 (nx360)) ;
    nor03_2x ix363 (.Y (nx362), .A0 (nx3087), .A1 (nx9691), .A2 (nx10179)) ;
    dffr gen_0_cmp_mRegCmp_reg_Q_15 (.Q (gen_0_cmp_mReg_15), .QB (nx3087), .D (
         window_0__15), .CLK (start), .R (rst)) ;
    nor03_2x ix361 (.Y (nx360), .A0 (gen_0_cmp_mReg_15), .A1 (nx10003), .A2 (
             nx10187)) ;
    nand02 ix385 (.Y (gen_0_cmp_BSCmp_op2_16), .A0 (nx3093), .A1 (nx3083)) ;
    nor02_2x ix3094 (.Y (nx3093), .A0 (nx380), .A1 (nx376)) ;
    nor03_2x ix381 (.Y (nx380), .A0 (gen_0_cmp_mReg_15), .A1 (nx9697), .A2 (
             nx10155)) ;
    nor03_2x ix377 (.Y (nx376), .A0 (nx3087), .A1 (nx10161), .A2 (nx10171)) ;
    nand02 ix453 (.Y (gen_1_cmp_BSCmp_op2_1), .A0 (nx3099), .A1 (nx3117)) ;
    nor02_2x ix3100 (.Y (nx3099), .A0 (nx448), .A1 (nx444)) ;
    nor03_2x ix449 (.Y (nx448), .A0 (gen_1_cmp_mReg_0), .A1 (nx9681), .A2 (
             nx10191)) ;
    dffr gen_1_cmp_mRegCmp_reg_Q_0 (.Q (gen_1_cmp_mReg_0), .QB (nx3103), .D (
         window_1__0), .CLK (start), .R (rst)) ;
    inv01 ix3108 (.Y (nx3107), .A (gen_1_cmp_pMux_0)) ;
    nor03_2x ix445 (.Y (nx444), .A0 (nx3103), .A1 (nx10197), .A2 (nx10207)) ;
    inv02 ix3116 (.Y (nx3115), .A (gen_1_cmp_pMux_2)) ;
    nor02_2x ix3118 (.Y (nx3117), .A0 (nx434), .A1 (nx432)) ;
    nor03_2x ix435 (.Y (nx434), .A0 (nx3121), .A1 (nx9675), .A2 (nx10215)) ;
    dffr gen_1_cmp_mRegCmp_reg_Q_1 (.Q (gen_1_cmp_mReg_1), .QB (nx3121), .D (
         window_1__1), .CLK (start), .R (rst)) ;
    nor03_2x ix433 (.Y (nx432), .A0 (gen_1_cmp_mReg_1), .A1 (nx10005), .A2 (
             nx10223)) ;
    nor03_2x ix393 (.Y (nx392), .A0 (nx9681), .A1 (nx3115), .A2 (
             gen_1_cmp_pMux_0)) ;
    nand02 ix475 (.Y (gen_1_cmp_BSCmp_op2_2), .A0 (nx3132), .A1 (nx3139)) ;
    nor02_2x ix3134 (.Y (nx3132), .A0 (nx470), .A1 (nx466)) ;
    nor03_2x ix471 (.Y (nx470), .A0 (gen_1_cmp_mReg_1), .A1 (nx9681), .A2 (
             nx10191)) ;
    nor03_2x ix467 (.Y (nx466), .A0 (nx3121), .A1 (nx10197), .A2 (nx10207)) ;
    nor02_2x ix3140 (.Y (nx3139), .A0 (nx462), .A1 (nx460)) ;
    nor03_2x ix463 (.Y (nx462), .A0 (nx3143), .A1 (nx9675), .A2 (nx10215)) ;
    dffr gen_1_cmp_mRegCmp_reg_Q_2 (.Q (gen_1_cmp_mReg_2), .QB (nx3143), .D (
         window_1__2), .CLK (start), .R (rst)) ;
    nor03_2x ix461 (.Y (nx460), .A0 (gen_1_cmp_mReg_2), .A1 (nx10005), .A2 (
             nx10223)) ;
    nand02 ix497 (.Y (gen_1_cmp_BSCmp_op2_3), .A0 (nx3149), .A1 (nx3155)) ;
    nor02_2x ix3150 (.Y (nx3149), .A0 (nx492), .A1 (nx488)) ;
    nor03_2x ix493 (.Y (nx492), .A0 (gen_1_cmp_mReg_2), .A1 (nx9681), .A2 (
             nx10191)) ;
    nor03_2x ix489 (.Y (nx488), .A0 (nx3143), .A1 (nx10197), .A2 (nx10207)) ;
    nor02_2x ix3156 (.Y (nx3155), .A0 (nx484), .A1 (nx482)) ;
    nor03_2x ix485 (.Y (nx484), .A0 (nx3158), .A1 (nx9675), .A2 (nx10215)) ;
    dffr gen_1_cmp_mRegCmp_reg_Q_3 (.Q (gen_1_cmp_mReg_3), .QB (nx3158), .D (
         window_1__3), .CLK (start), .R (rst)) ;
    nor03_2x ix483 (.Y (nx482), .A0 (gen_1_cmp_mReg_3), .A1 (nx10005), .A2 (
             nx10223)) ;
    nand02 ix519 (.Y (gen_1_cmp_BSCmp_op2_4), .A0 (nx3163), .A1 (nx3169)) ;
    nor02_2x ix3164 (.Y (nx3163), .A0 (nx514), .A1 (nx510)) ;
    nor03_2x ix515 (.Y (nx514), .A0 (gen_1_cmp_mReg_3), .A1 (nx9681), .A2 (
             nx10191)) ;
    nor03_2x ix511 (.Y (nx510), .A0 (nx3158), .A1 (nx10197), .A2 (nx10207)) ;
    nor02_2x ix3170 (.Y (nx3169), .A0 (nx506), .A1 (nx504)) ;
    nor03_2x ix507 (.Y (nx506), .A0 (nx3173), .A1 (nx9675), .A2 (nx10215)) ;
    dffr gen_1_cmp_mRegCmp_reg_Q_4 (.Q (gen_1_cmp_mReg_4), .QB (nx3173), .D (
         window_1__4), .CLK (start), .R (rst)) ;
    nor03_2x ix505 (.Y (nx504), .A0 (gen_1_cmp_mReg_4), .A1 (nx10005), .A2 (
             nx10223)) ;
    nand02 ix541 (.Y (gen_1_cmp_BSCmp_op2_5), .A0 (nx3179), .A1 (nx3183)) ;
    nor02_2x ix3180 (.Y (nx3179), .A0 (nx536), .A1 (nx532)) ;
    nor03_2x ix537 (.Y (nx536), .A0 (gen_1_cmp_mReg_4), .A1 (nx9681), .A2 (
             nx10191)) ;
    nor03_2x ix533 (.Y (nx532), .A0 (nx3173), .A1 (nx10197), .A2 (nx10207)) ;
    nor02_2x ix3184 (.Y (nx3183), .A0 (nx528), .A1 (nx526)) ;
    nor03_2x ix529 (.Y (nx528), .A0 (nx3187), .A1 (nx9677), .A2 (nx10215)) ;
    dffr gen_1_cmp_mRegCmp_reg_Q_5 (.Q (gen_1_cmp_mReg_5), .QB (nx3187), .D (
         window_1__5), .CLK (start), .R (rst)) ;
    nor03_2x ix527 (.Y (nx526), .A0 (gen_1_cmp_mReg_5), .A1 (nx10005), .A2 (
             nx10223)) ;
    nand02 ix563 (.Y (gen_1_cmp_BSCmp_op2_6), .A0 (nx3193), .A1 (nx3199)) ;
    nor02_2x ix3194 (.Y (nx3193), .A0 (nx558), .A1 (nx554)) ;
    nor03_2x ix559 (.Y (nx558), .A0 (gen_1_cmp_mReg_5), .A1 (nx9683), .A2 (
             nx10191)) ;
    nor03_2x ix555 (.Y (nx554), .A0 (nx3187), .A1 (nx10197), .A2 (nx10207)) ;
    nor02_2x ix3200 (.Y (nx3199), .A0 (nx550), .A1 (nx548)) ;
    nor03_2x ix551 (.Y (nx550), .A0 (nx3202), .A1 (nx9677), .A2 (nx10215)) ;
    dffr gen_1_cmp_mRegCmp_reg_Q_6 (.Q (gen_1_cmp_mReg_6), .QB (nx3202), .D (
         window_1__6), .CLK (start), .R (rst)) ;
    nor03_2x ix549 (.Y (nx548), .A0 (gen_1_cmp_mReg_6), .A1 (nx10005), .A2 (
             nx10223)) ;
    nand02 ix585 (.Y (gen_1_cmp_BSCmp_op2_7), .A0 (nx3207), .A1 (nx3213)) ;
    nor02_2x ix3208 (.Y (nx3207), .A0 (nx580), .A1 (nx576)) ;
    nor03_2x ix581 (.Y (nx580), .A0 (gen_1_cmp_mReg_6), .A1 (nx9683), .A2 (
             nx10193)) ;
    nor03_2x ix577 (.Y (nx576), .A0 (nx3202), .A1 (nx10199), .A2 (nx10209)) ;
    nor02_2x ix3214 (.Y (nx3213), .A0 (nx572), .A1 (nx570)) ;
    nor03_2x ix573 (.Y (nx572), .A0 (nx3217), .A1 (nx9677), .A2 (nx10217)) ;
    dffr gen_1_cmp_mRegCmp_reg_Q_7 (.Q (gen_1_cmp_mReg_7), .QB (nx3217), .D (
         window_1__7), .CLK (start), .R (rst)) ;
    nor03_2x ix571 (.Y (nx570), .A0 (gen_1_cmp_mReg_7), .A1 (nx10005), .A2 (
             nx10225)) ;
    nand02 ix607 (.Y (gen_1_cmp_BSCmp_op2_8), .A0 (nx3223), .A1 (nx3227)) ;
    nor02_2x ix3224 (.Y (nx3223), .A0 (nx602), .A1 (nx598)) ;
    nor03_2x ix603 (.Y (nx602), .A0 (gen_1_cmp_mReg_7), .A1 (nx9683), .A2 (
             nx10193)) ;
    nor03_2x ix599 (.Y (nx598), .A0 (nx3217), .A1 (nx10199), .A2 (nx10209)) ;
    nor02_2x ix3228 (.Y (nx3227), .A0 (nx594), .A1 (nx592)) ;
    nor03_2x ix595 (.Y (nx594), .A0 (nx3231), .A1 (nx9677), .A2 (nx10217)) ;
    dffr gen_1_cmp_mRegCmp_reg_Q_8 (.Q (gen_1_cmp_mReg_8), .QB (nx3231), .D (
         window_1__8), .CLK (start), .R (rst)) ;
    nor03_2x ix593 (.Y (nx592), .A0 (gen_1_cmp_mReg_8), .A1 (nx10007), .A2 (
             nx10225)) ;
    nand02 ix629 (.Y (gen_1_cmp_BSCmp_op2_9), .A0 (nx3237), .A1 (nx3243)) ;
    nor02_2x ix3238 (.Y (nx3237), .A0 (nx624), .A1 (nx620)) ;
    nor03_2x ix625 (.Y (nx624), .A0 (gen_1_cmp_mReg_8), .A1 (nx9683), .A2 (
             nx10193)) ;
    nor03_2x ix621 (.Y (nx620), .A0 (nx3231), .A1 (nx10199), .A2 (nx10209)) ;
    nor02_2x ix3244 (.Y (nx3243), .A0 (nx616), .A1 (nx614)) ;
    nor03_2x ix617 (.Y (nx616), .A0 (nx3246), .A1 (nx9677), .A2 (nx10217)) ;
    dffr gen_1_cmp_mRegCmp_reg_Q_9 (.Q (gen_1_cmp_mReg_9), .QB (nx3246), .D (
         window_1__9), .CLK (start), .R (rst)) ;
    nor03_2x ix615 (.Y (nx614), .A0 (gen_1_cmp_mReg_9), .A1 (nx10007), .A2 (
             nx10225)) ;
    nand02 ix651 (.Y (gen_1_cmp_BSCmp_op2_10), .A0 (nx3251), .A1 (nx3257)) ;
    nor02_2x ix3252 (.Y (nx3251), .A0 (nx646), .A1 (nx642)) ;
    nor03_2x ix647 (.Y (nx646), .A0 (gen_1_cmp_mReg_9), .A1 (nx9683), .A2 (
             nx10193)) ;
    nor03_2x ix643 (.Y (nx642), .A0 (nx3246), .A1 (nx10199), .A2 (nx10209)) ;
    nor02_2x ix3258 (.Y (nx3257), .A0 (nx638), .A1 (nx636)) ;
    nor03_2x ix639 (.Y (nx638), .A0 (nx3261), .A1 (nx9677), .A2 (nx10217)) ;
    dffr gen_1_cmp_mRegCmp_reg_Q_10 (.Q (gen_1_cmp_mReg_10), .QB (nx3261), .D (
         window_1__10), .CLK (start), .R (rst)) ;
    nor03_2x ix637 (.Y (nx636), .A0 (gen_1_cmp_mReg_10), .A1 (nx10007), .A2 (
             nx10225)) ;
    nand02 ix673 (.Y (gen_1_cmp_BSCmp_op2_11), .A0 (nx3267), .A1 (nx3271)) ;
    nor02_2x ix3268 (.Y (nx3267), .A0 (nx668), .A1 (nx664)) ;
    nor03_2x ix669 (.Y (nx668), .A0 (gen_1_cmp_mReg_10), .A1 (nx9683), .A2 (
             nx10193)) ;
    nor03_2x ix665 (.Y (nx664), .A0 (nx3261), .A1 (nx10199), .A2 (nx10209)) ;
    nor02_2x ix3272 (.Y (nx3271), .A0 (nx660), .A1 (nx658)) ;
    nor03_2x ix661 (.Y (nx660), .A0 (nx3275), .A1 (nx9677), .A2 (nx10217)) ;
    dffr gen_1_cmp_mRegCmp_reg_Q_11 (.Q (gen_1_cmp_mReg_11), .QB (nx3275), .D (
         window_1__11), .CLK (start), .R (rst)) ;
    nor03_2x ix659 (.Y (nx658), .A0 (gen_1_cmp_mReg_11), .A1 (nx10007), .A2 (
             nx10225)) ;
    nand02 ix695 (.Y (gen_1_cmp_BSCmp_op2_12), .A0 (nx3281), .A1 (nx3287)) ;
    nor02_2x ix3282 (.Y (nx3281), .A0 (nx690), .A1 (nx686)) ;
    nor03_2x ix691 (.Y (nx690), .A0 (gen_1_cmp_mReg_11), .A1 (nx9683), .A2 (
             nx10193)) ;
    nor03_2x ix687 (.Y (nx686), .A0 (nx3275), .A1 (nx10199), .A2 (nx10209)) ;
    nor02_2x ix3288 (.Y (nx3287), .A0 (nx682), .A1 (nx680)) ;
    nor03_2x ix683 (.Y (nx682), .A0 (nx3290), .A1 (nx9679), .A2 (nx10217)) ;
    dffr gen_1_cmp_mRegCmp_reg_Q_12 (.Q (gen_1_cmp_mReg_12), .QB (nx3290), .D (
         window_1__12), .CLK (start), .R (rst)) ;
    nor03_2x ix681 (.Y (nx680), .A0 (gen_1_cmp_mReg_12), .A1 (nx10007), .A2 (
             nx10225)) ;
    nand02 ix717 (.Y (gen_1_cmp_BSCmp_op2_13), .A0 (nx3295), .A1 (nx3301)) ;
    nor02_2x ix3296 (.Y (nx3295), .A0 (nx712), .A1 (nx708)) ;
    nor03_2x ix713 (.Y (nx712), .A0 (gen_1_cmp_mReg_12), .A1 (nx9685), .A2 (
             nx10195)) ;
    nor03_2x ix709 (.Y (nx708), .A0 (nx3290), .A1 (nx10199), .A2 (nx10211)) ;
    nor02_2x ix3302 (.Y (nx3301), .A0 (nx704), .A1 (nx702)) ;
    nor03_2x ix705 (.Y (nx704), .A0 (nx3305), .A1 (nx9679), .A2 (nx10219)) ;
    dffr gen_1_cmp_mRegCmp_reg_Q_13 (.Q (gen_1_cmp_mReg_13), .QB (nx3305), .D (
         window_1__13), .CLK (start), .R (rst)) ;
    nor03_2x ix703 (.Y (nx702), .A0 (gen_1_cmp_mReg_13), .A1 (nx10007), .A2 (
             nx10227)) ;
    nand02 ix739 (.Y (gen_1_cmp_BSCmp_op2_14), .A0 (nx3311), .A1 (nx3315)) ;
    nor02_2x ix3312 (.Y (nx3311), .A0 (nx734), .A1 (nx730)) ;
    nor03_2x ix735 (.Y (nx734), .A0 (gen_1_cmp_mReg_13), .A1 (nx9685), .A2 (
             nx10195)) ;
    nor03_2x ix731 (.Y (nx730), .A0 (nx3305), .A1 (nx10201), .A2 (nx10211)) ;
    nor02_2x ix3316 (.Y (nx3315), .A0 (nx726), .A1 (nx724)) ;
    nor03_2x ix727 (.Y (nx726), .A0 (nx3319), .A1 (nx9679), .A2 (nx10219)) ;
    dffr gen_1_cmp_mRegCmp_reg_Q_14 (.Q (gen_1_cmp_mReg_14), .QB (nx3319), .D (
         window_1__14), .CLK (start), .R (rst)) ;
    nor03_2x ix725 (.Y (nx724), .A0 (gen_1_cmp_mReg_14), .A1 (nx10007), .A2 (
             nx10227)) ;
    nand02 ix761 (.Y (gen_1_cmp_BSCmp_op2_15), .A0 (nx3325), .A1 (nx3331)) ;
    nor02_2x ix3326 (.Y (nx3325), .A0 (nx756), .A1 (nx752)) ;
    nor03_2x ix757 (.Y (nx756), .A0 (gen_1_cmp_mReg_14), .A1 (nx9685), .A2 (
             nx10195)) ;
    nor03_2x ix753 (.Y (nx752), .A0 (nx3319), .A1 (nx10201), .A2 (nx10211)) ;
    nor02_2x ix3332 (.Y (nx3331), .A0 (nx748), .A1 (nx746)) ;
    nor03_2x ix749 (.Y (nx748), .A0 (nx3334), .A1 (nx9679), .A2 (nx10219)) ;
    dffr gen_1_cmp_mRegCmp_reg_Q_15 (.Q (gen_1_cmp_mReg_15), .QB (nx3334), .D (
         window_1__15), .CLK (start), .R (rst)) ;
    nor03_2x ix747 (.Y (nx746), .A0 (gen_1_cmp_mReg_15), .A1 (nx10009), .A2 (
             nx10227)) ;
    nand02 ix771 (.Y (gen_1_cmp_BSCmp_op2_16), .A0 (nx3339), .A1 (nx3331)) ;
    nor02_2x ix3340 (.Y (nx3339), .A0 (nx766), .A1 (nx762)) ;
    nor03_2x ix767 (.Y (nx766), .A0 (gen_1_cmp_mReg_15), .A1 (nx9685), .A2 (
             nx10195)) ;
    nor03_2x ix763 (.Y (nx762), .A0 (nx3334), .A1 (nx10201), .A2 (nx10211)) ;
    nand02 ix839 (.Y (gen_2_cmp_BSCmp_op2_1), .A0 (nx3347), .A1 (nx3365)) ;
    nor02_2x ix3348 (.Y (nx3347), .A0 (nx834), .A1 (nx830)) ;
    nor03_2x ix835 (.Y (nx834), .A0 (gen_2_cmp_mReg_0), .A1 (nx9669), .A2 (
             nx10231)) ;
    dffr gen_2_cmp_mRegCmp_reg_Q_0 (.Q (gen_2_cmp_mReg_0), .QB (nx3353), .D (
         window_2__0), .CLK (start), .R (rst)) ;
    inv01 ix3357 (.Y (nx3356), .A (gen_2_cmp_pMux_0)) ;
    nor03_2x ix831 (.Y (nx830), .A0 (nx3353), .A1 (nx10237), .A2 (nx10247)) ;
    inv02 ix3364 (.Y (nx3363), .A (gen_2_cmp_pMux_2)) ;
    nor02_2x ix3366 (.Y (nx3365), .A0 (nx820), .A1 (nx818)) ;
    nor03_2x ix821 (.Y (nx820), .A0 (nx3369), .A1 (nx9663), .A2 (nx10255)) ;
    dffr gen_2_cmp_mRegCmp_reg_Q_1 (.Q (gen_2_cmp_mReg_1), .QB (nx3369), .D (
         window_2__1), .CLK (start), .R (rst)) ;
    nor03_2x ix819 (.Y (nx818), .A0 (gen_2_cmp_mReg_1), .A1 (nx10011), .A2 (
             nx10263)) ;
    nor03_2x ix779 (.Y (nx778), .A0 (nx9669), .A1 (nx3363), .A2 (
             gen_2_cmp_pMux_0)) ;
    nand02 ix861 (.Y (gen_2_cmp_BSCmp_op2_2), .A0 (nx3380), .A1 (nx3387)) ;
    nor02_2x ix3382 (.Y (nx3380), .A0 (nx856), .A1 (nx852)) ;
    nor03_2x ix857 (.Y (nx856), .A0 (gen_2_cmp_mReg_1), .A1 (nx9669), .A2 (
             nx10231)) ;
    nor03_2x ix853 (.Y (nx852), .A0 (nx3369), .A1 (nx10237), .A2 (nx10247)) ;
    nor02_2x ix3388 (.Y (nx3387), .A0 (nx848), .A1 (nx846)) ;
    nor03_2x ix849 (.Y (nx848), .A0 (nx3391), .A1 (nx9663), .A2 (nx10255)) ;
    dffr gen_2_cmp_mRegCmp_reg_Q_2 (.Q (gen_2_cmp_mReg_2), .QB (nx3391), .D (
         window_2__2), .CLK (start), .R (rst)) ;
    nor03_2x ix847 (.Y (nx846), .A0 (gen_2_cmp_mReg_2), .A1 (nx10011), .A2 (
             nx10263)) ;
    nand02 ix883 (.Y (gen_2_cmp_BSCmp_op2_3), .A0 (nx3397), .A1 (nx3401)) ;
    nor02_2x ix3398 (.Y (nx3397), .A0 (nx878), .A1 (nx874)) ;
    nor03_2x ix879 (.Y (nx878), .A0 (gen_2_cmp_mReg_2), .A1 (nx9669), .A2 (
             nx10231)) ;
    nor03_2x ix875 (.Y (nx874), .A0 (nx3391), .A1 (nx10237), .A2 (nx10247)) ;
    nor02_2x ix3402 (.Y (nx3401), .A0 (nx870), .A1 (nx868)) ;
    nor03_2x ix871 (.Y (nx870), .A0 (nx3405), .A1 (nx9663), .A2 (nx10255)) ;
    dffr gen_2_cmp_mRegCmp_reg_Q_3 (.Q (gen_2_cmp_mReg_3), .QB (nx3405), .D (
         window_2__3), .CLK (start), .R (rst)) ;
    nor03_2x ix869 (.Y (nx868), .A0 (gen_2_cmp_mReg_3), .A1 (nx10011), .A2 (
             nx10263)) ;
    nand02 ix905 (.Y (gen_2_cmp_BSCmp_op2_4), .A0 (nx3411), .A1 (nx3415)) ;
    nor02_2x ix3412 (.Y (nx3411), .A0 (nx900), .A1 (nx896)) ;
    nor03_2x ix901 (.Y (nx900), .A0 (gen_2_cmp_mReg_3), .A1 (nx9669), .A2 (
             nx10231)) ;
    nor03_2x ix897 (.Y (nx896), .A0 (nx3405), .A1 (nx10237), .A2 (nx10247)) ;
    nor02_2x ix3416 (.Y (nx3415), .A0 (nx892), .A1 (nx890)) ;
    nor03_2x ix893 (.Y (nx892), .A0 (nx3419), .A1 (nx9663), .A2 (nx10255)) ;
    dffr gen_2_cmp_mRegCmp_reg_Q_4 (.Q (gen_2_cmp_mReg_4), .QB (nx3419), .D (
         window_2__4), .CLK (start), .R (rst)) ;
    nor03_2x ix891 (.Y (nx890), .A0 (gen_2_cmp_mReg_4), .A1 (nx10011), .A2 (
             nx10263)) ;
    nand02 ix927 (.Y (gen_2_cmp_BSCmp_op2_5), .A0 (nx3423), .A1 (nx3429)) ;
    nor02_2x ix3424 (.Y (nx3423), .A0 (nx922), .A1 (nx918)) ;
    nor03_2x ix923 (.Y (nx922), .A0 (gen_2_cmp_mReg_4), .A1 (nx9669), .A2 (
             nx10231)) ;
    nor03_2x ix919 (.Y (nx918), .A0 (nx3419), .A1 (nx10237), .A2 (nx10247)) ;
    nor02_2x ix3430 (.Y (nx3429), .A0 (nx914), .A1 (nx912)) ;
    nor03_2x ix915 (.Y (nx914), .A0 (nx3433), .A1 (nx9665), .A2 (nx10255)) ;
    dffr gen_2_cmp_mRegCmp_reg_Q_5 (.Q (gen_2_cmp_mReg_5), .QB (nx3433), .D (
         window_2__5), .CLK (start), .R (rst)) ;
    nor03_2x ix913 (.Y (nx912), .A0 (gen_2_cmp_mReg_5), .A1 (nx10011), .A2 (
             nx10263)) ;
    nand02 ix949 (.Y (gen_2_cmp_BSCmp_op2_6), .A0 (nx3437), .A1 (nx3443)) ;
    nor02_2x ix3438 (.Y (nx3437), .A0 (nx944), .A1 (nx940)) ;
    nor03_2x ix945 (.Y (nx944), .A0 (gen_2_cmp_mReg_5), .A1 (nx9671), .A2 (
             nx10231)) ;
    nor03_2x ix941 (.Y (nx940), .A0 (nx3433), .A1 (nx10237), .A2 (nx10247)) ;
    nor02_2x ix3444 (.Y (nx3443), .A0 (nx936), .A1 (nx934)) ;
    nor03_2x ix937 (.Y (nx936), .A0 (nx3446), .A1 (nx9665), .A2 (nx10255)) ;
    dffr gen_2_cmp_mRegCmp_reg_Q_6 (.Q (gen_2_cmp_mReg_6), .QB (nx3446), .D (
         window_2__6), .CLK (start), .R (rst)) ;
    nor03_2x ix935 (.Y (nx934), .A0 (gen_2_cmp_mReg_6), .A1 (nx10011), .A2 (
             nx10263)) ;
    nand02 ix971 (.Y (gen_2_cmp_BSCmp_op2_7), .A0 (nx3453), .A1 (nx3459)) ;
    nor02_2x ix3454 (.Y (nx3453), .A0 (nx966), .A1 (nx962)) ;
    nor03_2x ix967 (.Y (nx966), .A0 (gen_2_cmp_mReg_6), .A1 (nx9671), .A2 (
             nx10233)) ;
    nor03_2x ix963 (.Y (nx962), .A0 (nx3446), .A1 (nx10239), .A2 (nx10249)) ;
    nor02_2x ix3460 (.Y (nx3459), .A0 (nx958), .A1 (nx956)) ;
    nor03_2x ix959 (.Y (nx958), .A0 (nx3463), .A1 (nx9665), .A2 (nx10257)) ;
    dffr gen_2_cmp_mRegCmp_reg_Q_7 (.Q (gen_2_cmp_mReg_7), .QB (nx3463), .D (
         window_2__7), .CLK (start), .R (rst)) ;
    nor03_2x ix957 (.Y (nx956), .A0 (gen_2_cmp_mReg_7), .A1 (nx10011), .A2 (
             nx10265)) ;
    nand02 ix993 (.Y (gen_2_cmp_BSCmp_op2_8), .A0 (nx3469), .A1 (nx3475)) ;
    nor02_2x ix3470 (.Y (nx3469), .A0 (nx988), .A1 (nx984)) ;
    nor03_2x ix989 (.Y (nx988), .A0 (gen_2_cmp_mReg_7), .A1 (nx9671), .A2 (
             nx10233)) ;
    nor03_2x ix985 (.Y (nx984), .A0 (nx3463), .A1 (nx10239), .A2 (nx10249)) ;
    nor02_2x ix3476 (.Y (nx3475), .A0 (nx980), .A1 (nx978)) ;
    nor03_2x ix981 (.Y (nx980), .A0 (nx3479), .A1 (nx9665), .A2 (nx10257)) ;
    dffr gen_2_cmp_mRegCmp_reg_Q_8 (.Q (gen_2_cmp_mReg_8), .QB (nx3479), .D (
         window_2__8), .CLK (start), .R (rst)) ;
    nor03_2x ix979 (.Y (nx978), .A0 (gen_2_cmp_mReg_8), .A1 (nx10013), .A2 (
             nx10265)) ;
    nand02 ix1015 (.Y (gen_2_cmp_BSCmp_op2_9), .A0 (nx3484), .A1 (nx3488)) ;
    nor02_2x ix3485 (.Y (nx3484), .A0 (nx1010), .A1 (nx1006)) ;
    nor03_2x ix1011 (.Y (nx1010), .A0 (gen_2_cmp_mReg_8), .A1 (nx9671), .A2 (
             nx10233)) ;
    nor03_2x ix1007 (.Y (nx1006), .A0 (nx3479), .A1 (nx10239), .A2 (nx10249)) ;
    nor02_2x ix3489 (.Y (nx3488), .A0 (nx1002), .A1 (nx1000)) ;
    nor03_2x ix1003 (.Y (nx1002), .A0 (nx3491), .A1 (nx9665), .A2 (nx10257)) ;
    dffr gen_2_cmp_mRegCmp_reg_Q_9 (.Q (gen_2_cmp_mReg_9), .QB (nx3491), .D (
         window_2__9), .CLK (start), .R (rst)) ;
    nor03_2x ix1001 (.Y (nx1000), .A0 (gen_2_cmp_mReg_9), .A1 (nx10013), .A2 (
             nx10265)) ;
    nand02 ix1037 (.Y (gen_2_cmp_BSCmp_op2_10), .A0 (nx3497), .A1 (nx3503)) ;
    nor02_2x ix3498 (.Y (nx3497), .A0 (nx1032), .A1 (nx1028)) ;
    nor03_2x ix1033 (.Y (nx1032), .A0 (gen_2_cmp_mReg_9), .A1 (nx9671), .A2 (
             nx10233)) ;
    nor03_2x ix1029 (.Y (nx1028), .A0 (nx3491), .A1 (nx10239), .A2 (nx10249)) ;
    nor02_2x ix3504 (.Y (nx3503), .A0 (nx1024), .A1 (nx1022)) ;
    nor03_2x ix1025 (.Y (nx1024), .A0 (nx3507), .A1 (nx9665), .A2 (nx10257)) ;
    dffr gen_2_cmp_mRegCmp_reg_Q_10 (.Q (gen_2_cmp_mReg_10), .QB (nx3507), .D (
         window_2__10), .CLK (start), .R (rst)) ;
    nor03_2x ix1023 (.Y (nx1022), .A0 (gen_2_cmp_mReg_10), .A1 (nx10013), .A2 (
             nx10265)) ;
    nand02 ix1059 (.Y (gen_2_cmp_BSCmp_op2_11), .A0 (nx3513), .A1 (nx3517)) ;
    nor02_2x ix3514 (.Y (nx3513), .A0 (nx1054), .A1 (nx1050)) ;
    nor03_2x ix1055 (.Y (nx1054), .A0 (gen_2_cmp_mReg_10), .A1 (nx9671), .A2 (
             nx10233)) ;
    nor03_2x ix1051 (.Y (nx1050), .A0 (nx3507), .A1 (nx10239), .A2 (nx10249)) ;
    nor02_2x ix3518 (.Y (nx3517), .A0 (nx1046), .A1 (nx1044)) ;
    nor03_2x ix1047 (.Y (nx1046), .A0 (nx3521), .A1 (nx9665), .A2 (nx10257)) ;
    dffr gen_2_cmp_mRegCmp_reg_Q_11 (.Q (gen_2_cmp_mReg_11), .QB (nx3521), .D (
         window_2__11), .CLK (start), .R (rst)) ;
    nor03_2x ix1045 (.Y (nx1044), .A0 (gen_2_cmp_mReg_11), .A1 (nx10013), .A2 (
             nx10265)) ;
    nand02 ix1081 (.Y (gen_2_cmp_BSCmp_op2_12), .A0 (nx3527), .A1 (nx3533)) ;
    nor02_2x ix3528 (.Y (nx3527), .A0 (nx1076), .A1 (nx1072)) ;
    nor03_2x ix1077 (.Y (nx1076), .A0 (gen_2_cmp_mReg_11), .A1 (nx9671), .A2 (
             nx10233)) ;
    nor03_2x ix1073 (.Y (nx1072), .A0 (nx3521), .A1 (nx10239), .A2 (nx10249)) ;
    nor02_2x ix3534 (.Y (nx3533), .A0 (nx1068), .A1 (nx1066)) ;
    nor03_2x ix1069 (.Y (nx1068), .A0 (nx3537), .A1 (nx9667), .A2 (nx10257)) ;
    dffr gen_2_cmp_mRegCmp_reg_Q_12 (.Q (gen_2_cmp_mReg_12), .QB (nx3537), .D (
         window_2__12), .CLK (start), .R (rst)) ;
    nor03_2x ix1067 (.Y (nx1066), .A0 (gen_2_cmp_mReg_12), .A1 (nx10013), .A2 (
             nx10265)) ;
    nand02 ix1103 (.Y (gen_2_cmp_BSCmp_op2_13), .A0 (nx3543), .A1 (nx3547)) ;
    nor02_2x ix3544 (.Y (nx3543), .A0 (nx1098), .A1 (nx1094)) ;
    nor03_2x ix1099 (.Y (nx1098), .A0 (gen_2_cmp_mReg_12), .A1 (nx9673), .A2 (
             nx10235)) ;
    nor03_2x ix1095 (.Y (nx1094), .A0 (nx3537), .A1 (nx10239), .A2 (nx10251)) ;
    nor02_2x ix3548 (.Y (nx3547), .A0 (nx1090), .A1 (nx1088)) ;
    nor03_2x ix1091 (.Y (nx1090), .A0 (nx3551), .A1 (nx9667), .A2 (nx10259)) ;
    dffr gen_2_cmp_mRegCmp_reg_Q_13 (.Q (gen_2_cmp_mReg_13), .QB (nx3551), .D (
         window_2__13), .CLK (start), .R (rst)) ;
    nor03_2x ix1089 (.Y (nx1088), .A0 (gen_2_cmp_mReg_13), .A1 (nx10013), .A2 (
             nx10267)) ;
    nand02 ix1125 (.Y (gen_2_cmp_BSCmp_op2_14), .A0 (nx3557), .A1 (nx3563)) ;
    nor02_2x ix3558 (.Y (nx3557), .A0 (nx1120), .A1 (nx1116)) ;
    nor03_2x ix1121 (.Y (nx1120), .A0 (gen_2_cmp_mReg_13), .A1 (nx9673), .A2 (
             nx10235)) ;
    nor03_2x ix1117 (.Y (nx1116), .A0 (nx3551), .A1 (nx10241), .A2 (nx10251)) ;
    nor02_2x ix3564 (.Y (nx3563), .A0 (nx1112), .A1 (nx1110)) ;
    nor03_2x ix1113 (.Y (nx1112), .A0 (nx3566), .A1 (nx9667), .A2 (nx10259)) ;
    dffr gen_2_cmp_mRegCmp_reg_Q_14 (.Q (gen_2_cmp_mReg_14), .QB (nx3566), .D (
         window_2__14), .CLK (start), .R (rst)) ;
    nor03_2x ix1111 (.Y (nx1110), .A0 (gen_2_cmp_mReg_14), .A1 (nx10013), .A2 (
             nx10267)) ;
    nand02 ix1147 (.Y (gen_2_cmp_BSCmp_op2_15), .A0 (nx3571), .A1 (nx3577)) ;
    nor02_2x ix3572 (.Y (nx3571), .A0 (nx1142), .A1 (nx1138)) ;
    nor03_2x ix1143 (.Y (nx1142), .A0 (gen_2_cmp_mReg_14), .A1 (nx9673), .A2 (
             nx10235)) ;
    nor03_2x ix1139 (.Y (nx1138), .A0 (nx3566), .A1 (nx10241), .A2 (nx10251)) ;
    nor02_2x ix3578 (.Y (nx3577), .A0 (nx1134), .A1 (nx1132)) ;
    nor03_2x ix1135 (.Y (nx1134), .A0 (nx3581), .A1 (nx9667), .A2 (nx10259)) ;
    dffr gen_2_cmp_mRegCmp_reg_Q_15 (.Q (gen_2_cmp_mReg_15), .QB (nx3581), .D (
         window_2__15), .CLK (start), .R (rst)) ;
    nor03_2x ix1133 (.Y (nx1132), .A0 (gen_2_cmp_mReg_15), .A1 (nx10015), .A2 (
             nx10267)) ;
    nand02 ix1157 (.Y (gen_2_cmp_BSCmp_op2_16), .A0 (nx3587), .A1 (nx3577)) ;
    nor02_2x ix3588 (.Y (nx3587), .A0 (nx1152), .A1 (nx1148)) ;
    nor03_2x ix1153 (.Y (nx1152), .A0 (gen_2_cmp_mReg_15), .A1 (nx9673), .A2 (
             nx10235)) ;
    nor03_2x ix1149 (.Y (nx1148), .A0 (nx3581), .A1 (nx10241), .A2 (nx10251)) ;
    nand02 ix1225 (.Y (gen_3_cmp_BSCmp_op2_1), .A0 (nx3593), .A1 (nx3613)) ;
    nor02_2x ix3594 (.Y (nx3593), .A0 (nx1220), .A1 (nx1216)) ;
    nor03_2x ix1221 (.Y (nx1220), .A0 (gen_3_cmp_mReg_0), .A1 (nx9657), .A2 (
             nx10271)) ;
    dffr gen_3_cmp_mRegCmp_reg_Q_0 (.Q (gen_3_cmp_mReg_0), .QB (nx3599), .D (
         window_3__0), .CLK (start), .R (rst)) ;
    inv01 ix3604 (.Y (nx3603), .A (gen_3_cmp_pMux_0)) ;
    nor03_2x ix1217 (.Y (nx1216), .A0 (nx3599), .A1 (nx10277), .A2 (nx10287)) ;
    inv02 ix3612 (.Y (nx3611), .A (gen_3_cmp_pMux_2)) ;
    nor02_2x ix3614 (.Y (nx3613), .A0 (nx1206), .A1 (nx1204)) ;
    nor03_2x ix1207 (.Y (nx1206), .A0 (nx3617), .A1 (nx9651), .A2 (nx10295)) ;
    dffr gen_3_cmp_mRegCmp_reg_Q_1 (.Q (gen_3_cmp_mReg_1), .QB (nx3617), .D (
         window_3__1), .CLK (start), .R (rst)) ;
    nor03_2x ix1205 (.Y (nx1204), .A0 (gen_3_cmp_mReg_1), .A1 (nx10017), .A2 (
             nx10303)) ;
    nor03_2x ix1165 (.Y (nx1164), .A0 (nx9657), .A1 (nx3611), .A2 (
             gen_3_cmp_pMux_0)) ;
    nand02 ix1247 (.Y (gen_3_cmp_BSCmp_op2_2), .A0 (nx3629), .A1 (nx3633)) ;
    nor02_2x ix3630 (.Y (nx3629), .A0 (nx1242), .A1 (nx1238)) ;
    nor03_2x ix1243 (.Y (nx1242), .A0 (gen_3_cmp_mReg_1), .A1 (nx9657), .A2 (
             nx10271)) ;
    nor03_2x ix1239 (.Y (nx1238), .A0 (nx3617), .A1 (nx10277), .A2 (nx10287)) ;
    nor02_2x ix3634 (.Y (nx3633), .A0 (nx1234), .A1 (nx1232)) ;
    nor03_2x ix1235 (.Y (nx1234), .A0 (nx3637), .A1 (nx9651), .A2 (nx10295)) ;
    dffr gen_3_cmp_mRegCmp_reg_Q_2 (.Q (gen_3_cmp_mReg_2), .QB (nx3637), .D (
         window_3__2), .CLK (start), .R (rst)) ;
    nor03_2x ix1233 (.Y (nx1232), .A0 (gen_3_cmp_mReg_2), .A1 (nx10017), .A2 (
             nx10303)) ;
    nand02 ix1269 (.Y (gen_3_cmp_BSCmp_op2_3), .A0 (nx3643), .A1 (nx3647)) ;
    nor02_2x ix3644 (.Y (nx3643), .A0 (nx1264), .A1 (nx1260)) ;
    nor03_2x ix1265 (.Y (nx1264), .A0 (gen_3_cmp_mReg_2), .A1 (nx9657), .A2 (
             nx10271)) ;
    nor03_2x ix1261 (.Y (nx1260), .A0 (nx3637), .A1 (nx10277), .A2 (nx10287)) ;
    nor02_2x ix3648 (.Y (nx3647), .A0 (nx1256), .A1 (nx1254)) ;
    nor03_2x ix1257 (.Y (nx1256), .A0 (nx3651), .A1 (nx9651), .A2 (nx10295)) ;
    dffr gen_3_cmp_mRegCmp_reg_Q_3 (.Q (gen_3_cmp_mReg_3), .QB (nx3651), .D (
         window_3__3), .CLK (start), .R (rst)) ;
    nor03_2x ix1255 (.Y (nx1254), .A0 (gen_3_cmp_mReg_3), .A1 (nx10017), .A2 (
             nx10303)) ;
    nand02 ix1291 (.Y (gen_3_cmp_BSCmp_op2_4), .A0 (nx3655), .A1 (nx3661)) ;
    nor02_2x ix3656 (.Y (nx3655), .A0 (nx1286), .A1 (nx1282)) ;
    nor03_2x ix1287 (.Y (nx1286), .A0 (gen_3_cmp_mReg_3), .A1 (nx9657), .A2 (
             nx10271)) ;
    nor03_2x ix1283 (.Y (nx1282), .A0 (nx3651), .A1 (nx10277), .A2 (nx10287)) ;
    nor02_2x ix3662 (.Y (nx3661), .A0 (nx1278), .A1 (nx1276)) ;
    nor03_2x ix1279 (.Y (nx1278), .A0 (nx3665), .A1 (nx9651), .A2 (nx10295)) ;
    dffr gen_3_cmp_mRegCmp_reg_Q_4 (.Q (gen_3_cmp_mReg_4), .QB (nx3665), .D (
         window_3__4), .CLK (start), .R (rst)) ;
    nor03_2x ix1277 (.Y (nx1276), .A0 (gen_3_cmp_mReg_4), .A1 (nx10017), .A2 (
             nx10303)) ;
    nand02 ix1313 (.Y (gen_3_cmp_BSCmp_op2_5), .A0 (nx3669), .A1 (nx3675)) ;
    nor02_2x ix3670 (.Y (nx3669), .A0 (nx1308), .A1 (nx1304)) ;
    nor03_2x ix1309 (.Y (nx1308), .A0 (gen_3_cmp_mReg_4), .A1 (nx9657), .A2 (
             nx10271)) ;
    nor03_2x ix1305 (.Y (nx1304), .A0 (nx3665), .A1 (nx10277), .A2 (nx10287)) ;
    nor02_2x ix3676 (.Y (nx3675), .A0 (nx1300), .A1 (nx1298)) ;
    nor03_2x ix1301 (.Y (nx1300), .A0 (nx3678), .A1 (nx9653), .A2 (nx10295)) ;
    dffr gen_3_cmp_mRegCmp_reg_Q_5 (.Q (gen_3_cmp_mReg_5), .QB (nx3678), .D (
         window_3__5), .CLK (start), .R (rst)) ;
    nor03_2x ix1299 (.Y (nx1298), .A0 (gen_3_cmp_mReg_5), .A1 (nx10017), .A2 (
             nx10303)) ;
    nand02 ix1335 (.Y (gen_3_cmp_BSCmp_op2_6), .A0 (nx3685), .A1 (nx3691)) ;
    nor02_2x ix3686 (.Y (nx3685), .A0 (nx1330), .A1 (nx1326)) ;
    nor03_2x ix1331 (.Y (nx1330), .A0 (gen_3_cmp_mReg_5), .A1 (nx9659), .A2 (
             nx10271)) ;
    nor03_2x ix1327 (.Y (nx1326), .A0 (nx3678), .A1 (nx10277), .A2 (nx10287)) ;
    nor02_2x ix3692 (.Y (nx3691), .A0 (nx1322), .A1 (nx1320)) ;
    nor03_2x ix1323 (.Y (nx1322), .A0 (nx3695), .A1 (nx9653), .A2 (nx10295)) ;
    dffr gen_3_cmp_mRegCmp_reg_Q_6 (.Q (gen_3_cmp_mReg_6), .QB (nx3695), .D (
         window_3__6), .CLK (start), .R (rst)) ;
    nor03_2x ix1321 (.Y (nx1320), .A0 (gen_3_cmp_mReg_6), .A1 (nx10017), .A2 (
             nx10303)) ;
    nand02 ix1357 (.Y (gen_3_cmp_BSCmp_op2_7), .A0 (nx3699), .A1 (nx3705)) ;
    nor02_2x ix3700 (.Y (nx3699), .A0 (nx1352), .A1 (nx1348)) ;
    nor03_2x ix1353 (.Y (nx1352), .A0 (gen_3_cmp_mReg_6), .A1 (nx9659), .A2 (
             nx10273)) ;
    nor03_2x ix1349 (.Y (nx1348), .A0 (nx3695), .A1 (nx10279), .A2 (nx10289)) ;
    nor02_2x ix3706 (.Y (nx3705), .A0 (nx1344), .A1 (nx1342)) ;
    nor03_2x ix1345 (.Y (nx1344), .A0 (nx3709), .A1 (nx9653), .A2 (nx10297)) ;
    dffr gen_3_cmp_mRegCmp_reg_Q_7 (.Q (gen_3_cmp_mReg_7), .QB (nx3709), .D (
         window_3__7), .CLK (start), .R (rst)) ;
    nor03_2x ix1343 (.Y (nx1342), .A0 (gen_3_cmp_mReg_7), .A1 (nx10017), .A2 (
             nx10305)) ;
    nand02 ix1379 (.Y (gen_3_cmp_BSCmp_op2_8), .A0 (nx3713), .A1 (nx3719)) ;
    nor02_2x ix3714 (.Y (nx3713), .A0 (nx1374), .A1 (nx1370)) ;
    nor03_2x ix1375 (.Y (nx1374), .A0 (gen_3_cmp_mReg_7), .A1 (nx9659), .A2 (
             nx10273)) ;
    nor03_2x ix1371 (.Y (nx1370), .A0 (nx3709), .A1 (nx10279), .A2 (nx10289)) ;
    nor02_2x ix3720 (.Y (nx3719), .A0 (nx1366), .A1 (nx1364)) ;
    nor03_2x ix1367 (.Y (nx1366), .A0 (nx3722), .A1 (nx9653), .A2 (nx10297)) ;
    dffr gen_3_cmp_mRegCmp_reg_Q_8 (.Q (gen_3_cmp_mReg_8), .QB (nx3722), .D (
         window_3__8), .CLK (start), .R (rst)) ;
    nor03_2x ix1365 (.Y (nx1364), .A0 (gen_3_cmp_mReg_8), .A1 (nx10019), .A2 (
             nx10305)) ;
    nand02 ix1401 (.Y (gen_3_cmp_BSCmp_op2_9), .A0 (nx3729), .A1 (nx3735)) ;
    nor02_2x ix3730 (.Y (nx3729), .A0 (nx1396), .A1 (nx1392)) ;
    nor03_2x ix1397 (.Y (nx1396), .A0 (gen_3_cmp_mReg_8), .A1 (nx9659), .A2 (
             nx10273)) ;
    nor03_2x ix1393 (.Y (nx1392), .A0 (nx3722), .A1 (nx10279), .A2 (nx10289)) ;
    nor02_2x ix3736 (.Y (nx3735), .A0 (nx1388), .A1 (nx1386)) ;
    nor03_2x ix1389 (.Y (nx1388), .A0 (nx3739), .A1 (nx9653), .A2 (nx10297)) ;
    dffr gen_3_cmp_mRegCmp_reg_Q_9 (.Q (gen_3_cmp_mReg_9), .QB (nx3739), .D (
         window_3__9), .CLK (start), .R (rst)) ;
    nor03_2x ix1387 (.Y (nx1386), .A0 (gen_3_cmp_mReg_9), .A1 (nx10019), .A2 (
             nx10305)) ;
    nand02 ix1423 (.Y (gen_3_cmp_BSCmp_op2_10), .A0 (nx3743), .A1 (nx3749)) ;
    nor02_2x ix3744 (.Y (nx3743), .A0 (nx1418), .A1 (nx1414)) ;
    nor03_2x ix1419 (.Y (nx1418), .A0 (gen_3_cmp_mReg_9), .A1 (nx9659), .A2 (
             nx10273)) ;
    nor03_2x ix1415 (.Y (nx1414), .A0 (nx3739), .A1 (nx10279), .A2 (nx10289)) ;
    nor02_2x ix3750 (.Y (nx3749), .A0 (nx1410), .A1 (nx1408)) ;
    nor03_2x ix1411 (.Y (nx1410), .A0 (nx3753), .A1 (nx9653), .A2 (nx10297)) ;
    dffr gen_3_cmp_mRegCmp_reg_Q_10 (.Q (gen_3_cmp_mReg_10), .QB (nx3753), .D (
         window_3__10), .CLK (start), .R (rst)) ;
    nor03_2x ix1409 (.Y (nx1408), .A0 (gen_3_cmp_mReg_10), .A1 (nx10019), .A2 (
             nx10305)) ;
    nand02 ix1445 (.Y (gen_3_cmp_BSCmp_op2_11), .A0 (nx3757), .A1 (nx3763)) ;
    nor02_2x ix3758 (.Y (nx3757), .A0 (nx1440), .A1 (nx1436)) ;
    nor03_2x ix1441 (.Y (nx1440), .A0 (gen_3_cmp_mReg_10), .A1 (nx9659), .A2 (
             nx10273)) ;
    nor03_2x ix1437 (.Y (nx1436), .A0 (nx3753), .A1 (nx10279), .A2 (nx10289)) ;
    nor02_2x ix3764 (.Y (nx3763), .A0 (nx1432), .A1 (nx1430)) ;
    nor03_2x ix1433 (.Y (nx1432), .A0 (nx3766), .A1 (nx9653), .A2 (nx10297)) ;
    dffr gen_3_cmp_mRegCmp_reg_Q_11 (.Q (gen_3_cmp_mReg_11), .QB (nx3766), .D (
         window_3__11), .CLK (start), .R (rst)) ;
    nor03_2x ix1431 (.Y (nx1430), .A0 (gen_3_cmp_mReg_11), .A1 (nx10019), .A2 (
             nx10305)) ;
    nand02 ix1467 (.Y (gen_3_cmp_BSCmp_op2_12), .A0 (nx3773), .A1 (nx3779)) ;
    nor02_2x ix3774 (.Y (nx3773), .A0 (nx1462), .A1 (nx1458)) ;
    nor03_2x ix1463 (.Y (nx1462), .A0 (gen_3_cmp_mReg_11), .A1 (nx9659), .A2 (
             nx10273)) ;
    nor03_2x ix1459 (.Y (nx1458), .A0 (nx3766), .A1 (nx10279), .A2 (nx10289)) ;
    nor02_2x ix3780 (.Y (nx3779), .A0 (nx1454), .A1 (nx1452)) ;
    nor03_2x ix1455 (.Y (nx1454), .A0 (nx3783), .A1 (nx9655), .A2 (nx10297)) ;
    dffr gen_3_cmp_mRegCmp_reg_Q_12 (.Q (gen_3_cmp_mReg_12), .QB (nx3783), .D (
         window_3__12), .CLK (start), .R (rst)) ;
    nor03_2x ix1453 (.Y (nx1452), .A0 (gen_3_cmp_mReg_12), .A1 (nx10019), .A2 (
             nx10305)) ;
    nand02 ix1489 (.Y (gen_3_cmp_BSCmp_op2_13), .A0 (nx3787), .A1 (nx3793)) ;
    nor02_2x ix3788 (.Y (nx3787), .A0 (nx1484), .A1 (nx1480)) ;
    nor03_2x ix1485 (.Y (nx1484), .A0 (gen_3_cmp_mReg_12), .A1 (nx9661), .A2 (
             nx10275)) ;
    nor03_2x ix1481 (.Y (nx1480), .A0 (nx3783), .A1 (nx10279), .A2 (nx10291)) ;
    nor02_2x ix3794 (.Y (nx3793), .A0 (nx1476), .A1 (nx1474)) ;
    nor03_2x ix1477 (.Y (nx1476), .A0 (nx3797), .A1 (nx9655), .A2 (nx10299)) ;
    dffr gen_3_cmp_mRegCmp_reg_Q_13 (.Q (gen_3_cmp_mReg_13), .QB (nx3797), .D (
         window_3__13), .CLK (start), .R (rst)) ;
    nor03_2x ix1475 (.Y (nx1474), .A0 (gen_3_cmp_mReg_13), .A1 (nx10019), .A2 (
             nx10307)) ;
    nand02 ix1511 (.Y (gen_3_cmp_BSCmp_op2_14), .A0 (nx3801), .A1 (nx3807)) ;
    nor02_2x ix3802 (.Y (nx3801), .A0 (nx1506), .A1 (nx1502)) ;
    nor03_2x ix1507 (.Y (nx1506), .A0 (gen_3_cmp_mReg_13), .A1 (nx9661), .A2 (
             nx10275)) ;
    nor03_2x ix1503 (.Y (nx1502), .A0 (nx3797), .A1 (nx10281), .A2 (nx10291)) ;
    nor02_2x ix3808 (.Y (nx3807), .A0 (nx1498), .A1 (nx1496)) ;
    nor03_2x ix1499 (.Y (nx1498), .A0 (nx3810), .A1 (nx9655), .A2 (nx10299)) ;
    dffr gen_3_cmp_mRegCmp_reg_Q_14 (.Q (gen_3_cmp_mReg_14), .QB (nx3810), .D (
         window_3__14), .CLK (start), .R (rst)) ;
    nor03_2x ix1497 (.Y (nx1496), .A0 (gen_3_cmp_mReg_14), .A1 (nx10019), .A2 (
             nx10307)) ;
    nand02 ix1533 (.Y (gen_3_cmp_BSCmp_op2_15), .A0 (nx3817), .A1 (nx3823)) ;
    nor02_2x ix3818 (.Y (nx3817), .A0 (nx1528), .A1 (nx1524)) ;
    nor03_2x ix1529 (.Y (nx1528), .A0 (gen_3_cmp_mReg_14), .A1 (nx9661), .A2 (
             nx10275)) ;
    nor03_2x ix1525 (.Y (nx1524), .A0 (nx3810), .A1 (nx10281), .A2 (nx10291)) ;
    nor02_2x ix3824 (.Y (nx3823), .A0 (nx1520), .A1 (nx1518)) ;
    nor03_2x ix1521 (.Y (nx1520), .A0 (nx3827), .A1 (nx9655), .A2 (nx10299)) ;
    dffr gen_3_cmp_mRegCmp_reg_Q_15 (.Q (gen_3_cmp_mReg_15), .QB (nx3827), .D (
         window_3__15), .CLK (start), .R (rst)) ;
    nor03_2x ix1519 (.Y (nx1518), .A0 (gen_3_cmp_mReg_15), .A1 (nx10021), .A2 (
             nx10307)) ;
    nand02 ix1543 (.Y (gen_3_cmp_BSCmp_op2_16), .A0 (nx3831), .A1 (nx3823)) ;
    nor02_2x ix3832 (.Y (nx3831), .A0 (nx1538), .A1 (nx1534)) ;
    nor03_2x ix1539 (.Y (nx1538), .A0 (gen_3_cmp_mReg_15), .A1 (nx9661), .A2 (
             nx10275)) ;
    nor03_2x ix1535 (.Y (nx1534), .A0 (nx3827), .A1 (nx10281), .A2 (nx10291)) ;
    nand02 ix1611 (.Y (gen_4_cmp_BSCmp_op2_1), .A0 (nx3839), .A1 (nx3859)) ;
    nor02_2x ix3840 (.Y (nx3839), .A0 (nx1606), .A1 (nx1602)) ;
    nor03_2x ix1607 (.Y (nx1606), .A0 (gen_4_cmp_mReg_0), .A1 (nx9645), .A2 (
             nx10311)) ;
    dffr gen_4_cmp_mRegCmp_reg_Q_0 (.Q (gen_4_cmp_mReg_0), .QB (nx3845), .D (
         window_4__0), .CLK (start), .R (rst)) ;
    inv01 ix3850 (.Y (nx3849), .A (gen_4_cmp_pMux_0)) ;
    nor03_2x ix1603 (.Y (nx1602), .A0 (nx3845), .A1 (nx10317), .A2 (nx10327)) ;
    inv02 ix3858 (.Y (nx3857), .A (gen_4_cmp_pMux_2)) ;
    nor02_2x ix3860 (.Y (nx3859), .A0 (nx1592), .A1 (nx1590)) ;
    nor03_2x ix1593 (.Y (nx1592), .A0 (nx3863), .A1 (nx9639), .A2 (nx10335)) ;
    dffr gen_4_cmp_mRegCmp_reg_Q_1 (.Q (gen_4_cmp_mReg_1), .QB (nx3863), .D (
         window_4__1), .CLK (start), .R (rst)) ;
    nor03_2x ix1591 (.Y (nx1590), .A0 (gen_4_cmp_mReg_1), .A1 (nx10023), .A2 (
             nx10343)) ;
    nor03_2x ix1551 (.Y (nx1550), .A0 (nx9645), .A1 (nx3857), .A2 (
             gen_4_cmp_pMux_0)) ;
    nand02 ix1633 (.Y (gen_4_cmp_BSCmp_op2_2), .A0 (nx3873), .A1 (nx3877)) ;
    nor02_2x ix3874 (.Y (nx3873), .A0 (nx1628), .A1 (nx1624)) ;
    nor03_2x ix1629 (.Y (nx1628), .A0 (gen_4_cmp_mReg_1), .A1 (nx9645), .A2 (
             nx10311)) ;
    nor03_2x ix1625 (.Y (nx1624), .A0 (nx3863), .A1 (nx10317), .A2 (nx10327)) ;
    nor02_2x ix3878 (.Y (nx3877), .A0 (nx1620), .A1 (nx1618)) ;
    nor03_2x ix1621 (.Y (nx1620), .A0 (nx3881), .A1 (nx9639), .A2 (nx10335)) ;
    dffr gen_4_cmp_mRegCmp_reg_Q_2 (.Q (gen_4_cmp_mReg_2), .QB (nx3881), .D (
         window_4__2), .CLK (start), .R (rst)) ;
    nor03_2x ix1619 (.Y (nx1618), .A0 (gen_4_cmp_mReg_2), .A1 (nx10023), .A2 (
             nx10343)) ;
    nand02 ix1655 (.Y (gen_4_cmp_BSCmp_op2_3), .A0 (nx3887), .A1 (nx3893)) ;
    nor02_2x ix3888 (.Y (nx3887), .A0 (nx1650), .A1 (nx1646)) ;
    nor03_2x ix1651 (.Y (nx1650), .A0 (gen_4_cmp_mReg_2), .A1 (nx9645), .A2 (
             nx10311)) ;
    nor03_2x ix1647 (.Y (nx1646), .A0 (nx3881), .A1 (nx10317), .A2 (nx10327)) ;
    nor02_2x ix3894 (.Y (nx3893), .A0 (nx1642), .A1 (nx1640)) ;
    nor03_2x ix1643 (.Y (nx1642), .A0 (nx3897), .A1 (nx9639), .A2 (nx10335)) ;
    dffr gen_4_cmp_mRegCmp_reg_Q_3 (.Q (gen_4_cmp_mReg_3), .QB (nx3897), .D (
         window_4__3), .CLK (start), .R (rst)) ;
    nor03_2x ix1641 (.Y (nx1640), .A0 (gen_4_cmp_mReg_3), .A1 (nx10023), .A2 (
             nx10343)) ;
    nand02 ix1677 (.Y (gen_4_cmp_BSCmp_op2_4), .A0 (nx3902), .A1 (nx3907)) ;
    nor02_2x ix3903 (.Y (nx3902), .A0 (nx1672), .A1 (nx1668)) ;
    nor03_2x ix1673 (.Y (nx1672), .A0 (gen_4_cmp_mReg_3), .A1 (nx9645), .A2 (
             nx10311)) ;
    nor03_2x ix1669 (.Y (nx1668), .A0 (nx3897), .A1 (nx10317), .A2 (nx10327)) ;
    nor02_2x ix3908 (.Y (nx3907), .A0 (nx1664), .A1 (nx1662)) ;
    nor03_2x ix1665 (.Y (nx1664), .A0 (nx3911), .A1 (nx9639), .A2 (nx10335)) ;
    dffr gen_4_cmp_mRegCmp_reg_Q_4 (.Q (gen_4_cmp_mReg_4), .QB (nx3911), .D (
         window_4__4), .CLK (start), .R (rst)) ;
    nor03_2x ix1663 (.Y (nx1662), .A0 (gen_4_cmp_mReg_4), .A1 (nx10023), .A2 (
             nx10343)) ;
    nand02 ix1699 (.Y (gen_4_cmp_BSCmp_op2_5), .A0 (nx3915), .A1 (nx3921)) ;
    nor02_2x ix3916 (.Y (nx3915), .A0 (nx1694), .A1 (nx1690)) ;
    nor03_2x ix1695 (.Y (nx1694), .A0 (gen_4_cmp_mReg_4), .A1 (nx9645), .A2 (
             nx10311)) ;
    nor03_2x ix1691 (.Y (nx1690), .A0 (nx3911), .A1 (nx10317), .A2 (nx10327)) ;
    nor02_2x ix3922 (.Y (nx3921), .A0 (nx1686), .A1 (nx1684)) ;
    nor03_2x ix1687 (.Y (nx1686), .A0 (nx3925), .A1 (nx9641), .A2 (nx10335)) ;
    dffr gen_4_cmp_mRegCmp_reg_Q_5 (.Q (gen_4_cmp_mReg_5), .QB (nx3925), .D (
         window_4__5), .CLK (start), .R (rst)) ;
    nor03_2x ix1685 (.Y (nx1684), .A0 (gen_4_cmp_mReg_5), .A1 (nx10023), .A2 (
             nx10343)) ;
    nand02 ix1721 (.Y (gen_4_cmp_BSCmp_op2_6), .A0 (nx3930), .A1 (nx3935)) ;
    nor02_2x ix3931 (.Y (nx3930), .A0 (nx1716), .A1 (nx1712)) ;
    nor03_2x ix1717 (.Y (nx1716), .A0 (gen_4_cmp_mReg_5), .A1 (nx9647), .A2 (
             nx10311)) ;
    nor03_2x ix1713 (.Y (nx1712), .A0 (nx3925), .A1 (nx10317), .A2 (nx10327)) ;
    nor02_2x ix3936 (.Y (nx3935), .A0 (nx1708), .A1 (nx1706)) ;
    nor03_2x ix1709 (.Y (nx1708), .A0 (nx3939), .A1 (nx9641), .A2 (nx10335)) ;
    dffr gen_4_cmp_mRegCmp_reg_Q_6 (.Q (gen_4_cmp_mReg_6), .QB (nx3939), .D (
         window_4__6), .CLK (start), .R (rst)) ;
    nor03_2x ix1707 (.Y (nx1706), .A0 (gen_4_cmp_mReg_6), .A1 (nx10023), .A2 (
             nx10343)) ;
    nand02 ix1743 (.Y (gen_4_cmp_BSCmp_op2_7), .A0 (nx3945), .A1 (nx3951)) ;
    nor02_2x ix3946 (.Y (nx3945), .A0 (nx1738), .A1 (nx1734)) ;
    nor03_2x ix1739 (.Y (nx1738), .A0 (gen_4_cmp_mReg_6), .A1 (nx9647), .A2 (
             nx10313)) ;
    nor03_2x ix1735 (.Y (nx1734), .A0 (nx3939), .A1 (nx10319), .A2 (nx10329)) ;
    nor02_2x ix3952 (.Y (nx3951), .A0 (nx1730), .A1 (nx1728)) ;
    nor03_2x ix1731 (.Y (nx1730), .A0 (nx3954), .A1 (nx9641), .A2 (nx10337)) ;
    dffr gen_4_cmp_mRegCmp_reg_Q_7 (.Q (gen_4_cmp_mReg_7), .QB (nx3954), .D (
         window_4__7), .CLK (start), .R (rst)) ;
    nor03_2x ix1729 (.Y (nx1728), .A0 (gen_4_cmp_mReg_7), .A1 (nx10023), .A2 (
             nx10345)) ;
    nand02 ix1765 (.Y (gen_4_cmp_BSCmp_op2_8), .A0 (nx3961), .A1 (nx3967)) ;
    nor02_2x ix3962 (.Y (nx3961), .A0 (nx1760), .A1 (nx1756)) ;
    nor03_2x ix1761 (.Y (nx1760), .A0 (gen_4_cmp_mReg_7), .A1 (nx9647), .A2 (
             nx10313)) ;
    nor03_2x ix1757 (.Y (nx1756), .A0 (nx3954), .A1 (nx10319), .A2 (nx10329)) ;
    nor02_2x ix3968 (.Y (nx3967), .A0 (nx1752), .A1 (nx1750)) ;
    nor03_2x ix1753 (.Y (nx1752), .A0 (nx3971), .A1 (nx9641), .A2 (nx10337)) ;
    dffr gen_4_cmp_mRegCmp_reg_Q_8 (.Q (gen_4_cmp_mReg_8), .QB (nx3971), .D (
         window_4__8), .CLK (start), .R (rst)) ;
    nor03_2x ix1751 (.Y (nx1750), .A0 (gen_4_cmp_mReg_8), .A1 (nx10025), .A2 (
             nx10345)) ;
    nand02 ix1787 (.Y (gen_4_cmp_BSCmp_op2_9), .A0 (nx3975), .A1 (nx3981)) ;
    nor02_2x ix3976 (.Y (nx3975), .A0 (nx1782), .A1 (nx1778)) ;
    nor03_2x ix1783 (.Y (nx1782), .A0 (gen_4_cmp_mReg_8), .A1 (nx9647), .A2 (
             nx10313)) ;
    nor03_2x ix1779 (.Y (nx1778), .A0 (nx3971), .A1 (nx10319), .A2 (nx10329)) ;
    nor02_2x ix3982 (.Y (nx3981), .A0 (nx1774), .A1 (nx1772)) ;
    nor03_2x ix1775 (.Y (nx1774), .A0 (nx3985), .A1 (nx9641), .A2 (nx10337)) ;
    dffr gen_4_cmp_mRegCmp_reg_Q_9 (.Q (gen_4_cmp_mReg_9), .QB (nx3985), .D (
         window_4__9), .CLK (start), .R (rst)) ;
    nor03_2x ix1773 (.Y (nx1772), .A0 (gen_4_cmp_mReg_9), .A1 (nx10025), .A2 (
             nx10345)) ;
    nand02 ix1809 (.Y (gen_4_cmp_BSCmp_op2_10), .A0 (nx3989), .A1 (nx3995)) ;
    nor02_2x ix3990 (.Y (nx3989), .A0 (nx1804), .A1 (nx1800)) ;
    nor03_2x ix1805 (.Y (nx1804), .A0 (gen_4_cmp_mReg_9), .A1 (nx9647), .A2 (
             nx10313)) ;
    nor03_2x ix1801 (.Y (nx1800), .A0 (nx3985), .A1 (nx10319), .A2 (nx10329)) ;
    nor02_2x ix3996 (.Y (nx3995), .A0 (nx1796), .A1 (nx1794)) ;
    nor03_2x ix1797 (.Y (nx1796), .A0 (nx3998), .A1 (nx9641), .A2 (nx10337)) ;
    dffr gen_4_cmp_mRegCmp_reg_Q_10 (.Q (gen_4_cmp_mReg_10), .QB (nx3998), .D (
         window_4__10), .CLK (start), .R (rst)) ;
    nor03_2x ix1795 (.Y (nx1794), .A0 (gen_4_cmp_mReg_10), .A1 (nx10025), .A2 (
             nx10345)) ;
    nand02 ix1831 (.Y (gen_4_cmp_BSCmp_op2_11), .A0 (nx4005), .A1 (nx4011)) ;
    nor02_2x ix4006 (.Y (nx4005), .A0 (nx1826), .A1 (nx1822)) ;
    nor03_2x ix1827 (.Y (nx1826), .A0 (gen_4_cmp_mReg_10), .A1 (nx9647), .A2 (
             nx10313)) ;
    nor03_2x ix1823 (.Y (nx1822), .A0 (nx3998), .A1 (nx10319), .A2 (nx10329)) ;
    nor02_2x ix4012 (.Y (nx4011), .A0 (nx1818), .A1 (nx1816)) ;
    nor03_2x ix1819 (.Y (nx1818), .A0 (nx4015), .A1 (nx9641), .A2 (nx10337)) ;
    dffr gen_4_cmp_mRegCmp_reg_Q_11 (.Q (gen_4_cmp_mReg_11), .QB (nx4015), .D (
         window_4__11), .CLK (start), .R (rst)) ;
    nor03_2x ix1817 (.Y (nx1816), .A0 (gen_4_cmp_mReg_11), .A1 (nx10025), .A2 (
             nx10345)) ;
    nand02 ix1853 (.Y (gen_4_cmp_BSCmp_op2_12), .A0 (nx4019), .A1 (nx4025)) ;
    nor02_2x ix4020 (.Y (nx4019), .A0 (nx1848), .A1 (nx1844)) ;
    nor03_2x ix1849 (.Y (nx1848), .A0 (gen_4_cmp_mReg_11), .A1 (nx9647), .A2 (
             nx10313)) ;
    nor03_2x ix1845 (.Y (nx1844), .A0 (nx4015), .A1 (nx10319), .A2 (nx10329)) ;
    nor02_2x ix4026 (.Y (nx4025), .A0 (nx1840), .A1 (nx1838)) ;
    nor03_2x ix1841 (.Y (nx1840), .A0 (nx4029), .A1 (nx9643), .A2 (nx10337)) ;
    dffr gen_4_cmp_mRegCmp_reg_Q_12 (.Q (gen_4_cmp_mReg_12), .QB (nx4029), .D (
         window_4__12), .CLK (start), .R (rst)) ;
    nor03_2x ix1839 (.Y (nx1838), .A0 (gen_4_cmp_mReg_12), .A1 (nx10025), .A2 (
             nx10345)) ;
    nand02 ix1875 (.Y (gen_4_cmp_BSCmp_op2_13), .A0 (nx4033), .A1 (nx4039)) ;
    nor02_2x ix4034 (.Y (nx4033), .A0 (nx1870), .A1 (nx1866)) ;
    nor03_2x ix1871 (.Y (nx1870), .A0 (gen_4_cmp_mReg_12), .A1 (nx9649), .A2 (
             nx10315)) ;
    nor03_2x ix1867 (.Y (nx1866), .A0 (nx4029), .A1 (nx10319), .A2 (nx10331)) ;
    nor02_2x ix4040 (.Y (nx4039), .A0 (nx1862), .A1 (nx1860)) ;
    nor03_2x ix1863 (.Y (nx1862), .A0 (nx4042), .A1 (nx9643), .A2 (nx10339)) ;
    dffr gen_4_cmp_mRegCmp_reg_Q_13 (.Q (gen_4_cmp_mReg_13), .QB (nx4042), .D (
         window_4__13), .CLK (start), .R (rst)) ;
    nor03_2x ix1861 (.Y (nx1860), .A0 (gen_4_cmp_mReg_13), .A1 (nx10025), .A2 (
             nx10347)) ;
    nand02 ix1897 (.Y (gen_4_cmp_BSCmp_op2_14), .A0 (nx4049), .A1 (nx4055)) ;
    nor02_2x ix4050 (.Y (nx4049), .A0 (nx1892), .A1 (nx1888)) ;
    nor03_2x ix1893 (.Y (nx1892), .A0 (gen_4_cmp_mReg_13), .A1 (nx9649), .A2 (
             nx10315)) ;
    nor03_2x ix1889 (.Y (nx1888), .A0 (nx4042), .A1 (nx10321), .A2 (nx10331)) ;
    nor02_2x ix4056 (.Y (nx4055), .A0 (nx1884), .A1 (nx1882)) ;
    nor03_2x ix1885 (.Y (nx1884), .A0 (nx4059), .A1 (nx9643), .A2 (nx10339)) ;
    dffr gen_4_cmp_mRegCmp_reg_Q_14 (.Q (gen_4_cmp_mReg_14), .QB (nx4059), .D (
         window_4__14), .CLK (start), .R (rst)) ;
    nor03_2x ix1883 (.Y (nx1882), .A0 (gen_4_cmp_mReg_14), .A1 (nx10025), .A2 (
             nx10347)) ;
    nand02 ix1919 (.Y (gen_4_cmp_BSCmp_op2_15), .A0 (nx4063), .A1 (nx4069)) ;
    nor02_2x ix4064 (.Y (nx4063), .A0 (nx1914), .A1 (nx1910)) ;
    nor03_2x ix1915 (.Y (nx1914), .A0 (gen_4_cmp_mReg_14), .A1 (nx9649), .A2 (
             nx10315)) ;
    nor03_2x ix1911 (.Y (nx1910), .A0 (nx4059), .A1 (nx10321), .A2 (nx10331)) ;
    nor02_2x ix4070 (.Y (nx4069), .A0 (nx1906), .A1 (nx1904)) ;
    nor03_2x ix1907 (.Y (nx1906), .A0 (nx4073), .A1 (nx9643), .A2 (nx10339)) ;
    dffr gen_4_cmp_mRegCmp_reg_Q_15 (.Q (gen_4_cmp_mReg_15), .QB (nx4073), .D (
         window_4__15), .CLK (start), .R (rst)) ;
    nor03_2x ix1905 (.Y (nx1904), .A0 (gen_4_cmp_mReg_15), .A1 (nx10027), .A2 (
             nx10347)) ;
    nand02 ix1929 (.Y (gen_4_cmp_BSCmp_op2_16), .A0 (nx4077), .A1 (nx4069)) ;
    nor02_2x ix4078 (.Y (nx4077), .A0 (nx1924), .A1 (nx1920)) ;
    nor03_2x ix1925 (.Y (nx1924), .A0 (gen_4_cmp_mReg_15), .A1 (nx9649), .A2 (
             nx10315)) ;
    nor03_2x ix1921 (.Y (nx1920), .A0 (nx4073), .A1 (nx10321), .A2 (nx10331)) ;
    nand02 ix1997 (.Y (gen_5_cmp_BSCmp_op2_1), .A0 (nx4084), .A1 (nx4103)) ;
    nor02_2x ix4085 (.Y (nx4084), .A0 (nx1992), .A1 (nx1988)) ;
    nor03_2x ix1993 (.Y (nx1992), .A0 (gen_5_cmp_mReg_0), .A1 (nx9633), .A2 (
             nx10351)) ;
    dffr gen_5_cmp_mRegCmp_reg_Q_0 (.Q (gen_5_cmp_mReg_0), .QB (nx4089), .D (
         window_5__0), .CLK (start), .R (rst)) ;
    inv01 ix4094 (.Y (nx4093), .A (gen_5_cmp_pMux_0)) ;
    nor03_2x ix1989 (.Y (nx1988), .A0 (nx4089), .A1 (nx10357), .A2 (nx10367)) ;
    inv02 ix4102 (.Y (nx4101), .A (gen_5_cmp_pMux_2)) ;
    nor02_2x ix4104 (.Y (nx4103), .A0 (nx1978), .A1 (nx1976)) ;
    nor03_2x ix1979 (.Y (nx1978), .A0 (nx4106), .A1 (nx9627), .A2 (nx10375)) ;
    dffr gen_5_cmp_mRegCmp_reg_Q_1 (.Q (gen_5_cmp_mReg_1), .QB (nx4106), .D (
         window_5__1), .CLK (start), .R (rst)) ;
    nor03_2x ix1977 (.Y (nx1976), .A0 (gen_5_cmp_mReg_1), .A1 (nx10029), .A2 (
             nx10383)) ;
    nor03_2x ix1937 (.Y (nx1936), .A0 (nx9633), .A1 (nx4101), .A2 (
             gen_5_cmp_pMux_0)) ;
    nand02 ix2019 (.Y (gen_5_cmp_BSCmp_op2_2), .A0 (nx4119), .A1 (nx4125)) ;
    nor02_2x ix4120 (.Y (nx4119), .A0 (nx2014), .A1 (nx2010)) ;
    nor03_2x ix2015 (.Y (nx2014), .A0 (gen_5_cmp_mReg_1), .A1 (nx9633), .A2 (
             nx10351)) ;
    nor03_2x ix2011 (.Y (nx2010), .A0 (nx4106), .A1 (nx10357), .A2 (nx10367)) ;
    nor02_2x ix4126 (.Y (nx4125), .A0 (nx2006), .A1 (nx2004)) ;
    nor03_2x ix2007 (.Y (nx2006), .A0 (nx4128), .A1 (nx9627), .A2 (nx10375)) ;
    dffr gen_5_cmp_mRegCmp_reg_Q_2 (.Q (gen_5_cmp_mReg_2), .QB (nx4128), .D (
         window_5__2), .CLK (start), .R (rst)) ;
    nor03_2x ix2005 (.Y (nx2004), .A0 (gen_5_cmp_mReg_2), .A1 (nx10029), .A2 (
             nx10383)) ;
    nand02 ix2041 (.Y (gen_5_cmp_BSCmp_op2_3), .A0 (nx4133), .A1 (nx4139)) ;
    nor02_2x ix4134 (.Y (nx4133), .A0 (nx2036), .A1 (nx2032)) ;
    nor03_2x ix2037 (.Y (nx2036), .A0 (gen_5_cmp_mReg_2), .A1 (nx9633), .A2 (
             nx10351)) ;
    nor03_2x ix2033 (.Y (nx2032), .A0 (nx4128), .A1 (nx10357), .A2 (nx10367)) ;
    nor02_2x ix4140 (.Y (nx4139), .A0 (nx2028), .A1 (nx2026)) ;
    nor03_2x ix2029 (.Y (nx2028), .A0 (nx4143), .A1 (nx9627), .A2 (nx10375)) ;
    dffr gen_5_cmp_mRegCmp_reg_Q_3 (.Q (gen_5_cmp_mReg_3), .QB (nx4143), .D (
         window_5__3), .CLK (start), .R (rst)) ;
    nor03_2x ix2027 (.Y (nx2026), .A0 (gen_5_cmp_mReg_3), .A1 (nx10029), .A2 (
             nx10383)) ;
    nand02 ix2063 (.Y (gen_5_cmp_BSCmp_op2_4), .A0 (nx4149), .A1 (nx4153)) ;
    nor02_2x ix4150 (.Y (nx4149), .A0 (nx2058), .A1 (nx2054)) ;
    nor03_2x ix2059 (.Y (nx2058), .A0 (gen_5_cmp_mReg_3), .A1 (nx9633), .A2 (
             nx10351)) ;
    nor03_2x ix2055 (.Y (nx2054), .A0 (nx4143), .A1 (nx10357), .A2 (nx10367)) ;
    nor02_2x ix4154 (.Y (nx4153), .A0 (nx2050), .A1 (nx2048)) ;
    nor03_2x ix2051 (.Y (nx2050), .A0 (nx4157), .A1 (nx9627), .A2 (nx10375)) ;
    dffr gen_5_cmp_mRegCmp_reg_Q_4 (.Q (gen_5_cmp_mReg_4), .QB (nx4157), .D (
         window_5__4), .CLK (start), .R (rst)) ;
    nor03_2x ix2049 (.Y (nx2048), .A0 (gen_5_cmp_mReg_4), .A1 (nx10029), .A2 (
             nx10383)) ;
    nand02 ix2085 (.Y (gen_5_cmp_BSCmp_op2_5), .A0 (nx4163), .A1 (nx4169)) ;
    nor02_2x ix4164 (.Y (nx4163), .A0 (nx2080), .A1 (nx2076)) ;
    nor03_2x ix2081 (.Y (nx2080), .A0 (gen_5_cmp_mReg_4), .A1 (nx9633), .A2 (
             nx10351)) ;
    nor03_2x ix2077 (.Y (nx2076), .A0 (nx4157), .A1 (nx10357), .A2 (nx10367)) ;
    nor02_2x ix4170 (.Y (nx4169), .A0 (nx2072), .A1 (nx2070)) ;
    nor03_2x ix2073 (.Y (nx2072), .A0 (nx4172), .A1 (nx9629), .A2 (nx10375)) ;
    dffr gen_5_cmp_mRegCmp_reg_Q_5 (.Q (gen_5_cmp_mReg_5), .QB (nx4172), .D (
         window_5__5), .CLK (start), .R (rst)) ;
    nor03_2x ix2071 (.Y (nx2070), .A0 (gen_5_cmp_mReg_5), .A1 (nx10029), .A2 (
             nx10383)) ;
    nand02 ix2107 (.Y (gen_5_cmp_BSCmp_op2_6), .A0 (nx4177), .A1 (nx4183)) ;
    nor02_2x ix4178 (.Y (nx4177), .A0 (nx2102), .A1 (nx2098)) ;
    nor03_2x ix2103 (.Y (nx2102), .A0 (gen_5_cmp_mReg_5), .A1 (nx9635), .A2 (
             nx10351)) ;
    nor03_2x ix2099 (.Y (nx2098), .A0 (nx4172), .A1 (nx10357), .A2 (nx10367)) ;
    nor02_2x ix4184 (.Y (nx4183), .A0 (nx2094), .A1 (nx2092)) ;
    nor03_2x ix2095 (.Y (nx2094), .A0 (nx4187), .A1 (nx9629), .A2 (nx10375)) ;
    dffr gen_5_cmp_mRegCmp_reg_Q_6 (.Q (gen_5_cmp_mReg_6), .QB (nx4187), .D (
         window_5__6), .CLK (start), .R (rst)) ;
    nor03_2x ix2093 (.Y (nx2092), .A0 (gen_5_cmp_mReg_6), .A1 (nx10029), .A2 (
             nx10383)) ;
    nand02 ix2129 (.Y (gen_5_cmp_BSCmp_op2_7), .A0 (nx4193), .A1 (nx4197)) ;
    nor02_2x ix4194 (.Y (nx4193), .A0 (nx2124), .A1 (nx2120)) ;
    nor03_2x ix2125 (.Y (nx2124), .A0 (gen_5_cmp_mReg_6), .A1 (nx9635), .A2 (
             nx10353)) ;
    nor03_2x ix2121 (.Y (nx2120), .A0 (nx4187), .A1 (nx10359), .A2 (nx10369)) ;
    nor02_2x ix4198 (.Y (nx4197), .A0 (nx2116), .A1 (nx2114)) ;
    nor03_2x ix2117 (.Y (nx2116), .A0 (nx4201), .A1 (nx9629), .A2 (nx10377)) ;
    dffr gen_5_cmp_mRegCmp_reg_Q_7 (.Q (gen_5_cmp_mReg_7), .QB (nx4201), .D (
         window_5__7), .CLK (start), .R (rst)) ;
    nor03_2x ix2115 (.Y (nx2114), .A0 (gen_5_cmp_mReg_7), .A1 (nx10029), .A2 (
             nx10385)) ;
    nand02 ix2151 (.Y (gen_5_cmp_BSCmp_op2_8), .A0 (nx4207), .A1 (nx4213)) ;
    nor02_2x ix4208 (.Y (nx4207), .A0 (nx2146), .A1 (nx2142)) ;
    nor03_2x ix2147 (.Y (nx2146), .A0 (gen_5_cmp_mReg_7), .A1 (nx9635), .A2 (
             nx10353)) ;
    nor03_2x ix2143 (.Y (nx2142), .A0 (nx4201), .A1 (nx10359), .A2 (nx10369)) ;
    nor02_2x ix4214 (.Y (nx4213), .A0 (nx2138), .A1 (nx2136)) ;
    nor03_2x ix2139 (.Y (nx2138), .A0 (nx4216), .A1 (nx9629), .A2 (nx10377)) ;
    dffr gen_5_cmp_mRegCmp_reg_Q_8 (.Q (gen_5_cmp_mReg_8), .QB (nx4216), .D (
         window_5__8), .CLK (start), .R (rst)) ;
    nor03_2x ix2137 (.Y (nx2136), .A0 (gen_5_cmp_mReg_8), .A1 (nx10031), .A2 (
             nx10385)) ;
    nand02 ix2173 (.Y (gen_5_cmp_BSCmp_op2_9), .A0 (nx4221), .A1 (nx4227)) ;
    nor02_2x ix4222 (.Y (nx4221), .A0 (nx2168), .A1 (nx2164)) ;
    nor03_2x ix2169 (.Y (nx2168), .A0 (gen_5_cmp_mReg_8), .A1 (nx9635), .A2 (
             nx10353)) ;
    nor03_2x ix2165 (.Y (nx2164), .A0 (nx4216), .A1 (nx10359), .A2 (nx10369)) ;
    nor02_2x ix4228 (.Y (nx4227), .A0 (nx2160), .A1 (nx2158)) ;
    nor03_2x ix2161 (.Y (nx2160), .A0 (nx4231), .A1 (nx9629), .A2 (nx10377)) ;
    dffr gen_5_cmp_mRegCmp_reg_Q_9 (.Q (gen_5_cmp_mReg_9), .QB (nx4231), .D (
         window_5__9), .CLK (start), .R (rst)) ;
    nor03_2x ix2159 (.Y (nx2158), .A0 (gen_5_cmp_mReg_9), .A1 (nx10031), .A2 (
             nx10385)) ;
    nand02 ix2195 (.Y (gen_5_cmp_BSCmp_op2_10), .A0 (nx4237), .A1 (nx4241)) ;
    nor02_2x ix4238 (.Y (nx4237), .A0 (nx2190), .A1 (nx2186)) ;
    nor03_2x ix2191 (.Y (nx2190), .A0 (gen_5_cmp_mReg_9), .A1 (nx9635), .A2 (
             nx10353)) ;
    nor03_2x ix2187 (.Y (nx2186), .A0 (nx4231), .A1 (nx10359), .A2 (nx10369)) ;
    nor02_2x ix4242 (.Y (nx4241), .A0 (nx2182), .A1 (nx2180)) ;
    nor03_2x ix2183 (.Y (nx2182), .A0 (nx4245), .A1 (nx9629), .A2 (nx10377)) ;
    dffr gen_5_cmp_mRegCmp_reg_Q_10 (.Q (gen_5_cmp_mReg_10), .QB (nx4245), .D (
         window_5__10), .CLK (start), .R (rst)) ;
    nor03_2x ix2181 (.Y (nx2180), .A0 (gen_5_cmp_mReg_10), .A1 (nx10031), .A2 (
             nx10385)) ;
    nand02 ix2217 (.Y (gen_5_cmp_BSCmp_op2_11), .A0 (nx4251), .A1 (nx4256)) ;
    nor02_2x ix4252 (.Y (nx4251), .A0 (nx2212), .A1 (nx2208)) ;
    nor03_2x ix2213 (.Y (nx2212), .A0 (gen_5_cmp_mReg_10), .A1 (nx9635), .A2 (
             nx10353)) ;
    nor03_2x ix2209 (.Y (nx2208), .A0 (nx4245), .A1 (nx10359), .A2 (nx10369)) ;
    nor02_2x ix4257 (.Y (nx4256), .A0 (nx2204), .A1 (nx2202)) ;
    nor03_2x ix2205 (.Y (nx2204), .A0 (nx4259), .A1 (nx9629), .A2 (nx10377)) ;
    dffr gen_5_cmp_mRegCmp_reg_Q_11 (.Q (gen_5_cmp_mReg_11), .QB (nx4259), .D (
         window_5__11), .CLK (start), .R (rst)) ;
    nor03_2x ix2203 (.Y (nx2202), .A0 (gen_5_cmp_mReg_11), .A1 (nx10031), .A2 (
             nx10385)) ;
    nand02 ix2239 (.Y (gen_5_cmp_BSCmp_op2_12), .A0 (nx4263), .A1 (nx4269)) ;
    nor02_2x ix4264 (.Y (nx4263), .A0 (nx2234), .A1 (nx2230)) ;
    nor03_2x ix2235 (.Y (nx2234), .A0 (gen_5_cmp_mReg_11), .A1 (nx9635), .A2 (
             nx10353)) ;
    nor03_2x ix2231 (.Y (nx2230), .A0 (nx4259), .A1 (nx10359), .A2 (nx10369)) ;
    nor02_2x ix4270 (.Y (nx4269), .A0 (nx2226), .A1 (nx2224)) ;
    nor03_2x ix2227 (.Y (nx2226), .A0 (nx4273), .A1 (nx9631), .A2 (nx10377)) ;
    dffr gen_5_cmp_mRegCmp_reg_Q_12 (.Q (gen_5_cmp_mReg_12), .QB (nx4273), .D (
         window_5__12), .CLK (start), .R (rst)) ;
    nor03_2x ix2225 (.Y (nx2224), .A0 (gen_5_cmp_mReg_12), .A1 (nx10031), .A2 (
             nx10385)) ;
    nand02 ix2261 (.Y (gen_5_cmp_BSCmp_op2_13), .A0 (nx4279), .A1 (nx4285)) ;
    nor02_2x ix4280 (.Y (nx4279), .A0 (nx2256), .A1 (nx2252)) ;
    nor03_2x ix2257 (.Y (nx2256), .A0 (gen_5_cmp_mReg_12), .A1 (nx9637), .A2 (
             nx10355)) ;
    nor03_2x ix2253 (.Y (nx2252), .A0 (nx4273), .A1 (nx10359), .A2 (nx10371)) ;
    nor02_2x ix4286 (.Y (nx4285), .A0 (nx2248), .A1 (nx2246)) ;
    nor03_2x ix2249 (.Y (nx2248), .A0 (nx4288), .A1 (nx9631), .A2 (nx10379)) ;
    dffr gen_5_cmp_mRegCmp_reg_Q_13 (.Q (gen_5_cmp_mReg_13), .QB (nx4288), .D (
         window_5__13), .CLK (start), .R (rst)) ;
    nor03_2x ix2247 (.Y (nx2246), .A0 (gen_5_cmp_mReg_13), .A1 (nx10031), .A2 (
             nx10387)) ;
    nand02 ix2283 (.Y (gen_5_cmp_BSCmp_op2_14), .A0 (nx4293), .A1 (nx4299)) ;
    nor02_2x ix4294 (.Y (nx4293), .A0 (nx2278), .A1 (nx2274)) ;
    nor03_2x ix2279 (.Y (nx2278), .A0 (gen_5_cmp_mReg_13), .A1 (nx9637), .A2 (
             nx10355)) ;
    nor03_2x ix2275 (.Y (nx2274), .A0 (nx4288), .A1 (nx10361), .A2 (nx10371)) ;
    nor02_2x ix4300 (.Y (nx4299), .A0 (nx2270), .A1 (nx2268)) ;
    nor03_2x ix2271 (.Y (nx2270), .A0 (nx4303), .A1 (nx9631), .A2 (nx10379)) ;
    dffr gen_5_cmp_mRegCmp_reg_Q_14 (.Q (gen_5_cmp_mReg_14), .QB (nx4303), .D (
         window_5__14), .CLK (start), .R (rst)) ;
    nor03_2x ix2269 (.Y (nx2268), .A0 (gen_5_cmp_mReg_14), .A1 (nx10031), .A2 (
             nx10387)) ;
    nand02 ix2305 (.Y (gen_5_cmp_BSCmp_op2_15), .A0 (nx4309), .A1 (nx4315)) ;
    nor02_2x ix4310 (.Y (nx4309), .A0 (nx2300), .A1 (nx2296)) ;
    nor03_2x ix2301 (.Y (nx2300), .A0 (gen_5_cmp_mReg_14), .A1 (nx9637), .A2 (
             nx10355)) ;
    nor03_2x ix2297 (.Y (nx2296), .A0 (nx4303), .A1 (nx10361), .A2 (nx10371)) ;
    nor02_2x ix4316 (.Y (nx4315), .A0 (nx2292), .A1 (nx2290)) ;
    nor03_2x ix2293 (.Y (nx2292), .A0 (nx4318), .A1 (nx9631), .A2 (nx10379)) ;
    dffr gen_5_cmp_mRegCmp_reg_Q_15 (.Q (gen_5_cmp_mReg_15), .QB (nx4318), .D (
         window_5__15), .CLK (start), .R (rst)) ;
    nor03_2x ix2291 (.Y (nx2290), .A0 (gen_5_cmp_mReg_15), .A1 (nx10033), .A2 (
             nx10387)) ;
    nand02 ix2315 (.Y (gen_5_cmp_BSCmp_op2_16), .A0 (nx4325), .A1 (nx4315)) ;
    nor02_2x ix4326 (.Y (nx4325), .A0 (nx2310), .A1 (nx2306)) ;
    nor03_2x ix2311 (.Y (nx2310), .A0 (gen_5_cmp_mReg_15), .A1 (nx9637), .A2 (
             nx10355)) ;
    nor03_2x ix2307 (.Y (nx2306), .A0 (nx4318), .A1 (nx10361), .A2 (nx10371)) ;
    nand02 ix2383 (.Y (gen_6_cmp_BSCmp_op2_1), .A0 (nx4331), .A1 (nx4351)) ;
    nor02_2x ix4332 (.Y (nx4331), .A0 (nx2378), .A1 (nx2374)) ;
    nor03_2x ix2379 (.Y (nx2378), .A0 (gen_6_cmp_mReg_0), .A1 (nx9621), .A2 (
             nx10391)) ;
    dffr gen_6_cmp_mRegCmp_reg_Q_0 (.Q (gen_6_cmp_mReg_0), .QB (nx4337), .D (
         window_6__0), .CLK (start), .R (rst)) ;
    inv01 ix4342 (.Y (nx4340), .A (gen_6_cmp_pMux_0)) ;
    nor03_2x ix2375 (.Y (nx2374), .A0 (nx4337), .A1 (nx10397), .A2 (nx10407)) ;
    inv02 ix4350 (.Y (nx4349), .A (gen_6_cmp_pMux_2)) ;
    nor02_2x ix4352 (.Y (nx4351), .A0 (nx2364), .A1 (nx2362)) ;
    nor03_2x ix2365 (.Y (nx2364), .A0 (nx4355), .A1 (nx9615), .A2 (nx10415)) ;
    dffr gen_6_cmp_mRegCmp_reg_Q_1 (.Q (gen_6_cmp_mReg_1), .QB (nx4355), .D (
         window_6__1), .CLK (start), .R (rst)) ;
    nor03_2x ix2363 (.Y (nx2362), .A0 (gen_6_cmp_mReg_1), .A1 (nx10035), .A2 (
             nx10423)) ;
    nor03_2x ix2326 (.Y (nx2322), .A0 (nx9621), .A1 (nx4349), .A2 (
             gen_6_cmp_pMux_0)) ;
    nand02 ix2405 (.Y (gen_6_cmp_BSCmp_op2_2), .A0 (nx4365), .A1 (nx4371)) ;
    nor02_2x ix4366 (.Y (nx4365), .A0 (nx2400), .A1 (nx2396)) ;
    nor03_2x ix2401 (.Y (nx2400), .A0 (gen_6_cmp_mReg_1), .A1 (nx9621), .A2 (
             nx10391)) ;
    nor03_2x ix2397 (.Y (nx2396), .A0 (nx4355), .A1 (nx10397), .A2 (nx10407)) ;
    nor02_2x ix4372 (.Y (nx4371), .A0 (nx2392), .A1 (nx2390)) ;
    nor03_2x ix2393 (.Y (nx2392), .A0 (nx4375), .A1 (nx9615), .A2 (nx10415)) ;
    dffr gen_6_cmp_mRegCmp_reg_Q_2 (.Q (gen_6_cmp_mReg_2), .QB (nx4375), .D (
         window_6__2), .CLK (start), .R (rst)) ;
    nor03_2x ix2391 (.Y (nx2390), .A0 (gen_6_cmp_mReg_2), .A1 (nx10035), .A2 (
             nx10423)) ;
    nand02 ix2427 (.Y (gen_6_cmp_BSCmp_op2_3), .A0 (nx4381), .A1 (nx4385)) ;
    nor02_2x ix4382 (.Y (nx4381), .A0 (nx2422), .A1 (nx2418)) ;
    nor03_2x ix2423 (.Y (nx2422), .A0 (gen_6_cmp_mReg_2), .A1 (nx9621), .A2 (
             nx10391)) ;
    nor03_2x ix2419 (.Y (nx2418), .A0 (nx4375), .A1 (nx10397), .A2 (nx10407)) ;
    nor02_2x ix4386 (.Y (nx4385), .A0 (nx2414), .A1 (nx2412)) ;
    nor03_2x ix2415 (.Y (nx2414), .A0 (nx4389), .A1 (nx9615), .A2 (nx10415)) ;
    dffr gen_6_cmp_mRegCmp_reg_Q_3 (.Q (gen_6_cmp_mReg_3), .QB (nx4389), .D (
         window_6__3), .CLK (start), .R (rst)) ;
    nor03_2x ix2413 (.Y (nx2412), .A0 (gen_6_cmp_mReg_3), .A1 (nx10035), .A2 (
             nx10423)) ;
    nand02 ix2449 (.Y (gen_6_cmp_BSCmp_op2_4), .A0 (nx4395), .A1 (nx4401)) ;
    nor02_2x ix4396 (.Y (nx4395), .A0 (nx2444), .A1 (nx2440)) ;
    nor03_2x ix2445 (.Y (nx2444), .A0 (gen_6_cmp_mReg_3), .A1 (nx9621), .A2 (
             nx10391)) ;
    nor03_2x ix2441 (.Y (nx2440), .A0 (nx4389), .A1 (nx10397), .A2 (nx10407)) ;
    nor02_2x ix4402 (.Y (nx4401), .A0 (nx2436), .A1 (nx2434)) ;
    nor03_2x ix2437 (.Y (nx2436), .A0 (nx4404), .A1 (nx9615), .A2 (nx10415)) ;
    dffr gen_6_cmp_mRegCmp_reg_Q_4 (.Q (gen_6_cmp_mReg_4), .QB (nx4404), .D (
         window_6__4), .CLK (start), .R (rst)) ;
    nor03_2x ix2435 (.Y (nx2434), .A0 (gen_6_cmp_mReg_4), .A1 (nx10035), .A2 (
             nx10423)) ;
    nand02 ix2471 (.Y (gen_6_cmp_BSCmp_op2_5), .A0 (nx4409), .A1 (nx4415)) ;
    nor02_2x ix4410 (.Y (nx4409), .A0 (nx2466), .A1 (nx2462)) ;
    nor03_2x ix2467 (.Y (nx2466), .A0 (gen_6_cmp_mReg_4), .A1 (nx9621), .A2 (
             nx10391)) ;
    nor03_2x ix2463 (.Y (nx2462), .A0 (nx4404), .A1 (nx10397), .A2 (nx10407)) ;
    nor02_2x ix4416 (.Y (nx4415), .A0 (nx2458), .A1 (nx2456)) ;
    nor03_2x ix2459 (.Y (nx2458), .A0 (nx4419), .A1 (nx9617), .A2 (nx10415)) ;
    dffr gen_6_cmp_mRegCmp_reg_Q_5 (.Q (gen_6_cmp_mReg_5), .QB (nx4419), .D (
         window_6__5), .CLK (start), .R (rst)) ;
    nor03_2x ix2457 (.Y (nx2456), .A0 (gen_6_cmp_mReg_5), .A1 (nx10035), .A2 (
             nx10423)) ;
    nand02 ix2493 (.Y (gen_6_cmp_BSCmp_op2_6), .A0 (nx4425), .A1 (nx4429)) ;
    nor02_2x ix4426 (.Y (nx4425), .A0 (nx2488), .A1 (nx2484)) ;
    nor03_2x ix2489 (.Y (nx2488), .A0 (gen_6_cmp_mReg_5), .A1 (nx9623), .A2 (
             nx10391)) ;
    nor03_2x ix2485 (.Y (nx2484), .A0 (nx4419), .A1 (nx10397), .A2 (nx10407)) ;
    nor02_2x ix4430 (.Y (nx4429), .A0 (nx2480), .A1 (nx2478)) ;
    nor03_2x ix2481 (.Y (nx2480), .A0 (nx4433), .A1 (nx9617), .A2 (nx10415)) ;
    dffr gen_6_cmp_mRegCmp_reg_Q_6 (.Q (gen_6_cmp_mReg_6), .QB (nx4433), .D (
         window_6__6), .CLK (start), .R (rst)) ;
    nor03_2x ix2479 (.Y (nx2478), .A0 (gen_6_cmp_mReg_6), .A1 (nx10035), .A2 (
             nx10423)) ;
    nand02 ix2515 (.Y (gen_6_cmp_BSCmp_op2_7), .A0 (nx4439), .A1 (nx4445)) ;
    nor02_2x ix4440 (.Y (nx4439), .A0 (nx2510), .A1 (nx2506)) ;
    nor03_2x ix2511 (.Y (nx2510), .A0 (gen_6_cmp_mReg_6), .A1 (nx9623), .A2 (
             nx10393)) ;
    nor03_2x ix2507 (.Y (nx2506), .A0 (nx4433), .A1 (nx10399), .A2 (nx10409)) ;
    nor02_2x ix4446 (.Y (nx4445), .A0 (nx2502), .A1 (nx2500)) ;
    nor03_2x ix2503 (.Y (nx2502), .A0 (nx4448), .A1 (nx9617), .A2 (nx10417)) ;
    dffr gen_6_cmp_mRegCmp_reg_Q_7 (.Q (gen_6_cmp_mReg_7), .QB (nx4448), .D (
         window_6__7), .CLK (start), .R (rst)) ;
    nor03_2x ix2501 (.Y (nx2500), .A0 (gen_6_cmp_mReg_7), .A1 (nx10035), .A2 (
             nx10425)) ;
    nand02 ix2537 (.Y (gen_6_cmp_BSCmp_op2_8), .A0 (nx4453), .A1 (nx4459)) ;
    nor02_2x ix4454 (.Y (nx4453), .A0 (nx2532), .A1 (nx2528)) ;
    nor03_2x ix2533 (.Y (nx2532), .A0 (gen_6_cmp_mReg_7), .A1 (nx9623), .A2 (
             nx10393)) ;
    nor03_2x ix2529 (.Y (nx2528), .A0 (nx4448), .A1 (nx10399), .A2 (nx10409)) ;
    nor02_2x ix4460 (.Y (nx4459), .A0 (nx2524), .A1 (nx2522)) ;
    nor03_2x ix2525 (.Y (nx2524), .A0 (nx4463), .A1 (nx9617), .A2 (nx10417)) ;
    dffr gen_6_cmp_mRegCmp_reg_Q_8 (.Q (gen_6_cmp_mReg_8), .QB (nx4463), .D (
         window_6__8), .CLK (start), .R (rst)) ;
    nor03_2x ix2523 (.Y (nx2522), .A0 (gen_6_cmp_mReg_8), .A1 (nx10037), .A2 (
             nx10425)) ;
    nand02 ix2559 (.Y (gen_6_cmp_BSCmp_op2_9), .A0 (nx4469), .A1 (nx4473)) ;
    nor02_2x ix4470 (.Y (nx4469), .A0 (nx2554), .A1 (nx2550)) ;
    nor03_2x ix2555 (.Y (nx2554), .A0 (gen_6_cmp_mReg_8), .A1 (nx9623), .A2 (
             nx10393)) ;
    nor03_2x ix2551 (.Y (nx2550), .A0 (nx4463), .A1 (nx10399), .A2 (nx10409)) ;
    nor02_2x ix4474 (.Y (nx4473), .A0 (nx2546), .A1 (nx2544)) ;
    nor03_2x ix2547 (.Y (nx2546), .A0 (nx4477), .A1 (nx9617), .A2 (nx10417)) ;
    dffr gen_6_cmp_mRegCmp_reg_Q_9 (.Q (gen_6_cmp_mReg_9), .QB (nx4477), .D (
         window_6__9), .CLK (start), .R (rst)) ;
    nor03_2x ix2545 (.Y (nx2544), .A0 (gen_6_cmp_mReg_9), .A1 (nx10037), .A2 (
             nx10425)) ;
    nand02 ix2581 (.Y (gen_6_cmp_BSCmp_op2_10), .A0 (nx4483), .A1 (nx4489)) ;
    nor02_2x ix4484 (.Y (nx4483), .A0 (nx2576), .A1 (nx2572)) ;
    nor03_2x ix2577 (.Y (nx2576), .A0 (gen_6_cmp_mReg_9), .A1 (nx9623), .A2 (
             nx10393)) ;
    nor03_2x ix2573 (.Y (nx2572), .A0 (nx4477), .A1 (nx10399), .A2 (nx10409)) ;
    nor02_2x ix4490 (.Y (nx4489), .A0 (nx2568), .A1 (nx2566)) ;
    nor03_2x ix2569 (.Y (nx2568), .A0 (nx4492), .A1 (nx9617), .A2 (nx10417)) ;
    dffr gen_6_cmp_mRegCmp_reg_Q_10 (.Q (gen_6_cmp_mReg_10), .QB (nx4492), .D (
         window_6__10), .CLK (start), .R (rst)) ;
    nor03_2x ix2567 (.Y (nx2566), .A0 (gen_6_cmp_mReg_10), .A1 (nx10037), .A2 (
             nx10425)) ;
    nand02 ix2603 (.Y (gen_6_cmp_BSCmp_op2_11), .A0 (nx4497), .A1 (nx4503)) ;
    nor02_2x ix4498 (.Y (nx4497), .A0 (nx2598), .A1 (nx2594)) ;
    nor03_2x ix2599 (.Y (nx2598), .A0 (gen_6_cmp_mReg_10), .A1 (nx9623), .A2 (
             nx10393)) ;
    nor03_2x ix2595 (.Y (nx2594), .A0 (nx4492), .A1 (nx10399), .A2 (nx10409)) ;
    nor02_2x ix4504 (.Y (nx4503), .A0 (nx2590), .A1 (nx2588)) ;
    nor03_2x ix2591 (.Y (nx2590), .A0 (nx4507), .A1 (nx9617), .A2 (nx10417)) ;
    dffr gen_6_cmp_mRegCmp_reg_Q_11 (.Q (gen_6_cmp_mReg_11), .QB (nx4507), .D (
         window_6__11), .CLK (start), .R (rst)) ;
    nor03_2x ix2589 (.Y (nx2588), .A0 (gen_6_cmp_mReg_11), .A1 (nx10037), .A2 (
             nx10425)) ;
    nand02 ix2625 (.Y (gen_6_cmp_BSCmp_op2_12), .A0 (nx4513), .A1 (nx4517)) ;
    nor02_2x ix4514 (.Y (nx4513), .A0 (nx2620), .A1 (nx2616)) ;
    nor03_2x ix2621 (.Y (nx2620), .A0 (gen_6_cmp_mReg_11), .A1 (nx9623), .A2 (
             nx10393)) ;
    nor03_2x ix2617 (.Y (nx2616), .A0 (nx4507), .A1 (nx10399), .A2 (nx10409)) ;
    nor02_2x ix4518 (.Y (nx4517), .A0 (nx2612), .A1 (nx2610)) ;
    nor03_2x ix2613 (.Y (nx2612), .A0 (nx4521), .A1 (nx9619), .A2 (nx10417)) ;
    dffr gen_6_cmp_mRegCmp_reg_Q_12 (.Q (gen_6_cmp_mReg_12), .QB (nx4521), .D (
         window_6__12), .CLK (start), .R (rst)) ;
    nor03_2x ix2611 (.Y (nx2610), .A0 (gen_6_cmp_mReg_12), .A1 (nx10037), .A2 (
             nx10425)) ;
    nand02 ix2647 (.Y (gen_6_cmp_BSCmp_op2_13), .A0 (nx4527), .A1 (nx4533)) ;
    nor02_2x ix4528 (.Y (nx4527), .A0 (nx2642), .A1 (nx2638)) ;
    nor03_2x ix2643 (.Y (nx2642), .A0 (gen_6_cmp_mReg_12), .A1 (nx9625), .A2 (
             nx10395)) ;
    nor03_2x ix2639 (.Y (nx2638), .A0 (nx4521), .A1 (nx10399), .A2 (nx10411)) ;
    nor02_2x ix4534 (.Y (nx4533), .A0 (nx2634), .A1 (nx2632)) ;
    nor03_2x ix2635 (.Y (nx2634), .A0 (nx4536), .A1 (nx9619), .A2 (nx10419)) ;
    dffr gen_6_cmp_mRegCmp_reg_Q_13 (.Q (gen_6_cmp_mReg_13), .QB (nx4536), .D (
         window_6__13), .CLK (start), .R (rst)) ;
    nor03_2x ix2633 (.Y (nx2632), .A0 (gen_6_cmp_mReg_13), .A1 (nx10037), .A2 (
             nx10427)) ;
    nand02 ix2669 (.Y (gen_6_cmp_BSCmp_op2_14), .A0 (nx4541), .A1 (nx4547)) ;
    nor02_2x ix4542 (.Y (nx4541), .A0 (nx2664), .A1 (nx2660)) ;
    nor03_2x ix2665 (.Y (nx2664), .A0 (gen_6_cmp_mReg_13), .A1 (nx9625), .A2 (
             nx10395)) ;
    nor03_2x ix2661 (.Y (nx2660), .A0 (nx4536), .A1 (nx10401), .A2 (nx10411)) ;
    nor02_2x ix4548 (.Y (nx4547), .A0 (nx2656), .A1 (nx2654)) ;
    nor03_2x ix2657 (.Y (nx2656), .A0 (nx4551), .A1 (nx9619), .A2 (nx10419)) ;
    dffr gen_6_cmp_mRegCmp_reg_Q_14 (.Q (gen_6_cmp_mReg_14), .QB (nx4551), .D (
         window_6__14), .CLK (start), .R (rst)) ;
    nor03_2x ix2655 (.Y (nx2654), .A0 (gen_6_cmp_mReg_14), .A1 (nx10037), .A2 (
             nx10427)) ;
    nand02 ix2691 (.Y (gen_6_cmp_BSCmp_op2_15), .A0 (nx4557), .A1 (nx4561)) ;
    nor02_2x ix4558 (.Y (nx4557), .A0 (nx2686), .A1 (nx2682)) ;
    nor03_2x ix2687 (.Y (nx2686), .A0 (gen_6_cmp_mReg_14), .A1 (nx9625), .A2 (
             nx10395)) ;
    nor03_2x ix2683 (.Y (nx2682), .A0 (nx4551), .A1 (nx10401), .A2 (nx10411)) ;
    nor02_2x ix4562 (.Y (nx4561), .A0 (nx2678), .A1 (nx2676)) ;
    nor03_2x ix2679 (.Y (nx2678), .A0 (nx4565), .A1 (nx9619), .A2 (nx10419)) ;
    dffr gen_6_cmp_mRegCmp_reg_Q_15 (.Q (gen_6_cmp_mReg_15), .QB (nx4565), .D (
         window_6__15), .CLK (start), .R (rst)) ;
    nor03_2x ix2677 (.Y (nx2676), .A0 (gen_6_cmp_mReg_15), .A1 (nx10039), .A2 (
             nx10427)) ;
    nand02 ix2701 (.Y (gen_6_cmp_BSCmp_op2_16), .A0 (nx4571), .A1 (nx4561)) ;
    nor02_2x ix4572 (.Y (nx4571), .A0 (nx2696), .A1 (nx2692)) ;
    nor03_2x ix2697 (.Y (nx2696), .A0 (gen_6_cmp_mReg_15), .A1 (nx9625), .A2 (
             nx10395)) ;
    nor03_2x ix2693 (.Y (nx2692), .A0 (nx4565), .A1 (nx10401), .A2 (nx10411)) ;
    nand02 ix2769 (.Y (gen_7_cmp_BSCmp_op2_1), .A0 (nx4579), .A1 (nx4597)) ;
    nor02_2x ix4580 (.Y (nx4579), .A0 (nx2764), .A1 (nx2760)) ;
    nor03_2x ix2765 (.Y (nx2764), .A0 (gen_7_cmp_mReg_0), .A1 (nx9609), .A2 (
             nx10431)) ;
    dffr gen_7_cmp_mRegCmp_reg_Q_0 (.Q (gen_7_cmp_mReg_0), .QB (nx4583), .D (
         window_7__0), .CLK (start), .R (rst)) ;
    inv01 ix4588 (.Y (nx4587), .A (gen_7_cmp_pMux_0)) ;
    nor03_2x ix2761 (.Y (nx2760), .A0 (nx4583), .A1 (nx10437), .A2 (nx10447)) ;
    inv02 ix4596 (.Y (nx4595), .A (gen_7_cmp_pMux_2)) ;
    nor02_2x ix4598 (.Y (nx4597), .A0 (nx2750), .A1 (nx2748)) ;
    nor03_2x ix2751 (.Y (nx2750), .A0 (nx4601), .A1 (nx9603), .A2 (nx10455)) ;
    dffr gen_7_cmp_mRegCmp_reg_Q_1 (.Q (gen_7_cmp_mReg_1), .QB (nx4601), .D (
         window_7__1), .CLK (start), .R (rst)) ;
    nor03_2x ix2749 (.Y (nx2748), .A0 (gen_7_cmp_mReg_1), .A1 (nx10041), .A2 (
             nx10463)) ;
    nor03_2x ix2709 (.Y (nx2708), .A0 (nx9609), .A1 (nx4595), .A2 (
             gen_7_cmp_pMux_0)) ;
    nand02 ix2791 (.Y (gen_7_cmp_BSCmp_op2_2), .A0 (nx4613), .A1 (nx4617)) ;
    nor02_2x ix4614 (.Y (nx4613), .A0 (nx2786), .A1 (nx2782)) ;
    nor03_2x ix2787 (.Y (nx2786), .A0 (gen_7_cmp_mReg_1), .A1 (nx9609), .A2 (
             nx10431)) ;
    nor03_2x ix2783 (.Y (nx2782), .A0 (nx4601), .A1 (nx10437), .A2 (nx10447)) ;
    nor02_2x ix4618 (.Y (nx4617), .A0 (nx2778), .A1 (nx2776)) ;
    nor03_2x ix2779 (.Y (nx2778), .A0 (nx4621), .A1 (nx9603), .A2 (nx10455)) ;
    dffr gen_7_cmp_mRegCmp_reg_Q_2 (.Q (gen_7_cmp_mReg_2), .QB (nx4621), .D (
         window_7__2), .CLK (start), .R (rst)) ;
    nor03_2x ix2777 (.Y (nx2776), .A0 (gen_7_cmp_mReg_2), .A1 (nx10041), .A2 (
             nx10463)) ;
    nand02 ix2813 (.Y (gen_7_cmp_BSCmp_op2_3), .A0 (nx4627), .A1 (nx4633)) ;
    nor02_2x ix4628 (.Y (nx4627), .A0 (nx2808), .A1 (nx2804)) ;
    nor03_2x ix2809 (.Y (nx2808), .A0 (gen_7_cmp_mReg_2), .A1 (nx9609), .A2 (
             nx10431)) ;
    nor03_2x ix2805 (.Y (nx2804), .A0 (nx4621), .A1 (nx10437), .A2 (nx10447)) ;
    nor02_2x ix4634 (.Y (nx4633), .A0 (nx2800), .A1 (nx2798)) ;
    nor03_2x ix2801 (.Y (nx2800), .A0 (nx4637), .A1 (nx9603), .A2 (nx10455)) ;
    dffr gen_7_cmp_mRegCmp_reg_Q_3 (.Q (gen_7_cmp_mReg_3), .QB (nx4637), .D (
         window_7__3), .CLK (start), .R (rst)) ;
    nor03_2x ix2799 (.Y (nx2798), .A0 (gen_7_cmp_mReg_3), .A1 (nx10041), .A2 (
             nx10463)) ;
    nand02 ix2835 (.Y (gen_7_cmp_BSCmp_op2_4), .A0 (nx4642), .A1 (nx4646)) ;
    nor02_2x ix4643 (.Y (nx4642), .A0 (nx2830), .A1 (nx2826)) ;
    nor03_2x ix2831 (.Y (nx2830), .A0 (gen_7_cmp_mReg_3), .A1 (nx9609), .A2 (
             nx10431)) ;
    nor03_2x ix2827 (.Y (nx2826), .A0 (nx4637), .A1 (nx10437), .A2 (nx10447)) ;
    nor02_2x ix4647 (.Y (nx4646), .A0 (nx2822), .A1 (nx2820)) ;
    nor03_2x ix2823 (.Y (nx2822), .A0 (nx4649), .A1 (nx9603), .A2 (nx10455)) ;
    dffr gen_7_cmp_mRegCmp_reg_Q_4 (.Q (gen_7_cmp_mReg_4), .QB (nx4649), .D (
         window_7__4), .CLK (start), .R (rst)) ;
    nor03_2x ix2821 (.Y (nx2820), .A0 (gen_7_cmp_mReg_4), .A1 (nx10041), .A2 (
             nx10463)) ;
    nand02 ix2857 (.Y (gen_7_cmp_BSCmp_op2_5), .A0 (nx4655), .A1 (nx4661)) ;
    nor02_2x ix4656 (.Y (nx4655), .A0 (nx2852), .A1 (nx2848)) ;
    nor03_2x ix2853 (.Y (nx2852), .A0 (gen_7_cmp_mReg_4), .A1 (nx9609), .A2 (
             nx10431)) ;
    nor03_2x ix2849 (.Y (nx2848), .A0 (nx4649), .A1 (nx10437), .A2 (nx10447)) ;
    nor02_2x ix4662 (.Y (nx4661), .A0 (nx2844), .A1 (nx2842)) ;
    nor03_2x ix2845 (.Y (nx2844), .A0 (nx4665), .A1 (nx9605), .A2 (nx10455)) ;
    dffr gen_7_cmp_mRegCmp_reg_Q_5 (.Q (gen_7_cmp_mReg_5), .QB (nx4665), .D (
         window_7__5), .CLK (start), .R (rst)) ;
    nor03_2x ix2843 (.Y (nx2842), .A0 (gen_7_cmp_mReg_5), .A1 (nx10041), .A2 (
             nx10463)) ;
    nand02 ix2879 (.Y (gen_7_cmp_BSCmp_op2_6), .A0 (nx4671), .A1 (nx4675)) ;
    nor02_2x ix4672 (.Y (nx4671), .A0 (nx2874), .A1 (nx2870)) ;
    nor03_2x ix2875 (.Y (nx2874), .A0 (gen_7_cmp_mReg_5), .A1 (nx9611), .A2 (
             nx10431)) ;
    nor03_2x ix2871 (.Y (nx2870), .A0 (nx4665), .A1 (nx10437), .A2 (nx10447)) ;
    nor02_2x ix4676 (.Y (nx4675), .A0 (nx2866), .A1 (nx2864)) ;
    nor03_2x ix2867 (.Y (nx2866), .A0 (nx4679), .A1 (nx9605), .A2 (nx10455)) ;
    dffr gen_7_cmp_mRegCmp_reg_Q_6 (.Q (gen_7_cmp_mReg_6), .QB (nx4679), .D (
         window_7__6), .CLK (start), .R (rst)) ;
    nor03_2x ix2865 (.Y (nx2864), .A0 (gen_7_cmp_mReg_6), .A1 (nx10041), .A2 (
             nx10463)) ;
    nand02 ix2901 (.Y (gen_7_cmp_BSCmp_op2_7), .A0 (nx4685), .A1 (nx4691)) ;
    nor02_2x ix4686 (.Y (nx4685), .A0 (nx2896), .A1 (nx2892)) ;
    nor03_2x ix2897 (.Y (nx2896), .A0 (gen_7_cmp_mReg_6), .A1 (nx9611), .A2 (
             nx10433)) ;
    nor03_2x ix2893 (.Y (nx2892), .A0 (nx4679), .A1 (nx10439), .A2 (nx10449)) ;
    nor02_2x ix4692 (.Y (nx4691), .A0 (nx2888), .A1 (nx2886)) ;
    nor03_2x ix2889 (.Y (nx2888), .A0 (nx4695), .A1 (nx9605), .A2 (nx10457)) ;
    dffr gen_7_cmp_mRegCmp_reg_Q_7 (.Q (gen_7_cmp_mReg_7), .QB (nx4695), .D (
         window_7__7), .CLK (start), .R (rst)) ;
    nor03_2x ix2887 (.Y (nx2886), .A0 (gen_7_cmp_mReg_7), .A1 (nx10041), .A2 (
             nx10465)) ;
    nand02 ix2923 (.Y (gen_7_cmp_BSCmp_op2_8), .A0 (nx4701), .A1 (nx4705)) ;
    nor02_2x ix4702 (.Y (nx4701), .A0 (nx2918), .A1 (nx2914)) ;
    nor03_2x ix2919 (.Y (nx2918), .A0 (gen_7_cmp_mReg_7), .A1 (nx9611), .A2 (
             nx10433)) ;
    nor03_2x ix2915 (.Y (nx2914), .A0 (nx4695), .A1 (nx10439), .A2 (nx10449)) ;
    nor02_2x ix4706 (.Y (nx4705), .A0 (nx2910), .A1 (nx2908)) ;
    nor03_2x ix2911 (.Y (nx2910), .A0 (nx4709), .A1 (nx9605), .A2 (nx10457)) ;
    dffr gen_7_cmp_mRegCmp_reg_Q_8 (.Q (gen_7_cmp_mReg_8), .QB (nx4709), .D (
         window_7__8), .CLK (start), .R (rst)) ;
    nor03_2x ix2909 (.Y (nx2908), .A0 (gen_7_cmp_mReg_8), .A1 (nx10043), .A2 (
             nx10465)) ;
    nand02 ix2945 (.Y (gen_7_cmp_BSCmp_op2_9), .A0 (nx4715), .A1 (nx4721)) ;
    nor02_2x ix4716 (.Y (nx4715), .A0 (nx2940), .A1 (nx2936)) ;
    nor03_2x ix2941 (.Y (nx2940), .A0 (gen_7_cmp_mReg_8), .A1 (nx9611), .A2 (
             nx10433)) ;
    nor03_2x ix2937 (.Y (nx2936), .A0 (nx4709), .A1 (nx10439), .A2 (nx10449)) ;
    nor02_2x ix4722 (.Y (nx4721), .A0 (nx2932), .A1 (nx2930)) ;
    nor03_2x ix2933 (.Y (nx2932), .A0 (nx4724), .A1 (nx9605), .A2 (nx10457)) ;
    dffr gen_7_cmp_mRegCmp_reg_Q_9 (.Q (gen_7_cmp_mReg_9), .QB (nx4724), .D (
         window_7__9), .CLK (start), .R (rst)) ;
    nor03_2x ix2931 (.Y (nx2930), .A0 (gen_7_cmp_mReg_9), .A1 (nx10043), .A2 (
             nx10465)) ;
    nand02 ix2967 (.Y (gen_7_cmp_BSCmp_op2_10), .A0 (nx4729), .A1 (nx4735)) ;
    nor02_2x ix4730 (.Y (nx4729), .A0 (nx2962), .A1 (nx2958)) ;
    nor03_2x ix2963 (.Y (nx2962), .A0 (gen_7_cmp_mReg_9), .A1 (nx9611), .A2 (
             nx10433)) ;
    nor03_2x ix2959 (.Y (nx2958), .A0 (nx4724), .A1 (nx10439), .A2 (nx10449)) ;
    nor02_2x ix4736 (.Y (nx4735), .A0 (nx2954), .A1 (nx2952)) ;
    nor03_2x ix2955 (.Y (nx2954), .A0 (nx4739), .A1 (nx9605), .A2 (nx10457)) ;
    dffr gen_7_cmp_mRegCmp_reg_Q_10 (.Q (gen_7_cmp_mReg_10), .QB (nx4739), .D (
         window_7__10), .CLK (start), .R (rst)) ;
    nor03_2x ix2953 (.Y (nx2952), .A0 (gen_7_cmp_mReg_10), .A1 (nx10043), .A2 (
             nx10465)) ;
    nand02 ix2989 (.Y (gen_7_cmp_BSCmp_op2_11), .A0 (nx4745), .A1 (nx4749)) ;
    nor02_2x ix4746 (.Y (nx4745), .A0 (nx2984), .A1 (nx2980)) ;
    nor03_2x ix2985 (.Y (nx2984), .A0 (gen_7_cmp_mReg_10), .A1 (nx9611), .A2 (
             nx10433)) ;
    nor03_2x ix2981 (.Y (nx2980), .A0 (nx4739), .A1 (nx10439), .A2 (nx10449)) ;
    nor02_2x ix4750 (.Y (nx4749), .A0 (nx2976), .A1 (nx2974)) ;
    nor03_2x ix2977 (.Y (nx2976), .A0 (nx4753), .A1 (nx9605), .A2 (nx10457)) ;
    dffr gen_7_cmp_mRegCmp_reg_Q_11 (.Q (gen_7_cmp_mReg_11), .QB (nx4753), .D (
         window_7__11), .CLK (start), .R (rst)) ;
    nor03_2x ix2975 (.Y (nx2974), .A0 (gen_7_cmp_mReg_11), .A1 (nx10043), .A2 (
             nx10465)) ;
    nand02 ix3011 (.Y (gen_7_cmp_BSCmp_op2_12), .A0 (nx4759), .A1 (nx4765)) ;
    nor02_2x ix4760 (.Y (nx4759), .A0 (nx3006), .A1 (nx3002)) ;
    nor03_2x ix3007 (.Y (nx3006), .A0 (gen_7_cmp_mReg_11), .A1 (nx9611), .A2 (
             nx10433)) ;
    nor03_2x ix3003 (.Y (nx3002), .A0 (nx4753), .A1 (nx10439), .A2 (nx10449)) ;
    nor02_2x ix4766 (.Y (nx4765), .A0 (nx2998), .A1 (nx2996)) ;
    nor03_2x ix2999 (.Y (nx2998), .A0 (nx4768), .A1 (nx9607), .A2 (nx10457)) ;
    dffr gen_7_cmp_mRegCmp_reg_Q_12 (.Q (gen_7_cmp_mReg_12), .QB (nx4768), .D (
         window_7__12), .CLK (start), .R (rst)) ;
    nor03_2x ix2997 (.Y (nx2996), .A0 (gen_7_cmp_mReg_12), .A1 (nx10043), .A2 (
             nx10465)) ;
    nand02 ix3033 (.Y (gen_7_cmp_BSCmp_op2_13), .A0 (nx4773), .A1 (nx4779)) ;
    nor02_2x ix4774 (.Y (nx4773), .A0 (nx3028), .A1 (nx3024)) ;
    nor03_2x ix3029 (.Y (nx3028), .A0 (gen_7_cmp_mReg_12), .A1 (nx9613), .A2 (
             nx10435)) ;
    nor03_2x ix3025 (.Y (nx3024), .A0 (nx4768), .A1 (nx10439), .A2 (nx10451)) ;
    nor02_2x ix4780 (.Y (nx4779), .A0 (nx3020), .A1 (nx3018)) ;
    nor03_2x ix3021 (.Y (nx3020), .A0 (nx4783), .A1 (nx9607), .A2 (nx10459)) ;
    dffr gen_7_cmp_mRegCmp_reg_Q_13 (.Q (gen_7_cmp_mReg_13), .QB (nx4783), .D (
         window_7__13), .CLK (start), .R (rst)) ;
    nor03_2x ix3019 (.Y (nx3018), .A0 (gen_7_cmp_mReg_13), .A1 (nx10043), .A2 (
             nx10467)) ;
    nand02 ix3055 (.Y (gen_7_cmp_BSCmp_op2_14), .A0 (nx4789), .A1 (nx4793)) ;
    nor02_2x ix4790 (.Y (nx4789), .A0 (nx3050), .A1 (nx3046)) ;
    nor03_2x ix3051 (.Y (nx3050), .A0 (gen_7_cmp_mReg_13), .A1 (nx9613), .A2 (
             nx10435)) ;
    nor03_2x ix3047 (.Y (nx3046), .A0 (nx4783), .A1 (nx10441), .A2 (nx10451)) ;
    nor02_2x ix4794 (.Y (nx4793), .A0 (nx3042), .A1 (nx3040)) ;
    nor03_2x ix3043 (.Y (nx3042), .A0 (nx4797), .A1 (nx9607), .A2 (nx10459)) ;
    dffr gen_7_cmp_mRegCmp_reg_Q_14 (.Q (gen_7_cmp_mReg_14), .QB (nx4797), .D (
         window_7__14), .CLK (start), .R (rst)) ;
    nor03_2x ix3041 (.Y (nx3040), .A0 (gen_7_cmp_mReg_14), .A1 (nx10043), .A2 (
             nx10467)) ;
    nand02 ix3077 (.Y (gen_7_cmp_BSCmp_op2_15), .A0 (nx4803), .A1 (nx4809)) ;
    nor02_2x ix4804 (.Y (nx4803), .A0 (nx3072), .A1 (nx3068)) ;
    nor03_2x ix3073 (.Y (nx3072), .A0 (gen_7_cmp_mReg_14), .A1 (nx9613), .A2 (
             nx10435)) ;
    nor03_2x ix3069 (.Y (nx3068), .A0 (nx4797), .A1 (nx10441), .A2 (nx10451)) ;
    nor02_2x ix4810 (.Y (nx4809), .A0 (nx3064), .A1 (nx3062)) ;
    nor03_2x ix3065 (.Y (nx3064), .A0 (nx4812), .A1 (nx9607), .A2 (nx10459)) ;
    dffr gen_7_cmp_mRegCmp_reg_Q_15 (.Q (gen_7_cmp_mReg_15), .QB (nx4812), .D (
         window_7__15), .CLK (start), .R (rst)) ;
    nor03_2x ix3063 (.Y (nx3062), .A0 (gen_7_cmp_mReg_15), .A1 (nx10045), .A2 (
             nx10467)) ;
    nand02 ix3087 (.Y (gen_7_cmp_BSCmp_op2_16), .A0 (nx4817), .A1 (nx4809)) ;
    nor02_2x ix4818 (.Y (nx4817), .A0 (nx3082), .A1 (nx3078)) ;
    nor03_2x ix3083 (.Y (nx3082), .A0 (gen_7_cmp_mReg_15), .A1 (nx9613), .A2 (
             nx10435)) ;
    nor03_2x ix3079 (.Y (nx3078), .A0 (nx4812), .A1 (nx10441), .A2 (nx10451)) ;
    nand02 ix3155 (.Y (gen_8_cmp_BSCmp_op2_1), .A0 (nx4825), .A1 (nx4843)) ;
    nor02_2x ix4826 (.Y (nx4825), .A0 (nx3150), .A1 (nx3146)) ;
    nor03_2x ix3151 (.Y (nx3150), .A0 (gen_8_cmp_mReg_0), .A1 (nx9597), .A2 (
             nx10471)) ;
    dffr gen_8_cmp_mRegCmp_reg_Q_0 (.Q (gen_8_cmp_mReg_0), .QB (nx4831), .D (
         window_8__0), .CLK (start), .R (rst)) ;
    inv01 ix4835 (.Y (nx4834), .A (gen_8_cmp_pMux_0)) ;
    nor03_2x ix3147 (.Y (nx3146), .A0 (nx4831), .A1 (nx10477), .A2 (nx10487)) ;
    inv02 ix4842 (.Y (nx4841), .A (gen_8_cmp_pMux_2)) ;
    nor02_2x ix4844 (.Y (nx4843), .A0 (nx3136), .A1 (nx3134)) ;
    nor03_2x ix3137 (.Y (nx3136), .A0 (nx4847), .A1 (nx9591), .A2 (nx10495)) ;
    dffr gen_8_cmp_mRegCmp_reg_Q_1 (.Q (gen_8_cmp_mReg_1), .QB (nx4847), .D (
         window_8__1), .CLK (start), .R (rst)) ;
    nor03_2x ix3135 (.Y (nx3134), .A0 (gen_8_cmp_mReg_1), .A1 (nx10047), .A2 (
             nx10503)) ;
    nor03_2x ix3095 (.Y (nx3094), .A0 (nx9597), .A1 (nx4841), .A2 (
             gen_8_cmp_pMux_0)) ;
    nand02 ix3177 (.Y (gen_8_cmp_BSCmp_op2_2), .A0 (nx4858), .A1 (nx4865)) ;
    nor02_2x ix4860 (.Y (nx4858), .A0 (nx3172), .A1 (nx3168)) ;
    nor03_2x ix3173 (.Y (nx3172), .A0 (gen_8_cmp_mReg_1), .A1 (nx9597), .A2 (
             nx10471)) ;
    nor03_2x ix3169 (.Y (nx3168), .A0 (nx4847), .A1 (nx10477), .A2 (nx10487)) ;
    nor02_2x ix4866 (.Y (nx4865), .A0 (nx3164), .A1 (nx3162)) ;
    nor03_2x ix3165 (.Y (nx3164), .A0 (nx4869), .A1 (nx9591), .A2 (nx10495)) ;
    dffr gen_8_cmp_mRegCmp_reg_Q_2 (.Q (gen_8_cmp_mReg_2), .QB (nx4869), .D (
         window_8__2), .CLK (start), .R (rst)) ;
    nor03_2x ix3163 (.Y (nx3162), .A0 (gen_8_cmp_mReg_2), .A1 (nx10047), .A2 (
             nx10503)) ;
    nand02 ix3199 (.Y (gen_8_cmp_BSCmp_op2_3), .A0 (nx4875), .A1 (nx4879)) ;
    nor02_2x ix4876 (.Y (nx4875), .A0 (nx3194), .A1 (nx3190)) ;
    nor03_2x ix3195 (.Y (nx3194), .A0 (gen_8_cmp_mReg_2), .A1 (nx9597), .A2 (
             nx10471)) ;
    nor03_2x ix3191 (.Y (nx3190), .A0 (nx4869), .A1 (nx10477), .A2 (nx10487)) ;
    nor02_2x ix4880 (.Y (nx4879), .A0 (nx3186), .A1 (nx3184)) ;
    nor03_2x ix3187 (.Y (nx3186), .A0 (nx4883), .A1 (nx9591), .A2 (nx10495)) ;
    dffr gen_8_cmp_mRegCmp_reg_Q_3 (.Q (gen_8_cmp_mReg_3), .QB (nx4883), .D (
         window_8__3), .CLK (start), .R (rst)) ;
    nor03_2x ix3185 (.Y (nx3184), .A0 (gen_8_cmp_mReg_3), .A1 (nx10047), .A2 (
             nx10503)) ;
    nand02 ix3221 (.Y (gen_8_cmp_BSCmp_op2_4), .A0 (nx4889), .A1 (nx4893)) ;
    nor02_2x ix4890 (.Y (nx4889), .A0 (nx3216), .A1 (nx3212)) ;
    nor03_2x ix3217 (.Y (nx3216), .A0 (gen_8_cmp_mReg_3), .A1 (nx9597), .A2 (
             nx10471)) ;
    nor03_2x ix3213 (.Y (nx3212), .A0 (nx4883), .A1 (nx10477), .A2 (nx10487)) ;
    nor02_2x ix4894 (.Y (nx4893), .A0 (nx3208), .A1 (nx3206)) ;
    nor03_2x ix3209 (.Y (nx3208), .A0 (nx4897), .A1 (nx9591), .A2 (nx10495)) ;
    dffr gen_8_cmp_mRegCmp_reg_Q_4 (.Q (gen_8_cmp_mReg_4), .QB (nx4897), .D (
         window_8__4), .CLK (start), .R (rst)) ;
    nor03_2x ix3207 (.Y (nx3206), .A0 (gen_8_cmp_mReg_4), .A1 (nx10047), .A2 (
             nx10503)) ;
    nand02 ix3243 (.Y (gen_8_cmp_BSCmp_op2_5), .A0 (nx4901), .A1 (nx4907)) ;
    nor02_2x ix4902 (.Y (nx4901), .A0 (nx3238), .A1 (nx3234)) ;
    nor03_2x ix3239 (.Y (nx3238), .A0 (gen_8_cmp_mReg_4), .A1 (nx9597), .A2 (
             nx10471)) ;
    nor03_2x ix3235 (.Y (nx3234), .A0 (nx4897), .A1 (nx10477), .A2 (nx10487)) ;
    nor02_2x ix4908 (.Y (nx4907), .A0 (nx3230), .A1 (nx3228)) ;
    nor03_2x ix3231 (.Y (nx3230), .A0 (nx4911), .A1 (nx9593), .A2 (nx10495)) ;
    dffr gen_8_cmp_mRegCmp_reg_Q_5 (.Q (gen_8_cmp_mReg_5), .QB (nx4911), .D (
         window_8__5), .CLK (start), .R (rst)) ;
    nor03_2x ix3229 (.Y (nx3228), .A0 (gen_8_cmp_mReg_5), .A1 (nx10047), .A2 (
             nx10503)) ;
    nand02 ix3265 (.Y (gen_8_cmp_BSCmp_op2_6), .A0 (nx4915), .A1 (nx4921)) ;
    nor02_2x ix4916 (.Y (nx4915), .A0 (nx3260), .A1 (nx3256)) ;
    nor03_2x ix3261 (.Y (nx3260), .A0 (gen_8_cmp_mReg_5), .A1 (nx9599), .A2 (
             nx10471)) ;
    nor03_2x ix3257 (.Y (nx3256), .A0 (nx4911), .A1 (nx10477), .A2 (nx10487)) ;
    nor02_2x ix4922 (.Y (nx4921), .A0 (nx3252), .A1 (nx3250)) ;
    nor03_2x ix3253 (.Y (nx3252), .A0 (nx4924), .A1 (nx9593), .A2 (nx10495)) ;
    dffr gen_8_cmp_mRegCmp_reg_Q_6 (.Q (gen_8_cmp_mReg_6), .QB (nx4924), .D (
         window_8__6), .CLK (start), .R (rst)) ;
    nor03_2x ix3251 (.Y (nx3250), .A0 (gen_8_cmp_mReg_6), .A1 (nx10047), .A2 (
             nx10503)) ;
    nand02 ix3287 (.Y (gen_8_cmp_BSCmp_op2_7), .A0 (nx4931), .A1 (nx4937)) ;
    nor02_2x ix4932 (.Y (nx4931), .A0 (nx3282), .A1 (nx3278)) ;
    nor03_2x ix3283 (.Y (nx3282), .A0 (gen_8_cmp_mReg_6), .A1 (nx9599), .A2 (
             nx10473)) ;
    nor03_2x ix3279 (.Y (nx3278), .A0 (nx4924), .A1 (nx10479), .A2 (nx10489)) ;
    nor02_2x ix4938 (.Y (nx4937), .A0 (nx3274), .A1 (nx3272)) ;
    nor03_2x ix3275 (.Y (nx3274), .A0 (nx4941), .A1 (nx9593), .A2 (nx10497)) ;
    dffr gen_8_cmp_mRegCmp_reg_Q_7 (.Q (gen_8_cmp_mReg_7), .QB (nx4941), .D (
         window_8__7), .CLK (start), .R (rst)) ;
    nor03_2x ix3273 (.Y (nx3272), .A0 (gen_8_cmp_mReg_7), .A1 (nx10047), .A2 (
             nx10505)) ;
    nand02 ix3309 (.Y (gen_8_cmp_BSCmp_op2_8), .A0 (nx4945), .A1 (nx4951)) ;
    nor02_2x ix4946 (.Y (nx4945), .A0 (nx3304), .A1 (nx3300)) ;
    nor03_2x ix3305 (.Y (nx3304), .A0 (gen_8_cmp_mReg_7), .A1 (nx9599), .A2 (
             nx10473)) ;
    nor03_2x ix3301 (.Y (nx3300), .A0 (nx4941), .A1 (nx10479), .A2 (nx10489)) ;
    nor02_2x ix4952 (.Y (nx4951), .A0 (nx3296), .A1 (nx3294)) ;
    nor03_2x ix3297 (.Y (nx3296), .A0 (nx4955), .A1 (nx9593), .A2 (nx10497)) ;
    dffr gen_8_cmp_mRegCmp_reg_Q_8 (.Q (gen_8_cmp_mReg_8), .QB (nx4955), .D (
         window_8__8), .CLK (start), .R (rst)) ;
    nor03_2x ix3295 (.Y (nx3294), .A0 (gen_8_cmp_mReg_8), .A1 (nx10049), .A2 (
             nx10505)) ;
    nand02 ix3331 (.Y (gen_8_cmp_BSCmp_op2_9), .A0 (nx4959), .A1 (nx4965)) ;
    nor02_2x ix4960 (.Y (nx4959), .A0 (nx3326), .A1 (nx3322)) ;
    nor03_2x ix3327 (.Y (nx3326), .A0 (gen_8_cmp_mReg_8), .A1 (nx9599), .A2 (
             nx10473)) ;
    nor03_2x ix3323 (.Y (nx3322), .A0 (nx4955), .A1 (nx10479), .A2 (nx10489)) ;
    nor02_2x ix4966 (.Y (nx4965), .A0 (nx3318), .A1 (nx3316)) ;
    nor03_2x ix3319 (.Y (nx3318), .A0 (nx4968), .A1 (nx9593), .A2 (nx10497)) ;
    dffr gen_8_cmp_mRegCmp_reg_Q_9 (.Q (gen_8_cmp_mReg_9), .QB (nx4968), .D (
         window_8__9), .CLK (start), .R (rst)) ;
    nor03_2x ix3317 (.Y (nx3316), .A0 (gen_8_cmp_mReg_9), .A1 (nx10049), .A2 (
             nx10505)) ;
    nand02 ix3353 (.Y (gen_8_cmp_BSCmp_op2_10), .A0 (nx4975), .A1 (nx4981)) ;
    nor02_2x ix4976 (.Y (nx4975), .A0 (nx3348), .A1 (nx3344)) ;
    nor03_2x ix3349 (.Y (nx3348), .A0 (gen_8_cmp_mReg_9), .A1 (nx9599), .A2 (
             nx10473)) ;
    nor03_2x ix3345 (.Y (nx3344), .A0 (nx4968), .A1 (nx10479), .A2 (nx10489)) ;
    nor02_2x ix4982 (.Y (nx4981), .A0 (nx3340), .A1 (nx3338)) ;
    nor03_2x ix3341 (.Y (nx3340), .A0 (nx4985), .A1 (nx9593), .A2 (nx10497)) ;
    dffr gen_8_cmp_mRegCmp_reg_Q_10 (.Q (gen_8_cmp_mReg_10), .QB (nx4985), .D (
         window_8__10), .CLK (start), .R (rst)) ;
    nor03_2x ix3339 (.Y (nx3338), .A0 (gen_8_cmp_mReg_10), .A1 (nx10049), .A2 (
             nx10505)) ;
    nand02 ix3375 (.Y (gen_8_cmp_BSCmp_op2_11), .A0 (nx4989), .A1 (nx4995)) ;
    nor02_2x ix4990 (.Y (nx4989), .A0 (nx3370), .A1 (nx3366)) ;
    nor03_2x ix3371 (.Y (nx3370), .A0 (gen_8_cmp_mReg_10), .A1 (nx9599), .A2 (
             nx10473)) ;
    nor03_2x ix3367 (.Y (nx3366), .A0 (nx4985), .A1 (nx10479), .A2 (nx10489)) ;
    nor02_2x ix4996 (.Y (nx4995), .A0 (nx3362), .A1 (nx3360)) ;
    nor03_2x ix3363 (.Y (nx3362), .A0 (nx4999), .A1 (nx9593), .A2 (nx10497)) ;
    dffr gen_8_cmp_mRegCmp_reg_Q_11 (.Q (gen_8_cmp_mReg_11), .QB (nx4999), .D (
         window_8__11), .CLK (start), .R (rst)) ;
    nor03_2x ix3361 (.Y (nx3360), .A0 (gen_8_cmp_mReg_11), .A1 (nx10049), .A2 (
             nx10505)) ;
    nand02 ix3397 (.Y (gen_8_cmp_BSCmp_op2_12), .A0 (nx5003), .A1 (nx5009)) ;
    nor02_2x ix5004 (.Y (nx5003), .A0 (nx3392), .A1 (nx3388)) ;
    nor03_2x ix3393 (.Y (nx3392), .A0 (gen_8_cmp_mReg_11), .A1 (nx9599), .A2 (
             nx10473)) ;
    nor03_2x ix3389 (.Y (nx3388), .A0 (nx4999), .A1 (nx10479), .A2 (nx10489)) ;
    nor02_2x ix5010 (.Y (nx5009), .A0 (nx3384), .A1 (nx3382)) ;
    nor03_2x ix3385 (.Y (nx3384), .A0 (nx5013), .A1 (nx9595), .A2 (nx10497)) ;
    dffr gen_8_cmp_mRegCmp_reg_Q_12 (.Q (gen_8_cmp_mReg_12), .QB (nx5013), .D (
         window_8__12), .CLK (start), .R (rst)) ;
    nor03_2x ix3383 (.Y (nx3382), .A0 (gen_8_cmp_mReg_12), .A1 (nx10049), .A2 (
             nx10505)) ;
    nand02 ix3419 (.Y (gen_8_cmp_BSCmp_op2_13), .A0 (nx5019), .A1 (nx5025)) ;
    nor02_2x ix5020 (.Y (nx5019), .A0 (nx3414), .A1 (nx3410)) ;
    nor03_2x ix3415 (.Y (nx3414), .A0 (gen_8_cmp_mReg_12), .A1 (nx9601), .A2 (
             nx10475)) ;
    nor03_2x ix3411 (.Y (nx3410), .A0 (nx5013), .A1 (nx10479), .A2 (nx10491)) ;
    nor02_2x ix5026 (.Y (nx5025), .A0 (nx3406), .A1 (nx3404)) ;
    nor03_2x ix3407 (.Y (nx3406), .A0 (nx5028), .A1 (nx9595), .A2 (nx10499)) ;
    dffr gen_8_cmp_mRegCmp_reg_Q_13 (.Q (gen_8_cmp_mReg_13), .QB (nx5028), .D (
         window_8__13), .CLK (start), .R (rst)) ;
    nor03_2x ix3405 (.Y (nx3404), .A0 (gen_8_cmp_mReg_13), .A1 (nx10049), .A2 (
             nx10507)) ;
    nand02 ix3441 (.Y (gen_8_cmp_BSCmp_op2_14), .A0 (nx5032), .A1 (nx5037)) ;
    nor02_2x ix5033 (.Y (nx5032), .A0 (nx3436), .A1 (nx3432)) ;
    nor03_2x ix3437 (.Y (nx3436), .A0 (gen_8_cmp_mReg_13), .A1 (nx9601), .A2 (
             nx10475)) ;
    nor03_2x ix3433 (.Y (nx3432), .A0 (nx5028), .A1 (nx10481), .A2 (nx10491)) ;
    nor02_2x ix5038 (.Y (nx5037), .A0 (nx3428), .A1 (nx3426)) ;
    nor03_2x ix3429 (.Y (nx3428), .A0 (nx5041), .A1 (nx9595), .A2 (nx10499)) ;
    dffr gen_8_cmp_mRegCmp_reg_Q_14 (.Q (gen_8_cmp_mReg_14), .QB (nx5041), .D (
         window_8__14), .CLK (start), .R (rst)) ;
    nor03_2x ix3427 (.Y (nx3426), .A0 (gen_8_cmp_mReg_14), .A1 (nx10049), .A2 (
             nx10507)) ;
    nand02 ix3463 (.Y (gen_8_cmp_BSCmp_op2_15), .A0 (nx5047), .A1 (nx5053)) ;
    nor02_2x ix5048 (.Y (nx5047), .A0 (nx3458), .A1 (nx3454)) ;
    nor03_2x ix3459 (.Y (nx3458), .A0 (gen_8_cmp_mReg_14), .A1 (nx9601), .A2 (
             nx10475)) ;
    nor03_2x ix3455 (.Y (nx3454), .A0 (nx5041), .A1 (nx10481), .A2 (nx10491)) ;
    nor02_2x ix5054 (.Y (nx5053), .A0 (nx3450), .A1 (nx3448)) ;
    nor03_2x ix3451 (.Y (nx3450), .A0 (nx5057), .A1 (nx9595), .A2 (nx10499)) ;
    dffr gen_8_cmp_mRegCmp_reg_Q_15 (.Q (gen_8_cmp_mReg_15), .QB (nx5057), .D (
         window_8__15), .CLK (start), .R (rst)) ;
    nor03_2x ix3449 (.Y (nx3448), .A0 (gen_8_cmp_mReg_15), .A1 (nx10051), .A2 (
             nx10507)) ;
    nand02 ix3473 (.Y (gen_8_cmp_BSCmp_op2_16), .A0 (nx5061), .A1 (nx5053)) ;
    nor02_2x ix5062 (.Y (nx5061), .A0 (nx3468), .A1 (nx3464)) ;
    nor03_2x ix3469 (.Y (nx3468), .A0 (gen_8_cmp_mReg_15), .A1 (nx9601), .A2 (
             nx10475)) ;
    nor03_2x ix3465 (.Y (nx3464), .A0 (nx5057), .A1 (nx10481), .A2 (nx10491)) ;
    nand02 ix3541 (.Y (gen_9_cmp_BSCmp_op2_1), .A0 (nx5069), .A1 (nx5087)) ;
    nor02_2x ix5070 (.Y (nx5069), .A0 (nx3536), .A1 (nx3532)) ;
    nor03_2x ix3537 (.Y (nx3536), .A0 (gen_9_cmp_mReg_0), .A1 (nx9585), .A2 (
             nx10511)) ;
    dffr gen_9_cmp_mRegCmp_reg_Q_0 (.Q (gen_9_cmp_mReg_0), .QB (nx5073), .D (
         window_9__0), .CLK (start), .R (rst)) ;
    inv01 ix5078 (.Y (nx5077), .A (gen_9_cmp_pMux_0)) ;
    nor03_2x ix3533 (.Y (nx3532), .A0 (nx5073), .A1 (nx10517), .A2 (nx10527)) ;
    inv02 ix5086 (.Y (nx5085), .A (gen_9_cmp_pMux_2)) ;
    nor02_2x ix5088 (.Y (nx5087), .A0 (nx3522), .A1 (nx3520)) ;
    nor03_2x ix3523 (.Y (nx3522), .A0 (nx5090), .A1 (nx9579), .A2 (nx10535)) ;
    dffr gen_9_cmp_mRegCmp_reg_Q_1 (.Q (gen_9_cmp_mReg_1), .QB (nx5090), .D (
         window_9__1), .CLK (start), .R (rst)) ;
    nor03_2x ix3521 (.Y (nx3520), .A0 (gen_9_cmp_mReg_1), .A1 (nx10053), .A2 (
             nx10543)) ;
    nor03_2x ix3481 (.Y (nx3480), .A0 (nx9585), .A1 (nx5085), .A2 (
             gen_9_cmp_pMux_0)) ;
    nand02 ix3563 (.Y (gen_9_cmp_BSCmp_op2_2), .A0 (nx5103), .A1 (nx5109)) ;
    nor02_2x ix5104 (.Y (nx5103), .A0 (nx3558), .A1 (nx3554)) ;
    nor03_2x ix3559 (.Y (nx3558), .A0 (gen_9_cmp_mReg_1), .A1 (nx9585), .A2 (
             nx10511)) ;
    nor03_2x ix3555 (.Y (nx3554), .A0 (nx5090), .A1 (nx10517), .A2 (nx10527)) ;
    nor02_2x ix5110 (.Y (nx5109), .A0 (nx3550), .A1 (nx3548)) ;
    nor03_2x ix3551 (.Y (nx3550), .A0 (nx5112), .A1 (nx9579), .A2 (nx10535)) ;
    dffr gen_9_cmp_mRegCmp_reg_Q_2 (.Q (gen_9_cmp_mReg_2), .QB (nx5112), .D (
         window_9__2), .CLK (start), .R (rst)) ;
    nor03_2x ix3549 (.Y (nx3548), .A0 (gen_9_cmp_mReg_2), .A1 (nx10053), .A2 (
             nx10543)) ;
    nand02 ix3585 (.Y (gen_9_cmp_BSCmp_op2_3), .A0 (nx5119), .A1 (nx5125)) ;
    nor02_2x ix5120 (.Y (nx5119), .A0 (nx3580), .A1 (nx3576)) ;
    nor03_2x ix3581 (.Y (nx3580), .A0 (gen_9_cmp_mReg_2), .A1 (nx9585), .A2 (
             nx10511)) ;
    nor03_2x ix3577 (.Y (nx3576), .A0 (nx5112), .A1 (nx10517), .A2 (nx10527)) ;
    nor02_2x ix5126 (.Y (nx5125), .A0 (nx3572), .A1 (nx3570)) ;
    nor03_2x ix3573 (.Y (nx3572), .A0 (nx5129), .A1 (nx9579), .A2 (nx10535)) ;
    dffr gen_9_cmp_mRegCmp_reg_Q_3 (.Q (gen_9_cmp_mReg_3), .QB (nx5129), .D (
         window_9__3), .CLK (start), .R (rst)) ;
    nor03_2x ix3571 (.Y (nx3570), .A0 (gen_9_cmp_mReg_3), .A1 (nx10053), .A2 (
             nx10543)) ;
    nand02 ix3607 (.Y (gen_9_cmp_BSCmp_op2_4), .A0 (nx5133), .A1 (nx5139)) ;
    nor02_2x ix5134 (.Y (nx5133), .A0 (nx3602), .A1 (nx3598)) ;
    nor03_2x ix3603 (.Y (nx3602), .A0 (gen_9_cmp_mReg_3), .A1 (nx9585), .A2 (
             nx10511)) ;
    nor03_2x ix3599 (.Y (nx3598), .A0 (nx5129), .A1 (nx10517), .A2 (nx10527)) ;
    nor02_2x ix5140 (.Y (nx5139), .A0 (nx3594), .A1 (nx3592)) ;
    nor03_2x ix3595 (.Y (nx3594), .A0 (nx5143), .A1 (nx9579), .A2 (nx10535)) ;
    dffr gen_9_cmp_mRegCmp_reg_Q_4 (.Q (gen_9_cmp_mReg_4), .QB (nx5143), .D (
         window_9__4), .CLK (start), .R (rst)) ;
    nor03_2x ix3593 (.Y (nx3592), .A0 (gen_9_cmp_mReg_4), .A1 (nx10053), .A2 (
             nx10543)) ;
    nand02 ix3629 (.Y (gen_9_cmp_BSCmp_op2_5), .A0 (nx5147), .A1 (nx5153)) ;
    nor02_2x ix5148 (.Y (nx5147), .A0 (nx3624), .A1 (nx3620)) ;
    nor03_2x ix3625 (.Y (nx3624), .A0 (gen_9_cmp_mReg_4), .A1 (nx9585), .A2 (
             nx10511)) ;
    nor03_2x ix3621 (.Y (nx3620), .A0 (nx5143), .A1 (nx10517), .A2 (nx10527)) ;
    nor02_2x ix5154 (.Y (nx5153), .A0 (nx3616), .A1 (nx3614)) ;
    nor03_2x ix3617 (.Y (nx3616), .A0 (nx5156), .A1 (nx9581), .A2 (nx10535)) ;
    dffr gen_9_cmp_mRegCmp_reg_Q_5 (.Q (gen_9_cmp_mReg_5), .QB (nx5156), .D (
         window_9__5), .CLK (start), .R (rst)) ;
    nor03_2x ix3615 (.Y (nx3614), .A0 (gen_9_cmp_mReg_5), .A1 (nx10053), .A2 (
             nx10543)) ;
    nand02 ix3651 (.Y (gen_9_cmp_BSCmp_op2_6), .A0 (nx5163), .A1 (nx5169)) ;
    nor02_2x ix5164 (.Y (nx5163), .A0 (nx3646), .A1 (nx3642)) ;
    nor03_2x ix3647 (.Y (nx3646), .A0 (gen_9_cmp_mReg_5), .A1 (nx9587), .A2 (
             nx10511)) ;
    nor03_2x ix3643 (.Y (nx3642), .A0 (nx5156), .A1 (nx10517), .A2 (nx10527)) ;
    nor02_2x ix5170 (.Y (nx5169), .A0 (nx3638), .A1 (nx3636)) ;
    nor03_2x ix3639 (.Y (nx3638), .A0 (nx5173), .A1 (nx9581), .A2 (nx10535)) ;
    dffr gen_9_cmp_mRegCmp_reg_Q_6 (.Q (gen_9_cmp_mReg_6), .QB (nx5173), .D (
         window_9__6), .CLK (start), .R (rst)) ;
    nor03_2x ix3637 (.Y (nx3636), .A0 (gen_9_cmp_mReg_6), .A1 (nx10053), .A2 (
             nx10543)) ;
    nand02 ix3673 (.Y (gen_9_cmp_BSCmp_op2_7), .A0 (nx5177), .A1 (nx5183)) ;
    nor02_2x ix5178 (.Y (nx5177), .A0 (nx3668), .A1 (nx3664)) ;
    nor03_2x ix3669 (.Y (nx3668), .A0 (gen_9_cmp_mReg_6), .A1 (nx9587), .A2 (
             nx10513)) ;
    nor03_2x ix3665 (.Y (nx3664), .A0 (nx5173), .A1 (nx10519), .A2 (nx10529)) ;
    nor02_2x ix5184 (.Y (nx5183), .A0 (nx3660), .A1 (nx3658)) ;
    nor03_2x ix3661 (.Y (nx3660), .A0 (nx5187), .A1 (nx9581), .A2 (nx10537)) ;
    dffr gen_9_cmp_mRegCmp_reg_Q_7 (.Q (gen_9_cmp_mReg_7), .QB (nx5187), .D (
         window_9__7), .CLK (start), .R (rst)) ;
    nor03_2x ix3659 (.Y (nx3658), .A0 (gen_9_cmp_mReg_7), .A1 (nx10053), .A2 (
             nx10545)) ;
    nand02 ix3695 (.Y (gen_9_cmp_BSCmp_op2_8), .A0 (nx5191), .A1 (nx5197)) ;
    nor02_2x ix5192 (.Y (nx5191), .A0 (nx3690), .A1 (nx3686)) ;
    nor03_2x ix3691 (.Y (nx3690), .A0 (gen_9_cmp_mReg_7), .A1 (nx9587), .A2 (
             nx10513)) ;
    nor03_2x ix3687 (.Y (nx3686), .A0 (nx5187), .A1 (nx10519), .A2 (nx10529)) ;
    nor02_2x ix5198 (.Y (nx5197), .A0 (nx3682), .A1 (nx3680)) ;
    nor03_2x ix3683 (.Y (nx3682), .A0 (nx5200), .A1 (nx9581), .A2 (nx10537)) ;
    dffr gen_9_cmp_mRegCmp_reg_Q_8 (.Q (gen_9_cmp_mReg_8), .QB (nx5200), .D (
         window_9__8), .CLK (start), .R (rst)) ;
    nor03_2x ix3681 (.Y (nx3680), .A0 (gen_9_cmp_mReg_8), .A1 (nx10055), .A2 (
             nx10545)) ;
    nand02 ix3717 (.Y (gen_9_cmp_BSCmp_op2_9), .A0 (nx5207), .A1 (nx5213)) ;
    nor02_2x ix5208 (.Y (nx5207), .A0 (nx3712), .A1 (nx3708)) ;
    nor03_2x ix3713 (.Y (nx3712), .A0 (gen_9_cmp_mReg_8), .A1 (nx9587), .A2 (
             nx10513)) ;
    nor03_2x ix3709 (.Y (nx3708), .A0 (nx5200), .A1 (nx10519), .A2 (nx10529)) ;
    nor02_2x ix5214 (.Y (nx5213), .A0 (nx3704), .A1 (nx3702)) ;
    nor03_2x ix3705 (.Y (nx3704), .A0 (nx5217), .A1 (nx9581), .A2 (nx10537)) ;
    dffr gen_9_cmp_mRegCmp_reg_Q_9 (.Q (gen_9_cmp_mReg_9), .QB (nx5217), .D (
         window_9__9), .CLK (start), .R (rst)) ;
    nor03_2x ix3703 (.Y (nx3702), .A0 (gen_9_cmp_mReg_9), .A1 (nx10055), .A2 (
             nx10545)) ;
    nand02 ix3739 (.Y (gen_9_cmp_BSCmp_op2_10), .A0 (nx5221), .A1 (nx5227)) ;
    nor02_2x ix5222 (.Y (nx5221), .A0 (nx3734), .A1 (nx3730)) ;
    nor03_2x ix3735 (.Y (nx3734), .A0 (gen_9_cmp_mReg_9), .A1 (nx9587), .A2 (
             nx10513)) ;
    nor03_2x ix3731 (.Y (nx3730), .A0 (nx5217), .A1 (nx10519), .A2 (nx10529)) ;
    nor02_2x ix5228 (.Y (nx5227), .A0 (nx3726), .A1 (nx3724)) ;
    nor03_2x ix3727 (.Y (nx3726), .A0 (nx5231), .A1 (nx9581), .A2 (nx10537)) ;
    dffr gen_9_cmp_mRegCmp_reg_Q_10 (.Q (gen_9_cmp_mReg_10), .QB (nx5231), .D (
         window_9__10), .CLK (start), .R (rst)) ;
    nor03_2x ix3725 (.Y (nx3724), .A0 (gen_9_cmp_mReg_10), .A1 (nx10055), .A2 (
             nx10545)) ;
    nand02 ix3761 (.Y (gen_9_cmp_BSCmp_op2_11), .A0 (nx5235), .A1 (nx5241)) ;
    nor02_2x ix5236 (.Y (nx5235), .A0 (nx3756), .A1 (nx3752)) ;
    nor03_2x ix3757 (.Y (nx3756), .A0 (gen_9_cmp_mReg_10), .A1 (nx9587), .A2 (
             nx10513)) ;
    nor03_2x ix3753 (.Y (nx3752), .A0 (nx5231), .A1 (nx10519), .A2 (nx10529)) ;
    nor02_2x ix5242 (.Y (nx5241), .A0 (nx3748), .A1 (nx3746)) ;
    nor03_2x ix3749 (.Y (nx3748), .A0 (nx5244), .A1 (nx9581), .A2 (nx10537)) ;
    dffr gen_9_cmp_mRegCmp_reg_Q_11 (.Q (gen_9_cmp_mReg_11), .QB (nx5244), .D (
         window_9__11), .CLK (start), .R (rst)) ;
    nor03_2x ix3747 (.Y (nx3746), .A0 (gen_9_cmp_mReg_11), .A1 (nx10055), .A2 (
             nx10545)) ;
    nand02 ix3783 (.Y (gen_9_cmp_BSCmp_op2_12), .A0 (nx5251), .A1 (nx5257)) ;
    nor02_2x ix5252 (.Y (nx5251), .A0 (nx3778), .A1 (nx3774)) ;
    nor03_2x ix3779 (.Y (nx3778), .A0 (gen_9_cmp_mReg_11), .A1 (nx9587), .A2 (
             nx10513)) ;
    nor03_2x ix3775 (.Y (nx3774), .A0 (nx5244), .A1 (nx10519), .A2 (nx10529)) ;
    nor02_2x ix5258 (.Y (nx5257), .A0 (nx3770), .A1 (nx3768)) ;
    nor03_2x ix3771 (.Y (nx3770), .A0 (nx5261), .A1 (nx9583), .A2 (nx10537)) ;
    dffr gen_9_cmp_mRegCmp_reg_Q_12 (.Q (gen_9_cmp_mReg_12), .QB (nx5261), .D (
         window_9__12), .CLK (start), .R (rst)) ;
    nor03_2x ix3769 (.Y (nx3768), .A0 (gen_9_cmp_mReg_12), .A1 (nx10055), .A2 (
             nx10545)) ;
    nand02 ix3805 (.Y (gen_9_cmp_BSCmp_op2_13), .A0 (nx5265), .A1 (nx5271)) ;
    nor02_2x ix5266 (.Y (nx5265), .A0 (nx3800), .A1 (nx3796)) ;
    nor03_2x ix3801 (.Y (nx3800), .A0 (gen_9_cmp_mReg_12), .A1 (nx9589), .A2 (
             nx10515)) ;
    nor03_2x ix3797 (.Y (nx3796), .A0 (nx5261), .A1 (nx10519), .A2 (nx10531)) ;
    nor02_2x ix5272 (.Y (nx5271), .A0 (nx3792), .A1 (nx3790)) ;
    nor03_2x ix3793 (.Y (nx3792), .A0 (nx5275), .A1 (nx9583), .A2 (nx10539)) ;
    dffr gen_9_cmp_mRegCmp_reg_Q_13 (.Q (gen_9_cmp_mReg_13), .QB (nx5275), .D (
         window_9__13), .CLK (start), .R (rst)) ;
    nor03_2x ix3791 (.Y (nx3790), .A0 (gen_9_cmp_mReg_13), .A1 (nx10055), .A2 (
             nx10547)) ;
    nand02 ix3827 (.Y (gen_9_cmp_BSCmp_op2_14), .A0 (nx5279), .A1 (nx5285)) ;
    nor02_2x ix5280 (.Y (nx5279), .A0 (nx3822), .A1 (nx3818)) ;
    nor03_2x ix3823 (.Y (nx3822), .A0 (gen_9_cmp_mReg_13), .A1 (nx9589), .A2 (
             nx10515)) ;
    nor03_2x ix3819 (.Y (nx3818), .A0 (nx5275), .A1 (nx10521), .A2 (nx10531)) ;
    nor02_2x ix5286 (.Y (nx5285), .A0 (nx3814), .A1 (nx3812)) ;
    nor03_2x ix3815 (.Y (nx3814), .A0 (nx5288), .A1 (nx9583), .A2 (nx10539)) ;
    dffr gen_9_cmp_mRegCmp_reg_Q_14 (.Q (gen_9_cmp_mReg_14), .QB (nx5288), .D (
         window_9__14), .CLK (start), .R (rst)) ;
    nor03_2x ix3813 (.Y (nx3812), .A0 (gen_9_cmp_mReg_14), .A1 (nx10055), .A2 (
             nx10547)) ;
    nand02 ix3849 (.Y (gen_9_cmp_BSCmp_op2_15), .A0 (nx5295), .A1 (nx5301)) ;
    nor02_2x ix5296 (.Y (nx5295), .A0 (nx3844), .A1 (nx3840)) ;
    nor03_2x ix3845 (.Y (nx3844), .A0 (gen_9_cmp_mReg_14), .A1 (nx9589), .A2 (
             nx10515)) ;
    nor03_2x ix3841 (.Y (nx3840), .A0 (nx5288), .A1 (nx10521), .A2 (nx10531)) ;
    nor02_2x ix5302 (.Y (nx5301), .A0 (nx3836), .A1 (nx3834)) ;
    nor03_2x ix3837 (.Y (nx3836), .A0 (nx5305), .A1 (nx9583), .A2 (nx10539)) ;
    dffr gen_9_cmp_mRegCmp_reg_Q_15 (.Q (gen_9_cmp_mReg_15), .QB (nx5305), .D (
         window_9__15), .CLK (start), .R (rst)) ;
    nor03_2x ix3835 (.Y (nx3834), .A0 (gen_9_cmp_mReg_15), .A1 (nx10057), .A2 (
             nx10547)) ;
    nand02 ix3859 (.Y (gen_9_cmp_BSCmp_op2_16), .A0 (nx5309), .A1 (nx5301)) ;
    nor02_2x ix5310 (.Y (nx5309), .A0 (nx3854), .A1 (nx3850)) ;
    nor03_2x ix3855 (.Y (nx3854), .A0 (gen_9_cmp_mReg_15), .A1 (nx9589), .A2 (
             nx10515)) ;
    nor03_2x ix3851 (.Y (nx3850), .A0 (nx5305), .A1 (nx10521), .A2 (nx10531)) ;
    nand02 ix3927 (.Y (gen_10_cmp_BSCmp_op2_1), .A0 (nx5317), .A1 (nx5337)) ;
    nor02_2x ix5318 (.Y (nx5317), .A0 (nx3922), .A1 (nx3918)) ;
    nor03_2x ix3923 (.Y (nx3922), .A0 (gen_10_cmp_mReg_0), .A1 (nx9573), .A2 (
             nx10551)) ;
    dffr gen_10_cmp_mRegCmp_reg_Q_0 (.Q (gen_10_cmp_mReg_0), .QB (nx5323), .D (
         window_10__0), .CLK (start), .R (rst)) ;
    inv01 ix5328 (.Y (nx5327), .A (gen_10_cmp_pMux_0)) ;
    nor03_2x ix3919 (.Y (nx3918), .A0 (nx5323), .A1 (nx10557), .A2 (nx10567)) ;
    inv02 ix5336 (.Y (nx5335), .A (gen_10_cmp_pMux_2)) ;
    nor02_2x ix5338 (.Y (nx5337), .A0 (nx3908), .A1 (nx3906)) ;
    nor03_2x ix3909 (.Y (nx3908), .A0 (nx5341), .A1 (nx9567), .A2 (nx10575)) ;
    dffr gen_10_cmp_mRegCmp_reg_Q_1 (.Q (gen_10_cmp_mReg_1), .QB (nx5341), .D (
         window_10__1), .CLK (start), .R (rst)) ;
    nor03_2x ix3907 (.Y (nx3906), .A0 (gen_10_cmp_mReg_1), .A1 (nx10059), .A2 (
             nx10583)) ;
    nor03_2x ix3867 (.Y (nx3866), .A0 (nx9573), .A1 (nx5335), .A2 (
             gen_10_cmp_pMux_0)) ;
    nand02 ix3949 (.Y (gen_10_cmp_BSCmp_op2_2), .A0 (nx5352), .A1 (nx5357)) ;
    nor02_2x ix5353 (.Y (nx5352), .A0 (nx3944), .A1 (nx3940)) ;
    nor03_2x ix3945 (.Y (nx3944), .A0 (gen_10_cmp_mReg_1), .A1 (nx9573), .A2 (
             nx10551)) ;
    nor03_2x ix3941 (.Y (nx3940), .A0 (nx5341), .A1 (nx10557), .A2 (nx10567)) ;
    nor02_2x ix5358 (.Y (nx5357), .A0 (nx3936), .A1 (nx3934)) ;
    nor03_2x ix3937 (.Y (nx3936), .A0 (nx5361), .A1 (nx9567), .A2 (nx10575)) ;
    dffr gen_10_cmp_mRegCmp_reg_Q_2 (.Q (gen_10_cmp_mReg_2), .QB (nx5361), .D (
         window_10__2), .CLK (start), .R (rst)) ;
    nor03_2x ix3935 (.Y (nx3934), .A0 (gen_10_cmp_mReg_2), .A1 (nx10059), .A2 (
             nx10583)) ;
    nand02 ix3971 (.Y (gen_10_cmp_BSCmp_op2_3), .A0 (nx5367), .A1 (nx5373)) ;
    nor02_2x ix5368 (.Y (nx5367), .A0 (nx3966), .A1 (nx3962)) ;
    nor03_2x ix3967 (.Y (nx3966), .A0 (gen_10_cmp_mReg_2), .A1 (nx9573), .A2 (
             nx10551)) ;
    nor03_2x ix3963 (.Y (nx3962), .A0 (nx5361), .A1 (nx10557), .A2 (nx10567)) ;
    nor02_2x ix5374 (.Y (nx5373), .A0 (nx3958), .A1 (nx3956)) ;
    nor03_2x ix3959 (.Y (nx3958), .A0 (nx5376), .A1 (nx9567), .A2 (nx10575)) ;
    dffr gen_10_cmp_mRegCmp_reg_Q_3 (.Q (gen_10_cmp_mReg_3), .QB (nx5376), .D (
         window_10__3), .CLK (start), .R (rst)) ;
    nor03_2x ix3957 (.Y (nx3956), .A0 (gen_10_cmp_mReg_3), .A1 (nx10059), .A2 (
             nx10583)) ;
    nand02 ix3993 (.Y (gen_10_cmp_BSCmp_op2_4), .A0 (nx5383), .A1 (nx5389)) ;
    nor02_2x ix5384 (.Y (nx5383), .A0 (nx3988), .A1 (nx3984)) ;
    nor03_2x ix3989 (.Y (nx3988), .A0 (gen_10_cmp_mReg_3), .A1 (nx9573), .A2 (
             nx10551)) ;
    nor03_2x ix3985 (.Y (nx3984), .A0 (nx5376), .A1 (nx10557), .A2 (nx10567)) ;
    nor02_2x ix5390 (.Y (nx5389), .A0 (nx3980), .A1 (nx3978)) ;
    nor03_2x ix3981 (.Y (nx3980), .A0 (nx5393), .A1 (nx9567), .A2 (nx10575)) ;
    dffr gen_10_cmp_mRegCmp_reg_Q_4 (.Q (gen_10_cmp_mReg_4), .QB (nx5393), .D (
         window_10__4), .CLK (start), .R (rst)) ;
    nor03_2x ix3979 (.Y (nx3978), .A0 (gen_10_cmp_mReg_4), .A1 (nx10059), .A2 (
             nx10583)) ;
    nand02 ix4015 (.Y (gen_10_cmp_BSCmp_op2_5), .A0 (nx5399), .A1 (nx5405)) ;
    nor02_2x ix5400 (.Y (nx5399), .A0 (nx4010), .A1 (nx4006)) ;
    nor03_2x ix4011 (.Y (nx4010), .A0 (gen_10_cmp_mReg_4), .A1 (nx9573), .A2 (
             nx10551)) ;
    nor03_2x ix4007 (.Y (nx4006), .A0 (nx5393), .A1 (nx10557), .A2 (nx10567)) ;
    nor02_2x ix5406 (.Y (nx5405), .A0 (nx4002), .A1 (nx4000)) ;
    nor03_2x ix4003 (.Y (nx4002), .A0 (nx5409), .A1 (nx9569), .A2 (nx10575)) ;
    dffr gen_10_cmp_mRegCmp_reg_Q_5 (.Q (gen_10_cmp_mReg_5), .QB (nx5409), .D (
         window_10__5), .CLK (start), .R (rst)) ;
    nor03_2x ix4001 (.Y (nx4000), .A0 (gen_10_cmp_mReg_5), .A1 (nx10059), .A2 (
             nx10583)) ;
    nand02 ix4037 (.Y (gen_10_cmp_BSCmp_op2_6), .A0 (nx5414), .A1 (nx5418)) ;
    nor02_2x ix5415 (.Y (nx5414), .A0 (nx4032), .A1 (nx4028)) ;
    nor03_2x ix4033 (.Y (nx4032), .A0 (gen_10_cmp_mReg_5), .A1 (nx9575), .A2 (
             nx10551)) ;
    nor03_2x ix4029 (.Y (nx4028), .A0 (nx5409), .A1 (nx10557), .A2 (nx10567)) ;
    nor02_2x ix5419 (.Y (nx5418), .A0 (nx4024), .A1 (nx4022)) ;
    nor03_2x ix4025 (.Y (nx4024), .A0 (nx5421), .A1 (nx9569), .A2 (nx10575)) ;
    dffr gen_10_cmp_mRegCmp_reg_Q_6 (.Q (gen_10_cmp_mReg_6), .QB (nx5421), .D (
         window_10__6), .CLK (start), .R (rst)) ;
    nor03_2x ix4023 (.Y (nx4022), .A0 (gen_10_cmp_mReg_6), .A1 (nx10059), .A2 (
             nx10583)) ;
    nand02 ix4059 (.Y (gen_10_cmp_BSCmp_op2_7), .A0 (nx5427), .A1 (nx5433)) ;
    nor02_2x ix5428 (.Y (nx5427), .A0 (nx4054), .A1 (nx4050)) ;
    nor03_2x ix4055 (.Y (nx4054), .A0 (gen_10_cmp_mReg_6), .A1 (nx9575), .A2 (
             nx10553)) ;
    nor03_2x ix4051 (.Y (nx4050), .A0 (nx5421), .A1 (nx10559), .A2 (nx10569)) ;
    nor02_2x ix5434 (.Y (nx5433), .A0 (nx4046), .A1 (nx4044)) ;
    nor03_2x ix4047 (.Y (nx4046), .A0 (nx5437), .A1 (nx9569), .A2 (nx10577)) ;
    dffr gen_10_cmp_mRegCmp_reg_Q_7 (.Q (gen_10_cmp_mReg_7), .QB (nx5437), .D (
         window_10__7), .CLK (start), .R (rst)) ;
    nor03_2x ix4045 (.Y (nx4044), .A0 (gen_10_cmp_mReg_7), .A1 (nx10059), .A2 (
             nx10585)) ;
    nand02 ix4081 (.Y (gen_10_cmp_BSCmp_op2_8), .A0 (nx5443), .A1 (nx5447)) ;
    nor02_2x ix5444 (.Y (nx5443), .A0 (nx4076), .A1 (nx4072)) ;
    nor03_2x ix4077 (.Y (nx4076), .A0 (gen_10_cmp_mReg_7), .A1 (nx9575), .A2 (
             nx10553)) ;
    nor03_2x ix4073 (.Y (nx4072), .A0 (nx5437), .A1 (nx10559), .A2 (nx10569)) ;
    nor02_2x ix5448 (.Y (nx5447), .A0 (nx4068), .A1 (nx4066)) ;
    nor03_2x ix4069 (.Y (nx4068), .A0 (nx5451), .A1 (nx9569), .A2 (nx10577)) ;
    dffr gen_10_cmp_mRegCmp_reg_Q_8 (.Q (gen_10_cmp_mReg_8), .QB (nx5451), .D (
         window_10__8), .CLK (start), .R (rst)) ;
    nor03_2x ix4067 (.Y (nx4066), .A0 (gen_10_cmp_mReg_8), .A1 (nx10061), .A2 (
             nx10585)) ;
    nand02 ix4103 (.Y (gen_10_cmp_BSCmp_op2_9), .A0 (nx5457), .A1 (nx5463)) ;
    nor02_2x ix5458 (.Y (nx5457), .A0 (nx4098), .A1 (nx4094)) ;
    nor03_2x ix4099 (.Y (nx4098), .A0 (gen_10_cmp_mReg_8), .A1 (nx9575), .A2 (
             nx10553)) ;
    nor03_2x ix4095 (.Y (nx4094), .A0 (nx5451), .A1 (nx10559), .A2 (nx10569)) ;
    nor02_2x ix5464 (.Y (nx5463), .A0 (nx4090), .A1 (nx4088)) ;
    nor03_2x ix4091 (.Y (nx4090), .A0 (nx5467), .A1 (nx9569), .A2 (nx10577)) ;
    dffr gen_10_cmp_mRegCmp_reg_Q_9 (.Q (gen_10_cmp_mReg_9), .QB (nx5467), .D (
         window_10__9), .CLK (start), .R (rst)) ;
    nor03_2x ix4089 (.Y (nx4088), .A0 (gen_10_cmp_mReg_9), .A1 (nx10061), .A2 (
             nx10585)) ;
    nand02 ix4125 (.Y (gen_10_cmp_BSCmp_op2_10), .A0 (nx5473), .A1 (nx5477)) ;
    nor02_2x ix5474 (.Y (nx5473), .A0 (nx4120), .A1 (nx4116)) ;
    nor03_2x ix4121 (.Y (nx4120), .A0 (gen_10_cmp_mReg_9), .A1 (nx9575), .A2 (
             nx10553)) ;
    nor03_2x ix4117 (.Y (nx4116), .A0 (nx5467), .A1 (nx10559), .A2 (nx10569)) ;
    nor02_2x ix5478 (.Y (nx5477), .A0 (nx4112), .A1 (nx4110)) ;
    nor03_2x ix4113 (.Y (nx4112), .A0 (nx5481), .A1 (nx9569), .A2 (nx10577)) ;
    dffr gen_10_cmp_mRegCmp_reg_Q_10 (.Q (gen_10_cmp_mReg_10), .QB (nx5481), .D (
         window_10__10), .CLK (start), .R (rst)) ;
    nor03_2x ix4111 (.Y (nx4110), .A0 (gen_10_cmp_mReg_10), .A1 (nx10061), .A2 (
             nx10585)) ;
    nand02 ix4147 (.Y (gen_10_cmp_BSCmp_op2_11), .A0 (nx5487), .A1 (nx5493)) ;
    nor02_2x ix5488 (.Y (nx5487), .A0 (nx4142), .A1 (nx4138)) ;
    nor03_2x ix4143 (.Y (nx4142), .A0 (gen_10_cmp_mReg_10), .A1 (nx9575), .A2 (
             nx10553)) ;
    nor03_2x ix4139 (.Y (nx4138), .A0 (nx5481), .A1 (nx10559), .A2 (nx10569)) ;
    nor02_2x ix5494 (.Y (nx5493), .A0 (nx4134), .A1 (nx4132)) ;
    nor03_2x ix4135 (.Y (nx4134), .A0 (nx5496), .A1 (nx9569), .A2 (nx10577)) ;
    dffr gen_10_cmp_mRegCmp_reg_Q_11 (.Q (gen_10_cmp_mReg_11), .QB (nx5496), .D (
         window_10__11), .CLK (start), .R (rst)) ;
    nor03_2x ix4133 (.Y (nx4132), .A0 (gen_10_cmp_mReg_11), .A1 (nx10061), .A2 (
             nx10585)) ;
    nand02 ix4169 (.Y (gen_10_cmp_BSCmp_op2_12), .A0 (nx5501), .A1 (nx5507)) ;
    nor02_2x ix5502 (.Y (nx5501), .A0 (nx4164), .A1 (nx4160)) ;
    nor03_2x ix4165 (.Y (nx4164), .A0 (gen_10_cmp_mReg_11), .A1 (nx9575), .A2 (
             nx10553)) ;
    nor03_2x ix4161 (.Y (nx4160), .A0 (nx5496), .A1 (nx10559), .A2 (nx10569)) ;
    nor02_2x ix5508 (.Y (nx5507), .A0 (nx4156), .A1 (nx4154)) ;
    nor03_2x ix4157 (.Y (nx4156), .A0 (nx5511), .A1 (nx9571), .A2 (nx10577)) ;
    dffr gen_10_cmp_mRegCmp_reg_Q_12 (.Q (gen_10_cmp_mReg_12), .QB (nx5511), .D (
         window_10__12), .CLK (start), .R (rst)) ;
    nor03_2x ix4155 (.Y (nx4154), .A0 (gen_10_cmp_mReg_12), .A1 (nx10061), .A2 (
             nx10585)) ;
    nand02 ix4191 (.Y (gen_10_cmp_BSCmp_op2_13), .A0 (nx5517), .A1 (nx5521)) ;
    nor02_2x ix5518 (.Y (nx5517), .A0 (nx4186), .A1 (nx4182)) ;
    nor03_2x ix4187 (.Y (nx4186), .A0 (gen_10_cmp_mReg_12), .A1 (nx9577), .A2 (
             nx10555)) ;
    nor03_2x ix4183 (.Y (nx4182), .A0 (nx5511), .A1 (nx10559), .A2 (nx10571)) ;
    nor02_2x ix5522 (.Y (nx5521), .A0 (nx4178), .A1 (nx4176)) ;
    nor03_2x ix4179 (.Y (nx4178), .A0 (nx5525), .A1 (nx9571), .A2 (nx10579)) ;
    dffr gen_10_cmp_mRegCmp_reg_Q_13 (.Q (gen_10_cmp_mReg_13), .QB (nx5525), .D (
         window_10__13), .CLK (start), .R (rst)) ;
    nor03_2x ix4177 (.Y (nx4176), .A0 (gen_10_cmp_mReg_13), .A1 (nx10061), .A2 (
             nx10587)) ;
    nand02 ix4213 (.Y (gen_10_cmp_BSCmp_op2_14), .A0 (nx5531), .A1 (nx5537)) ;
    nor02_2x ix5532 (.Y (nx5531), .A0 (nx4208), .A1 (nx4204)) ;
    nor03_2x ix4209 (.Y (nx4208), .A0 (gen_10_cmp_mReg_13), .A1 (nx9577), .A2 (
             nx10555)) ;
    nor03_2x ix4205 (.Y (nx4204), .A0 (nx5525), .A1 (nx10561), .A2 (nx10571)) ;
    nor02_2x ix5538 (.Y (nx5537), .A0 (nx4200), .A1 (nx4198)) ;
    nor03_2x ix4201 (.Y (nx4200), .A0 (nx5540), .A1 (nx9571), .A2 (nx10579)) ;
    dffr gen_10_cmp_mRegCmp_reg_Q_14 (.Q (gen_10_cmp_mReg_14), .QB (nx5540), .D (
         window_10__14), .CLK (start), .R (rst)) ;
    nor03_2x ix4199 (.Y (nx4198), .A0 (gen_10_cmp_mReg_14), .A1 (nx10061), .A2 (
             nx10587)) ;
    nand02 ix4235 (.Y (gen_10_cmp_BSCmp_op2_15), .A0 (nx5545), .A1 (nx5551)) ;
    nor02_2x ix5546 (.Y (nx5545), .A0 (nx4230), .A1 (nx4226)) ;
    nor03_2x ix4231 (.Y (nx4230), .A0 (gen_10_cmp_mReg_14), .A1 (nx9577), .A2 (
             nx10555)) ;
    nor03_2x ix4227 (.Y (nx4226), .A0 (nx5540), .A1 (nx10561), .A2 (nx10571)) ;
    nor02_2x ix5552 (.Y (nx5551), .A0 (nx4222), .A1 (nx4220)) ;
    nor03_2x ix4223 (.Y (nx4222), .A0 (nx5555), .A1 (nx9571), .A2 (nx10579)) ;
    dffr gen_10_cmp_mRegCmp_reg_Q_15 (.Q (gen_10_cmp_mReg_15), .QB (nx5555), .D (
         window_10__15), .CLK (start), .R (rst)) ;
    nor03_2x ix4221 (.Y (nx4220), .A0 (gen_10_cmp_mReg_15), .A1 (nx10063), .A2 (
             nx10587)) ;
    nand02 ix4245 (.Y (gen_10_cmp_BSCmp_op2_16), .A0 (nx5561), .A1 (nx5551)) ;
    nor02_2x ix5562 (.Y (nx5561), .A0 (nx4240), .A1 (nx4236)) ;
    nor03_2x ix4241 (.Y (nx4240), .A0 (gen_10_cmp_mReg_15), .A1 (nx9577), .A2 (
             nx10555)) ;
    nor03_2x ix4237 (.Y (nx4236), .A0 (nx5555), .A1 (nx10561), .A2 (nx10571)) ;
    nand02 ix4313 (.Y (gen_11_cmp_BSCmp_op2_1), .A0 (nx5567), .A1 (nx5587)) ;
    nor02_2x ix5568 (.Y (nx5567), .A0 (nx4308), .A1 (nx4304)) ;
    nor03_2x ix4309 (.Y (nx4308), .A0 (gen_11_cmp_mReg_0), .A1 (nx9561), .A2 (
             nx10591)) ;
    dffr gen_11_cmp_mRegCmp_reg_Q_0 (.Q (gen_11_cmp_mReg_0), .QB (nx5573), .D (
         window_11__0), .CLK (start), .R (rst)) ;
    inv01 ix5578 (.Y (nx5577), .A (gen_11_cmp_pMux_0)) ;
    nor03_2x ix4305 (.Y (nx4304), .A0 (nx5573), .A1 (nx10597), .A2 (nx10607)) ;
    inv02 ix5586 (.Y (nx5585), .A (gen_11_cmp_pMux_2)) ;
    nor02_2x ix5588 (.Y (nx5587), .A0 (nx4294), .A1 (nx4292)) ;
    nor03_2x ix4295 (.Y (nx4294), .A0 (nx5591), .A1 (nx9555), .A2 (nx10615)) ;
    dffr gen_11_cmp_mRegCmp_reg_Q_1 (.Q (gen_11_cmp_mReg_1), .QB (nx5591), .D (
         window_11__1), .CLK (start), .R (rst)) ;
    nor03_2x ix4293 (.Y (nx4292), .A0 (gen_11_cmp_mReg_1), .A1 (nx10065), .A2 (
             nx10623)) ;
    nor03_2x ix4253 (.Y (nx4252), .A0 (nx9561), .A1 (nx5585), .A2 (
             gen_11_cmp_pMux_0)) ;
    nand02 ix4335 (.Y (gen_11_cmp_BSCmp_op2_2), .A0 (nx5603), .A1 (nx5607)) ;
    nor02_2x ix5604 (.Y (nx5603), .A0 (nx4330), .A1 (nx4326)) ;
    nor03_2x ix4331 (.Y (nx4330), .A0 (gen_11_cmp_mReg_1), .A1 (nx9561), .A2 (
             nx10591)) ;
    nor03_2x ix4327 (.Y (nx4326), .A0 (nx5591), .A1 (nx10597), .A2 (nx10607)) ;
    nor02_2x ix5608 (.Y (nx5607), .A0 (nx4322), .A1 (nx4320)) ;
    nor03_2x ix4323 (.Y (nx4322), .A0 (nx5611), .A1 (nx9555), .A2 (nx10615)) ;
    dffr gen_11_cmp_mRegCmp_reg_Q_2 (.Q (gen_11_cmp_mReg_2), .QB (nx5611), .D (
         window_11__2), .CLK (start), .R (rst)) ;
    nor03_2x ix4321 (.Y (nx4320), .A0 (gen_11_cmp_mReg_2), .A1 (nx10065), .A2 (
             nx10623)) ;
    nand02 ix4357 (.Y (gen_11_cmp_BSCmp_op2_3), .A0 (nx5617), .A1 (nx5621)) ;
    nor02_2x ix5618 (.Y (nx5617), .A0 (nx4352), .A1 (nx4348)) ;
    nor03_2x ix4353 (.Y (nx4352), .A0 (gen_11_cmp_mReg_2), .A1 (nx9561), .A2 (
             nx10591)) ;
    nor03_2x ix4349 (.Y (nx4348), .A0 (nx5611), .A1 (nx10597), .A2 (nx10607)) ;
    nor02_2x ix5622 (.Y (nx5621), .A0 (nx4344), .A1 (nx4342)) ;
    nor03_2x ix4345 (.Y (nx4344), .A0 (nx5625), .A1 (nx9555), .A2 (nx10615)) ;
    dffr gen_11_cmp_mRegCmp_reg_Q_3 (.Q (gen_11_cmp_mReg_3), .QB (nx5625), .D (
         window_11__3), .CLK (start), .R (rst)) ;
    nor03_2x ix4343 (.Y (nx4342), .A0 (gen_11_cmp_mReg_3), .A1 (nx10065), .A2 (
             nx10623)) ;
    nand02 ix4379 (.Y (gen_11_cmp_BSCmp_op2_4), .A0 (nx5629), .A1 (nx5635)) ;
    nor02_2x ix5630 (.Y (nx5629), .A0 (nx4374), .A1 (nx4370)) ;
    nor03_2x ix4375 (.Y (nx4374), .A0 (gen_11_cmp_mReg_3), .A1 (nx9561), .A2 (
             nx10591)) ;
    nor03_2x ix4371 (.Y (nx4370), .A0 (nx5625), .A1 (nx10597), .A2 (nx10607)) ;
    nor02_2x ix5636 (.Y (nx5635), .A0 (nx4366), .A1 (nx4364)) ;
    nor03_2x ix4367 (.Y (nx4366), .A0 (nx5639), .A1 (nx9555), .A2 (nx10615)) ;
    dffr gen_11_cmp_mRegCmp_reg_Q_4 (.Q (gen_11_cmp_mReg_4), .QB (nx5639), .D (
         window_11__4), .CLK (start), .R (rst)) ;
    nor03_2x ix4365 (.Y (nx4364), .A0 (gen_11_cmp_mReg_4), .A1 (nx10065), .A2 (
             nx10623)) ;
    nand02 ix4401 (.Y (gen_11_cmp_BSCmp_op2_5), .A0 (nx5643), .A1 (nx5649)) ;
    nor02_2x ix5644 (.Y (nx5643), .A0 (nx4396), .A1 (nx4392)) ;
    nor03_2x ix4397 (.Y (nx4396), .A0 (gen_11_cmp_mReg_4), .A1 (nx9561), .A2 (
             nx10591)) ;
    nor03_2x ix4393 (.Y (nx4392), .A0 (nx5639), .A1 (nx10597), .A2 (nx10607)) ;
    nor02_2x ix5650 (.Y (nx5649), .A0 (nx4388), .A1 (nx4386)) ;
    nor03_2x ix4389 (.Y (nx4388), .A0 (nx5652), .A1 (nx9557), .A2 (nx10615)) ;
    dffr gen_11_cmp_mRegCmp_reg_Q_5 (.Q (gen_11_cmp_mReg_5), .QB (nx5652), .D (
         window_11__5), .CLK (start), .R (rst)) ;
    nor03_2x ix4387 (.Y (nx4386), .A0 (gen_11_cmp_mReg_5), .A1 (nx10065), .A2 (
             nx10623)) ;
    nand02 ix4423 (.Y (gen_11_cmp_BSCmp_op2_6), .A0 (nx5659), .A1 (nx5665)) ;
    nor02_2x ix5660 (.Y (nx5659), .A0 (nx4418), .A1 (nx4414)) ;
    nor03_2x ix4419 (.Y (nx4418), .A0 (gen_11_cmp_mReg_5), .A1 (nx9563), .A2 (
             nx10591)) ;
    nor03_2x ix4415 (.Y (nx4414), .A0 (nx5652), .A1 (nx10597), .A2 (nx10607)) ;
    nor02_2x ix5666 (.Y (nx5665), .A0 (nx4410), .A1 (nx4408)) ;
    nor03_2x ix4411 (.Y (nx4410), .A0 (nx5669), .A1 (nx9557), .A2 (nx10615)) ;
    dffr gen_11_cmp_mRegCmp_reg_Q_6 (.Q (gen_11_cmp_mReg_6), .QB (nx5669), .D (
         window_11__6), .CLK (start), .R (rst)) ;
    nor03_2x ix4409 (.Y (nx4408), .A0 (gen_11_cmp_mReg_6), .A1 (nx10065), .A2 (
             nx10623)) ;
    nand02 ix4445 (.Y (gen_11_cmp_BSCmp_op2_7), .A0 (nx5673), .A1 (nx5679)) ;
    nor02_2x ix5674 (.Y (nx5673), .A0 (nx4440), .A1 (nx4436)) ;
    nor03_2x ix4441 (.Y (nx4440), .A0 (gen_11_cmp_mReg_6), .A1 (nx9563), .A2 (
             nx10593)) ;
    nor03_2x ix4437 (.Y (nx4436), .A0 (nx5669), .A1 (nx10599), .A2 (nx10609)) ;
    nor02_2x ix5680 (.Y (nx5679), .A0 (nx4432), .A1 (nx4430)) ;
    nor03_2x ix4433 (.Y (nx4432), .A0 (nx5683), .A1 (nx9557), .A2 (nx10617)) ;
    dffr gen_11_cmp_mRegCmp_reg_Q_7 (.Q (gen_11_cmp_mReg_7), .QB (nx5683), .D (
         window_11__7), .CLK (start), .R (rst)) ;
    nor03_2x ix4431 (.Y (nx4430), .A0 (gen_11_cmp_mReg_7), .A1 (nx10065), .A2 (
             nx10625)) ;
    nand02 ix4467 (.Y (gen_11_cmp_BSCmp_op2_8), .A0 (nx5687), .A1 (nx5693)) ;
    nor02_2x ix5688 (.Y (nx5687), .A0 (nx4462), .A1 (nx4458)) ;
    nor03_2x ix4463 (.Y (nx4462), .A0 (gen_11_cmp_mReg_7), .A1 (nx9563), .A2 (
             nx10593)) ;
    nor03_2x ix4459 (.Y (nx4458), .A0 (nx5683), .A1 (nx10599), .A2 (nx10609)) ;
    nor02_2x ix5694 (.Y (nx5693), .A0 (nx4454), .A1 (nx4452)) ;
    nor03_2x ix4455 (.Y (nx4454), .A0 (nx5696), .A1 (nx9557), .A2 (nx10617)) ;
    dffr gen_11_cmp_mRegCmp_reg_Q_8 (.Q (gen_11_cmp_mReg_8), .QB (nx5696), .D (
         window_11__8), .CLK (start), .R (rst)) ;
    nor03_2x ix4453 (.Y (nx4452), .A0 (gen_11_cmp_mReg_8), .A1 (nx10067), .A2 (
             nx10625)) ;
    nand02 ix4489 (.Y (gen_11_cmp_BSCmp_op2_9), .A0 (nx5703), .A1 (nx5709)) ;
    nor02_2x ix5704 (.Y (nx5703), .A0 (nx4484), .A1 (nx4480)) ;
    nor03_2x ix4485 (.Y (nx4484), .A0 (gen_11_cmp_mReg_8), .A1 (nx9563), .A2 (
             nx10593)) ;
    nor03_2x ix4481 (.Y (nx4480), .A0 (nx5696), .A1 (nx10599), .A2 (nx10609)) ;
    nor02_2x ix5710 (.Y (nx5709), .A0 (nx4476), .A1 (nx4474)) ;
    nor03_2x ix4477 (.Y (nx4476), .A0 (nx5713), .A1 (nx9557), .A2 (nx10617)) ;
    dffr gen_11_cmp_mRegCmp_reg_Q_9 (.Q (gen_11_cmp_mReg_9), .QB (nx5713), .D (
         window_11__9), .CLK (start), .R (rst)) ;
    nor03_2x ix4475 (.Y (nx4474), .A0 (gen_11_cmp_mReg_9), .A1 (nx10067), .A2 (
             nx10625)) ;
    nand02 ix4511 (.Y (gen_11_cmp_BSCmp_op2_10), .A0 (nx5717), .A1 (nx5723)) ;
    nor02_2x ix5718 (.Y (nx5717), .A0 (nx4506), .A1 (nx4502)) ;
    nor03_2x ix4507 (.Y (nx4506), .A0 (gen_11_cmp_mReg_9), .A1 (nx9563), .A2 (
             nx10593)) ;
    nor03_2x ix4503 (.Y (nx4502), .A0 (nx5713), .A1 (nx10599), .A2 (nx10609)) ;
    nor02_2x ix5724 (.Y (nx5723), .A0 (nx4498), .A1 (nx4496)) ;
    nor03_2x ix4499 (.Y (nx4498), .A0 (nx5727), .A1 (nx9557), .A2 (nx10617)) ;
    dffr gen_11_cmp_mRegCmp_reg_Q_10 (.Q (gen_11_cmp_mReg_10), .QB (nx5727), .D (
         window_11__10), .CLK (start), .R (rst)) ;
    nor03_2x ix4497 (.Y (nx4496), .A0 (gen_11_cmp_mReg_10), .A1 (nx10067), .A2 (
             nx10625)) ;
    nand02 ix4533 (.Y (gen_11_cmp_BSCmp_op2_11), .A0 (nx5731), .A1 (nx5737)) ;
    nor02_2x ix5732 (.Y (nx5731), .A0 (nx4528), .A1 (nx4524)) ;
    nor03_2x ix4529 (.Y (nx4528), .A0 (gen_11_cmp_mReg_10), .A1 (nx9563), .A2 (
             nx10593)) ;
    nor03_2x ix4525 (.Y (nx4524), .A0 (nx5727), .A1 (nx10599), .A2 (nx10609)) ;
    nor02_2x ix5738 (.Y (nx5737), .A0 (nx4520), .A1 (nx4518)) ;
    nor03_2x ix4521 (.Y (nx4520), .A0 (nx5740), .A1 (nx9557), .A2 (nx10617)) ;
    dffr gen_11_cmp_mRegCmp_reg_Q_11 (.Q (gen_11_cmp_mReg_11), .QB (nx5740), .D (
         window_11__11), .CLK (start), .R (rst)) ;
    nor03_2x ix4519 (.Y (nx4518), .A0 (gen_11_cmp_mReg_11), .A1 (nx10067), .A2 (
             nx10625)) ;
    nand02 ix4555 (.Y (gen_11_cmp_BSCmp_op2_12), .A0 (nx5747), .A1 (nx5753)) ;
    nor02_2x ix5748 (.Y (nx5747), .A0 (nx4550), .A1 (nx4546)) ;
    nor03_2x ix4551 (.Y (nx4550), .A0 (gen_11_cmp_mReg_11), .A1 (nx9563), .A2 (
             nx10593)) ;
    nor03_2x ix4547 (.Y (nx4546), .A0 (nx5740), .A1 (nx10599), .A2 (nx10609)) ;
    nor02_2x ix5754 (.Y (nx5753), .A0 (nx4542), .A1 (nx4540)) ;
    nor03_2x ix4543 (.Y (nx4542), .A0 (nx5757), .A1 (nx9559), .A2 (nx10617)) ;
    dffr gen_11_cmp_mRegCmp_reg_Q_12 (.Q (gen_11_cmp_mReg_12), .QB (nx5757), .D (
         window_11__12), .CLK (start), .R (rst)) ;
    nor03_2x ix4541 (.Y (nx4540), .A0 (gen_11_cmp_mReg_12), .A1 (nx10067), .A2 (
             nx10625)) ;
    nand02 ix4577 (.Y (gen_11_cmp_BSCmp_op2_13), .A0 (nx5761), .A1 (nx5767)) ;
    nor02_2x ix5762 (.Y (nx5761), .A0 (nx4572), .A1 (nx4568)) ;
    nor03_2x ix4573 (.Y (nx4572), .A0 (gen_11_cmp_mReg_12), .A1 (nx9565), .A2 (
             nx10595)) ;
    nor03_2x ix4569 (.Y (nx4568), .A0 (nx5757), .A1 (nx10599), .A2 (nx10611)) ;
    nor02_2x ix5768 (.Y (nx5767), .A0 (nx4564), .A1 (nx4562)) ;
    nor03_2x ix4565 (.Y (nx4564), .A0 (nx5771), .A1 (nx9559), .A2 (nx10619)) ;
    dffr gen_11_cmp_mRegCmp_reg_Q_13 (.Q (gen_11_cmp_mReg_13), .QB (nx5771), .D (
         window_11__13), .CLK (start), .R (rst)) ;
    nor03_2x ix4563 (.Y (nx4562), .A0 (gen_11_cmp_mReg_13), .A1 (nx10067), .A2 (
             nx10627)) ;
    nand02 ix4599 (.Y (gen_11_cmp_BSCmp_op2_14), .A0 (nx5775), .A1 (nx5781)) ;
    nor02_2x ix5776 (.Y (nx5775), .A0 (nx4594), .A1 (nx4590)) ;
    nor03_2x ix4595 (.Y (nx4594), .A0 (gen_11_cmp_mReg_13), .A1 (nx9565), .A2 (
             nx10595)) ;
    nor03_2x ix4591 (.Y (nx4590), .A0 (nx5771), .A1 (nx10601), .A2 (nx10611)) ;
    nor02_2x ix5782 (.Y (nx5781), .A0 (nx4586), .A1 (nx4584)) ;
    nor03_2x ix4587 (.Y (nx4586), .A0 (nx5785), .A1 (nx9559), .A2 (nx10619)) ;
    dffr gen_11_cmp_mRegCmp_reg_Q_14 (.Q (gen_11_cmp_mReg_14), .QB (nx5785), .D (
         window_11__14), .CLK (start), .R (rst)) ;
    nor03_2x ix4585 (.Y (nx4584), .A0 (gen_11_cmp_mReg_14), .A1 (nx10067), .A2 (
             nx10627)) ;
    nand02 ix4621 (.Y (gen_11_cmp_BSCmp_op2_15), .A0 (nx5791), .A1 (nx5797)) ;
    nor02_2x ix5792 (.Y (nx5791), .A0 (nx4616), .A1 (nx4612)) ;
    nor03_2x ix4617 (.Y (nx4616), .A0 (gen_11_cmp_mReg_14), .A1 (nx9565), .A2 (
             nx10595)) ;
    nor03_2x ix4613 (.Y (nx4612), .A0 (nx5785), .A1 (nx10601), .A2 (nx10611)) ;
    nor02_2x ix5798 (.Y (nx5797), .A0 (nx4608), .A1 (nx4606)) ;
    nor03_2x ix4609 (.Y (nx4608), .A0 (nx5800), .A1 (nx9559), .A2 (nx10619)) ;
    dffr gen_11_cmp_mRegCmp_reg_Q_15 (.Q (gen_11_cmp_mReg_15), .QB (nx5800), .D (
         window_11__15), .CLK (start), .R (rst)) ;
    nor03_2x ix4607 (.Y (nx4606), .A0 (gen_11_cmp_mReg_15), .A1 (nx10069), .A2 (
             nx10627)) ;
    nand02 ix4631 (.Y (gen_11_cmp_BSCmp_op2_16), .A0 (nx5804), .A1 (nx5797)) ;
    nor02_2x ix5805 (.Y (nx5804), .A0 (nx4626), .A1 (nx4622)) ;
    nor03_2x ix4627 (.Y (nx4626), .A0 (gen_11_cmp_mReg_15), .A1 (nx9565), .A2 (
             nx10595)) ;
    nor03_2x ix4623 (.Y (nx4622), .A0 (nx5800), .A1 (nx10601), .A2 (nx10611)) ;
    nand02 ix4699 (.Y (gen_12_cmp_BSCmp_op2_1), .A0 (nx5811), .A1 (nx5831)) ;
    nor02_2x ix5812 (.Y (nx5811), .A0 (nx4694), .A1 (nx4690)) ;
    nor03_2x ix4695 (.Y (nx4694), .A0 (gen_12_cmp_mReg_0), .A1 (nx9549), .A2 (
             nx10631)) ;
    dffr gen_12_cmp_mRegCmp_reg_Q_0 (.Q (gen_12_cmp_mReg_0), .QB (nx5817), .D (
         window_12__0), .CLK (start), .R (rst)) ;
    inv01 ix5822 (.Y (nx5821), .A (gen_12_cmp_pMux_0)) ;
    nor03_2x ix4691 (.Y (nx4690), .A0 (nx5817), .A1 (nx10637), .A2 (nx10647)) ;
    inv02 ix5830 (.Y (nx5829), .A (gen_12_cmp_pMux_2)) ;
    nor02_2x ix5832 (.Y (nx5831), .A0 (nx4680), .A1 (nx4678)) ;
    nor03_2x ix4681 (.Y (nx4680), .A0 (nx5834), .A1 (nx9543), .A2 (nx10655)) ;
    dffr gen_12_cmp_mRegCmp_reg_Q_1 (.Q (gen_12_cmp_mReg_1), .QB (nx5834), .D (
         window_12__1), .CLK (start), .R (rst)) ;
    nor03_2x ix4679 (.Y (nx4678), .A0 (gen_12_cmp_mReg_1), .A1 (nx10071), .A2 (
             nx10663)) ;
    nor03_2x ix4639 (.Y (nx4638), .A0 (nx9549), .A1 (nx5829), .A2 (
             gen_12_cmp_pMux_0)) ;
    nand02 ix4721 (.Y (gen_12_cmp_BSCmp_op2_2), .A0 (nx5847), .A1 (nx5853)) ;
    nor02_2x ix5848 (.Y (nx5847), .A0 (nx4716), .A1 (nx4712)) ;
    nor03_2x ix4717 (.Y (nx4716), .A0 (gen_12_cmp_mReg_1), .A1 (nx9549), .A2 (
             nx10631)) ;
    nor03_2x ix4713 (.Y (nx4712), .A0 (nx5834), .A1 (nx10637), .A2 (nx10647)) ;
    nor02_2x ix5854 (.Y (nx5853), .A0 (nx4708), .A1 (nx4706)) ;
    nor03_2x ix4709 (.Y (nx4708), .A0 (nx5857), .A1 (nx9543), .A2 (nx10655)) ;
    dffr gen_12_cmp_mRegCmp_reg_Q_2 (.Q (gen_12_cmp_mReg_2), .QB (nx5857), .D (
         window_12__2), .CLK (start), .R (rst)) ;
    nor03_2x ix4707 (.Y (nx4706), .A0 (gen_12_cmp_mReg_2), .A1 (nx10071), .A2 (
             nx10663)) ;
    nand02 ix4743 (.Y (gen_12_cmp_BSCmp_op2_3), .A0 (nx5861), .A1 (nx5867)) ;
    nor02_2x ix5862 (.Y (nx5861), .A0 (nx4738), .A1 (nx4734)) ;
    nor03_2x ix4739 (.Y (nx4738), .A0 (gen_12_cmp_mReg_2), .A1 (nx9549), .A2 (
             nx10631)) ;
    nor03_2x ix4735 (.Y (nx4734), .A0 (nx5857), .A1 (nx10637), .A2 (nx10647)) ;
    nor02_2x ix5868 (.Y (nx5867), .A0 (nx4730), .A1 (nx4728)) ;
    nor03_2x ix4731 (.Y (nx4730), .A0 (nx5871), .A1 (nx9543), .A2 (nx10655)) ;
    dffr gen_12_cmp_mRegCmp_reg_Q_3 (.Q (gen_12_cmp_mReg_3), .QB (nx5871), .D (
         window_12__3), .CLK (start), .R (rst)) ;
    nor03_2x ix4729 (.Y (nx4728), .A0 (gen_12_cmp_mReg_3), .A1 (nx10071), .A2 (
             nx10663)) ;
    nand02 ix4765 (.Y (gen_12_cmp_BSCmp_op2_4), .A0 (nx5875), .A1 (nx5881)) ;
    nor02_2x ix5876 (.Y (nx5875), .A0 (nx4760), .A1 (nx4756)) ;
    nor03_2x ix4761 (.Y (nx4760), .A0 (gen_12_cmp_mReg_3), .A1 (nx9549), .A2 (
             nx10631)) ;
    nor03_2x ix4757 (.Y (nx4756), .A0 (nx5871), .A1 (nx10637), .A2 (nx10647)) ;
    nor02_2x ix5882 (.Y (nx5881), .A0 (nx4752), .A1 (nx4750)) ;
    nor03_2x ix4753 (.Y (nx4752), .A0 (nx5884), .A1 (nx9543), .A2 (nx10655)) ;
    dffr gen_12_cmp_mRegCmp_reg_Q_4 (.Q (gen_12_cmp_mReg_4), .QB (nx5884), .D (
         window_12__4), .CLK (start), .R (rst)) ;
    nor03_2x ix4751 (.Y (nx4750), .A0 (gen_12_cmp_mReg_4), .A1 (nx10071), .A2 (
             nx10663)) ;
    nand02 ix4787 (.Y (gen_12_cmp_BSCmp_op2_5), .A0 (nx5891), .A1 (nx5897)) ;
    nor02_2x ix5892 (.Y (nx5891), .A0 (nx4782), .A1 (nx4778)) ;
    nor03_2x ix4783 (.Y (nx4782), .A0 (gen_12_cmp_mReg_4), .A1 (nx9549), .A2 (
             nx10631)) ;
    nor03_2x ix4779 (.Y (nx4778), .A0 (nx5884), .A1 (nx10637), .A2 (nx10647)) ;
    nor02_2x ix5898 (.Y (nx5897), .A0 (nx4774), .A1 (nx4772)) ;
    nor03_2x ix4775 (.Y (nx4774), .A0 (nx5901), .A1 (nx9545), .A2 (nx10655)) ;
    dffr gen_12_cmp_mRegCmp_reg_Q_5 (.Q (gen_12_cmp_mReg_5), .QB (nx5901), .D (
         window_12__5), .CLK (start), .R (rst)) ;
    nor03_2x ix4773 (.Y (nx4772), .A0 (gen_12_cmp_mReg_5), .A1 (nx10071), .A2 (
             nx10663)) ;
    nand02 ix4809 (.Y (gen_12_cmp_BSCmp_op2_6), .A0 (nx5905), .A1 (nx5911)) ;
    nor02_2x ix5906 (.Y (nx5905), .A0 (nx4804), .A1 (nx4800)) ;
    nor03_2x ix4805 (.Y (nx4804), .A0 (gen_12_cmp_mReg_5), .A1 (nx9551), .A2 (
             nx10631)) ;
    nor03_2x ix4801 (.Y (nx4800), .A0 (nx5901), .A1 (nx10637), .A2 (nx10647)) ;
    nor02_2x ix5912 (.Y (nx5911), .A0 (nx4796), .A1 (nx4794)) ;
    nor03_2x ix4797 (.Y (nx4796), .A0 (nx5915), .A1 (nx9545), .A2 (nx10655)) ;
    dffr gen_12_cmp_mRegCmp_reg_Q_6 (.Q (gen_12_cmp_mReg_6), .QB (nx5915), .D (
         window_12__6), .CLK (start), .R (rst)) ;
    nor03_2x ix4795 (.Y (nx4794), .A0 (gen_12_cmp_mReg_6), .A1 (nx10071), .A2 (
             nx10663)) ;
    nand02 ix4831 (.Y (gen_12_cmp_BSCmp_op2_7), .A0 (nx5919), .A1 (nx5925)) ;
    nor02_2x ix5920 (.Y (nx5919), .A0 (nx4826), .A1 (nx4822)) ;
    nor03_2x ix4827 (.Y (nx4826), .A0 (gen_12_cmp_mReg_6), .A1 (nx9551), .A2 (
             nx10633)) ;
    nor03_2x ix4823 (.Y (nx4822), .A0 (nx5915), .A1 (nx10639), .A2 (nx10649)) ;
    nor02_2x ix5926 (.Y (nx5925), .A0 (nx4818), .A1 (nx4816)) ;
    nor03_2x ix4819 (.Y (nx4818), .A0 (nx5928), .A1 (nx9545), .A2 (nx10657)) ;
    dffr gen_12_cmp_mRegCmp_reg_Q_7 (.Q (gen_12_cmp_mReg_7), .QB (nx5928), .D (
         window_12__7), .CLK (start), .R (rst)) ;
    nor03_2x ix4817 (.Y (nx4816), .A0 (gen_12_cmp_mReg_7), .A1 (nx10071), .A2 (
             nx10665)) ;
    nand02 ix4853 (.Y (gen_12_cmp_BSCmp_op2_8), .A0 (nx5935), .A1 (nx5941)) ;
    nor02_2x ix5936 (.Y (nx5935), .A0 (nx4848), .A1 (nx4844)) ;
    nor03_2x ix4849 (.Y (nx4848), .A0 (gen_12_cmp_mReg_7), .A1 (nx9551), .A2 (
             nx10633)) ;
    nor03_2x ix4845 (.Y (nx4844), .A0 (nx5928), .A1 (nx10639), .A2 (nx10649)) ;
    nor02_2x ix5942 (.Y (nx5941), .A0 (nx4840), .A1 (nx4838)) ;
    nor03_2x ix4841 (.Y (nx4840), .A0 (nx5945), .A1 (nx9545), .A2 (nx10657)) ;
    dffr gen_12_cmp_mRegCmp_reg_Q_8 (.Q (gen_12_cmp_mReg_8), .QB (nx5945), .D (
         window_12__8), .CLK (start), .R (rst)) ;
    nor03_2x ix4839 (.Y (nx4838), .A0 (gen_12_cmp_mReg_8), .A1 (nx10073), .A2 (
             nx10665)) ;
    nand02 ix4875 (.Y (gen_12_cmp_BSCmp_op2_9), .A0 (nx5949), .A1 (nx5955)) ;
    nor02_2x ix5950 (.Y (nx5949), .A0 (nx4870), .A1 (nx4866)) ;
    nor03_2x ix4871 (.Y (nx4870), .A0 (gen_12_cmp_mReg_8), .A1 (nx9551), .A2 (
             nx10633)) ;
    nor03_2x ix4867 (.Y (nx4866), .A0 (nx5945), .A1 (nx10639), .A2 (nx10649)) ;
    nor02_2x ix5956 (.Y (nx5955), .A0 (nx4862), .A1 (nx4860)) ;
    nor03_2x ix4863 (.Y (nx4862), .A0 (nx5959), .A1 (nx9545), .A2 (nx10657)) ;
    dffr gen_12_cmp_mRegCmp_reg_Q_9 (.Q (gen_12_cmp_mReg_9), .QB (nx5959), .D (
         window_12__9), .CLK (start), .R (rst)) ;
    nor03_2x ix4861 (.Y (nx4860), .A0 (gen_12_cmp_mReg_9), .A1 (nx10073), .A2 (
             nx10665)) ;
    nand02 ix4897 (.Y (gen_12_cmp_BSCmp_op2_10), .A0 (nx5963), .A1 (nx5969)) ;
    nor02_2x ix5964 (.Y (nx5963), .A0 (nx4892), .A1 (nx4888)) ;
    nor03_2x ix4893 (.Y (nx4892), .A0 (gen_12_cmp_mReg_9), .A1 (nx9551), .A2 (
             nx10633)) ;
    nor03_2x ix4889 (.Y (nx4888), .A0 (nx5959), .A1 (nx10639), .A2 (nx10649)) ;
    nor02_2x ix5970 (.Y (nx5969), .A0 (nx4884), .A1 (nx4882)) ;
    nor03_2x ix4885 (.Y (nx4884), .A0 (nx5972), .A1 (nx9545), .A2 (nx10657)) ;
    dffr gen_12_cmp_mRegCmp_reg_Q_10 (.Q (gen_12_cmp_mReg_10), .QB (nx5972), .D (
         window_12__10), .CLK (start), .R (rst)) ;
    nor03_2x ix4883 (.Y (nx4882), .A0 (gen_12_cmp_mReg_10), .A1 (nx10073), .A2 (
             nx10665)) ;
    nand02 ix4919 (.Y (gen_12_cmp_BSCmp_op2_11), .A0 (nx5979), .A1 (nx5985)) ;
    nor02_2x ix5980 (.Y (nx5979), .A0 (nx4914), .A1 (nx4910)) ;
    nor03_2x ix4915 (.Y (nx4914), .A0 (gen_12_cmp_mReg_10), .A1 (nx9551), .A2 (
             nx10633)) ;
    nor03_2x ix4911 (.Y (nx4910), .A0 (nx5972), .A1 (nx10639), .A2 (nx10649)) ;
    nor02_2x ix5986 (.Y (nx5985), .A0 (nx4906), .A1 (nx4904)) ;
    nor03_2x ix4907 (.Y (nx4906), .A0 (nx5989), .A1 (nx9545), .A2 (nx10657)) ;
    dffr gen_12_cmp_mRegCmp_reg_Q_11 (.Q (gen_12_cmp_mReg_11), .QB (nx5989), .D (
         window_12__11), .CLK (start), .R (rst)) ;
    nor03_2x ix4905 (.Y (nx4904), .A0 (gen_12_cmp_mReg_11), .A1 (nx10073), .A2 (
             nx10665)) ;
    nand02 ix4941 (.Y (gen_12_cmp_BSCmp_op2_12), .A0 (nx5993), .A1 (nx5999)) ;
    nor02_2x ix5994 (.Y (nx5993), .A0 (nx4936), .A1 (nx4932)) ;
    nor03_2x ix4937 (.Y (nx4936), .A0 (gen_12_cmp_mReg_11), .A1 (nx9551), .A2 (
             nx10633)) ;
    nor03_2x ix4933 (.Y (nx4932), .A0 (nx5989), .A1 (nx10639), .A2 (nx10649)) ;
    nor02_2x ix6000 (.Y (nx5999), .A0 (nx4928), .A1 (nx4926)) ;
    nor03_2x ix4929 (.Y (nx4928), .A0 (nx6003), .A1 (nx9547), .A2 (nx10657)) ;
    dffr gen_12_cmp_mRegCmp_reg_Q_12 (.Q (gen_12_cmp_mReg_12), .QB (nx6003), .D (
         window_12__12), .CLK (start), .R (rst)) ;
    nor03_2x ix4927 (.Y (nx4926), .A0 (gen_12_cmp_mReg_12), .A1 (nx10073), .A2 (
             nx10665)) ;
    nand02 ix4963 (.Y (gen_12_cmp_BSCmp_op2_13), .A0 (nx6007), .A1 (nx6013)) ;
    nor02_2x ix6008 (.Y (nx6007), .A0 (nx4958), .A1 (nx4954)) ;
    nor03_2x ix4959 (.Y (nx4958), .A0 (gen_12_cmp_mReg_12), .A1 (nx9553), .A2 (
             nx10635)) ;
    nor03_2x ix4955 (.Y (nx4954), .A0 (nx6003), .A1 (nx10639), .A2 (nx10651)) ;
    nor02_2x ix6014 (.Y (nx6013), .A0 (nx4950), .A1 (nx4948)) ;
    nor03_2x ix4951 (.Y (nx4950), .A0 (nx6016), .A1 (nx9547), .A2 (nx10659)) ;
    dffr gen_12_cmp_mRegCmp_reg_Q_13 (.Q (gen_12_cmp_mReg_13), .QB (nx6016), .D (
         window_12__13), .CLK (start), .R (rst)) ;
    nor03_2x ix4949 (.Y (nx4948), .A0 (gen_12_cmp_mReg_13), .A1 (nx10073), .A2 (
             nx10667)) ;
    nand02 ix4985 (.Y (gen_12_cmp_BSCmp_op2_14), .A0 (nx6023), .A1 (nx6029)) ;
    nor02_2x ix6024 (.Y (nx6023), .A0 (nx4980), .A1 (nx4976)) ;
    nor03_2x ix4981 (.Y (nx4980), .A0 (gen_12_cmp_mReg_13), .A1 (nx9553), .A2 (
             nx10635)) ;
    nor03_2x ix4977 (.Y (nx4976), .A0 (nx6016), .A1 (nx10641), .A2 (nx10651)) ;
    nor02_2x ix6030 (.Y (nx6029), .A0 (nx4972), .A1 (nx4970)) ;
    nor03_2x ix4973 (.Y (nx4972), .A0 (nx6033), .A1 (nx9547), .A2 (nx10659)) ;
    dffr gen_12_cmp_mRegCmp_reg_Q_14 (.Q (gen_12_cmp_mReg_14), .QB (nx6033), .D (
         window_12__14), .CLK (start), .R (rst)) ;
    nor03_2x ix4971 (.Y (nx4970), .A0 (gen_12_cmp_mReg_14), .A1 (nx10073), .A2 (
             nx10667)) ;
    nand02 ix5007 (.Y (gen_12_cmp_BSCmp_op2_15), .A0 (nx6037), .A1 (nx6043)) ;
    nor02_2x ix6038 (.Y (nx6037), .A0 (nx5002), .A1 (nx4998)) ;
    nor03_2x ix5003 (.Y (nx5002), .A0 (gen_12_cmp_mReg_14), .A1 (nx9553), .A2 (
             nx10635)) ;
    nor03_2x ix4999 (.Y (nx4998), .A0 (nx6033), .A1 (nx10641), .A2 (nx10651)) ;
    nor02_2x ix6044 (.Y (nx6043), .A0 (nx4994), .A1 (nx4992)) ;
    nor03_2x ix4995 (.Y (nx4994), .A0 (nx6047), .A1 (nx9547), .A2 (nx10659)) ;
    dffr gen_12_cmp_mRegCmp_reg_Q_15 (.Q (gen_12_cmp_mReg_15), .QB (nx6047), .D (
         window_12__15), .CLK (start), .R (rst)) ;
    nor03_2x ix4993 (.Y (nx4992), .A0 (gen_12_cmp_mReg_15), .A1 (nx10075), .A2 (
             nx10667)) ;
    nand02 ix5017 (.Y (gen_12_cmp_BSCmp_op2_16), .A0 (nx6051), .A1 (nx6043)) ;
    nor02_2x ix6052 (.Y (nx6051), .A0 (nx5012), .A1 (nx5008)) ;
    nor03_2x ix5013 (.Y (nx5012), .A0 (gen_12_cmp_mReg_15), .A1 (nx9553), .A2 (
             nx10635)) ;
    nor03_2x ix5009 (.Y (nx5008), .A0 (nx6047), .A1 (nx10641), .A2 (nx10651)) ;
    nand02 ix5085 (.Y (gen_13_cmp_BSCmp_op2_1), .A0 (nx6058), .A1 (nx6077)) ;
    nor02_2x ix6059 (.Y (nx6058), .A0 (nx5080), .A1 (nx5076)) ;
    nor03_2x ix5081 (.Y (nx5080), .A0 (gen_13_cmp_mReg_0), .A1 (nx9537), .A2 (
             nx10671)) ;
    dffr gen_13_cmp_mRegCmp_reg_Q_0 (.Q (gen_13_cmp_mReg_0), .QB (nx6063), .D (
         window_13__0), .CLK (start), .R (rst)) ;
    inv01 ix6068 (.Y (nx6067), .A (gen_13_cmp_pMux_0)) ;
    nor03_2x ix5077 (.Y (nx5076), .A0 (nx6063), .A1 (nx10677), .A2 (nx10687)) ;
    inv02 ix6076 (.Y (nx6075), .A (gen_13_cmp_pMux_2)) ;
    nor02_2x ix6078 (.Y (nx6077), .A0 (nx5066), .A1 (nx5064)) ;
    nor03_2x ix5067 (.Y (nx5066), .A0 (nx6080), .A1 (nx9531), .A2 (nx10695)) ;
    dffr gen_13_cmp_mRegCmp_reg_Q_1 (.Q (gen_13_cmp_mReg_1), .QB (nx6080), .D (
         window_13__1), .CLK (start), .R (rst)) ;
    nor03_2x ix5065 (.Y (nx5064), .A0 (gen_13_cmp_mReg_1), .A1 (nx10077), .A2 (
             nx10703)) ;
    nor03_2x ix5025 (.Y (nx5024), .A0 (nx9537), .A1 (nx6075), .A2 (
             gen_13_cmp_pMux_0)) ;
    nand02 ix5107 (.Y (gen_13_cmp_BSCmp_op2_2), .A0 (nx6093), .A1 (nx6099)) ;
    nor02_2x ix6094 (.Y (nx6093), .A0 (nx5102), .A1 (nx5098)) ;
    nor03_2x ix5103 (.Y (nx5102), .A0 (gen_13_cmp_mReg_1), .A1 (nx9537), .A2 (
             nx10671)) ;
    nor03_2x ix5099 (.Y (nx5098), .A0 (nx6080), .A1 (nx10677), .A2 (nx10687)) ;
    nor02_2x ix6100 (.Y (nx6099), .A0 (nx5094), .A1 (nx5092)) ;
    nor03_2x ix5095 (.Y (nx5094), .A0 (nx6102), .A1 (nx9531), .A2 (nx10695)) ;
    dffr gen_13_cmp_mRegCmp_reg_Q_2 (.Q (gen_13_cmp_mReg_2), .QB (nx6102), .D (
         window_13__2), .CLK (start), .R (rst)) ;
    nor03_2x ix5093 (.Y (nx5092), .A0 (gen_13_cmp_mReg_2), .A1 (nx10077), .A2 (
             nx10703)) ;
    nand02 ix5129 (.Y (gen_13_cmp_BSCmp_op2_3), .A0 (nx6107), .A1 (nx6113)) ;
    nor02_2x ix6108 (.Y (nx6107), .A0 (nx5124), .A1 (nx5120)) ;
    nor03_2x ix5125 (.Y (nx5124), .A0 (gen_13_cmp_mReg_2), .A1 (nx9537), .A2 (
             nx10671)) ;
    nor03_2x ix5121 (.Y (nx5120), .A0 (nx6102), .A1 (nx10677), .A2 (nx10687)) ;
    nor02_2x ix6114 (.Y (nx6113), .A0 (nx5116), .A1 (nx5114)) ;
    nor03_2x ix5117 (.Y (nx5116), .A0 (nx6117), .A1 (nx9531), .A2 (nx10695)) ;
    dffr gen_13_cmp_mRegCmp_reg_Q_3 (.Q (gen_13_cmp_mReg_3), .QB (nx6117), .D (
         window_13__3), .CLK (start), .R (rst)) ;
    nor03_2x ix5115 (.Y (nx5114), .A0 (gen_13_cmp_mReg_3), .A1 (nx10077), .A2 (
             nx10703)) ;
    nand02 ix5151 (.Y (gen_13_cmp_BSCmp_op2_4), .A0 (nx6123), .A1 (nx6127)) ;
    nor02_2x ix6124 (.Y (nx6123), .A0 (nx5146), .A1 (nx5142)) ;
    nor03_2x ix5147 (.Y (nx5146), .A0 (gen_13_cmp_mReg_3), .A1 (nx9537), .A2 (
             nx10671)) ;
    nor03_2x ix5143 (.Y (nx5142), .A0 (nx6117), .A1 (nx10677), .A2 (nx10687)) ;
    nor02_2x ix6128 (.Y (nx6127), .A0 (nx5138), .A1 (nx5136)) ;
    nor03_2x ix5139 (.Y (nx5138), .A0 (nx6131), .A1 (nx9531), .A2 (nx10695)) ;
    dffr gen_13_cmp_mRegCmp_reg_Q_4 (.Q (gen_13_cmp_mReg_4), .QB (nx6131), .D (
         window_13__4), .CLK (start), .R (rst)) ;
    nor03_2x ix5137 (.Y (nx5136), .A0 (gen_13_cmp_mReg_4), .A1 (nx10077), .A2 (
             nx10703)) ;
    nand02 ix5173 (.Y (gen_13_cmp_BSCmp_op2_5), .A0 (nx6137), .A1 (nx6143)) ;
    nor02_2x ix6138 (.Y (nx6137), .A0 (nx5168), .A1 (nx5164)) ;
    nor03_2x ix5169 (.Y (nx5168), .A0 (gen_13_cmp_mReg_4), .A1 (nx9537), .A2 (
             nx10671)) ;
    nor03_2x ix5165 (.Y (nx5164), .A0 (nx6131), .A1 (nx10677), .A2 (nx10687)) ;
    nor02_2x ix6144 (.Y (nx6143), .A0 (nx5160), .A1 (nx5158)) ;
    nor03_2x ix5161 (.Y (nx5160), .A0 (nx6146), .A1 (nx9533), .A2 (nx10695)) ;
    dffr gen_13_cmp_mRegCmp_reg_Q_5 (.Q (gen_13_cmp_mReg_5), .QB (nx6146), .D (
         window_13__5), .CLK (start), .R (rst)) ;
    nor03_2x ix5159 (.Y (nx5158), .A0 (gen_13_cmp_mReg_5), .A1 (nx10077), .A2 (
             nx10703)) ;
    nand02 ix5195 (.Y (gen_13_cmp_BSCmp_op2_6), .A0 (nx6151), .A1 (nx6157)) ;
    nor02_2x ix6152 (.Y (nx6151), .A0 (nx5190), .A1 (nx5186)) ;
    nor03_2x ix5191 (.Y (nx5190), .A0 (gen_13_cmp_mReg_5), .A1 (nx9539), .A2 (
             nx10671)) ;
    nor03_2x ix5187 (.Y (nx5186), .A0 (nx6146), .A1 (nx10677), .A2 (nx10687)) ;
    nor02_2x ix6158 (.Y (nx6157), .A0 (nx5182), .A1 (nx5180)) ;
    nor03_2x ix5183 (.Y (nx5182), .A0 (nx6161), .A1 (nx9533), .A2 (nx10695)) ;
    dffr gen_13_cmp_mRegCmp_reg_Q_6 (.Q (gen_13_cmp_mReg_6), .QB (nx6161), .D (
         window_13__6), .CLK (start), .R (rst)) ;
    nor03_2x ix5181 (.Y (nx5180), .A0 (gen_13_cmp_mReg_6), .A1 (nx10077), .A2 (
             nx10703)) ;
    nand02 ix5217 (.Y (gen_13_cmp_BSCmp_op2_7), .A0 (nx6167), .A1 (nx6171)) ;
    nor02_2x ix6168 (.Y (nx6167), .A0 (nx5212), .A1 (nx5208)) ;
    nor03_2x ix5213 (.Y (nx5212), .A0 (gen_13_cmp_mReg_6), .A1 (nx9539), .A2 (
             nx10673)) ;
    nor03_2x ix5209 (.Y (nx5208), .A0 (nx6161), .A1 (nx10679), .A2 (nx10689)) ;
    nor02_2x ix6172 (.Y (nx6171), .A0 (nx5204), .A1 (nx5202)) ;
    nor03_2x ix5205 (.Y (nx5204), .A0 (nx6175), .A1 (nx9533), .A2 (nx10697)) ;
    dffr gen_13_cmp_mRegCmp_reg_Q_7 (.Q (gen_13_cmp_mReg_7), .QB (nx6175), .D (
         window_13__7), .CLK (start), .R (rst)) ;
    nor03_2x ix5203 (.Y (nx5202), .A0 (gen_13_cmp_mReg_7), .A1 (nx10077), .A2 (
             nx10705)) ;
    nand02 ix5239 (.Y (gen_13_cmp_BSCmp_op2_8), .A0 (nx6181), .A1 (nx6186)) ;
    nor02_2x ix6182 (.Y (nx6181), .A0 (nx5234), .A1 (nx5230)) ;
    nor03_2x ix5235 (.Y (nx5234), .A0 (gen_13_cmp_mReg_7), .A1 (nx9539), .A2 (
             nx10673)) ;
    nor03_2x ix5231 (.Y (nx5230), .A0 (nx6175), .A1 (nx10679), .A2 (nx10689)) ;
    nor02_2x ix6187 (.Y (nx6186), .A0 (nx5226), .A1 (nx5224)) ;
    nor03_2x ix5227 (.Y (nx5226), .A0 (nx6189), .A1 (nx9533), .A2 (nx10697)) ;
    dffr gen_13_cmp_mRegCmp_reg_Q_8 (.Q (gen_13_cmp_mReg_8), .QB (nx6189), .D (
         window_13__8), .CLK (start), .R (rst)) ;
    nor03_2x ix5225 (.Y (nx5224), .A0 (gen_13_cmp_mReg_8), .A1 (nx10079), .A2 (
             nx10705)) ;
    nand02 ix5261 (.Y (gen_13_cmp_BSCmp_op2_9), .A0 (nx6193), .A1 (nx6199)) ;
    nor02_2x ix6194 (.Y (nx6193), .A0 (nx5256), .A1 (nx5252)) ;
    nor03_2x ix5257 (.Y (nx5256), .A0 (gen_13_cmp_mReg_8), .A1 (nx9539), .A2 (
             nx10673)) ;
    nor03_2x ix5253 (.Y (nx5252), .A0 (nx6189), .A1 (nx10679), .A2 (nx10689)) ;
    nor02_2x ix6200 (.Y (nx6199), .A0 (nx5248), .A1 (nx5246)) ;
    nor03_2x ix5249 (.Y (nx5248), .A0 (nx6203), .A1 (nx9533), .A2 (nx10697)) ;
    dffr gen_13_cmp_mRegCmp_reg_Q_9 (.Q (gen_13_cmp_mReg_9), .QB (nx6203), .D (
         window_13__9), .CLK (start), .R (rst)) ;
    nor03_2x ix5247 (.Y (nx5246), .A0 (gen_13_cmp_mReg_9), .A1 (nx10079), .A2 (
             nx10705)) ;
    nand02 ix5283 (.Y (gen_13_cmp_BSCmp_op2_10), .A0 (nx6209), .A1 (nx6215)) ;
    nor02_2x ix6210 (.Y (nx6209), .A0 (nx5278), .A1 (nx5274)) ;
    nor03_2x ix5279 (.Y (nx5278), .A0 (gen_13_cmp_mReg_9), .A1 (nx9539), .A2 (
             nx10673)) ;
    nor03_2x ix5275 (.Y (nx5274), .A0 (nx6203), .A1 (nx10679), .A2 (nx10689)) ;
    nor02_2x ix6216 (.Y (nx6215), .A0 (nx5270), .A1 (nx5268)) ;
    nor03_2x ix5271 (.Y (nx5270), .A0 (nx6218), .A1 (nx9533), .A2 (nx10697)) ;
    dffr gen_13_cmp_mRegCmp_reg_Q_10 (.Q (gen_13_cmp_mReg_10), .QB (nx6218), .D (
         window_13__10), .CLK (start), .R (rst)) ;
    nor03_2x ix5269 (.Y (nx5268), .A0 (gen_13_cmp_mReg_10), .A1 (nx10079), .A2 (
             nx10705)) ;
    nand02 ix5305 (.Y (gen_13_cmp_BSCmp_op2_11), .A0 (nx6223), .A1 (nx6229)) ;
    nor02_2x ix6224 (.Y (nx6223), .A0 (nx5300), .A1 (nx5296)) ;
    nor03_2x ix5301 (.Y (nx5300), .A0 (gen_13_cmp_mReg_10), .A1 (nx9539), .A2 (
             nx10673)) ;
    nor03_2x ix5297 (.Y (nx5296), .A0 (nx6218), .A1 (nx10679), .A2 (nx10689)) ;
    nor02_2x ix6230 (.Y (nx6229), .A0 (nx5292), .A1 (nx5290)) ;
    nor03_2x ix5293 (.Y (nx5292), .A0 (nx6233), .A1 (nx9533), .A2 (nx10697)) ;
    dffr gen_13_cmp_mRegCmp_reg_Q_11 (.Q (gen_13_cmp_mReg_11), .QB (nx6233), .D (
         window_13__11), .CLK (start), .R (rst)) ;
    nor03_2x ix5291 (.Y (nx5290), .A0 (gen_13_cmp_mReg_11), .A1 (nx10079), .A2 (
             nx10705)) ;
    nand02 ix5327 (.Y (gen_13_cmp_BSCmp_op2_12), .A0 (nx6239), .A1 (nx6245)) ;
    nor02_2x ix6240 (.Y (nx6239), .A0 (nx5322), .A1 (nx5318)) ;
    nor03_2x ix5323 (.Y (nx5322), .A0 (gen_13_cmp_mReg_11), .A1 (nx9539), .A2 (
             nx10673)) ;
    nor03_2x ix5319 (.Y (nx5318), .A0 (nx6233), .A1 (nx10679), .A2 (nx10689)) ;
    nor02_2x ix6246 (.Y (nx6245), .A0 (nx5314), .A1 (nx5312)) ;
    nor03_2x ix5315 (.Y (nx5314), .A0 (nx6248), .A1 (nx9535), .A2 (nx10697)) ;
    dffr gen_13_cmp_mRegCmp_reg_Q_12 (.Q (gen_13_cmp_mReg_12), .QB (nx6248), .D (
         window_13__12), .CLK (start), .R (rst)) ;
    nor03_2x ix5313 (.Y (nx5312), .A0 (gen_13_cmp_mReg_12), .A1 (nx10079), .A2 (
             nx10705)) ;
    nand02 ix5349 (.Y (gen_13_cmp_BSCmp_op2_13), .A0 (nx6255), .A1 (nx6261)) ;
    nor02_2x ix6256 (.Y (nx6255), .A0 (nx5344), .A1 (nx5340)) ;
    nor03_2x ix5345 (.Y (nx5344), .A0 (gen_13_cmp_mReg_12), .A1 (nx9541), .A2 (
             nx10675)) ;
    nor03_2x ix5341 (.Y (nx5340), .A0 (nx6248), .A1 (nx10679), .A2 (nx10691)) ;
    nor02_2x ix6262 (.Y (nx6261), .A0 (nx5336), .A1 (nx5334)) ;
    nor03_2x ix5337 (.Y (nx5336), .A0 (nx6265), .A1 (nx9535), .A2 (nx10699)) ;
    dffr gen_13_cmp_mRegCmp_reg_Q_13 (.Q (gen_13_cmp_mReg_13), .QB (nx6265), .D (
         window_13__13), .CLK (start), .R (rst)) ;
    nor03_2x ix5335 (.Y (nx5334), .A0 (gen_13_cmp_mReg_13), .A1 (nx10079), .A2 (
             nx10707)) ;
    nand02 ix5371 (.Y (gen_13_cmp_BSCmp_op2_14), .A0 (nx6269), .A1 (nx6275)) ;
    nor02_2x ix6270 (.Y (nx6269), .A0 (nx5366), .A1 (nx5362)) ;
    nor03_2x ix5367 (.Y (nx5366), .A0 (gen_13_cmp_mReg_13), .A1 (nx9541), .A2 (
             nx10675)) ;
    nor03_2x ix5363 (.Y (nx5362), .A0 (nx6265), .A1 (nx10681), .A2 (nx10691)) ;
    nor02_2x ix6276 (.Y (nx6275), .A0 (nx5358), .A1 (nx5356)) ;
    nor03_2x ix5359 (.Y (nx5358), .A0 (nx6279), .A1 (nx9535), .A2 (nx10699)) ;
    dffr gen_13_cmp_mRegCmp_reg_Q_14 (.Q (gen_13_cmp_mReg_14), .QB (nx6279), .D (
         window_13__14), .CLK (start), .R (rst)) ;
    nor03_2x ix5357 (.Y (nx5356), .A0 (gen_13_cmp_mReg_14), .A1 (nx10079), .A2 (
             nx10707)) ;
    nand02 ix5393 (.Y (gen_13_cmp_BSCmp_op2_15), .A0 (nx6283), .A1 (nx6289)) ;
    nor02_2x ix6284 (.Y (nx6283), .A0 (nx5388), .A1 (nx5384)) ;
    nor03_2x ix5389 (.Y (nx5388), .A0 (gen_13_cmp_mReg_14), .A1 (nx9541), .A2 (
             nx10675)) ;
    nor03_2x ix5385 (.Y (nx5384), .A0 (nx6279), .A1 (nx10681), .A2 (nx10691)) ;
    nor02_2x ix6290 (.Y (nx6289), .A0 (nx5380), .A1 (nx5378)) ;
    nor03_2x ix5381 (.Y (nx5380), .A0 (nx6292), .A1 (nx9535), .A2 (nx10699)) ;
    dffr gen_13_cmp_mRegCmp_reg_Q_15 (.Q (gen_13_cmp_mReg_15), .QB (nx6292), .D (
         window_13__15), .CLK (start), .R (rst)) ;
    nor03_2x ix5379 (.Y (nx5378), .A0 (gen_13_cmp_mReg_15), .A1 (nx10081), .A2 (
             nx10707)) ;
    nand02 ix5403 (.Y (gen_13_cmp_BSCmp_op2_16), .A0 (nx6299), .A1 (nx6289)) ;
    nor02_2x ix6300 (.Y (nx6299), .A0 (nx5398), .A1 (nx5394)) ;
    nor03_2x ix5399 (.Y (nx5398), .A0 (gen_13_cmp_mReg_15), .A1 (nx9541), .A2 (
             nx10675)) ;
    nor03_2x ix5395 (.Y (nx5394), .A0 (nx6292), .A1 (nx10681), .A2 (nx10691)) ;
    nand02 ix5471 (.Y (gen_14_cmp_BSCmp_op2_1), .A0 (nx6305), .A1 (nx6325)) ;
    nor02_2x ix6306 (.Y (nx6305), .A0 (nx5466), .A1 (nx5462)) ;
    nor03_2x ix5467 (.Y (nx5466), .A0 (gen_14_cmp_mReg_0), .A1 (nx9525), .A2 (
             nx10711)) ;
    dffr gen_14_cmp_mRegCmp_reg_Q_0 (.Q (gen_14_cmp_mReg_0), .QB (nx6311), .D (
         window_14__0), .CLK (start), .R (rst)) ;
    inv01 ix6316 (.Y (nx6314), .A (gen_14_cmp_pMux_0)) ;
    nor03_2x ix5463 (.Y (nx5462), .A0 (nx6311), .A1 (nx10717), .A2 (nx10727)) ;
    inv02 ix6324 (.Y (nx6323), .A (gen_14_cmp_pMux_2)) ;
    nor02_2x ix6326 (.Y (nx6325), .A0 (nx5452), .A1 (nx5450)) ;
    nor03_2x ix5453 (.Y (nx5452), .A0 (nx6329), .A1 (nx9519), .A2 (nx10735)) ;
    dffr gen_14_cmp_mRegCmp_reg_Q_1 (.Q (gen_14_cmp_mReg_1), .QB (nx6329), .D (
         window_14__1), .CLK (start), .R (rst)) ;
    nor03_2x ix5451 (.Y (nx5450), .A0 (gen_14_cmp_mReg_1), .A1 (nx10083), .A2 (
             nx10743)) ;
    nor03_2x ix5411 (.Y (nx5410), .A0 (nx9525), .A1 (nx6323), .A2 (
             gen_14_cmp_pMux_0)) ;
    nand02 ix5493 (.Y (gen_14_cmp_BSCmp_op2_2), .A0 (nx6339), .A1 (nx6345)) ;
    nor02_2x ix6340 (.Y (nx6339), .A0 (nx5488), .A1 (nx5484)) ;
    nor03_2x ix5489 (.Y (nx5488), .A0 (gen_14_cmp_mReg_1), .A1 (nx9525), .A2 (
             nx10711)) ;
    nor03_2x ix5485 (.Y (nx5484), .A0 (nx6329), .A1 (nx10717), .A2 (nx10727)) ;
    nor02_2x ix6346 (.Y (nx6345), .A0 (nx5480), .A1 (nx5478)) ;
    nor03_2x ix5481 (.Y (nx5480), .A0 (nx6349), .A1 (nx9519), .A2 (nx10735)) ;
    dffr gen_14_cmp_mRegCmp_reg_Q_2 (.Q (gen_14_cmp_mReg_2), .QB (nx6349), .D (
         window_14__2), .CLK (start), .R (rst)) ;
    nor03_2x ix5479 (.Y (nx5478), .A0 (gen_14_cmp_mReg_2), .A1 (nx10083), .A2 (
             nx10743)) ;
    nand02 ix5515 (.Y (gen_14_cmp_BSCmp_op2_3), .A0 (nx6355), .A1 (nx6359)) ;
    nor02_2x ix6356 (.Y (nx6355), .A0 (nx5510), .A1 (nx5506)) ;
    nor03_2x ix5511 (.Y (nx5510), .A0 (gen_14_cmp_mReg_2), .A1 (nx9525), .A2 (
             nx10711)) ;
    nor03_2x ix5507 (.Y (nx5506), .A0 (nx6349), .A1 (nx10717), .A2 (nx10727)) ;
    nor02_2x ix6360 (.Y (nx6359), .A0 (nx5502), .A1 (nx5500)) ;
    nor03_2x ix5503 (.Y (nx5502), .A0 (nx6363), .A1 (nx9519), .A2 (nx10735)) ;
    dffr gen_14_cmp_mRegCmp_reg_Q_3 (.Q (gen_14_cmp_mReg_3), .QB (nx6363), .D (
         window_14__3), .CLK (start), .R (rst)) ;
    nor03_2x ix5501 (.Y (nx5500), .A0 (gen_14_cmp_mReg_3), .A1 (nx10083), .A2 (
             nx10743)) ;
    nand02 ix5537 (.Y (gen_14_cmp_BSCmp_op2_4), .A0 (nx6369), .A1 (nx6375)) ;
    nor02_2x ix6370 (.Y (nx6369), .A0 (nx5532), .A1 (nx5528)) ;
    nor03_2x ix5533 (.Y (nx5532), .A0 (gen_14_cmp_mReg_3), .A1 (nx9525), .A2 (
             nx10711)) ;
    nor03_2x ix5529 (.Y (nx5528), .A0 (nx6363), .A1 (nx10717), .A2 (nx10727)) ;
    nor02_2x ix6376 (.Y (nx6375), .A0 (nx5524), .A1 (nx5522)) ;
    nor03_2x ix5525 (.Y (nx5524), .A0 (nx6378), .A1 (nx9519), .A2 (nx10735)) ;
    dffr gen_14_cmp_mRegCmp_reg_Q_4 (.Q (gen_14_cmp_mReg_4), .QB (nx6378), .D (
         window_14__4), .CLK (start), .R (rst)) ;
    nor03_2x ix5523 (.Y (nx5522), .A0 (gen_14_cmp_mReg_4), .A1 (nx10083), .A2 (
             nx10743)) ;
    nand02 ix5559 (.Y (gen_14_cmp_BSCmp_op2_5), .A0 (nx6383), .A1 (nx6389)) ;
    nor02_2x ix6384 (.Y (nx6383), .A0 (nx5554), .A1 (nx5550)) ;
    nor03_2x ix5555 (.Y (nx5554), .A0 (gen_14_cmp_mReg_4), .A1 (nx9525), .A2 (
             nx10711)) ;
    nor03_2x ix5551 (.Y (nx5550), .A0 (nx6378), .A1 (nx10717), .A2 (nx10727)) ;
    nor02_2x ix6390 (.Y (nx6389), .A0 (nx5546), .A1 (nx5544)) ;
    nor03_2x ix5547 (.Y (nx5546), .A0 (nx6393), .A1 (nx9521), .A2 (nx10735)) ;
    dffr gen_14_cmp_mRegCmp_reg_Q_5 (.Q (gen_14_cmp_mReg_5), .QB (nx6393), .D (
         window_14__5), .CLK (start), .R (rst)) ;
    nor03_2x ix5545 (.Y (nx5544), .A0 (gen_14_cmp_mReg_5), .A1 (nx10083), .A2 (
             nx10743)) ;
    nand02 ix5581 (.Y (gen_14_cmp_BSCmp_op2_6), .A0 (nx6399), .A1 (nx6403)) ;
    nor02_2x ix6400 (.Y (nx6399), .A0 (nx5576), .A1 (nx5572)) ;
    nor03_2x ix5577 (.Y (nx5576), .A0 (gen_14_cmp_mReg_5), .A1 (nx9527), .A2 (
             nx10711)) ;
    nor03_2x ix5573 (.Y (nx5572), .A0 (nx6393), .A1 (nx10717), .A2 (nx10727)) ;
    nor02_2x ix6404 (.Y (nx6403), .A0 (nx5568), .A1 (nx5566)) ;
    nor03_2x ix5569 (.Y (nx5568), .A0 (nx6407), .A1 (nx9521), .A2 (nx10735)) ;
    dffr gen_14_cmp_mRegCmp_reg_Q_6 (.Q (gen_14_cmp_mReg_6), .QB (nx6407), .D (
         window_14__6), .CLK (start), .R (rst)) ;
    nor03_2x ix5567 (.Y (nx5566), .A0 (gen_14_cmp_mReg_6), .A1 (nx10083), .A2 (
             nx10743)) ;
    nand02 ix5603 (.Y (gen_14_cmp_BSCmp_op2_7), .A0 (nx6413), .A1 (nx6419)) ;
    nor02_2x ix6414 (.Y (nx6413), .A0 (nx5598), .A1 (nx5594)) ;
    nor03_2x ix5599 (.Y (nx5598), .A0 (gen_14_cmp_mReg_6), .A1 (nx9527), .A2 (
             nx10713)) ;
    nor03_2x ix5595 (.Y (nx5594), .A0 (nx6407), .A1 (nx10719), .A2 (nx10729)) ;
    nor02_2x ix6420 (.Y (nx6419), .A0 (nx5590), .A1 (nx5588)) ;
    nor03_2x ix5591 (.Y (nx5590), .A0 (nx6422), .A1 (nx9521), .A2 (nx10737)) ;
    dffr gen_14_cmp_mRegCmp_reg_Q_7 (.Q (gen_14_cmp_mReg_7), .QB (nx6422), .D (
         window_14__7), .CLK (start), .R (rst)) ;
    nor03_2x ix5589 (.Y (nx5588), .A0 (gen_14_cmp_mReg_7), .A1 (nx10083), .A2 (
             nx10745)) ;
    nand02 ix5625 (.Y (gen_14_cmp_BSCmp_op2_8), .A0 (nx6427), .A1 (nx6433)) ;
    nor02_2x ix6428 (.Y (nx6427), .A0 (nx5620), .A1 (nx5616)) ;
    nor03_2x ix5621 (.Y (nx5620), .A0 (gen_14_cmp_mReg_7), .A1 (nx9527), .A2 (
             nx10713)) ;
    nor03_2x ix5617 (.Y (nx5616), .A0 (nx6422), .A1 (nx10719), .A2 (nx10729)) ;
    nor02_2x ix6434 (.Y (nx6433), .A0 (nx5612), .A1 (nx5610)) ;
    nor03_2x ix5613 (.Y (nx5612), .A0 (nx6437), .A1 (nx9521), .A2 (nx10737)) ;
    dffr gen_14_cmp_mRegCmp_reg_Q_8 (.Q (gen_14_cmp_mReg_8), .QB (nx6437), .D (
         window_14__8), .CLK (start), .R (rst)) ;
    nor03_2x ix5611 (.Y (nx5610), .A0 (gen_14_cmp_mReg_8), .A1 (nx10085), .A2 (
             nx10745)) ;
    nand02 ix5647 (.Y (gen_14_cmp_BSCmp_op2_9), .A0 (nx6443), .A1 (nx6447)) ;
    nor02_2x ix6444 (.Y (nx6443), .A0 (nx5642), .A1 (nx5638)) ;
    nor03_2x ix5643 (.Y (nx5642), .A0 (gen_14_cmp_mReg_8), .A1 (nx9527), .A2 (
             nx10713)) ;
    nor03_2x ix5639 (.Y (nx5638), .A0 (nx6437), .A1 (nx10719), .A2 (nx10729)) ;
    nor02_2x ix6448 (.Y (nx6447), .A0 (nx5634), .A1 (nx5632)) ;
    nor03_2x ix5635 (.Y (nx5634), .A0 (nx6451), .A1 (nx9521), .A2 (nx10737)) ;
    dffr gen_14_cmp_mRegCmp_reg_Q_9 (.Q (gen_14_cmp_mReg_9), .QB (nx6451), .D (
         window_14__9), .CLK (start), .R (rst)) ;
    nor03_2x ix5633 (.Y (nx5632), .A0 (gen_14_cmp_mReg_9), .A1 (nx10085), .A2 (
             nx10745)) ;
    nand02 ix5669 (.Y (gen_14_cmp_BSCmp_op2_10), .A0 (nx6457), .A1 (nx6463)) ;
    nor02_2x ix6458 (.Y (nx6457), .A0 (nx5664), .A1 (nx5660)) ;
    nor03_2x ix5665 (.Y (nx5664), .A0 (gen_14_cmp_mReg_9), .A1 (nx9527), .A2 (
             nx10713)) ;
    nor03_2x ix5661 (.Y (nx5660), .A0 (nx6451), .A1 (nx10719), .A2 (nx10729)) ;
    nor02_2x ix6464 (.Y (nx6463), .A0 (nx5656), .A1 (nx5654)) ;
    nor03_2x ix5657 (.Y (nx5656), .A0 (nx6466), .A1 (nx9521), .A2 (nx10737)) ;
    dffr gen_14_cmp_mRegCmp_reg_Q_10 (.Q (gen_14_cmp_mReg_10), .QB (nx6466), .D (
         window_14__10), .CLK (start), .R (rst)) ;
    nor03_2x ix5655 (.Y (nx5654), .A0 (gen_14_cmp_mReg_10), .A1 (nx10085), .A2 (
             nx10745)) ;
    nand02 ix5691 (.Y (gen_14_cmp_BSCmp_op2_11), .A0 (nx6471), .A1 (nx6477)) ;
    nor02_2x ix6472 (.Y (nx6471), .A0 (nx5686), .A1 (nx5682)) ;
    nor03_2x ix5687 (.Y (nx5686), .A0 (gen_14_cmp_mReg_10), .A1 (nx9527), .A2 (
             nx10713)) ;
    nor03_2x ix5683 (.Y (nx5682), .A0 (nx6466), .A1 (nx10719), .A2 (nx10729)) ;
    nor02_2x ix6478 (.Y (nx6477), .A0 (nx5678), .A1 (nx5676)) ;
    nor03_2x ix5679 (.Y (nx5678), .A0 (nx6481), .A1 (nx9521), .A2 (nx10737)) ;
    dffr gen_14_cmp_mRegCmp_reg_Q_11 (.Q (gen_14_cmp_mReg_11), .QB (nx6481), .D (
         window_14__11), .CLK (start), .R (rst)) ;
    nor03_2x ix5677 (.Y (nx5676), .A0 (gen_14_cmp_mReg_11), .A1 (nx10085), .A2 (
             nx10745)) ;
    nand02 ix5713 (.Y (gen_14_cmp_BSCmp_op2_12), .A0 (nx6487), .A1 (nx6491)) ;
    nor02_2x ix6488 (.Y (nx6487), .A0 (nx5708), .A1 (nx5704)) ;
    nor03_2x ix5709 (.Y (nx5708), .A0 (gen_14_cmp_mReg_11), .A1 (nx9527), .A2 (
             nx10713)) ;
    nor03_2x ix5705 (.Y (nx5704), .A0 (nx6481), .A1 (nx10719), .A2 (nx10729)) ;
    nor02_2x ix6492 (.Y (nx6491), .A0 (nx5700), .A1 (nx5698)) ;
    nor03_2x ix5701 (.Y (nx5700), .A0 (nx6495), .A1 (nx9523), .A2 (nx10737)) ;
    dffr gen_14_cmp_mRegCmp_reg_Q_12 (.Q (gen_14_cmp_mReg_12), .QB (nx6495), .D (
         window_14__12), .CLK (start), .R (rst)) ;
    nor03_2x ix5699 (.Y (nx5698), .A0 (gen_14_cmp_mReg_12), .A1 (nx10085), .A2 (
             nx10745)) ;
    nand02 ix5735 (.Y (gen_14_cmp_BSCmp_op2_13), .A0 (nx6501), .A1 (nx6507)) ;
    nor02_2x ix6502 (.Y (nx6501), .A0 (nx5730), .A1 (nx5726)) ;
    nor03_2x ix5731 (.Y (nx5730), .A0 (gen_14_cmp_mReg_12), .A1 (nx9529), .A2 (
             nx10715)) ;
    nor03_2x ix5727 (.Y (nx5726), .A0 (nx6495), .A1 (nx10719), .A2 (nx10731)) ;
    nor02_2x ix6508 (.Y (nx6507), .A0 (nx5722), .A1 (nx5720)) ;
    nor03_2x ix5723 (.Y (nx5722), .A0 (nx6510), .A1 (nx9523), .A2 (nx10739)) ;
    dffr gen_14_cmp_mRegCmp_reg_Q_13 (.Q (gen_14_cmp_mReg_13), .QB (nx6510), .D (
         window_14__13), .CLK (start), .R (rst)) ;
    nor03_2x ix5721 (.Y (nx5720), .A0 (gen_14_cmp_mReg_13), .A1 (nx10085), .A2 (
             nx10747)) ;
    nand02 ix5757 (.Y (gen_14_cmp_BSCmp_op2_14), .A0 (nx6515), .A1 (nx6521)) ;
    nor02_2x ix6516 (.Y (nx6515), .A0 (nx5752), .A1 (nx5748)) ;
    nor03_2x ix5753 (.Y (nx5752), .A0 (gen_14_cmp_mReg_13), .A1 (nx9529), .A2 (
             nx10715)) ;
    nor03_2x ix5749 (.Y (nx5748), .A0 (nx6510), .A1 (nx10721), .A2 (nx10731)) ;
    nor02_2x ix6522 (.Y (nx6521), .A0 (nx5744), .A1 (nx5742)) ;
    nor03_2x ix5745 (.Y (nx5744), .A0 (nx6525), .A1 (nx9523), .A2 (nx10739)) ;
    dffr gen_14_cmp_mRegCmp_reg_Q_14 (.Q (gen_14_cmp_mReg_14), .QB (nx6525), .D (
         window_14__14), .CLK (start), .R (rst)) ;
    nor03_2x ix5743 (.Y (nx5742), .A0 (gen_14_cmp_mReg_14), .A1 (nx10085), .A2 (
             nx10747)) ;
    nand02 ix5779 (.Y (gen_14_cmp_BSCmp_op2_15), .A0 (nx6531), .A1 (nx6535)) ;
    nor02_2x ix6532 (.Y (nx6531), .A0 (nx5774), .A1 (nx5770)) ;
    nor03_2x ix5775 (.Y (nx5774), .A0 (gen_14_cmp_mReg_14), .A1 (nx9529), .A2 (
             nx10715)) ;
    nor03_2x ix5771 (.Y (nx5770), .A0 (nx6525), .A1 (nx10721), .A2 (nx10731)) ;
    nor02_2x ix6536 (.Y (nx6535), .A0 (nx5766), .A1 (nx5764)) ;
    nor03_2x ix5767 (.Y (nx5766), .A0 (nx6539), .A1 (nx9523), .A2 (nx10739)) ;
    dffr gen_14_cmp_mRegCmp_reg_Q_15 (.Q (gen_14_cmp_mReg_15), .QB (nx6539), .D (
         window_14__15), .CLK (start), .R (rst)) ;
    nor03_2x ix5765 (.Y (nx5764), .A0 (gen_14_cmp_mReg_15), .A1 (nx10087), .A2 (
             nx10747)) ;
    nand02 ix5789 (.Y (gen_14_cmp_BSCmp_op2_16), .A0 (nx6545), .A1 (nx6535)) ;
    nor02_2x ix6546 (.Y (nx6545), .A0 (nx5784), .A1 (nx5780)) ;
    nor03_2x ix5785 (.Y (nx5784), .A0 (gen_14_cmp_mReg_15), .A1 (nx9529), .A2 (
             nx10715)) ;
    nor03_2x ix5781 (.Y (nx5780), .A0 (nx6539), .A1 (nx10721), .A2 (nx10731)) ;
    nand02 ix5857 (.Y (gen_15_cmp_BSCmp_op2_1), .A0 (nx6553), .A1 (nx6571)) ;
    nor02_2x ix6554 (.Y (nx6553), .A0 (nx5852), .A1 (nx5848)) ;
    nor03_2x ix5853 (.Y (nx5852), .A0 (gen_15_cmp_mReg_0), .A1 (nx9513), .A2 (
             nx10751)) ;
    dffr gen_15_cmp_mRegCmp_reg_Q_0 (.Q (gen_15_cmp_mReg_0), .QB (nx6557), .D (
         window_15__0), .CLK (start), .R (rst)) ;
    inv01 ix6562 (.Y (nx6561), .A (gen_15_cmp_pMux_0)) ;
    nor03_2x ix5849 (.Y (nx5848), .A0 (nx6557), .A1 (nx10757), .A2 (nx10767)) ;
    inv02 ix6570 (.Y (nx6569), .A (gen_15_cmp_pMux_2)) ;
    nor02_2x ix6572 (.Y (nx6571), .A0 (nx5838), .A1 (nx5836)) ;
    nor03_2x ix5839 (.Y (nx5838), .A0 (nx6574), .A1 (nx9507), .A2 (nx10775)) ;
    dffr gen_15_cmp_mRegCmp_reg_Q_1 (.Q (gen_15_cmp_mReg_1), .QB (nx6574), .D (
         window_15__1), .CLK (start), .R (rst)) ;
    nor03_2x ix5837 (.Y (nx5836), .A0 (gen_15_cmp_mReg_1), .A1 (nx10089), .A2 (
             nx10783)) ;
    nor03_2x ix5797 (.Y (nx5796), .A0 (nx9513), .A1 (nx6569), .A2 (
             gen_15_cmp_pMux_0)) ;
    nand02 ix5879 (.Y (gen_15_cmp_BSCmp_op2_2), .A0 (nx6585), .A1 (nx6591)) ;
    nor02_2x ix6586 (.Y (nx6585), .A0 (nx5874), .A1 (nx5870)) ;
    nor03_2x ix5875 (.Y (nx5874), .A0 (gen_15_cmp_mReg_1), .A1 (nx9513), .A2 (
             nx10751)) ;
    nor03_2x ix5871 (.Y (nx5870), .A0 (nx6574), .A1 (nx10757), .A2 (nx10767)) ;
    nor02_2x ix6592 (.Y (nx6591), .A0 (nx5866), .A1 (nx5864)) ;
    nor03_2x ix5867 (.Y (nx5866), .A0 (nx6595), .A1 (nx9507), .A2 (nx10775)) ;
    dffr gen_15_cmp_mRegCmp_reg_Q_2 (.Q (gen_15_cmp_mReg_2), .QB (nx6595), .D (
         window_15__2), .CLK (start), .R (rst)) ;
    nor03_2x ix5865 (.Y (nx5864), .A0 (gen_15_cmp_mReg_2), .A1 (nx10089), .A2 (
             nx10783)) ;
    nand02 ix5901 (.Y (gen_15_cmp_BSCmp_op2_3), .A0 (nx6601), .A1 (nx6605)) ;
    nor02_2x ix6602 (.Y (nx6601), .A0 (nx5896), .A1 (nx5892)) ;
    nor03_2x ix5897 (.Y (nx5896), .A0 (gen_15_cmp_mReg_2), .A1 (nx9513), .A2 (
             nx10751)) ;
    nor03_2x ix5893 (.Y (nx5892), .A0 (nx6595), .A1 (nx10757), .A2 (nx10767)) ;
    nor02_2x ix6606 (.Y (nx6605), .A0 (nx5888), .A1 (nx5886)) ;
    nor03_2x ix5889 (.Y (nx5888), .A0 (nx6609), .A1 (nx9507), .A2 (nx10775)) ;
    dffr gen_15_cmp_mRegCmp_reg_Q_3 (.Q (gen_15_cmp_mReg_3), .QB (nx6609), .D (
         window_15__3), .CLK (start), .R (rst)) ;
    nor03_2x ix5887 (.Y (nx5886), .A0 (gen_15_cmp_mReg_3), .A1 (nx10089), .A2 (
             nx10783)) ;
    nand02 ix5923 (.Y (gen_15_cmp_BSCmp_op2_4), .A0 (nx6615), .A1 (nx6621)) ;
    nor02_2x ix6616 (.Y (nx6615), .A0 (nx5918), .A1 (nx5914)) ;
    nor03_2x ix5919 (.Y (nx5918), .A0 (gen_15_cmp_mReg_3), .A1 (nx9513), .A2 (
             nx10751)) ;
    nor03_2x ix5915 (.Y (nx5914), .A0 (nx6609), .A1 (nx10757), .A2 (nx10767)) ;
    nor02_2x ix6622 (.Y (nx6621), .A0 (nx5910), .A1 (nx5908)) ;
    nor03_2x ix5911 (.Y (nx5910), .A0 (nx6625), .A1 (nx9507), .A2 (nx10775)) ;
    dffr gen_15_cmp_mRegCmp_reg_Q_4 (.Q (gen_15_cmp_mReg_4), .QB (nx6625), .D (
         window_15__4), .CLK (start), .R (rst)) ;
    nor03_2x ix5909 (.Y (nx5908), .A0 (gen_15_cmp_mReg_4), .A1 (nx10089), .A2 (
             nx10783)) ;
    nand02 ix5945 (.Y (gen_15_cmp_BSCmp_op2_5), .A0 (nx6631), .A1 (nx6635)) ;
    nor02_2x ix6632 (.Y (nx6631), .A0 (nx5940), .A1 (nx5936)) ;
    nor03_2x ix5941 (.Y (nx5940), .A0 (gen_15_cmp_mReg_4), .A1 (nx9513), .A2 (
             nx10751)) ;
    nor03_2x ix5937 (.Y (nx5936), .A0 (nx6625), .A1 (nx10757), .A2 (nx10767)) ;
    nor02_2x ix6636 (.Y (nx6635), .A0 (nx5932), .A1 (nx5930)) ;
    nor03_2x ix5933 (.Y (nx5932), .A0 (nx6639), .A1 (nx9509), .A2 (nx10775)) ;
    dffr gen_15_cmp_mRegCmp_reg_Q_5 (.Q (gen_15_cmp_mReg_5), .QB (nx6639), .D (
         window_15__5), .CLK (start), .R (rst)) ;
    nor03_2x ix5931 (.Y (nx5930), .A0 (gen_15_cmp_mReg_5), .A1 (nx10089), .A2 (
             nx10783)) ;
    nand02 ix5967 (.Y (gen_15_cmp_BSCmp_op2_6), .A0 (nx6645), .A1 (nx6651)) ;
    nor02_2x ix6646 (.Y (nx6645), .A0 (nx5962), .A1 (nx5958)) ;
    nor03_2x ix5963 (.Y (nx5962), .A0 (gen_15_cmp_mReg_5), .A1 (nx9515), .A2 (
             nx10751)) ;
    nor03_2x ix5959 (.Y (nx5958), .A0 (nx6639), .A1 (nx10757), .A2 (nx10767)) ;
    nor02_2x ix6652 (.Y (nx6651), .A0 (nx5954), .A1 (nx5952)) ;
    nor03_2x ix5955 (.Y (nx5954), .A0 (nx6654), .A1 (nx9509), .A2 (nx10775)) ;
    dffr gen_15_cmp_mRegCmp_reg_Q_6 (.Q (gen_15_cmp_mReg_6), .QB (nx6654), .D (
         window_15__6), .CLK (start), .R (rst)) ;
    nor03_2x ix5953 (.Y (nx5952), .A0 (gen_15_cmp_mReg_6), .A1 (nx10089), .A2 (
             nx10783)) ;
    nand02 ix5989 (.Y (gen_15_cmp_BSCmp_op2_7), .A0 (nx6659), .A1 (nx6665)) ;
    nor02_2x ix6660 (.Y (nx6659), .A0 (nx5984), .A1 (nx5980)) ;
    nor03_2x ix5985 (.Y (nx5984), .A0 (gen_15_cmp_mReg_6), .A1 (nx9515), .A2 (
             nx10753)) ;
    nor03_2x ix5981 (.Y (nx5980), .A0 (nx6654), .A1 (nx10759), .A2 (nx10769)) ;
    nor02_2x ix6666 (.Y (nx6665), .A0 (nx5976), .A1 (nx5974)) ;
    nor03_2x ix5977 (.Y (nx5976), .A0 (nx6669), .A1 (nx9509), .A2 (nx10777)) ;
    dffr gen_15_cmp_mRegCmp_reg_Q_7 (.Q (gen_15_cmp_mReg_7), .QB (nx6669), .D (
         window_15__7), .CLK (start), .R (rst)) ;
    nor03_2x ix5975 (.Y (nx5974), .A0 (gen_15_cmp_mReg_7), .A1 (nx10089), .A2 (
             nx10785)) ;
    nand02 ix6011 (.Y (gen_15_cmp_BSCmp_op2_8), .A0 (nx6675), .A1 (nx6679)) ;
    nor02_2x ix6676 (.Y (nx6675), .A0 (nx6006), .A1 (nx6002)) ;
    nor03_2x ix6007 (.Y (nx6006), .A0 (gen_15_cmp_mReg_7), .A1 (nx9515), .A2 (
             nx10753)) ;
    nor03_2x ix6003 (.Y (nx6002), .A0 (nx6669), .A1 (nx10759), .A2 (nx10769)) ;
    nor02_2x ix6680 (.Y (nx6679), .A0 (nx5998), .A1 (nx5996)) ;
    nor03_2x ix5999 (.Y (nx5998), .A0 (nx6683), .A1 (nx9509), .A2 (nx10777)) ;
    dffr gen_15_cmp_mRegCmp_reg_Q_8 (.Q (gen_15_cmp_mReg_8), .QB (nx6683), .D (
         window_15__8), .CLK (start), .R (rst)) ;
    nor03_2x ix5997 (.Y (nx5996), .A0 (gen_15_cmp_mReg_8), .A1 (nx10091), .A2 (
             nx10785)) ;
    nand02 ix6033 (.Y (gen_15_cmp_BSCmp_op2_9), .A0 (nx6689), .A1 (nx6695)) ;
    nor02_2x ix6690 (.Y (nx6689), .A0 (nx6028), .A1 (nx6024)) ;
    nor03_2x ix6029 (.Y (nx6028), .A0 (gen_15_cmp_mReg_8), .A1 (nx9515), .A2 (
             nx10753)) ;
    nor03_2x ix6025 (.Y (nx6024), .A0 (nx6683), .A1 (nx10759), .A2 (nx10769)) ;
    nor02_2x ix6696 (.Y (nx6695), .A0 (nx6020), .A1 (nx6018)) ;
    nor03_2x ix6021 (.Y (nx6020), .A0 (nx6698), .A1 (nx9509), .A2 (nx10777)) ;
    dffr gen_15_cmp_mRegCmp_reg_Q_9 (.Q (gen_15_cmp_mReg_9), .QB (nx6698), .D (
         window_15__9), .CLK (start), .R (rst)) ;
    nor03_2x ix6019 (.Y (nx6018), .A0 (gen_15_cmp_mReg_9), .A1 (nx10091), .A2 (
             nx10785)) ;
    nand02 ix6055 (.Y (gen_15_cmp_BSCmp_op2_10), .A0 (nx6703), .A1 (nx6709)) ;
    nor02_2x ix6704 (.Y (nx6703), .A0 (nx6050), .A1 (nx6046)) ;
    nor03_2x ix6051 (.Y (nx6050), .A0 (gen_15_cmp_mReg_9), .A1 (nx9515), .A2 (
             nx10753)) ;
    nor03_2x ix6047 (.Y (nx6046), .A0 (nx6698), .A1 (nx10759), .A2 (nx10769)) ;
    nor02_2x ix6710 (.Y (nx6709), .A0 (nx6042), .A1 (nx6040)) ;
    nor03_2x ix6043 (.Y (nx6042), .A0 (nx6713), .A1 (nx9509), .A2 (nx10777)) ;
    dffr gen_15_cmp_mRegCmp_reg_Q_10 (.Q (gen_15_cmp_mReg_10), .QB (nx6713), .D (
         window_15__10), .CLK (start), .R (rst)) ;
    nor03_2x ix6041 (.Y (nx6040), .A0 (gen_15_cmp_mReg_10), .A1 (nx10091), .A2 (
             nx10785)) ;
    nand02 ix6077 (.Y (gen_15_cmp_BSCmp_op2_11), .A0 (nx6719), .A1 (nx6723)) ;
    nor02_2x ix6720 (.Y (nx6719), .A0 (nx6072), .A1 (nx6068)) ;
    nor03_2x ix6073 (.Y (nx6072), .A0 (gen_15_cmp_mReg_10), .A1 (nx9515), .A2 (
             nx10753)) ;
    nor03_2x ix6069 (.Y (nx6068), .A0 (nx6713), .A1 (nx10759), .A2 (nx10769)) ;
    nor02_2x ix6724 (.Y (nx6723), .A0 (nx6064), .A1 (nx6062)) ;
    nor03_2x ix6065 (.Y (nx6064), .A0 (nx6727), .A1 (nx9509), .A2 (nx10777)) ;
    dffr gen_15_cmp_mRegCmp_reg_Q_11 (.Q (gen_15_cmp_mReg_11), .QB (nx6727), .D (
         window_15__11), .CLK (start), .R (rst)) ;
    nor03_2x ix6063 (.Y (nx6062), .A0 (gen_15_cmp_mReg_11), .A1 (nx10091), .A2 (
             nx10785)) ;
    nand02 ix6099 (.Y (gen_15_cmp_BSCmp_op2_12), .A0 (nx6733), .A1 (nx6739)) ;
    nor02_2x ix6734 (.Y (nx6733), .A0 (nx6094), .A1 (nx6090)) ;
    nor03_2x ix6095 (.Y (nx6094), .A0 (gen_15_cmp_mReg_11), .A1 (nx9515), .A2 (
             nx10753)) ;
    nor03_2x ix6091 (.Y (nx6090), .A0 (nx6727), .A1 (nx10759), .A2 (nx10769)) ;
    nor02_2x ix6740 (.Y (nx6739), .A0 (nx6086), .A1 (nx6084)) ;
    nor03_2x ix6087 (.Y (nx6086), .A0 (nx6742), .A1 (nx9511), .A2 (nx10777)) ;
    dffr gen_15_cmp_mRegCmp_reg_Q_12 (.Q (gen_15_cmp_mReg_12), .QB (nx6742), .D (
         window_15__12), .CLK (start), .R (rst)) ;
    nor03_2x ix6085 (.Y (nx6084), .A0 (gen_15_cmp_mReg_12), .A1 (nx10091), .A2 (
             nx10785)) ;
    nand02 ix6121 (.Y (gen_15_cmp_BSCmp_op2_13), .A0 (nx6747), .A1 (nx6753)) ;
    nor02_2x ix6748 (.Y (nx6747), .A0 (nx6116), .A1 (nx6112)) ;
    nor03_2x ix6117 (.Y (nx6116), .A0 (gen_15_cmp_mReg_12), .A1 (nx9517), .A2 (
             nx10755)) ;
    nor03_2x ix6113 (.Y (nx6112), .A0 (nx6742), .A1 (nx10759), .A2 (nx10771)) ;
    nor02_2x ix6754 (.Y (nx6753), .A0 (nx6108), .A1 (nx6106)) ;
    nor03_2x ix6109 (.Y (nx6108), .A0 (nx6757), .A1 (nx9511), .A2 (nx10779)) ;
    dffr gen_15_cmp_mRegCmp_reg_Q_13 (.Q (gen_15_cmp_mReg_13), .QB (nx6757), .D (
         window_15__13), .CLK (start), .R (rst)) ;
    nor03_2x ix6107 (.Y (nx6106), .A0 (gen_15_cmp_mReg_13), .A1 (nx10091), .A2 (
             nx10787)) ;
    nand02 ix6143 (.Y (gen_15_cmp_BSCmp_op2_14), .A0 (nx6763), .A1 (nx6767)) ;
    nor02_2x ix6764 (.Y (nx6763), .A0 (nx6138), .A1 (nx6134)) ;
    nor03_2x ix6139 (.Y (nx6138), .A0 (gen_15_cmp_mReg_13), .A1 (nx9517), .A2 (
             nx10755)) ;
    nor03_2x ix6135 (.Y (nx6134), .A0 (nx6757), .A1 (nx10761), .A2 (nx10771)) ;
    nor02_2x ix6768 (.Y (nx6767), .A0 (nx6130), .A1 (nx6128)) ;
    nor03_2x ix6131 (.Y (nx6130), .A0 (nx6771), .A1 (nx9511), .A2 (nx10779)) ;
    dffr gen_15_cmp_mRegCmp_reg_Q_14 (.Q (gen_15_cmp_mReg_14), .QB (nx6771), .D (
         window_15__14), .CLK (start), .R (rst)) ;
    nor03_2x ix6129 (.Y (nx6128), .A0 (gen_15_cmp_mReg_14), .A1 (nx10091), .A2 (
             nx10787)) ;
    nand02 ix6165 (.Y (gen_15_cmp_BSCmp_op2_15), .A0 (nx6777), .A1 (nx6783)) ;
    nor02_2x ix6778 (.Y (nx6777), .A0 (nx6160), .A1 (nx6156)) ;
    nor03_2x ix6161 (.Y (nx6160), .A0 (gen_15_cmp_mReg_14), .A1 (nx9517), .A2 (
             nx10755)) ;
    nor03_2x ix6157 (.Y (nx6156), .A0 (nx6771), .A1 (nx10761), .A2 (nx10771)) ;
    nor02_2x ix6784 (.Y (nx6783), .A0 (nx6152), .A1 (nx6150)) ;
    nor03_2x ix6153 (.Y (nx6152), .A0 (nx6786), .A1 (nx9511), .A2 (nx10779)) ;
    dffr gen_15_cmp_mRegCmp_reg_Q_15 (.Q (gen_15_cmp_mReg_15), .QB (nx6786), .D (
         window_15__15), .CLK (start), .R (rst)) ;
    nor03_2x ix6151 (.Y (nx6150), .A0 (gen_15_cmp_mReg_15), .A1 (nx10093), .A2 (
             nx10787)) ;
    nand02 ix6175 (.Y (gen_15_cmp_BSCmp_op2_16), .A0 (nx6791), .A1 (nx6783)) ;
    nor02_2x ix6792 (.Y (nx6791), .A0 (nx6170), .A1 (nx6166)) ;
    nor03_2x ix6171 (.Y (nx6170), .A0 (gen_15_cmp_mReg_15), .A1 (nx9517), .A2 (
             nx10755)) ;
    nor03_2x ix6167 (.Y (nx6166), .A0 (nx6786), .A1 (nx10761), .A2 (nx10771)) ;
    nand02 ix6243 (.Y (gen_16_cmp_BSCmp_op2_1), .A0 (nx6799), .A1 (nx6817)) ;
    nor02_2x ix6800 (.Y (nx6799), .A0 (nx6238), .A1 (nx6234)) ;
    nor03_2x ix6239 (.Y (nx6238), .A0 (gen_16_cmp_mReg_0), .A1 (nx9501), .A2 (
             nx10791)) ;
    dffr gen_16_cmp_mRegCmp_reg_Q_0 (.Q (gen_16_cmp_mReg_0), .QB (nx6805), .D (
         window_16__0), .CLK (start), .R (rst)) ;
    inv01 ix6809 (.Y (nx6808), .A (gen_16_cmp_pMux_0)) ;
    nor03_2x ix6235 (.Y (nx6234), .A0 (nx6805), .A1 (nx10797), .A2 (nx10807)) ;
    inv02 ix6816 (.Y (nx6815), .A (gen_16_cmp_pMux_2)) ;
    nor02_2x ix6818 (.Y (nx6817), .A0 (nx6224), .A1 (nx6222)) ;
    nor03_2x ix6225 (.Y (nx6224), .A0 (nx6821), .A1 (nx9495), .A2 (nx10815)) ;
    dffr gen_16_cmp_mRegCmp_reg_Q_1 (.Q (gen_16_cmp_mReg_1), .QB (nx6821), .D (
         window_16__1), .CLK (start), .R (rst)) ;
    nor03_2x ix6223 (.Y (nx6222), .A0 (gen_16_cmp_mReg_1), .A1 (nx10095), .A2 (
             nx10823)) ;
    nor03_2x ix6183 (.Y (nx6182), .A0 (nx9501), .A1 (nx6815), .A2 (
             gen_16_cmp_pMux_0)) ;
    nand02 ix6265 (.Y (gen_16_cmp_BSCmp_op2_2), .A0 (nx6832), .A1 (nx6839)) ;
    nor02_2x ix6834 (.Y (nx6832), .A0 (nx6260), .A1 (nx6256)) ;
    nor03_2x ix6261 (.Y (nx6260), .A0 (gen_16_cmp_mReg_1), .A1 (nx9501), .A2 (
             nx10791)) ;
    nor03_2x ix6257 (.Y (nx6256), .A0 (nx6821), .A1 (nx10797), .A2 (nx10807)) ;
    nor02_2x ix6840 (.Y (nx6839), .A0 (nx6252), .A1 (nx6250)) ;
    nor03_2x ix6253 (.Y (nx6252), .A0 (nx6843), .A1 (nx9495), .A2 (nx10815)) ;
    dffr gen_16_cmp_mRegCmp_reg_Q_2 (.Q (gen_16_cmp_mReg_2), .QB (nx6843), .D (
         window_16__2), .CLK (start), .R (rst)) ;
    nor03_2x ix6251 (.Y (nx6250), .A0 (gen_16_cmp_mReg_2), .A1 (nx10095), .A2 (
             nx10823)) ;
    nand02 ix6287 (.Y (gen_16_cmp_BSCmp_op2_3), .A0 (nx6849), .A1 (nx6853)) ;
    nor02_2x ix6850 (.Y (nx6849), .A0 (nx6282), .A1 (nx6278)) ;
    nor03_2x ix6283 (.Y (nx6282), .A0 (gen_16_cmp_mReg_2), .A1 (nx9501), .A2 (
             nx10791)) ;
    nor03_2x ix6279 (.Y (nx6278), .A0 (nx6843), .A1 (nx10797), .A2 (nx10807)) ;
    nor02_2x ix6854 (.Y (nx6853), .A0 (nx6274), .A1 (nx6272)) ;
    nor03_2x ix6275 (.Y (nx6274), .A0 (nx6857), .A1 (nx9495), .A2 (nx10815)) ;
    dffr gen_16_cmp_mRegCmp_reg_Q_3 (.Q (gen_16_cmp_mReg_3), .QB (nx6857), .D (
         window_16__3), .CLK (start), .R (rst)) ;
    nor03_2x ix6273 (.Y (nx6272), .A0 (gen_16_cmp_mReg_3), .A1 (nx10095), .A2 (
             nx10823)) ;
    nand02 ix6309 (.Y (gen_16_cmp_BSCmp_op2_4), .A0 (nx6863), .A1 (nx6867)) ;
    nor02_2x ix6864 (.Y (nx6863), .A0 (nx6304), .A1 (nx6300)) ;
    nor03_2x ix6305 (.Y (nx6304), .A0 (gen_16_cmp_mReg_3), .A1 (nx9501), .A2 (
             nx10791)) ;
    nor03_2x ix6301 (.Y (nx6300), .A0 (nx6857), .A1 (nx10797), .A2 (nx10807)) ;
    nor02_2x ix6868 (.Y (nx6867), .A0 (nx6296), .A1 (nx6294)) ;
    nor03_2x ix6297 (.Y (nx6296), .A0 (nx6871), .A1 (nx9495), .A2 (nx10815)) ;
    dffr gen_16_cmp_mRegCmp_reg_Q_4 (.Q (gen_16_cmp_mReg_4), .QB (nx6871), .D (
         window_16__4), .CLK (start), .R (rst)) ;
    nor03_2x ix6295 (.Y (nx6294), .A0 (gen_16_cmp_mReg_4), .A1 (nx10095), .A2 (
             nx10823)) ;
    nand02 ix6331 (.Y (gen_16_cmp_BSCmp_op2_5), .A0 (nx6875), .A1 (nx6881)) ;
    nor02_2x ix6876 (.Y (nx6875), .A0 (nx6326), .A1 (nx6322)) ;
    nor03_2x ix6327 (.Y (nx6326), .A0 (gen_16_cmp_mReg_4), .A1 (nx9501), .A2 (
             nx10791)) ;
    nor03_2x ix6323 (.Y (nx6322), .A0 (nx6871), .A1 (nx10797), .A2 (nx10807)) ;
    nor02_2x ix6882 (.Y (nx6881), .A0 (nx6318), .A1 (nx6316)) ;
    nor03_2x ix6319 (.Y (nx6318), .A0 (nx6885), .A1 (nx9497), .A2 (nx10815)) ;
    dffr gen_16_cmp_mRegCmp_reg_Q_5 (.Q (gen_16_cmp_mReg_5), .QB (nx6885), .D (
         window_16__5), .CLK (start), .R (rst)) ;
    nor03_2x ix6317 (.Y (nx6316), .A0 (gen_16_cmp_mReg_5), .A1 (nx10095), .A2 (
             nx10823)) ;
    nand02 ix6353 (.Y (gen_16_cmp_BSCmp_op2_6), .A0 (nx6889), .A1 (nx6895)) ;
    nor02_2x ix6890 (.Y (nx6889), .A0 (nx6348), .A1 (nx6344)) ;
    nor03_2x ix6349 (.Y (nx6348), .A0 (gen_16_cmp_mReg_5), .A1 (nx9503), .A2 (
             nx10791)) ;
    nor03_2x ix6345 (.Y (nx6344), .A0 (nx6885), .A1 (nx10797), .A2 (nx10807)) ;
    nor02_2x ix6896 (.Y (nx6895), .A0 (nx6340), .A1 (nx6338)) ;
    nor03_2x ix6341 (.Y (nx6340), .A0 (nx6898), .A1 (nx9497), .A2 (nx10815)) ;
    dffr gen_16_cmp_mRegCmp_reg_Q_6 (.Q (gen_16_cmp_mReg_6), .QB (nx6898), .D (
         window_16__6), .CLK (start), .R (rst)) ;
    nor03_2x ix6339 (.Y (nx6338), .A0 (gen_16_cmp_mReg_6), .A1 (nx10095), .A2 (
             nx10823)) ;
    nand02 ix6375 (.Y (gen_16_cmp_BSCmp_op2_7), .A0 (nx6905), .A1 (nx6911)) ;
    nor02_2x ix6906 (.Y (nx6905), .A0 (nx6370), .A1 (nx6366)) ;
    nor03_2x ix6371 (.Y (nx6370), .A0 (gen_16_cmp_mReg_6), .A1 (nx9503), .A2 (
             nx10793)) ;
    nor03_2x ix6367 (.Y (nx6366), .A0 (nx6898), .A1 (nx10799), .A2 (nx10809)) ;
    nor02_2x ix6912 (.Y (nx6911), .A0 (nx6362), .A1 (nx6360)) ;
    nor03_2x ix6363 (.Y (nx6362), .A0 (nx6915), .A1 (nx9497), .A2 (nx10817)) ;
    dffr gen_16_cmp_mRegCmp_reg_Q_7 (.Q (gen_16_cmp_mReg_7), .QB (nx6915), .D (
         window_16__7), .CLK (start), .R (rst)) ;
    nor03_2x ix6361 (.Y (nx6360), .A0 (gen_16_cmp_mReg_7), .A1 (nx10095), .A2 (
             nx10825)) ;
    nand02 ix6397 (.Y (gen_16_cmp_BSCmp_op2_8), .A0 (nx6919), .A1 (nx6925)) ;
    nor02_2x ix6920 (.Y (nx6919), .A0 (nx6392), .A1 (nx6388)) ;
    nor03_2x ix6393 (.Y (nx6392), .A0 (gen_16_cmp_mReg_7), .A1 (nx9503), .A2 (
             nx10793)) ;
    nor03_2x ix6389 (.Y (nx6388), .A0 (nx6915), .A1 (nx10799), .A2 (nx10809)) ;
    nor02_2x ix6926 (.Y (nx6925), .A0 (nx6384), .A1 (nx6382)) ;
    nor03_2x ix6385 (.Y (nx6384), .A0 (nx6929), .A1 (nx9497), .A2 (nx10817)) ;
    dffr gen_16_cmp_mRegCmp_reg_Q_8 (.Q (gen_16_cmp_mReg_8), .QB (nx6929), .D (
         window_16__8), .CLK (start), .R (rst)) ;
    nor03_2x ix6383 (.Y (nx6382), .A0 (gen_16_cmp_mReg_8), .A1 (nx10097), .A2 (
             nx10825)) ;
    nand02 ix6419 (.Y (gen_16_cmp_BSCmp_op2_9), .A0 (nx6933), .A1 (nx6939)) ;
    nor02_2x ix6934 (.Y (nx6933), .A0 (nx6414), .A1 (nx6410)) ;
    nor03_2x ix6415 (.Y (nx6414), .A0 (gen_16_cmp_mReg_8), .A1 (nx9503), .A2 (
             nx10793)) ;
    nor03_2x ix6411 (.Y (nx6410), .A0 (nx6929), .A1 (nx10799), .A2 (nx10809)) ;
    nor02_2x ix6940 (.Y (nx6939), .A0 (nx6406), .A1 (nx6404)) ;
    nor03_2x ix6407 (.Y (nx6406), .A0 (nx6943), .A1 (nx9497), .A2 (nx10817)) ;
    dffr gen_16_cmp_mRegCmp_reg_Q_9 (.Q (gen_16_cmp_mReg_9), .QB (nx6943), .D (
         window_16__9), .CLK (start), .R (rst)) ;
    nor03_2x ix6405 (.Y (nx6404), .A0 (gen_16_cmp_mReg_9), .A1 (nx10097), .A2 (
             nx10825)) ;
    nand02 ix6441 (.Y (gen_16_cmp_BSCmp_op2_10), .A0 (nx6949), .A1 (nx6955)) ;
    nor02_2x ix6950 (.Y (nx6949), .A0 (nx6436), .A1 (nx6432)) ;
    nor03_2x ix6437 (.Y (nx6436), .A0 (gen_16_cmp_mReg_9), .A1 (nx9503), .A2 (
             nx10793)) ;
    nor03_2x ix6433 (.Y (nx6432), .A0 (nx6943), .A1 (nx10799), .A2 (nx10809)) ;
    nor02_2x ix6956 (.Y (nx6955), .A0 (nx6428), .A1 (nx6426)) ;
    nor03_2x ix6429 (.Y (nx6428), .A0 (nx6958), .A1 (nx9497), .A2 (nx10817)) ;
    dffr gen_16_cmp_mRegCmp_reg_Q_10 (.Q (gen_16_cmp_mReg_10), .QB (nx6958), .D (
         window_16__10), .CLK (start), .R (rst)) ;
    nor03_2x ix6427 (.Y (nx6426), .A0 (gen_16_cmp_mReg_10), .A1 (nx10097), .A2 (
             nx10825)) ;
    nand02 ix6463 (.Y (gen_16_cmp_BSCmp_op2_11), .A0 (nx6962), .A1 (nx6967)) ;
    nor02_2x ix6963 (.Y (nx6962), .A0 (nx6458), .A1 (nx6454)) ;
    nor03_2x ix6459 (.Y (nx6458), .A0 (gen_16_cmp_mReg_10), .A1 (nx9503), .A2 (
             nx10793)) ;
    nor03_2x ix6455 (.Y (nx6454), .A0 (nx6958), .A1 (nx10799), .A2 (nx10809)) ;
    nor02_2x ix6968 (.Y (nx6967), .A0 (nx6450), .A1 (nx6448)) ;
    nor03_2x ix6451 (.Y (nx6450), .A0 (nx6971), .A1 (nx9497), .A2 (nx10817)) ;
    dffr gen_16_cmp_mRegCmp_reg_Q_11 (.Q (gen_16_cmp_mReg_11), .QB (nx6971), .D (
         window_16__11), .CLK (start), .R (rst)) ;
    nor03_2x ix6449 (.Y (nx6448), .A0 (gen_16_cmp_mReg_11), .A1 (nx10097), .A2 (
             nx10825)) ;
    nand02 ix6485 (.Y (gen_16_cmp_BSCmp_op2_12), .A0 (nx6977), .A1 (nx6983)) ;
    nor02_2x ix6978 (.Y (nx6977), .A0 (nx6480), .A1 (nx6476)) ;
    nor03_2x ix6481 (.Y (nx6480), .A0 (gen_16_cmp_mReg_11), .A1 (nx9503), .A2 (
             nx10793)) ;
    nor03_2x ix6477 (.Y (nx6476), .A0 (nx6971), .A1 (nx10799), .A2 (nx10809)) ;
    nor02_2x ix6984 (.Y (nx6983), .A0 (nx6472), .A1 (nx6470)) ;
    nor03_2x ix6473 (.Y (nx6472), .A0 (nx6987), .A1 (nx9499), .A2 (nx10817)) ;
    dffr gen_16_cmp_mRegCmp_reg_Q_12 (.Q (gen_16_cmp_mReg_12), .QB (nx6987), .D (
         window_16__12), .CLK (start), .R (rst)) ;
    nor03_2x ix6471 (.Y (nx6470), .A0 (gen_16_cmp_mReg_12), .A1 (nx10097), .A2 (
             nx10825)) ;
    nand02 ix6507 (.Y (gen_16_cmp_BSCmp_op2_13), .A0 (nx6991), .A1 (nx6997)) ;
    nor02_2x ix6992 (.Y (nx6991), .A0 (nx6502), .A1 (nx6498)) ;
    nor03_2x ix6503 (.Y (nx6502), .A0 (gen_16_cmp_mReg_12), .A1 (nx9505), .A2 (
             nx10795)) ;
    nor03_2x ix6499 (.Y (nx6498), .A0 (nx6987), .A1 (nx10799), .A2 (nx10811)) ;
    nor02_2x ix6998 (.Y (nx6997), .A0 (nx6494), .A1 (nx6492)) ;
    nor03_2x ix6495 (.Y (nx6494), .A0 (nx7001), .A1 (nx9499), .A2 (nx10819)) ;
    dffr gen_16_cmp_mRegCmp_reg_Q_13 (.Q (gen_16_cmp_mReg_13), .QB (nx7001), .D (
         window_16__13), .CLK (start), .R (rst)) ;
    nor03_2x ix6493 (.Y (nx6492), .A0 (gen_16_cmp_mReg_13), .A1 (nx10097), .A2 (
             nx10827)) ;
    nand02 ix6529 (.Y (gen_16_cmp_BSCmp_op2_14), .A0 (nx7007), .A1 (nx7011)) ;
    nor02_2x ix7008 (.Y (nx7007), .A0 (nx6524), .A1 (nx6520)) ;
    nor03_2x ix6525 (.Y (nx6524), .A0 (gen_16_cmp_mReg_13), .A1 (nx9505), .A2 (
             nx10795)) ;
    nor03_2x ix6521 (.Y (nx6520), .A0 (nx7001), .A1 (nx10801), .A2 (nx10811)) ;
    nor02_2x ix7012 (.Y (nx7011), .A0 (nx6516), .A1 (nx6514)) ;
    nor03_2x ix6517 (.Y (nx6516), .A0 (nx7015), .A1 (nx9499), .A2 (nx10819)) ;
    dffr gen_16_cmp_mRegCmp_reg_Q_14 (.Q (gen_16_cmp_mReg_14), .QB (nx7015), .D (
         window_16__14), .CLK (start), .R (rst)) ;
    nor03_2x ix6515 (.Y (nx6514), .A0 (gen_16_cmp_mReg_14), .A1 (nx10097), .A2 (
             nx10827)) ;
    nand02 ix6551 (.Y (gen_16_cmp_BSCmp_op2_15), .A0 (nx7019), .A1 (nx7025)) ;
    nor02_2x ix7020 (.Y (nx7019), .A0 (nx6546), .A1 (nx6542)) ;
    nor03_2x ix6547 (.Y (nx6546), .A0 (gen_16_cmp_mReg_14), .A1 (nx9505), .A2 (
             nx10795)) ;
    nor03_2x ix6543 (.Y (nx6542), .A0 (nx7015), .A1 (nx10801), .A2 (nx10811)) ;
    nor02_2x ix7026 (.Y (nx7025), .A0 (nx6538), .A1 (nx6536)) ;
    nor03_2x ix6539 (.Y (nx6538), .A0 (nx7029), .A1 (nx9499), .A2 (nx10819)) ;
    dffr gen_16_cmp_mRegCmp_reg_Q_15 (.Q (gen_16_cmp_mReg_15), .QB (nx7029), .D (
         window_16__15), .CLK (start), .R (rst)) ;
    nor03_2x ix6537 (.Y (nx6536), .A0 (gen_16_cmp_mReg_15), .A1 (nx10099), .A2 (
             nx10827)) ;
    nand02 ix6561 (.Y (gen_16_cmp_BSCmp_op2_16), .A0 (nx7033), .A1 (nx7025)) ;
    nor02_2x ix7034 (.Y (nx7033), .A0 (nx6556), .A1 (nx6552)) ;
    nor03_2x ix6557 (.Y (nx6556), .A0 (gen_16_cmp_mReg_15), .A1 (nx9505), .A2 (
             nx10795)) ;
    nor03_2x ix6553 (.Y (nx6552), .A0 (nx7029), .A1 (nx10801), .A2 (nx10811)) ;
    nand02 ix6629 (.Y (gen_17_cmp_BSCmp_op2_1), .A0 (nx7040), .A1 (nx7059)) ;
    nor02_2x ix7041 (.Y (nx7040), .A0 (nx6624), .A1 (nx6620)) ;
    nor03_2x ix6625 (.Y (nx6624), .A0 (gen_17_cmp_mReg_0), .A1 (nx9489), .A2 (
             nx10831)) ;
    dffr gen_17_cmp_mRegCmp_reg_Q_0 (.Q (gen_17_cmp_mReg_0), .QB (nx7045), .D (
         window_17__0), .CLK (start), .R (rst)) ;
    inv01 ix7050 (.Y (nx7049), .A (gen_17_cmp_pMux_0)) ;
    nor03_2x ix6621 (.Y (nx6620), .A0 (nx7045), .A1 (nx10837), .A2 (nx10847)) ;
    inv02 ix7058 (.Y (nx7057), .A (gen_17_cmp_pMux_2)) ;
    nor02_2x ix7060 (.Y (nx7059), .A0 (nx6610), .A1 (nx6608)) ;
    nor03_2x ix6611 (.Y (nx6610), .A0 (nx7062), .A1 (nx9483), .A2 (nx10855)) ;
    dffr gen_17_cmp_mRegCmp_reg_Q_1 (.Q (gen_17_cmp_mReg_1), .QB (nx7062), .D (
         window_17__1), .CLK (start), .R (rst)) ;
    nor03_2x ix6609 (.Y (nx6608), .A0 (gen_17_cmp_mReg_1), .A1 (nx10101), .A2 (
             nx10863)) ;
    nor03_2x ix6569 (.Y (nx6568), .A0 (nx9489), .A1 (nx7057), .A2 (
             gen_17_cmp_pMux_0)) ;
    nand02 ix6651 (.Y (gen_17_cmp_BSCmp_op2_2), .A0 (nx7075), .A1 (nx7081)) ;
    nor02_2x ix7076 (.Y (nx7075), .A0 (nx6646), .A1 (nx6642)) ;
    nor03_2x ix6647 (.Y (nx6646), .A0 (gen_17_cmp_mReg_1), .A1 (nx9489), .A2 (
             nx10831)) ;
    nor03_2x ix6643 (.Y (nx6642), .A0 (nx7062), .A1 (nx10837), .A2 (nx10847)) ;
    nor02_2x ix7082 (.Y (nx7081), .A0 (nx6638), .A1 (nx6636)) ;
    nor03_2x ix6639 (.Y (nx6638), .A0 (nx7084), .A1 (nx9483), .A2 (nx10855)) ;
    dffr gen_17_cmp_mRegCmp_reg_Q_2 (.Q (gen_17_cmp_mReg_2), .QB (nx7084), .D (
         window_17__2), .CLK (start), .R (rst)) ;
    nor03_2x ix6637 (.Y (nx6636), .A0 (gen_17_cmp_mReg_2), .A1 (nx10101), .A2 (
             nx10863)) ;
    nand02 ix6673 (.Y (gen_17_cmp_BSCmp_op2_3), .A0 (nx7089), .A1 (nx7095)) ;
    nor02_2x ix7090 (.Y (nx7089), .A0 (nx6668), .A1 (nx6664)) ;
    nor03_2x ix6669 (.Y (nx6668), .A0 (gen_17_cmp_mReg_2), .A1 (nx9489), .A2 (
             nx10831)) ;
    nor03_2x ix6665 (.Y (nx6664), .A0 (nx7084), .A1 (nx10837), .A2 (nx10847)) ;
    nor02_2x ix7096 (.Y (nx7095), .A0 (nx6660), .A1 (nx6658)) ;
    nor03_2x ix6661 (.Y (nx6660), .A0 (nx7099), .A1 (nx9483), .A2 (nx10855)) ;
    dffr gen_17_cmp_mRegCmp_reg_Q_3 (.Q (gen_17_cmp_mReg_3), .QB (nx7099), .D (
         window_17__3), .CLK (start), .R (rst)) ;
    nor03_2x ix6659 (.Y (nx6658), .A0 (gen_17_cmp_mReg_3), .A1 (nx10101), .A2 (
             nx10863)) ;
    nand02 ix6695 (.Y (gen_17_cmp_BSCmp_op2_4), .A0 (nx7105), .A1 (nx7109)) ;
    nor02_2x ix7106 (.Y (nx7105), .A0 (nx6690), .A1 (nx6686)) ;
    nor03_2x ix6691 (.Y (nx6690), .A0 (gen_17_cmp_mReg_3), .A1 (nx9489), .A2 (
             nx10831)) ;
    nor03_2x ix6687 (.Y (nx6686), .A0 (nx7099), .A1 (nx10837), .A2 (nx10847)) ;
    nor02_2x ix7110 (.Y (nx7109), .A0 (nx6682), .A1 (nx6680)) ;
    nor03_2x ix6683 (.Y (nx6682), .A0 (nx7113), .A1 (nx9483), .A2 (nx10855)) ;
    dffr gen_17_cmp_mRegCmp_reg_Q_4 (.Q (gen_17_cmp_mReg_4), .QB (nx7113), .D (
         window_17__4), .CLK (start), .R (rst)) ;
    nor03_2x ix6681 (.Y (nx6680), .A0 (gen_17_cmp_mReg_4), .A1 (nx10101), .A2 (
             nx10863)) ;
    nand02 ix6717 (.Y (gen_17_cmp_BSCmp_op2_5), .A0 (nx7119), .A1 (nx7125)) ;
    nor02_2x ix7120 (.Y (nx7119), .A0 (nx6712), .A1 (nx6708)) ;
    nor03_2x ix6713 (.Y (nx6712), .A0 (gen_17_cmp_mReg_4), .A1 (nx9489), .A2 (
             nx10831)) ;
    nor03_2x ix6709 (.Y (nx6708), .A0 (nx7113), .A1 (nx10837), .A2 (nx10847)) ;
    nor02_2x ix7126 (.Y (nx7125), .A0 (nx6704), .A1 (nx6702)) ;
    nor03_2x ix6705 (.Y (nx6704), .A0 (nx7128), .A1 (nx9485), .A2 (nx10855)) ;
    dffr gen_17_cmp_mRegCmp_reg_Q_5 (.Q (gen_17_cmp_mReg_5), .QB (nx7128), .D (
         window_17__5), .CLK (start), .R (rst)) ;
    nor03_2x ix6703 (.Y (nx6702), .A0 (gen_17_cmp_mReg_5), .A1 (nx10101), .A2 (
             nx10863)) ;
    nand02 ix6739 (.Y (gen_17_cmp_BSCmp_op2_6), .A0 (nx7133), .A1 (nx7139)) ;
    nor02_2x ix7134 (.Y (nx7133), .A0 (nx6734), .A1 (nx6730)) ;
    nor03_2x ix6735 (.Y (nx6734), .A0 (gen_17_cmp_mReg_5), .A1 (nx9491), .A2 (
             nx10831)) ;
    nor03_2x ix6731 (.Y (nx6730), .A0 (nx7128), .A1 (nx10837), .A2 (nx10847)) ;
    nor02_2x ix7140 (.Y (nx7139), .A0 (nx6726), .A1 (nx6724)) ;
    nor03_2x ix6727 (.Y (nx6726), .A0 (nx7143), .A1 (nx9485), .A2 (nx10855)) ;
    dffr gen_17_cmp_mRegCmp_reg_Q_6 (.Q (gen_17_cmp_mReg_6), .QB (nx7143), .D (
         window_17__6), .CLK (start), .R (rst)) ;
    nor03_2x ix6725 (.Y (nx6724), .A0 (gen_17_cmp_mReg_6), .A1 (nx10101), .A2 (
             nx10863)) ;
    nand02 ix6761 (.Y (gen_17_cmp_BSCmp_op2_7), .A0 (nx7149), .A1 (nx7153)) ;
    nor02_2x ix7150 (.Y (nx7149), .A0 (nx6756), .A1 (nx6752)) ;
    nor03_2x ix6757 (.Y (nx6756), .A0 (gen_17_cmp_mReg_6), .A1 (nx9491), .A2 (
             nx10833)) ;
    nor03_2x ix6753 (.Y (nx6752), .A0 (nx7143), .A1 (nx10839), .A2 (nx10849)) ;
    nor02_2x ix7154 (.Y (nx7153), .A0 (nx6748), .A1 (nx6746)) ;
    nor03_2x ix6749 (.Y (nx6748), .A0 (nx7157), .A1 (nx9485), .A2 (nx10857)) ;
    dffr gen_17_cmp_mRegCmp_reg_Q_7 (.Q (gen_17_cmp_mReg_7), .QB (nx7157), .D (
         window_17__7), .CLK (start), .R (rst)) ;
    nor03_2x ix6747 (.Y (nx6746), .A0 (gen_17_cmp_mReg_7), .A1 (nx10101), .A2 (
             nx10865)) ;
    nand02 ix6783 (.Y (gen_17_cmp_BSCmp_op2_8), .A0 (nx7163), .A1 (nx7169)) ;
    nor02_2x ix7164 (.Y (nx7163), .A0 (nx6778), .A1 (nx6774)) ;
    nor03_2x ix6779 (.Y (nx6778), .A0 (gen_17_cmp_mReg_7), .A1 (nx9491), .A2 (
             nx10833)) ;
    nor03_2x ix6775 (.Y (nx6774), .A0 (nx7157), .A1 (nx10839), .A2 (nx10849)) ;
    nor02_2x ix7170 (.Y (nx7169), .A0 (nx6770), .A1 (nx6768)) ;
    nor03_2x ix6771 (.Y (nx6770), .A0 (nx7172), .A1 (nx9485), .A2 (nx10857)) ;
    dffr gen_17_cmp_mRegCmp_reg_Q_8 (.Q (gen_17_cmp_mReg_8), .QB (nx7172), .D (
         window_17__8), .CLK (start), .R (rst)) ;
    nor03_2x ix6769 (.Y (nx6768), .A0 (gen_17_cmp_mReg_8), .A1 (nx10103), .A2 (
             nx10865)) ;
    nand02 ix6805 (.Y (gen_17_cmp_BSCmp_op2_9), .A0 (nx7177), .A1 (nx7183)) ;
    nor02_2x ix7178 (.Y (nx7177), .A0 (nx6800), .A1 (nx6796)) ;
    nor03_2x ix6801 (.Y (nx6800), .A0 (gen_17_cmp_mReg_8), .A1 (nx9491), .A2 (
             nx10833)) ;
    nor03_2x ix6797 (.Y (nx6796), .A0 (nx7172), .A1 (nx10839), .A2 (nx10849)) ;
    nor02_2x ix7184 (.Y (nx7183), .A0 (nx6792), .A1 (nx6790)) ;
    nor03_2x ix6793 (.Y (nx6792), .A0 (nx7187), .A1 (nx9485), .A2 (nx10857)) ;
    dffr gen_17_cmp_mRegCmp_reg_Q_9 (.Q (gen_17_cmp_mReg_9), .QB (nx7187), .D (
         window_17__9), .CLK (start), .R (rst)) ;
    nor03_2x ix6791 (.Y (nx6790), .A0 (gen_17_cmp_mReg_9), .A1 (nx10103), .A2 (
             nx10865)) ;
    nand02 ix6827 (.Y (gen_17_cmp_BSCmp_op2_10), .A0 (nx7193), .A1 (nx7197)) ;
    nor02_2x ix7194 (.Y (nx7193), .A0 (nx6822), .A1 (nx6818)) ;
    nor03_2x ix6823 (.Y (nx6822), .A0 (gen_17_cmp_mReg_9), .A1 (nx9491), .A2 (
             nx10833)) ;
    nor03_2x ix6819 (.Y (nx6818), .A0 (nx7187), .A1 (nx10839), .A2 (nx10849)) ;
    nor02_2x ix7198 (.Y (nx7197), .A0 (nx6814), .A1 (nx6812)) ;
    nor03_2x ix6815 (.Y (nx6814), .A0 (nx7201), .A1 (nx9485), .A2 (nx10857)) ;
    dffr gen_17_cmp_mRegCmp_reg_Q_10 (.Q (gen_17_cmp_mReg_10), .QB (nx7201), .D (
         window_17__10), .CLK (start), .R (rst)) ;
    nor03_2x ix6813 (.Y (nx6812), .A0 (gen_17_cmp_mReg_10), .A1 (nx10103), .A2 (
             nx10865)) ;
    nand02 ix6849 (.Y (gen_17_cmp_BSCmp_op2_11), .A0 (nx7207), .A1 (nx7213)) ;
    nor02_2x ix7208 (.Y (nx7207), .A0 (nx6844), .A1 (nx6840)) ;
    nor03_2x ix6845 (.Y (nx6844), .A0 (gen_17_cmp_mReg_10), .A1 (nx9491), .A2 (
             nx10833)) ;
    nor03_2x ix6841 (.Y (nx6840), .A0 (nx7201), .A1 (nx10839), .A2 (nx10849)) ;
    nor02_2x ix7214 (.Y (nx7213), .A0 (nx6836), .A1 (nx6834)) ;
    nor03_2x ix6837 (.Y (nx6836), .A0 (nx7216), .A1 (nx9485), .A2 (nx10857)) ;
    dffr gen_17_cmp_mRegCmp_reg_Q_11 (.Q (gen_17_cmp_mReg_11), .QB (nx7216), .D (
         window_17__11), .CLK (start), .R (rst)) ;
    nor03_2x ix6835 (.Y (nx6834), .A0 (gen_17_cmp_mReg_11), .A1 (nx10103), .A2 (
             nx10865)) ;
    nand02 ix6871 (.Y (gen_17_cmp_BSCmp_op2_12), .A0 (nx7221), .A1 (nx7227)) ;
    nor02_2x ix7222 (.Y (nx7221), .A0 (nx6866), .A1 (nx6862)) ;
    nor03_2x ix6867 (.Y (nx6866), .A0 (gen_17_cmp_mReg_11), .A1 (nx9491), .A2 (
             nx10833)) ;
    nor03_2x ix6863 (.Y (nx6862), .A0 (nx7216), .A1 (nx10839), .A2 (nx10849)) ;
    nor02_2x ix7228 (.Y (nx7227), .A0 (nx6858), .A1 (nx6856)) ;
    nor03_2x ix6859 (.Y (nx6858), .A0 (nx7231), .A1 (nx9487), .A2 (nx10857)) ;
    dffr gen_17_cmp_mRegCmp_reg_Q_12 (.Q (gen_17_cmp_mReg_12), .QB (nx7231), .D (
         window_17__12), .CLK (start), .R (rst)) ;
    nor03_2x ix6857 (.Y (nx6856), .A0 (gen_17_cmp_mReg_12), .A1 (nx10103), .A2 (
             nx10865)) ;
    nand02 ix6893 (.Y (gen_17_cmp_BSCmp_op2_13), .A0 (nx7237), .A1 (nx7241)) ;
    nor02_2x ix7238 (.Y (nx7237), .A0 (nx6888), .A1 (nx6884)) ;
    nor03_2x ix6889 (.Y (nx6888), .A0 (gen_17_cmp_mReg_12), .A1 (nx9493), .A2 (
             nx10835)) ;
    nor03_2x ix6885 (.Y (nx6884), .A0 (nx7231), .A1 (nx10839), .A2 (nx10851)) ;
    nor02_2x ix7242 (.Y (nx7241), .A0 (nx6880), .A1 (nx6878)) ;
    nor03_2x ix6881 (.Y (nx6880), .A0 (nx7245), .A1 (nx9487), .A2 (nx10859)) ;
    dffr gen_17_cmp_mRegCmp_reg_Q_13 (.Q (gen_17_cmp_mReg_13), .QB (nx7245), .D (
         window_17__13), .CLK (start), .R (rst)) ;
    nor03_2x ix6879 (.Y (nx6878), .A0 (gen_17_cmp_mReg_13), .A1 (nx10103), .A2 (
             nx10867)) ;
    nand02 ix6915 (.Y (gen_17_cmp_BSCmp_op2_14), .A0 (nx7251), .A1 (nx7257)) ;
    nor02_2x ix7252 (.Y (nx7251), .A0 (nx6910), .A1 (nx6906)) ;
    nor03_2x ix6911 (.Y (nx6910), .A0 (gen_17_cmp_mReg_13), .A1 (nx9493), .A2 (
             nx10835)) ;
    nor03_2x ix6907 (.Y (nx6906), .A0 (nx7245), .A1 (nx10841), .A2 (nx10851)) ;
    nor02_2x ix7258 (.Y (nx7257), .A0 (nx6902), .A1 (nx6900)) ;
    nor03_2x ix6903 (.Y (nx6902), .A0 (nx7260), .A1 (nx9487), .A2 (nx10859)) ;
    dffr gen_17_cmp_mRegCmp_reg_Q_14 (.Q (gen_17_cmp_mReg_14), .QB (nx7260), .D (
         window_17__14), .CLK (start), .R (rst)) ;
    nor03_2x ix6901 (.Y (nx6900), .A0 (gen_17_cmp_mReg_14), .A1 (nx10103), .A2 (
             nx10867)) ;
    nand02 ix6937 (.Y (gen_17_cmp_BSCmp_op2_15), .A0 (nx7265), .A1 (nx7271)) ;
    nor02_2x ix7266 (.Y (nx7265), .A0 (nx6932), .A1 (nx6928)) ;
    nor03_2x ix6933 (.Y (nx6932), .A0 (gen_17_cmp_mReg_14), .A1 (nx9493), .A2 (
             nx10835)) ;
    nor03_2x ix6929 (.Y (nx6928), .A0 (nx7260), .A1 (nx10841), .A2 (nx10851)) ;
    nor02_2x ix7272 (.Y (nx7271), .A0 (nx6924), .A1 (nx6922)) ;
    nor03_2x ix6925 (.Y (nx6924), .A0 (nx7275), .A1 (nx9487), .A2 (nx10859)) ;
    dffr gen_17_cmp_mRegCmp_reg_Q_15 (.Q (gen_17_cmp_mReg_15), .QB (nx7275), .D (
         window_17__15), .CLK (start), .R (rst)) ;
    nor03_2x ix6923 (.Y (nx6922), .A0 (gen_17_cmp_mReg_15), .A1 (nx10105), .A2 (
             nx10867)) ;
    nand02 ix6947 (.Y (gen_17_cmp_BSCmp_op2_16), .A0 (nx7281), .A1 (nx7271)) ;
    nor02_2x ix7282 (.Y (nx7281), .A0 (nx6942), .A1 (nx6938)) ;
    nor03_2x ix6943 (.Y (nx6942), .A0 (gen_17_cmp_mReg_15), .A1 (nx9493), .A2 (
             nx10835)) ;
    nor03_2x ix6939 (.Y (nx6938), .A0 (nx7275), .A1 (nx10841), .A2 (nx10851)) ;
    nand02 ix7015 (.Y (gen_18_cmp_BSCmp_op2_1), .A0 (nx7287), .A1 (nx7307)) ;
    nor02_2x ix7288 (.Y (nx7287), .A0 (nx7010), .A1 (nx7006)) ;
    nor03_2x ix7011 (.Y (nx7010), .A0 (gen_18_cmp_mReg_0), .A1 (nx9477), .A2 (
             nx10871)) ;
    dffr gen_18_cmp_mRegCmp_reg_Q_0 (.Q (gen_18_cmp_mReg_0), .QB (nx7293), .D (
         window_18__0), .CLK (start), .R (rst)) ;
    inv01 ix7298 (.Y (nx7297), .A (gen_18_cmp_pMux_0)) ;
    nor03_2x ix7007 (.Y (nx7006), .A0 (nx7293), .A1 (nx10877), .A2 (nx10887)) ;
    inv02 ix7306 (.Y (nx7305), .A (gen_18_cmp_pMux_2)) ;
    nor02_2x ix7308 (.Y (nx7307), .A0 (nx6996), .A1 (nx6994)) ;
    nor03_2x ix6997 (.Y (nx6996), .A0 (nx7311), .A1 (nx9471), .A2 (nx10895)) ;
    dffr gen_18_cmp_mRegCmp_reg_Q_1 (.Q (gen_18_cmp_mReg_1), .QB (nx7311), .D (
         window_18__1), .CLK (start), .R (rst)) ;
    nor03_2x ix6995 (.Y (nx6994), .A0 (gen_18_cmp_mReg_1), .A1 (nx10107), .A2 (
             nx10903)) ;
    nor03_2x ix6955 (.Y (nx6954), .A0 (nx9477), .A1 (nx7305), .A2 (
             gen_18_cmp_pMux_0)) ;
    nand02 ix7037 (.Y (gen_18_cmp_BSCmp_op2_2), .A0 (nx7323), .A1 (nx7329)) ;
    nor02_2x ix7324 (.Y (nx7323), .A0 (nx7032), .A1 (nx7028)) ;
    nor03_2x ix7033 (.Y (nx7032), .A0 (gen_18_cmp_mReg_1), .A1 (nx9477), .A2 (
             nx10871)) ;
    nor03_2x ix7029 (.Y (nx7028), .A0 (nx7311), .A1 (nx10877), .A2 (nx10887)) ;
    nor02_2x ix7330 (.Y (nx7329), .A0 (nx7024), .A1 (nx7022)) ;
    nor03_2x ix7025 (.Y (nx7024), .A0 (nx7333), .A1 (nx9471), .A2 (nx10895)) ;
    dffr gen_18_cmp_mRegCmp_reg_Q_2 (.Q (gen_18_cmp_mReg_2), .QB (nx7333), .D (
         window_18__2), .CLK (start), .R (rst)) ;
    nor03_2x ix7023 (.Y (nx7022), .A0 (gen_18_cmp_mReg_2), .A1 (nx10107), .A2 (
             nx10903)) ;
    nand02 ix7059 (.Y (gen_18_cmp_BSCmp_op2_3), .A0 (nx7339), .A1 (nx7344)) ;
    nor02_2x ix7340 (.Y (nx7339), .A0 (nx7054), .A1 (nx7050)) ;
    nor03_2x ix7055 (.Y (nx7054), .A0 (gen_18_cmp_mReg_2), .A1 (nx9477), .A2 (
             nx10871)) ;
    nor03_2x ix7051 (.Y (nx7050), .A0 (nx7333), .A1 (nx10877), .A2 (nx10887)) ;
    nor02_2x ix7345 (.Y (nx7344), .A0 (nx7046), .A1 (nx7044)) ;
    nor03_2x ix7047 (.Y (nx7046), .A0 (nx7347), .A1 (nx9471), .A2 (nx10895)) ;
    dffr gen_18_cmp_mRegCmp_reg_Q_3 (.Q (gen_18_cmp_mReg_3), .QB (nx7347), .D (
         window_18__3), .CLK (start), .R (rst)) ;
    nor03_2x ix7045 (.Y (nx7044), .A0 (gen_18_cmp_mReg_3), .A1 (nx10107), .A2 (
             nx10903)) ;
    nand02 ix7081 (.Y (gen_18_cmp_BSCmp_op2_4), .A0 (nx7351), .A1 (nx7357)) ;
    nor02_2x ix7352 (.Y (nx7351), .A0 (nx7076), .A1 (nx7072)) ;
    nor03_2x ix7077 (.Y (nx7076), .A0 (gen_18_cmp_mReg_3), .A1 (nx9477), .A2 (
             nx10871)) ;
    nor03_2x ix7073 (.Y (nx7072), .A0 (nx7347), .A1 (nx10877), .A2 (nx10887)) ;
    nor02_2x ix7358 (.Y (nx7357), .A0 (nx7068), .A1 (nx7066)) ;
    nor03_2x ix7069 (.Y (nx7068), .A0 (nx7361), .A1 (nx9471), .A2 (nx10895)) ;
    dffr gen_18_cmp_mRegCmp_reg_Q_4 (.Q (gen_18_cmp_mReg_4), .QB (nx7361), .D (
         window_18__4), .CLK (start), .R (rst)) ;
    nor03_2x ix7067 (.Y (nx7066), .A0 (gen_18_cmp_mReg_4), .A1 (nx10107), .A2 (
             nx10903)) ;
    nand02 ix7103 (.Y (gen_18_cmp_BSCmp_op2_5), .A0 (nx7367), .A1 (nx7373)) ;
    nor02_2x ix7368 (.Y (nx7367), .A0 (nx7098), .A1 (nx7094)) ;
    nor03_2x ix7099 (.Y (nx7098), .A0 (gen_18_cmp_mReg_4), .A1 (nx9477), .A2 (
             nx10871)) ;
    nor03_2x ix7095 (.Y (nx7094), .A0 (nx7361), .A1 (nx10877), .A2 (nx10887)) ;
    nor02_2x ix7374 (.Y (nx7373), .A0 (nx7090), .A1 (nx7088)) ;
    nor03_2x ix7091 (.Y (nx7090), .A0 (nx7376), .A1 (nx9473), .A2 (nx10895)) ;
    dffr gen_18_cmp_mRegCmp_reg_Q_5 (.Q (gen_18_cmp_mReg_5), .QB (nx7376), .D (
         window_18__5), .CLK (start), .R (rst)) ;
    nor03_2x ix7089 (.Y (nx7088), .A0 (gen_18_cmp_mReg_5), .A1 (nx10107), .A2 (
             nx10903)) ;
    nand02 ix7125 (.Y (gen_18_cmp_BSCmp_op2_6), .A0 (nx7381), .A1 (nx7387)) ;
    nor02_2x ix7382 (.Y (nx7381), .A0 (nx7120), .A1 (nx7116)) ;
    nor03_2x ix7121 (.Y (nx7120), .A0 (gen_18_cmp_mReg_5), .A1 (nx9479), .A2 (
             nx10871)) ;
    nor03_2x ix7117 (.Y (nx7116), .A0 (nx7376), .A1 (nx10877), .A2 (nx10887)) ;
    nor02_2x ix7388 (.Y (nx7387), .A0 (nx7112), .A1 (nx7110)) ;
    nor03_2x ix7113 (.Y (nx7112), .A0 (nx7391), .A1 (nx9473), .A2 (nx10895)) ;
    dffr gen_18_cmp_mRegCmp_reg_Q_6 (.Q (gen_18_cmp_mReg_6), .QB (nx7391), .D (
         window_18__6), .CLK (start), .R (rst)) ;
    nor03_2x ix7111 (.Y (nx7110), .A0 (gen_18_cmp_mReg_6), .A1 (nx10107), .A2 (
             nx10903)) ;
    nand02 ix7147 (.Y (gen_18_cmp_BSCmp_op2_7), .A0 (nx7397), .A1 (nx7403)) ;
    nor02_2x ix7398 (.Y (nx7397), .A0 (nx7142), .A1 (nx7138)) ;
    nor03_2x ix7143 (.Y (nx7142), .A0 (gen_18_cmp_mReg_6), .A1 (nx9479), .A2 (
             nx10873)) ;
    nor03_2x ix7139 (.Y (nx7138), .A0 (nx7391), .A1 (nx10879), .A2 (nx10889)) ;
    nor02_2x ix7404 (.Y (nx7403), .A0 (nx7134), .A1 (nx7132)) ;
    nor03_2x ix7135 (.Y (nx7134), .A0 (nx7406), .A1 (nx9473), .A2 (nx10897)) ;
    dffr gen_18_cmp_mRegCmp_reg_Q_7 (.Q (gen_18_cmp_mReg_7), .QB (nx7406), .D (
         window_18__7), .CLK (start), .R (rst)) ;
    nor03_2x ix7133 (.Y (nx7132), .A0 (gen_18_cmp_mReg_7), .A1 (nx10107), .A2 (
             nx10905)) ;
    nand02 ix7169 (.Y (gen_18_cmp_BSCmp_op2_8), .A0 (nx7413), .A1 (nx7419)) ;
    nor02_2x ix7414 (.Y (nx7413), .A0 (nx7164), .A1 (nx7160)) ;
    nor03_2x ix7165 (.Y (nx7164), .A0 (gen_18_cmp_mReg_7), .A1 (nx9479), .A2 (
             nx10873)) ;
    nor03_2x ix7161 (.Y (nx7160), .A0 (nx7406), .A1 (nx10879), .A2 (nx10889)) ;
    nor02_2x ix7420 (.Y (nx7419), .A0 (nx7156), .A1 (nx7154)) ;
    nor03_2x ix7157 (.Y (nx7156), .A0 (nx7423), .A1 (nx9473), .A2 (nx10897)) ;
    dffr gen_18_cmp_mRegCmp_reg_Q_8 (.Q (gen_18_cmp_mReg_8), .QB (nx7423), .D (
         window_18__8), .CLK (start), .R (rst)) ;
    nor03_2x ix7155 (.Y (nx7154), .A0 (gen_18_cmp_mReg_8), .A1 (nx10109), .A2 (
             nx10905)) ;
    nand02 ix7191 (.Y (gen_18_cmp_BSCmp_op2_9), .A0 (nx7427), .A1 (nx7433)) ;
    nor02_2x ix7428 (.Y (nx7427), .A0 (nx7186), .A1 (nx7182)) ;
    nor03_2x ix7187 (.Y (nx7186), .A0 (gen_18_cmp_mReg_8), .A1 (nx9479), .A2 (
             nx10873)) ;
    nor03_2x ix7183 (.Y (nx7182), .A0 (nx7423), .A1 (nx10879), .A2 (nx10889)) ;
    nor02_2x ix7434 (.Y (nx7433), .A0 (nx7178), .A1 (nx7176)) ;
    nor03_2x ix7179 (.Y (nx7178), .A0 (nx7437), .A1 (nx9473), .A2 (nx10897)) ;
    dffr gen_18_cmp_mRegCmp_reg_Q_9 (.Q (gen_18_cmp_mReg_9), .QB (nx7437), .D (
         window_18__9), .CLK (start), .R (rst)) ;
    nor03_2x ix7177 (.Y (nx7176), .A0 (gen_18_cmp_mReg_9), .A1 (nx10109), .A2 (
             nx10905)) ;
    nand02 ix7213 (.Y (gen_18_cmp_BSCmp_op2_10), .A0 (nx7441), .A1 (nx7447)) ;
    nor02_2x ix7442 (.Y (nx7441), .A0 (nx7208), .A1 (nx7204)) ;
    nor03_2x ix7209 (.Y (nx7208), .A0 (gen_18_cmp_mReg_9), .A1 (nx9479), .A2 (
             nx10873)) ;
    nor03_2x ix7205 (.Y (nx7204), .A0 (nx7437), .A1 (nx10879), .A2 (nx10889)) ;
    nor02_2x ix7448 (.Y (nx7447), .A0 (nx7200), .A1 (nx7198)) ;
    nor03_2x ix7201 (.Y (nx7200), .A0 (nx7450), .A1 (nx9473), .A2 (nx10897)) ;
    dffr gen_18_cmp_mRegCmp_reg_Q_10 (.Q (gen_18_cmp_mReg_10), .QB (nx7450), .D (
         window_18__10), .CLK (start), .R (rst)) ;
    nor03_2x ix7199 (.Y (nx7198), .A0 (gen_18_cmp_mReg_10), .A1 (nx10109), .A2 (
             nx10905)) ;
    nand02 ix7235 (.Y (gen_18_cmp_BSCmp_op2_11), .A0 (nx7457), .A1 (nx7463)) ;
    nor02_2x ix7458 (.Y (nx7457), .A0 (nx7230), .A1 (nx7226)) ;
    nor03_2x ix7231 (.Y (nx7230), .A0 (gen_18_cmp_mReg_10), .A1 (nx9479), .A2 (
             nx10873)) ;
    nor03_2x ix7227 (.Y (nx7226), .A0 (nx7450), .A1 (nx10879), .A2 (nx10889)) ;
    nor02_2x ix7464 (.Y (nx7463), .A0 (nx7222), .A1 (nx7220)) ;
    nor03_2x ix7223 (.Y (nx7222), .A0 (nx7467), .A1 (nx9473), .A2 (nx10897)) ;
    dffr gen_18_cmp_mRegCmp_reg_Q_11 (.Q (gen_18_cmp_mReg_11), .QB (nx7467), .D (
         window_18__11), .CLK (start), .R (rst)) ;
    nor03_2x ix7221 (.Y (nx7220), .A0 (gen_18_cmp_mReg_11), .A1 (nx10109), .A2 (
             nx10905)) ;
    nand02 ix7257 (.Y (gen_18_cmp_BSCmp_op2_12), .A0 (nx7471), .A1 (nx7477)) ;
    nor02_2x ix7472 (.Y (nx7471), .A0 (nx7252), .A1 (nx7248)) ;
    nor03_2x ix7253 (.Y (nx7252), .A0 (gen_18_cmp_mReg_11), .A1 (nx9479), .A2 (
             nx10873)) ;
    nor03_2x ix7249 (.Y (nx7248), .A0 (nx7467), .A1 (nx10879), .A2 (nx10889)) ;
    nor02_2x ix7478 (.Y (nx7477), .A0 (nx7244), .A1 (nx7242)) ;
    nor03_2x ix7245 (.Y (nx7244), .A0 (nx7481), .A1 (nx9475), .A2 (nx10897)) ;
    dffr gen_18_cmp_mRegCmp_reg_Q_12 (.Q (gen_18_cmp_mReg_12), .QB (nx7481), .D (
         window_18__12), .CLK (start), .R (rst)) ;
    nor03_2x ix7243 (.Y (nx7242), .A0 (gen_18_cmp_mReg_12), .A1 (nx10109), .A2 (
             nx10905)) ;
    nand02 ix7279 (.Y (gen_18_cmp_BSCmp_op2_13), .A0 (nx7485), .A1 (nx7491)) ;
    nor02_2x ix7486 (.Y (nx7485), .A0 (nx7274), .A1 (nx7270)) ;
    nor03_2x ix7275 (.Y (nx7274), .A0 (gen_18_cmp_mReg_12), .A1 (nx9481), .A2 (
             nx10875)) ;
    nor03_2x ix7271 (.Y (nx7270), .A0 (nx7481), .A1 (nx10879), .A2 (nx10891)) ;
    nor02_2x ix7492 (.Y (nx7491), .A0 (nx7266), .A1 (nx7264)) ;
    nor03_2x ix7267 (.Y (nx7266), .A0 (nx7494), .A1 (nx9475), .A2 (nx10899)) ;
    dffr gen_18_cmp_mRegCmp_reg_Q_13 (.Q (gen_18_cmp_mReg_13), .QB (nx7494), .D (
         window_18__13), .CLK (start), .R (rst)) ;
    nor03_2x ix7265 (.Y (nx7264), .A0 (gen_18_cmp_mReg_13), .A1 (nx10109), .A2 (
             nx10907)) ;
    nand02 ix7301 (.Y (gen_18_cmp_BSCmp_op2_14), .A0 (nx7501), .A1 (nx7507)) ;
    nor02_2x ix7502 (.Y (nx7501), .A0 (nx7296), .A1 (nx7292)) ;
    nor03_2x ix7297 (.Y (nx7296), .A0 (gen_18_cmp_mReg_13), .A1 (nx9481), .A2 (
             nx10875)) ;
    nor03_2x ix7293 (.Y (nx7292), .A0 (nx7494), .A1 (nx10881), .A2 (nx10891)) ;
    nor02_2x ix7508 (.Y (nx7507), .A0 (nx7288), .A1 (nx7286)) ;
    nor03_2x ix7289 (.Y (nx7288), .A0 (nx7511), .A1 (nx9475), .A2 (nx10899)) ;
    dffr gen_18_cmp_mRegCmp_reg_Q_14 (.Q (gen_18_cmp_mReg_14), .QB (nx7511), .D (
         window_18__14), .CLK (start), .R (rst)) ;
    nor03_2x ix7287 (.Y (nx7286), .A0 (gen_18_cmp_mReg_14), .A1 (nx10109), .A2 (
             nx10907)) ;
    nand02 ix7323 (.Y (gen_18_cmp_BSCmp_op2_15), .A0 (nx7515), .A1 (nx7521)) ;
    nor02_2x ix7516 (.Y (nx7515), .A0 (nx7318), .A1 (nx7314)) ;
    nor03_2x ix7319 (.Y (nx7318), .A0 (gen_18_cmp_mReg_14), .A1 (nx9481), .A2 (
             nx10875)) ;
    nor03_2x ix7315 (.Y (nx7314), .A0 (nx7511), .A1 (nx10881), .A2 (nx10891)) ;
    nor02_2x ix7522 (.Y (nx7521), .A0 (nx7310), .A1 (nx7308)) ;
    nor03_2x ix7311 (.Y (nx7310), .A0 (nx7525), .A1 (nx9475), .A2 (nx10899)) ;
    dffr gen_18_cmp_mRegCmp_reg_Q_15 (.Q (gen_18_cmp_mReg_15), .QB (nx7525), .D (
         window_18__15), .CLK (start), .R (rst)) ;
    nor03_2x ix7309 (.Y (nx7308), .A0 (gen_18_cmp_mReg_15), .A1 (nx10111), .A2 (
             nx10907)) ;
    nand02 ix7333 (.Y (gen_18_cmp_BSCmp_op2_16), .A0 (nx7529), .A1 (nx7521)) ;
    nor02_2x ix7530 (.Y (nx7529), .A0 (nx7328), .A1 (nx7324)) ;
    nor03_2x ix7329 (.Y (nx7328), .A0 (gen_18_cmp_mReg_15), .A1 (nx9481), .A2 (
             nx10875)) ;
    nor03_2x ix7325 (.Y (nx7324), .A0 (nx7525), .A1 (nx10881), .A2 (nx10891)) ;
    nand02 ix7401 (.Y (gen_19_cmp_BSCmp_op2_1), .A0 (nx7536), .A1 (nx7555)) ;
    nor02_2x ix7537 (.Y (nx7536), .A0 (nx7396), .A1 (nx7392)) ;
    nor03_2x ix7397 (.Y (nx7396), .A0 (gen_19_cmp_mReg_0), .A1 (nx9465), .A2 (
             nx10911)) ;
    dffr gen_19_cmp_mRegCmp_reg_Q_0 (.Q (gen_19_cmp_mReg_0), .QB (nx7541), .D (
         window_19__0), .CLK (start), .R (rst)) ;
    inv01 ix7546 (.Y (nx7545), .A (gen_19_cmp_pMux_0)) ;
    nor03_2x ix7393 (.Y (nx7392), .A0 (nx7541), .A1 (nx10917), .A2 (nx10927)) ;
    inv02 ix7554 (.Y (nx7553), .A (gen_19_cmp_pMux_2)) ;
    nor02_2x ix7556 (.Y (nx7555), .A0 (nx7382), .A1 (nx7380)) ;
    nor03_2x ix7383 (.Y (nx7382), .A0 (nx7558), .A1 (nx9459), .A2 (nx10935)) ;
    dffr gen_19_cmp_mRegCmp_reg_Q_1 (.Q (gen_19_cmp_mReg_1), .QB (nx7558), .D (
         window_19__1), .CLK (start), .R (rst)) ;
    nor03_2x ix7381 (.Y (nx7380), .A0 (gen_19_cmp_mReg_1), .A1 (nx10113), .A2 (
             nx10943)) ;
    nor03_2x ix7341 (.Y (nx7340), .A0 (nx9465), .A1 (nx7553), .A2 (
             gen_19_cmp_pMux_0)) ;
    nand02 ix7423 (.Y (gen_19_cmp_BSCmp_op2_2), .A0 (nx7571), .A1 (nx7577)) ;
    nor02_2x ix7572 (.Y (nx7571), .A0 (nx7418), .A1 (nx7414)) ;
    nor03_2x ix7419 (.Y (nx7418), .A0 (gen_19_cmp_mReg_1), .A1 (nx9465), .A2 (
             nx10911)) ;
    nor03_2x ix7415 (.Y (nx7414), .A0 (nx7558), .A1 (nx10917), .A2 (nx10927)) ;
    nor02_2x ix7578 (.Y (nx7577), .A0 (nx7410), .A1 (nx7408)) ;
    nor03_2x ix7411 (.Y (nx7410), .A0 (nx7580), .A1 (nx9459), .A2 (nx10935)) ;
    dffr gen_19_cmp_mRegCmp_reg_Q_2 (.Q (gen_19_cmp_mReg_2), .QB (nx7580), .D (
         window_19__2), .CLK (start), .R (rst)) ;
    nor03_2x ix7409 (.Y (nx7408), .A0 (gen_19_cmp_mReg_2), .A1 (nx10113), .A2 (
             nx10943)) ;
    nand02 ix7445 (.Y (gen_19_cmp_BSCmp_op2_3), .A0 (nx7585), .A1 (nx7591)) ;
    nor02_2x ix7586 (.Y (nx7585), .A0 (nx7440), .A1 (nx7436)) ;
    nor03_2x ix7441 (.Y (nx7440), .A0 (gen_19_cmp_mReg_2), .A1 (nx9465), .A2 (
             nx10911)) ;
    nor03_2x ix7437 (.Y (nx7436), .A0 (nx7580), .A1 (nx10917), .A2 (nx10927)) ;
    nor02_2x ix7592 (.Y (nx7591), .A0 (nx7432), .A1 (nx7430)) ;
    nor03_2x ix7433 (.Y (nx7432), .A0 (nx7595), .A1 (nx9459), .A2 (nx10935)) ;
    dffr gen_19_cmp_mRegCmp_reg_Q_3 (.Q (gen_19_cmp_mReg_3), .QB (nx7595), .D (
         window_19__3), .CLK (start), .R (rst)) ;
    nor03_2x ix7431 (.Y (nx7430), .A0 (gen_19_cmp_mReg_3), .A1 (nx10113), .A2 (
             nx10943)) ;
    nand02 ix7467 (.Y (gen_19_cmp_BSCmp_op2_4), .A0 (nx7601), .A1 (nx7605)) ;
    nor02_2x ix7602 (.Y (nx7601), .A0 (nx7462), .A1 (nx7458)) ;
    nor03_2x ix7463 (.Y (nx7462), .A0 (gen_19_cmp_mReg_3), .A1 (nx9465), .A2 (
             nx10911)) ;
    nor03_2x ix7459 (.Y (nx7458), .A0 (nx7595), .A1 (nx10917), .A2 (nx10927)) ;
    nor02_2x ix7606 (.Y (nx7605), .A0 (nx7454), .A1 (nx7452)) ;
    nor03_2x ix7455 (.Y (nx7454), .A0 (nx7609), .A1 (nx9459), .A2 (nx10935)) ;
    dffr gen_19_cmp_mRegCmp_reg_Q_4 (.Q (gen_19_cmp_mReg_4), .QB (nx7609), .D (
         window_19__4), .CLK (start), .R (rst)) ;
    nor03_2x ix7453 (.Y (nx7452), .A0 (gen_19_cmp_mReg_4), .A1 (nx10113), .A2 (
             nx10943)) ;
    nand02 ix7489 (.Y (gen_19_cmp_BSCmp_op2_5), .A0 (nx7615), .A1 (nx7621)) ;
    nor02_2x ix7616 (.Y (nx7615), .A0 (nx7484), .A1 (nx7480)) ;
    nor03_2x ix7485 (.Y (nx7484), .A0 (gen_19_cmp_mReg_4), .A1 (nx9465), .A2 (
             nx10911)) ;
    nor03_2x ix7481 (.Y (nx7480), .A0 (nx7609), .A1 (nx10917), .A2 (nx10927)) ;
    nor02_2x ix7622 (.Y (nx7621), .A0 (nx7476), .A1 (nx7474)) ;
    nor03_2x ix7477 (.Y (nx7476), .A0 (nx7624), .A1 (nx9461), .A2 (nx10935)) ;
    dffr gen_19_cmp_mRegCmp_reg_Q_5 (.Q (gen_19_cmp_mReg_5), .QB (nx7624), .D (
         window_19__5), .CLK (start), .R (rst)) ;
    nor03_2x ix7475 (.Y (nx7474), .A0 (gen_19_cmp_mReg_5), .A1 (nx10113), .A2 (
             nx10943)) ;
    nand02 ix7511 (.Y (gen_19_cmp_BSCmp_op2_6), .A0 (nx7629), .A1 (nx7635)) ;
    nor02_2x ix7630 (.Y (nx7629), .A0 (nx7506), .A1 (nx7502)) ;
    nor03_2x ix7507 (.Y (nx7506), .A0 (gen_19_cmp_mReg_5), .A1 (nx9467), .A2 (
             nx10911)) ;
    nor03_2x ix7503 (.Y (nx7502), .A0 (nx7624), .A1 (nx10917), .A2 (nx10927)) ;
    nor02_2x ix7636 (.Y (nx7635), .A0 (nx7498), .A1 (nx7496)) ;
    nor03_2x ix7499 (.Y (nx7498), .A0 (nx7639), .A1 (nx9461), .A2 (nx10935)) ;
    dffr gen_19_cmp_mRegCmp_reg_Q_6 (.Q (gen_19_cmp_mReg_6), .QB (nx7639), .D (
         window_19__6), .CLK (start), .R (rst)) ;
    nor03_2x ix7497 (.Y (nx7496), .A0 (gen_19_cmp_mReg_6), .A1 (nx10113), .A2 (
             nx10943)) ;
    nand02 ix7533 (.Y (gen_19_cmp_BSCmp_op2_7), .A0 (nx7645), .A1 (nx7649)) ;
    nor02_2x ix7646 (.Y (nx7645), .A0 (nx7528), .A1 (nx7524)) ;
    nor03_2x ix7529 (.Y (nx7528), .A0 (gen_19_cmp_mReg_6), .A1 (nx9467), .A2 (
             nx10913)) ;
    nor03_2x ix7525 (.Y (nx7524), .A0 (nx7639), .A1 (nx10919), .A2 (nx10929)) ;
    nor02_2x ix7650 (.Y (nx7649), .A0 (nx7520), .A1 (nx7518)) ;
    nor03_2x ix7521 (.Y (nx7520), .A0 (nx7653), .A1 (nx9461), .A2 (nx10937)) ;
    dffr gen_19_cmp_mRegCmp_reg_Q_7 (.Q (gen_19_cmp_mReg_7), .QB (nx7653), .D (
         window_19__7), .CLK (start), .R (rst)) ;
    nor03_2x ix7519 (.Y (nx7518), .A0 (gen_19_cmp_mReg_7), .A1 (nx10113), .A2 (
             nx10945)) ;
    nand02 ix7555 (.Y (gen_19_cmp_BSCmp_op2_8), .A0 (nx7659), .A1 (nx7665)) ;
    nor02_2x ix7660 (.Y (nx7659), .A0 (nx7550), .A1 (nx7546)) ;
    nor03_2x ix7551 (.Y (nx7550), .A0 (gen_19_cmp_mReg_7), .A1 (nx9467), .A2 (
             nx10913)) ;
    nor03_2x ix7547 (.Y (nx7546), .A0 (nx7653), .A1 (nx10919), .A2 (nx10929)) ;
    nor02_2x ix7666 (.Y (nx7665), .A0 (nx7542), .A1 (nx7540)) ;
    nor03_2x ix7543 (.Y (nx7542), .A0 (nx7668), .A1 (nx9461), .A2 (nx10937)) ;
    dffr gen_19_cmp_mRegCmp_reg_Q_8 (.Q (gen_19_cmp_mReg_8), .QB (nx7668), .D (
         window_19__8), .CLK (start), .R (rst)) ;
    nor03_2x ix7541 (.Y (nx7540), .A0 (gen_19_cmp_mReg_8), .A1 (nx10115), .A2 (
             nx10945)) ;
    nand02 ix7577 (.Y (gen_19_cmp_BSCmp_op2_9), .A0 (nx7673), .A1 (nx7679)) ;
    nor02_2x ix7674 (.Y (nx7673), .A0 (nx7572), .A1 (nx7568)) ;
    nor03_2x ix7573 (.Y (nx7572), .A0 (gen_19_cmp_mReg_8), .A1 (nx9467), .A2 (
             nx10913)) ;
    nor03_2x ix7569 (.Y (nx7568), .A0 (nx7668), .A1 (nx10919), .A2 (nx10929)) ;
    nor02_2x ix7680 (.Y (nx7679), .A0 (nx7564), .A1 (nx7562)) ;
    nor03_2x ix7565 (.Y (nx7564), .A0 (nx7683), .A1 (nx9461), .A2 (nx10937)) ;
    dffr gen_19_cmp_mRegCmp_reg_Q_9 (.Q (gen_19_cmp_mReg_9), .QB (nx7683), .D (
         window_19__9), .CLK (start), .R (rst)) ;
    nor03_2x ix7563 (.Y (nx7562), .A0 (gen_19_cmp_mReg_9), .A1 (nx10115), .A2 (
             nx10945)) ;
    nand02 ix7599 (.Y (gen_19_cmp_BSCmp_op2_10), .A0 (nx7689), .A1 (nx7693)) ;
    nor02_2x ix7690 (.Y (nx7689), .A0 (nx7594), .A1 (nx7590)) ;
    nor03_2x ix7595 (.Y (nx7594), .A0 (gen_19_cmp_mReg_9), .A1 (nx9467), .A2 (
             nx10913)) ;
    nor03_2x ix7591 (.Y (nx7590), .A0 (nx7683), .A1 (nx10919), .A2 (nx10929)) ;
    nor02_2x ix7694 (.Y (nx7693), .A0 (nx7586), .A1 (nx7584)) ;
    nor03_2x ix7587 (.Y (nx7586), .A0 (nx7697), .A1 (nx9461), .A2 (nx10937)) ;
    dffr gen_19_cmp_mRegCmp_reg_Q_10 (.Q (gen_19_cmp_mReg_10), .QB (nx7697), .D (
         window_19__10), .CLK (start), .R (rst)) ;
    nor03_2x ix7585 (.Y (nx7584), .A0 (gen_19_cmp_mReg_10), .A1 (nx10115), .A2 (
             nx10945)) ;
    nand02 ix7621 (.Y (gen_19_cmp_BSCmp_op2_11), .A0 (nx7703), .A1 (nx7709)) ;
    nor02_2x ix7704 (.Y (nx7703), .A0 (nx7616), .A1 (nx7612)) ;
    nor03_2x ix7617 (.Y (nx7616), .A0 (gen_19_cmp_mReg_10), .A1 (nx9467), .A2 (
             nx10913)) ;
    nor03_2x ix7613 (.Y (nx7612), .A0 (nx7697), .A1 (nx10919), .A2 (nx10929)) ;
    nor02_2x ix7710 (.Y (nx7709), .A0 (nx7608), .A1 (nx7606)) ;
    nor03_2x ix7609 (.Y (nx7608), .A0 (nx7713), .A1 (nx9461), .A2 (nx10937)) ;
    dffr gen_19_cmp_mRegCmp_reg_Q_11 (.Q (gen_19_cmp_mReg_11), .QB (nx7713), .D (
         window_19__11), .CLK (start), .R (rst)) ;
    nor03_2x ix7607 (.Y (nx7606), .A0 (gen_19_cmp_mReg_11), .A1 (nx10115), .A2 (
             nx10945)) ;
    nand02 ix7643 (.Y (gen_19_cmp_BSCmp_op2_12), .A0 (nx7719), .A1 (nx7725)) ;
    nor02_2x ix7720 (.Y (nx7719), .A0 (nx7638), .A1 (nx7634)) ;
    nor03_2x ix7639 (.Y (nx7638), .A0 (gen_19_cmp_mReg_11), .A1 (nx9467), .A2 (
             nx10913)) ;
    nor03_2x ix7635 (.Y (nx7634), .A0 (nx7713), .A1 (nx10919), .A2 (nx10929)) ;
    nor02_2x ix7726 (.Y (nx7725), .A0 (nx7630), .A1 (nx7628)) ;
    nor03_2x ix7631 (.Y (nx7630), .A0 (nx7729), .A1 (nx9463), .A2 (nx10937)) ;
    dffr gen_19_cmp_mRegCmp_reg_Q_12 (.Q (gen_19_cmp_mReg_12), .QB (nx7729), .D (
         window_19__12), .CLK (start), .R (rst)) ;
    nor03_2x ix7629 (.Y (nx7628), .A0 (gen_19_cmp_mReg_12), .A1 (nx10115), .A2 (
             nx10945)) ;
    nand02 ix7665 (.Y (gen_19_cmp_BSCmp_op2_13), .A0 (nx7733), .A1 (nx7737)) ;
    nor02_2x ix7734 (.Y (nx7733), .A0 (nx7660), .A1 (nx7656)) ;
    nor03_2x ix7661 (.Y (nx7660), .A0 (gen_19_cmp_mReg_12), .A1 (nx9469), .A2 (
             nx10915)) ;
    nor03_2x ix7657 (.Y (nx7656), .A0 (nx7729), .A1 (nx10919), .A2 (nx10931)) ;
    nor02_2x ix7738 (.Y (nx7737), .A0 (nx7652), .A1 (nx7650)) ;
    nor03_2x ix7653 (.Y (nx7652), .A0 (nx7741), .A1 (nx9463), .A2 (nx10939)) ;
    dffr gen_19_cmp_mRegCmp_reg_Q_13 (.Q (gen_19_cmp_mReg_13), .QB (nx7741), .D (
         window_19__13), .CLK (start), .R (rst)) ;
    nor03_2x ix7651 (.Y (nx7650), .A0 (gen_19_cmp_mReg_13), .A1 (nx10115), .A2 (
             nx10947)) ;
    nand02 ix7687 (.Y (gen_19_cmp_BSCmp_op2_14), .A0 (nx7747), .A1 (nx7753)) ;
    nor02_2x ix7748 (.Y (nx7747), .A0 (nx7682), .A1 (nx7678)) ;
    nor03_2x ix7683 (.Y (nx7682), .A0 (gen_19_cmp_mReg_13), .A1 (nx9469), .A2 (
             nx10915)) ;
    nor03_2x ix7679 (.Y (nx7678), .A0 (nx7741), .A1 (nx10921), .A2 (nx10931)) ;
    nor02_2x ix7754 (.Y (nx7753), .A0 (nx7674), .A1 (nx7672)) ;
    nor03_2x ix7675 (.Y (nx7674), .A0 (nx7757), .A1 (nx9463), .A2 (nx10939)) ;
    dffr gen_19_cmp_mRegCmp_reg_Q_14 (.Q (gen_19_cmp_mReg_14), .QB (nx7757), .D (
         window_19__14), .CLK (start), .R (rst)) ;
    nor03_2x ix7673 (.Y (nx7672), .A0 (gen_19_cmp_mReg_14), .A1 (nx10115), .A2 (
             nx10947)) ;
    nand02 ix7709 (.Y (gen_19_cmp_BSCmp_op2_15), .A0 (nx7762), .A1 (nx7767)) ;
    nor02_2x ix7763 (.Y (nx7762), .A0 (nx7704), .A1 (nx7700)) ;
    nor03_2x ix7705 (.Y (nx7704), .A0 (gen_19_cmp_mReg_14), .A1 (nx9469), .A2 (
             nx10915)) ;
    nor03_2x ix7701 (.Y (nx7700), .A0 (nx7757), .A1 (nx10921), .A2 (nx10931)) ;
    nor02_2x ix7768 (.Y (nx7767), .A0 (nx7696), .A1 (nx7694)) ;
    nor03_2x ix7697 (.Y (nx7696), .A0 (nx7771), .A1 (nx9463), .A2 (nx10939)) ;
    dffr gen_19_cmp_mRegCmp_reg_Q_15 (.Q (gen_19_cmp_mReg_15), .QB (nx7771), .D (
         window_19__15), .CLK (start), .R (rst)) ;
    nor03_2x ix7695 (.Y (nx7694), .A0 (gen_19_cmp_mReg_15), .A1 (nx10117), .A2 (
             nx10947)) ;
    nand02 ix7719 (.Y (gen_19_cmp_BSCmp_op2_16), .A0 (nx7775), .A1 (nx7767)) ;
    nor02_2x ix7776 (.Y (nx7775), .A0 (nx7714), .A1 (nx7710)) ;
    nor03_2x ix7715 (.Y (nx7714), .A0 (gen_19_cmp_mReg_15), .A1 (nx9469), .A2 (
             nx10915)) ;
    nor03_2x ix7711 (.Y (nx7710), .A0 (nx7771), .A1 (nx10921), .A2 (nx10931)) ;
    nand02 ix7787 (.Y (gen_20_cmp_BSCmp_op2_1), .A0 (nx7783), .A1 (nx7803)) ;
    nor02_2x ix7784 (.Y (nx7783), .A0 (nx7782), .A1 (nx7778)) ;
    nor03_2x ix7783 (.Y (nx7782), .A0 (gen_20_cmp_mReg_0), .A1 (nx9453), .A2 (
             nx10951)) ;
    dffr gen_20_cmp_mRegCmp_reg_Q_0 (.Q (gen_20_cmp_mReg_0), .QB (nx7789), .D (
         window_20__0), .CLK (start), .R (rst)) ;
    inv01 ix7794 (.Y (nx7792), .A (gen_20_cmp_pMux_0)) ;
    nor03_2x ix7779 (.Y (nx7778), .A0 (nx7789), .A1 (nx10957), .A2 (nx10967)) ;
    inv02 ix7802 (.Y (nx7801), .A (gen_20_cmp_pMux_2)) ;
    nor02_2x ix7804 (.Y (nx7803), .A0 (nx7768), .A1 (nx7766)) ;
    nor03_2x ix7769 (.Y (nx7768), .A0 (nx7807), .A1 (nx9447), .A2 (nx10975)) ;
    dffr gen_20_cmp_mRegCmp_reg_Q_1 (.Q (gen_20_cmp_mReg_1), .QB (nx7807), .D (
         window_20__1), .CLK (start), .R (rst)) ;
    nor03_2x ix7767 (.Y (nx7766), .A0 (gen_20_cmp_mReg_1), .A1 (nx10119), .A2 (
             nx10983)) ;
    nor03_2x ix7727 (.Y (nx7726), .A0 (nx9453), .A1 (nx7801), .A2 (
             gen_20_cmp_pMux_0)) ;
    nand02 ix7809 (.Y (gen_20_cmp_BSCmp_op2_2), .A0 (nx7817), .A1 (nx7823)) ;
    nor02_2x ix7818 (.Y (nx7817), .A0 (nx7804), .A1 (nx7800)) ;
    nor03_2x ix7805 (.Y (nx7804), .A0 (gen_20_cmp_mReg_1), .A1 (nx9453), .A2 (
             nx10951)) ;
    nor03_2x ix7801 (.Y (nx7800), .A0 (nx7807), .A1 (nx10957), .A2 (nx10967)) ;
    nor02_2x ix7824 (.Y (nx7823), .A0 (nx7796), .A1 (nx7794)) ;
    nor03_2x ix7797 (.Y (nx7796), .A0 (nx7827), .A1 (nx9447), .A2 (nx10975)) ;
    dffr gen_20_cmp_mRegCmp_reg_Q_2 (.Q (gen_20_cmp_mReg_2), .QB (nx7827), .D (
         window_20__2), .CLK (start), .R (rst)) ;
    nor03_2x ix7795 (.Y (nx7794), .A0 (gen_20_cmp_mReg_2), .A1 (nx10119), .A2 (
             nx10983)) ;
    nand02 ix7831 (.Y (gen_20_cmp_BSCmp_op2_3), .A0 (nx7833), .A1 (nx7837)) ;
    nor02_2x ix7834 (.Y (nx7833), .A0 (nx7826), .A1 (nx7822)) ;
    nor03_2x ix7827 (.Y (nx7826), .A0 (gen_20_cmp_mReg_2), .A1 (nx9453), .A2 (
             nx10951)) ;
    nor03_2x ix7823 (.Y (nx7822), .A0 (nx7827), .A1 (nx10957), .A2 (nx10967)) ;
    nor02_2x ix7838 (.Y (nx7837), .A0 (nx7818), .A1 (nx7816)) ;
    nor03_2x ix7819 (.Y (nx7818), .A0 (nx7841), .A1 (nx9447), .A2 (nx10975)) ;
    dffr gen_20_cmp_mRegCmp_reg_Q_3 (.Q (gen_20_cmp_mReg_3), .QB (nx7841), .D (
         window_20__3), .CLK (start), .R (rst)) ;
    nor03_2x ix7817 (.Y (nx7816), .A0 (gen_20_cmp_mReg_3), .A1 (nx10119), .A2 (
             nx10983)) ;
    nand02 ix7853 (.Y (gen_20_cmp_BSCmp_op2_4), .A0 (nx7847), .A1 (nx7853)) ;
    nor02_2x ix7848 (.Y (nx7847), .A0 (nx7848), .A1 (nx7844)) ;
    nor03_2x ix7849 (.Y (nx7848), .A0 (gen_20_cmp_mReg_3), .A1 (nx9453), .A2 (
             nx10951)) ;
    nor03_2x ix7845 (.Y (nx7844), .A0 (nx7841), .A1 (nx10957), .A2 (nx10967)) ;
    nor02_2x ix7854 (.Y (nx7853), .A0 (nx7840), .A1 (nx7838)) ;
    nor03_2x ix7841 (.Y (nx7840), .A0 (nx7856), .A1 (nx9447), .A2 (nx10975)) ;
    dffr gen_20_cmp_mRegCmp_reg_Q_4 (.Q (gen_20_cmp_mReg_4), .QB (nx7856), .D (
         window_20__4), .CLK (start), .R (rst)) ;
    nor03_2x ix7839 (.Y (nx7838), .A0 (gen_20_cmp_mReg_4), .A1 (nx10119), .A2 (
             nx10983)) ;
    nand02 ix7875 (.Y (gen_20_cmp_BSCmp_op2_5), .A0 (nx7861), .A1 (nx7867)) ;
    nor02_2x ix7862 (.Y (nx7861), .A0 (nx7870), .A1 (nx7866)) ;
    nor03_2x ix7871 (.Y (nx7870), .A0 (gen_20_cmp_mReg_4), .A1 (nx9453), .A2 (
             nx10951)) ;
    nor03_2x ix7867 (.Y (nx7866), .A0 (nx7856), .A1 (nx10957), .A2 (nx10967)) ;
    nor02_2x ix7868 (.Y (nx7867), .A0 (nx7862), .A1 (nx7860)) ;
    nor03_2x ix7863 (.Y (nx7862), .A0 (nx7871), .A1 (nx9449), .A2 (nx10975)) ;
    dffr gen_20_cmp_mRegCmp_reg_Q_5 (.Q (gen_20_cmp_mReg_5), .QB (nx7871), .D (
         window_20__5), .CLK (start), .R (rst)) ;
    nor03_2x ix7861 (.Y (nx7860), .A0 (gen_20_cmp_mReg_5), .A1 (nx10119), .A2 (
             nx10983)) ;
    nand02 ix7897 (.Y (gen_20_cmp_BSCmp_op2_6), .A0 (nx7877), .A1 (nx7881)) ;
    nor02_2x ix7878 (.Y (nx7877), .A0 (nx7892), .A1 (nx7888)) ;
    nor03_2x ix7893 (.Y (nx7892), .A0 (gen_20_cmp_mReg_5), .A1 (nx9455), .A2 (
             nx10951)) ;
    nor03_2x ix7889 (.Y (nx7888), .A0 (nx7871), .A1 (nx10957), .A2 (nx10967)) ;
    nor02_2x ix7882 (.Y (nx7881), .A0 (nx7884), .A1 (nx7882)) ;
    nor03_2x ix7885 (.Y (nx7884), .A0 (nx7885), .A1 (nx9449), .A2 (nx10975)) ;
    dffr gen_20_cmp_mRegCmp_reg_Q_6 (.Q (gen_20_cmp_mReg_6), .QB (nx7885), .D (
         window_20__6), .CLK (start), .R (rst)) ;
    nor03_2x ix7883 (.Y (nx7882), .A0 (gen_20_cmp_mReg_6), .A1 (nx10119), .A2 (
             nx10983)) ;
    nand02 ix7919 (.Y (gen_20_cmp_BSCmp_op2_7), .A0 (nx7891), .A1 (nx7897)) ;
    nor02_2x ix7892 (.Y (nx7891), .A0 (nx7914), .A1 (nx7910)) ;
    nor03_2x ix7915 (.Y (nx7914), .A0 (gen_20_cmp_mReg_6), .A1 (nx9455), .A2 (
             nx10953)) ;
    nor03_2x ix7911 (.Y (nx7910), .A0 (nx7885), .A1 (nx10959), .A2 (nx10969)) ;
    nor02_2x ix7898 (.Y (nx7897), .A0 (nx7906), .A1 (nx7904)) ;
    nor03_2x ix7907 (.Y (nx7906), .A0 (nx7900), .A1 (nx9449), .A2 (nx10977)) ;
    dffr gen_20_cmp_mRegCmp_reg_Q_7 (.Q (gen_20_cmp_mReg_7), .QB (nx7900), .D (
         window_20__7), .CLK (start), .R (rst)) ;
    nor03_2x ix7905 (.Y (nx7904), .A0 (gen_20_cmp_mReg_7), .A1 (nx10119), .A2 (
             nx10985)) ;
    nand02 ix7941 (.Y (gen_20_cmp_BSCmp_op2_8), .A0 (nx7905), .A1 (nx7911)) ;
    nor02_2x ix7906 (.Y (nx7905), .A0 (nx7936), .A1 (nx7932)) ;
    nor03_2x ix7937 (.Y (nx7936), .A0 (gen_20_cmp_mReg_7), .A1 (nx9455), .A2 (
             nx10953)) ;
    nor03_2x ix7933 (.Y (nx7932), .A0 (nx7900), .A1 (nx10959), .A2 (nx10969)) ;
    nor02_2x ix7912 (.Y (nx7911), .A0 (nx7928), .A1 (nx7926)) ;
    nor03_2x ix7929 (.Y (nx7928), .A0 (nx7915), .A1 (nx9449), .A2 (nx10977)) ;
    dffr gen_20_cmp_mRegCmp_reg_Q_8 (.Q (gen_20_cmp_mReg_8), .QB (nx7915), .D (
         window_20__8), .CLK (start), .R (rst)) ;
    nor03_2x ix7927 (.Y (nx7926), .A0 (gen_20_cmp_mReg_8), .A1 (nx10121), .A2 (
             nx10985)) ;
    nand02 ix7963 (.Y (gen_20_cmp_BSCmp_op2_9), .A0 (nx7921), .A1 (nx7925)) ;
    nor02_2x ix7922 (.Y (nx7921), .A0 (nx7958), .A1 (nx7954)) ;
    nor03_2x ix7959 (.Y (nx7958), .A0 (gen_20_cmp_mReg_8), .A1 (nx9455), .A2 (
             nx10953)) ;
    nor03_2x ix7955 (.Y (nx7954), .A0 (nx7915), .A1 (nx10959), .A2 (nx10969)) ;
    nor02_2x ix7926 (.Y (nx7925), .A0 (nx7950), .A1 (nx7948)) ;
    nor03_2x ix7951 (.Y (nx7950), .A0 (nx7929), .A1 (nx9449), .A2 (nx10977)) ;
    dffr gen_20_cmp_mRegCmp_reg_Q_9 (.Q (gen_20_cmp_mReg_9), .QB (nx7929), .D (
         window_20__9), .CLK (start), .R (rst)) ;
    nor03_2x ix7949 (.Y (nx7948), .A0 (gen_20_cmp_mReg_9), .A1 (nx10121), .A2 (
             nx10985)) ;
    nand02 ix7985 (.Y (gen_20_cmp_BSCmp_op2_10), .A0 (nx7935), .A1 (nx7941)) ;
    nor02_2x ix7936 (.Y (nx7935), .A0 (nx7980), .A1 (nx7976)) ;
    nor03_2x ix7981 (.Y (nx7980), .A0 (gen_20_cmp_mReg_9), .A1 (nx9455), .A2 (
             nx10953)) ;
    nor03_2x ix7977 (.Y (nx7976), .A0 (nx7929), .A1 (nx10959), .A2 (nx10969)) ;
    nor02_2x ix7942 (.Y (nx7941), .A0 (nx7972), .A1 (nx7970)) ;
    nor03_2x ix7973 (.Y (nx7972), .A0 (nx7944), .A1 (nx9449), .A2 (nx10977)) ;
    dffr gen_20_cmp_mRegCmp_reg_Q_10 (.Q (gen_20_cmp_mReg_10), .QB (nx7944), .D (
         window_20__10), .CLK (start), .R (rst)) ;
    nor03_2x ix7971 (.Y (nx7970), .A0 (gen_20_cmp_mReg_10), .A1 (nx10121), .A2 (
             nx10985)) ;
    nand02 ix8007 (.Y (gen_20_cmp_BSCmp_op2_11), .A0 (nx7949), .A1 (nx7955)) ;
    nor02_2x ix7950 (.Y (nx7949), .A0 (nx8002), .A1 (nx7998)) ;
    nor03_2x ix8003 (.Y (nx8002), .A0 (gen_20_cmp_mReg_10), .A1 (nx9455), .A2 (
             nx10953)) ;
    nor03_2x ix7999 (.Y (nx7998), .A0 (nx7944), .A1 (nx10959), .A2 (nx10969)) ;
    nor02_2x ix7956 (.Y (nx7955), .A0 (nx7994), .A1 (nx7992)) ;
    nor03_2x ix7995 (.Y (nx7994), .A0 (nx7959), .A1 (nx9449), .A2 (nx10977)) ;
    dffr gen_20_cmp_mRegCmp_reg_Q_11 (.Q (gen_20_cmp_mReg_11), .QB (nx7959), .D (
         window_20__11), .CLK (start), .R (rst)) ;
    nor03_2x ix7993 (.Y (nx7992), .A0 (gen_20_cmp_mReg_11), .A1 (nx10121), .A2 (
             nx10985)) ;
    nand02 ix8029 (.Y (gen_20_cmp_BSCmp_op2_12), .A0 (nx7965), .A1 (nx7969)) ;
    nor02_2x ix7966 (.Y (nx7965), .A0 (nx8024), .A1 (nx8020)) ;
    nor03_2x ix8025 (.Y (nx8024), .A0 (gen_20_cmp_mReg_11), .A1 (nx9455), .A2 (
             nx10953)) ;
    nor03_2x ix8021 (.Y (nx8020), .A0 (nx7959), .A1 (nx10959), .A2 (nx10969)) ;
    nor02_2x ix7970 (.Y (nx7969), .A0 (nx8016), .A1 (nx8014)) ;
    nor03_2x ix8017 (.Y (nx8016), .A0 (nx7973), .A1 (nx9451), .A2 (nx10977)) ;
    dffr gen_20_cmp_mRegCmp_reg_Q_12 (.Q (gen_20_cmp_mReg_12), .QB (nx7973), .D (
         window_20__12), .CLK (start), .R (rst)) ;
    nor03_2x ix8015 (.Y (nx8014), .A0 (gen_20_cmp_mReg_12), .A1 (nx10121), .A2 (
             nx10985)) ;
    nand02 ix8051 (.Y (gen_20_cmp_BSCmp_op2_13), .A0 (nx7979), .A1 (nx7985)) ;
    nor02_2x ix7980 (.Y (nx7979), .A0 (nx8046), .A1 (nx8042)) ;
    nor03_2x ix8047 (.Y (nx8046), .A0 (gen_20_cmp_mReg_12), .A1 (nx9457), .A2 (
             nx10955)) ;
    nor03_2x ix8043 (.Y (nx8042), .A0 (nx7973), .A1 (nx10959), .A2 (nx10971)) ;
    nor02_2x ix7986 (.Y (nx7985), .A0 (nx8038), .A1 (nx8036)) ;
    nor03_2x ix8039 (.Y (nx8038), .A0 (nx7988), .A1 (nx9451), .A2 (nx10979)) ;
    dffr gen_20_cmp_mRegCmp_reg_Q_13 (.Q (gen_20_cmp_mReg_13), .QB (nx7988), .D (
         window_20__13), .CLK (start), .R (rst)) ;
    nor03_2x ix8037 (.Y (nx8036), .A0 (gen_20_cmp_mReg_13), .A1 (nx10121), .A2 (
             nx10987)) ;
    nand02 ix8073 (.Y (gen_20_cmp_BSCmp_op2_14), .A0 (nx7993), .A1 (nx7999)) ;
    nor02_2x ix7994 (.Y (nx7993), .A0 (nx8068), .A1 (nx8064)) ;
    nor03_2x ix8069 (.Y (nx8068), .A0 (gen_20_cmp_mReg_13), .A1 (nx9457), .A2 (
             nx10955)) ;
    nor03_2x ix8065 (.Y (nx8064), .A0 (nx7988), .A1 (nx10961), .A2 (nx10971)) ;
    nor02_2x ix8000 (.Y (nx7999), .A0 (nx8060), .A1 (nx8058)) ;
    nor03_2x ix8061 (.Y (nx8060), .A0 (nx8003), .A1 (nx9451), .A2 (nx10979)) ;
    dffr gen_20_cmp_mRegCmp_reg_Q_14 (.Q (gen_20_cmp_mReg_14), .QB (nx8003), .D (
         window_20__14), .CLK (start), .R (rst)) ;
    nor03_2x ix8059 (.Y (nx8058), .A0 (gen_20_cmp_mReg_14), .A1 (nx10121), .A2 (
             nx10987)) ;
    nand02 ix8095 (.Y (gen_20_cmp_BSCmp_op2_15), .A0 (nx8009), .A1 (nx8013)) ;
    nor02_2x ix8010 (.Y (nx8009), .A0 (nx8090), .A1 (nx8086)) ;
    nor03_2x ix8091 (.Y (nx8090), .A0 (gen_20_cmp_mReg_14), .A1 (nx9457), .A2 (
             nx10955)) ;
    nor03_2x ix8087 (.Y (nx8086), .A0 (nx8003), .A1 (nx10961), .A2 (nx10971)) ;
    nor02_2x ix8014 (.Y (nx8013), .A0 (nx8082), .A1 (nx8080)) ;
    nor03_2x ix8083 (.Y (nx8082), .A0 (nx8017), .A1 (nx9451), .A2 (nx10979)) ;
    dffr gen_20_cmp_mRegCmp_reg_Q_15 (.Q (gen_20_cmp_mReg_15), .QB (nx8017), .D (
         window_20__15), .CLK (start), .R (rst)) ;
    nor03_2x ix8081 (.Y (nx8080), .A0 (gen_20_cmp_mReg_15), .A1 (nx10123), .A2 (
             nx10987)) ;
    nand02 ix8105 (.Y (gen_20_cmp_BSCmp_op2_16), .A0 (nx8023), .A1 (nx8013)) ;
    nor02_2x ix8024 (.Y (nx8023), .A0 (nx8100), .A1 (nx8096)) ;
    nor03_2x ix8101 (.Y (nx8100), .A0 (gen_20_cmp_mReg_15), .A1 (nx9457), .A2 (
             nx10955)) ;
    nor03_2x ix8097 (.Y (nx8096), .A0 (nx8017), .A1 (nx10961), .A2 (nx10971)) ;
    nand02 ix8173 (.Y (gen_21_cmp_BSCmp_op2_1), .A0 (nx8031), .A1 (nx8049)) ;
    nor02_2x ix8032 (.Y (nx8031), .A0 (nx8168), .A1 (nx8164)) ;
    nor03_2x ix8169 (.Y (nx8168), .A0 (gen_21_cmp_mReg_0), .A1 (nx9441), .A2 (
             nx10991)) ;
    dffr gen_21_cmp_mRegCmp_reg_Q_0 (.Q (gen_21_cmp_mReg_0), .QB (nx8035), .D (
         window_21__0), .CLK (start), .R (rst)) ;
    inv01 ix8040 (.Y (nx8039), .A (gen_21_cmp_pMux_0)) ;
    nor03_2x ix8165 (.Y (nx8164), .A0 (nx8035), .A1 (nx10997), .A2 (nx11007)) ;
    inv02 ix8048 (.Y (nx8047), .A (gen_21_cmp_pMux_2)) ;
    nor02_2x ix8050 (.Y (nx8049), .A0 (nx8154), .A1 (nx8152)) ;
    nor03_2x ix8155 (.Y (nx8154), .A0 (nx8053), .A1 (nx9435), .A2 (nx11015)) ;
    dffr gen_21_cmp_mRegCmp_reg_Q_1 (.Q (gen_21_cmp_mReg_1), .QB (nx8053), .D (
         window_21__1), .CLK (start), .R (rst)) ;
    nor03_2x ix8153 (.Y (nx8152), .A0 (gen_21_cmp_mReg_1), .A1 (nx10125), .A2 (
             nx11023)) ;
    nor03_2x ix8113 (.Y (nx8112), .A0 (nx9441), .A1 (nx8047), .A2 (
             gen_21_cmp_pMux_0)) ;
    nand02 ix8195 (.Y (gen_21_cmp_BSCmp_op2_2), .A0 (nx8065), .A1 (nx8069)) ;
    nor02_2x ix8066 (.Y (nx8065), .A0 (nx8190), .A1 (nx8186)) ;
    nor03_2x ix8191 (.Y (nx8190), .A0 (gen_21_cmp_mReg_1), .A1 (nx9441), .A2 (
             nx10991)) ;
    nor03_2x ix8187 (.Y (nx8186), .A0 (nx8053), .A1 (nx10997), .A2 (nx11007)) ;
    nor02_2x ix8070 (.Y (nx8069), .A0 (nx8182), .A1 (nx8180)) ;
    nor03_2x ix8183 (.Y (nx8182), .A0 (nx8073), .A1 (nx9435), .A2 (nx11015)) ;
    dffr gen_21_cmp_mRegCmp_reg_Q_2 (.Q (gen_21_cmp_mReg_2), .QB (nx8073), .D (
         window_21__2), .CLK (start), .R (rst)) ;
    nor03_2x ix8181 (.Y (nx8180), .A0 (gen_21_cmp_mReg_2), .A1 (nx10125), .A2 (
             nx11023)) ;
    nand02 ix8217 (.Y (gen_21_cmp_BSCmp_op2_3), .A0 (nx8077), .A1 (nx8083)) ;
    nor02_2x ix8078 (.Y (nx8077), .A0 (nx8212), .A1 (nx8208)) ;
    nor03_2x ix8213 (.Y (nx8212), .A0 (gen_21_cmp_mReg_2), .A1 (nx9441), .A2 (
             nx10991)) ;
    nor03_2x ix8209 (.Y (nx8208), .A0 (nx8073), .A1 (nx10997), .A2 (nx11007)) ;
    nor02_2x ix8084 (.Y (nx8083), .A0 (nx8204), .A1 (nx8202)) ;
    nor03_2x ix8205 (.Y (nx8204), .A0 (nx8087), .A1 (nx9435), .A2 (nx11015)) ;
    dffr gen_21_cmp_mRegCmp_reg_Q_3 (.Q (gen_21_cmp_mReg_3), .QB (nx8087), .D (
         window_21__3), .CLK (start), .R (rst)) ;
    nor03_2x ix8203 (.Y (nx8202), .A0 (gen_21_cmp_mReg_3), .A1 (nx10125), .A2 (
             nx11023)) ;
    nand02 ix8239 (.Y (gen_21_cmp_BSCmp_op2_4), .A0 (nx8091), .A1 (nx8097)) ;
    nor02_2x ix8092 (.Y (nx8091), .A0 (nx8234), .A1 (nx8230)) ;
    nor03_2x ix8235 (.Y (nx8234), .A0 (gen_21_cmp_mReg_3), .A1 (nx9441), .A2 (
             nx10991)) ;
    nor03_2x ix8231 (.Y (nx8230), .A0 (nx8087), .A1 (nx10997), .A2 (nx11007)) ;
    nor02_2x ix8098 (.Y (nx8097), .A0 (nx8226), .A1 (nx8224)) ;
    nor03_2x ix8227 (.Y (nx8226), .A0 (nx8101), .A1 (nx9435), .A2 (nx11015)) ;
    dffr gen_21_cmp_mRegCmp_reg_Q_4 (.Q (gen_21_cmp_mReg_4), .QB (nx8101), .D (
         window_21__4), .CLK (start), .R (rst)) ;
    nor03_2x ix8225 (.Y (nx8224), .A0 (gen_21_cmp_mReg_4), .A1 (nx10125), .A2 (
             nx11023)) ;
    nand02 ix8261 (.Y (gen_21_cmp_BSCmp_op2_5), .A0 (nx8107), .A1 (nx8113)) ;
    nor02_2x ix8108 (.Y (nx8107), .A0 (nx8256), .A1 (nx8252)) ;
    nor03_2x ix8257 (.Y (nx8256), .A0 (gen_21_cmp_mReg_4), .A1 (nx9441), .A2 (
             nx10991)) ;
    nor03_2x ix8253 (.Y (nx8252), .A0 (nx8101), .A1 (nx10997), .A2 (nx11007)) ;
    nor02_2x ix8114 (.Y (nx8113), .A0 (nx8248), .A1 (nx8246)) ;
    nor03_2x ix8249 (.Y (nx8248), .A0 (nx8116), .A1 (nx9437), .A2 (nx11015)) ;
    dffr gen_21_cmp_mRegCmp_reg_Q_5 (.Q (gen_21_cmp_mReg_5), .QB (nx8116), .D (
         window_21__5), .CLK (start), .R (rst)) ;
    nor03_2x ix8247 (.Y (nx8246), .A0 (gen_21_cmp_mReg_5), .A1 (nx10125), .A2 (
             nx11023)) ;
    nand02 ix8283 (.Y (gen_21_cmp_BSCmp_op2_6), .A0 (nx8120), .A1 (nx8125)) ;
    nor02_2x ix8121 (.Y (nx8120), .A0 (nx8278), .A1 (nx8274)) ;
    nor03_2x ix8279 (.Y (nx8278), .A0 (gen_21_cmp_mReg_5), .A1 (nx9443), .A2 (
             nx10991)) ;
    nor03_2x ix8275 (.Y (nx8274), .A0 (nx8116), .A1 (nx10997), .A2 (nx11007)) ;
    nor02_2x ix8126 (.Y (nx8125), .A0 (nx8270), .A1 (nx8268)) ;
    nor03_2x ix8271 (.Y (nx8270), .A0 (nx8129), .A1 (nx9437), .A2 (nx11015)) ;
    dffr gen_21_cmp_mRegCmp_reg_Q_6 (.Q (gen_21_cmp_mReg_6), .QB (nx8129), .D (
         window_21__6), .CLK (start), .R (rst)) ;
    nor03_2x ix8269 (.Y (nx8268), .A0 (gen_21_cmp_mReg_6), .A1 (nx10125), .A2 (
             nx11023)) ;
    nand02 ix8305 (.Y (gen_21_cmp_BSCmp_op2_7), .A0 (nx8135), .A1 (nx8141)) ;
    nor02_2x ix8136 (.Y (nx8135), .A0 (nx8300), .A1 (nx8296)) ;
    nor03_2x ix8301 (.Y (nx8300), .A0 (gen_21_cmp_mReg_6), .A1 (nx9443), .A2 (
             nx10993)) ;
    nor03_2x ix8297 (.Y (nx8296), .A0 (nx8129), .A1 (nx10999), .A2 (nx11009)) ;
    nor02_2x ix8142 (.Y (nx8141), .A0 (nx8292), .A1 (nx8290)) ;
    nor03_2x ix8293 (.Y (nx8292), .A0 (nx8145), .A1 (nx9437), .A2 (nx11017)) ;
    dffr gen_21_cmp_mRegCmp_reg_Q_7 (.Q (gen_21_cmp_mReg_7), .QB (nx8145), .D (
         window_21__7), .CLK (start), .R (rst)) ;
    nor03_2x ix8291 (.Y (nx8290), .A0 (gen_21_cmp_mReg_7), .A1 (nx10125), .A2 (
             nx11025)) ;
    nand02 ix8327 (.Y (gen_21_cmp_BSCmp_op2_8), .A0 (nx8149), .A1 (nx8155)) ;
    nor02_2x ix8150 (.Y (nx8149), .A0 (nx8322), .A1 (nx8318)) ;
    nor03_2x ix8323 (.Y (nx8322), .A0 (gen_21_cmp_mReg_7), .A1 (nx9443), .A2 (
             nx10993)) ;
    nor03_2x ix8319 (.Y (nx8318), .A0 (nx8145), .A1 (nx10999), .A2 (nx11009)) ;
    nor02_2x ix8156 (.Y (nx8155), .A0 (nx8314), .A1 (nx8312)) ;
    nor03_2x ix8315 (.Y (nx8314), .A0 (nx8159), .A1 (nx9437), .A2 (nx11017)) ;
    dffr gen_21_cmp_mRegCmp_reg_Q_8 (.Q (gen_21_cmp_mReg_8), .QB (nx8159), .D (
         window_21__8), .CLK (start), .R (rst)) ;
    nor03_2x ix8313 (.Y (nx8312), .A0 (gen_21_cmp_mReg_8), .A1 (nx10127), .A2 (
             nx11025)) ;
    nand02 ix8349 (.Y (gen_21_cmp_BSCmp_op2_9), .A0 (nx8165), .A1 (nx8169)) ;
    nor02_2x ix8166 (.Y (nx8165), .A0 (nx8344), .A1 (nx8340)) ;
    nor03_2x ix8345 (.Y (nx8344), .A0 (gen_21_cmp_mReg_8), .A1 (nx9443), .A2 (
             nx10993)) ;
    nor03_2x ix8341 (.Y (nx8340), .A0 (nx8159), .A1 (nx10999), .A2 (nx11009)) ;
    nor02_2x ix8170 (.Y (nx8169), .A0 (nx8336), .A1 (nx8334)) ;
    nor03_2x ix8337 (.Y (nx8336), .A0 (nx8173), .A1 (nx9437), .A2 (nx11017)) ;
    dffr gen_21_cmp_mRegCmp_reg_Q_9 (.Q (gen_21_cmp_mReg_9), .QB (nx8173), .D (
         window_21__9), .CLK (start), .R (rst)) ;
    nor03_2x ix8335 (.Y (nx8334), .A0 (gen_21_cmp_mReg_9), .A1 (nx10127), .A2 (
             nx11025)) ;
    nand02 ix8371 (.Y (gen_21_cmp_BSCmp_op2_10), .A0 (nx8177), .A1 (nx8183)) ;
    nor02_2x ix8178 (.Y (nx8177), .A0 (nx8366), .A1 (nx8362)) ;
    nor03_2x ix8367 (.Y (nx8366), .A0 (gen_21_cmp_mReg_9), .A1 (nx9443), .A2 (
             nx10993)) ;
    nor03_2x ix8363 (.Y (nx8362), .A0 (nx8173), .A1 (nx10999), .A2 (nx11009)) ;
    nor02_2x ix8184 (.Y (nx8183), .A0 (nx8358), .A1 (nx8356)) ;
    nor03_2x ix8359 (.Y (nx8358), .A0 (nx8187), .A1 (nx9437), .A2 (nx11017)) ;
    dffr gen_21_cmp_mRegCmp_reg_Q_10 (.Q (gen_21_cmp_mReg_10), .QB (nx8187), .D (
         window_21__10), .CLK (start), .R (rst)) ;
    nor03_2x ix8357 (.Y (nx8356), .A0 (gen_21_cmp_mReg_10), .A1 (nx10127), .A2 (
             nx11025)) ;
    nand02 ix8393 (.Y (gen_21_cmp_BSCmp_op2_11), .A0 (nx8191), .A1 (nx8197)) ;
    nor02_2x ix8192 (.Y (nx8191), .A0 (nx8388), .A1 (nx8384)) ;
    nor03_2x ix8389 (.Y (nx8388), .A0 (gen_21_cmp_mReg_10), .A1 (nx9443), .A2 (
             nx10993)) ;
    nor03_2x ix8385 (.Y (nx8384), .A0 (nx8187), .A1 (nx10999), .A2 (nx11009)) ;
    nor02_2x ix8198 (.Y (nx8197), .A0 (nx8380), .A1 (nx8378)) ;
    nor03_2x ix8381 (.Y (nx8380), .A0 (nx8200), .A1 (nx9437), .A2 (nx11017)) ;
    dffr gen_21_cmp_mRegCmp_reg_Q_11 (.Q (gen_21_cmp_mReg_11), .QB (nx8200), .D (
         window_21__11), .CLK (start), .R (rst)) ;
    nor03_2x ix8379 (.Y (nx8378), .A0 (gen_21_cmp_mReg_11), .A1 (nx10127), .A2 (
             nx11025)) ;
    nand02 ix8415 (.Y (gen_21_cmp_BSCmp_op2_12), .A0 (nx8207), .A1 (nx8213)) ;
    nor02_2x ix8208 (.Y (nx8207), .A0 (nx8410), .A1 (nx8406)) ;
    nor03_2x ix8411 (.Y (nx8410), .A0 (gen_21_cmp_mReg_11), .A1 (nx9443), .A2 (
             nx10993)) ;
    nor03_2x ix8407 (.Y (nx8406), .A0 (nx8200), .A1 (nx10999), .A2 (nx11009)) ;
    nor02_2x ix8214 (.Y (nx8213), .A0 (nx8402), .A1 (nx8400)) ;
    nor03_2x ix8403 (.Y (nx8402), .A0 (nx8217), .A1 (nx9439), .A2 (nx11017)) ;
    dffr gen_21_cmp_mRegCmp_reg_Q_12 (.Q (gen_21_cmp_mReg_12), .QB (nx8217), .D (
         window_21__12), .CLK (start), .R (rst)) ;
    nor03_2x ix8401 (.Y (nx8400), .A0 (gen_21_cmp_mReg_12), .A1 (nx10127), .A2 (
             nx11025)) ;
    nand02 ix8437 (.Y (gen_21_cmp_BSCmp_op2_13), .A0 (nx8221), .A1 (nx8227)) ;
    nor02_2x ix8222 (.Y (nx8221), .A0 (nx8432), .A1 (nx8428)) ;
    nor03_2x ix8433 (.Y (nx8432), .A0 (gen_21_cmp_mReg_12), .A1 (nx9445), .A2 (
             nx10995)) ;
    nor03_2x ix8429 (.Y (nx8428), .A0 (nx8217), .A1 (nx10999), .A2 (nx11011)) ;
    nor02_2x ix8228 (.Y (nx8227), .A0 (nx8424), .A1 (nx8422)) ;
    nor03_2x ix8425 (.Y (nx8424), .A0 (nx8231), .A1 (nx9439), .A2 (nx11019)) ;
    dffr gen_21_cmp_mRegCmp_reg_Q_13 (.Q (gen_21_cmp_mReg_13), .QB (nx8231), .D (
         window_21__13), .CLK (start), .R (rst)) ;
    nor03_2x ix8423 (.Y (nx8422), .A0 (gen_21_cmp_mReg_13), .A1 (nx10127), .A2 (
             nx11027)) ;
    nand02 ix8459 (.Y (gen_21_cmp_BSCmp_op2_14), .A0 (nx8235), .A1 (nx8241)) ;
    nor02_2x ix8236 (.Y (nx8235), .A0 (nx8454), .A1 (nx8450)) ;
    nor03_2x ix8455 (.Y (nx8454), .A0 (gen_21_cmp_mReg_13), .A1 (nx9445), .A2 (
             nx10995)) ;
    nor03_2x ix8451 (.Y (nx8450), .A0 (nx8231), .A1 (nx11001), .A2 (nx11011)) ;
    nor02_2x ix8242 (.Y (nx8241), .A0 (nx8446), .A1 (nx8444)) ;
    nor03_2x ix8447 (.Y (nx8446), .A0 (nx8244), .A1 (nx9439), .A2 (nx11019)) ;
    dffr gen_21_cmp_mRegCmp_reg_Q_14 (.Q (gen_21_cmp_mReg_14), .QB (nx8244), .D (
         window_21__14), .CLK (start), .R (rst)) ;
    nor03_2x ix8445 (.Y (nx8444), .A0 (gen_21_cmp_mReg_14), .A1 (nx10127), .A2 (
             nx11027)) ;
    nand02 ix8481 (.Y (gen_21_cmp_BSCmp_op2_15), .A0 (nx8251), .A1 (nx8257)) ;
    nor02_2x ix8252 (.Y (nx8251), .A0 (nx8476), .A1 (nx8472)) ;
    nor03_2x ix8477 (.Y (nx8476), .A0 (gen_21_cmp_mReg_14), .A1 (nx9445), .A2 (
             nx10995)) ;
    nor03_2x ix8473 (.Y (nx8472), .A0 (nx8244), .A1 (nx11001), .A2 (nx11011)) ;
    nor02_2x ix8258 (.Y (nx8257), .A0 (nx8468), .A1 (nx8466)) ;
    nor03_2x ix8469 (.Y (nx8468), .A0 (nx8261), .A1 (nx9439), .A2 (nx11019)) ;
    dffr gen_21_cmp_mRegCmp_reg_Q_15 (.Q (gen_21_cmp_mReg_15), .QB (nx8261), .D (
         window_21__15), .CLK (start), .R (rst)) ;
    nor03_2x ix8467 (.Y (nx8466), .A0 (gen_21_cmp_mReg_15), .A1 (nx10129), .A2 (
             nx11027)) ;
    nand02 ix8491 (.Y (gen_21_cmp_BSCmp_op2_16), .A0 (nx8265), .A1 (nx8257)) ;
    nor02_2x ix8266 (.Y (nx8265), .A0 (nx8486), .A1 (nx8482)) ;
    nor03_2x ix8487 (.Y (nx8486), .A0 (gen_21_cmp_mReg_15), .A1 (nx9445), .A2 (
             nx10995)) ;
    nor03_2x ix8483 (.Y (nx8482), .A0 (nx8261), .A1 (nx11001), .A2 (nx11011)) ;
    nand02 ix8559 (.Y (gen_22_cmp_BSCmp_op2_1), .A0 (nx8273), .A1 (nx8293)) ;
    nor02_2x ix8274 (.Y (nx8273), .A0 (nx8554), .A1 (nx8550)) ;
    nor03_2x ix8555 (.Y (nx8554), .A0 (gen_22_cmp_mReg_0), .A1 (nx9429), .A2 (
             nx11031)) ;
    dffr gen_22_cmp_mRegCmp_reg_Q_0 (.Q (gen_22_cmp_mReg_0), .QB (nx8279), .D (
         window_22__0), .CLK (start), .R (rst)) ;
    inv01 ix8284 (.Y (nx8283), .A (gen_22_cmp_pMux_0)) ;
    nor03_2x ix8551 (.Y (nx8550), .A0 (nx8279), .A1 (nx11037), .A2 (nx11047)) ;
    inv02 ix8292 (.Y (nx8291), .A (gen_22_cmp_pMux_2)) ;
    nor02_2x ix8294 (.Y (nx8293), .A0 (nx8540), .A1 (nx8538)) ;
    nor03_2x ix8541 (.Y (nx8540), .A0 (nx8297), .A1 (nx9423), .A2 (nx11055)) ;
    dffr gen_22_cmp_mRegCmp_reg_Q_1 (.Q (gen_22_cmp_mReg_1), .QB (nx8297), .D (
         window_22__1), .CLK (start), .R (rst)) ;
    nor03_2x ix8539 (.Y (nx8538), .A0 (gen_22_cmp_mReg_1), .A1 (nx10131), .A2 (
             nx11063)) ;
    nor03_2x ix8499 (.Y (nx8498), .A0 (nx9429), .A1 (nx8291), .A2 (
             gen_22_cmp_pMux_0)) ;
    nand02 ix8581 (.Y (gen_22_cmp_BSCmp_op2_2), .A0 (nx8308), .A1 (nx8313)) ;
    nor02_2x ix8309 (.Y (nx8308), .A0 (nx8576), .A1 (nx8572)) ;
    nor03_2x ix8577 (.Y (nx8576), .A0 (gen_22_cmp_mReg_1), .A1 (nx9429), .A2 (
             nx11031)) ;
    nor03_2x ix8573 (.Y (nx8572), .A0 (nx8297), .A1 (nx11037), .A2 (nx11047)) ;
    nor02_2x ix8314 (.Y (nx8313), .A0 (nx8568), .A1 (nx8566)) ;
    nor03_2x ix8569 (.Y (nx8568), .A0 (nx8317), .A1 (nx9423), .A2 (nx11055)) ;
    dffr gen_22_cmp_mRegCmp_reg_Q_2 (.Q (gen_22_cmp_mReg_2), .QB (nx8317), .D (
         window_22__2), .CLK (start), .R (rst)) ;
    nor03_2x ix8567 (.Y (nx8566), .A0 (gen_22_cmp_mReg_2), .A1 (nx10131), .A2 (
             nx11063)) ;
    nand02 ix8603 (.Y (gen_22_cmp_BSCmp_op2_3), .A0 (nx8323), .A1 (nx8329)) ;
    nor02_2x ix8324 (.Y (nx8323), .A0 (nx8598), .A1 (nx8594)) ;
    nor03_2x ix8599 (.Y (nx8598), .A0 (gen_22_cmp_mReg_2), .A1 (nx9429), .A2 (
             nx11031)) ;
    nor03_2x ix8595 (.Y (nx8594), .A0 (nx8317), .A1 (nx11037), .A2 (nx11047)) ;
    nor02_2x ix8330 (.Y (nx8329), .A0 (nx8590), .A1 (nx8588)) ;
    nor03_2x ix8591 (.Y (nx8590), .A0 (nx8332), .A1 (nx9423), .A2 (nx11055)) ;
    dffr gen_22_cmp_mRegCmp_reg_Q_3 (.Q (gen_22_cmp_mReg_3), .QB (nx8332), .D (
         window_22__3), .CLK (start), .R (rst)) ;
    nor03_2x ix8589 (.Y (nx8588), .A0 (gen_22_cmp_mReg_3), .A1 (nx10131), .A2 (
             nx11063)) ;
    nand02 ix8625 (.Y (gen_22_cmp_BSCmp_op2_4), .A0 (nx8339), .A1 (nx8345)) ;
    nor02_2x ix8340 (.Y (nx8339), .A0 (nx8620), .A1 (nx8616)) ;
    nor03_2x ix8621 (.Y (nx8620), .A0 (gen_22_cmp_mReg_3), .A1 (nx9429), .A2 (
             nx11031)) ;
    nor03_2x ix8617 (.Y (nx8616), .A0 (nx8332), .A1 (nx11037), .A2 (nx11047)) ;
    nor02_2x ix8346 (.Y (nx8345), .A0 (nx8612), .A1 (nx8610)) ;
    nor03_2x ix8613 (.Y (nx8612), .A0 (nx8349), .A1 (nx9423), .A2 (nx11055)) ;
    dffr gen_22_cmp_mRegCmp_reg_Q_4 (.Q (gen_22_cmp_mReg_4), .QB (nx8349), .D (
         window_22__4), .CLK (start), .R (rst)) ;
    nor03_2x ix8611 (.Y (nx8610), .A0 (gen_22_cmp_mReg_4), .A1 (nx10131), .A2 (
             nx11063)) ;
    nand02 ix8647 (.Y (gen_22_cmp_BSCmp_op2_5), .A0 (nx8353), .A1 (nx8359)) ;
    nor02_2x ix8354 (.Y (nx8353), .A0 (nx8642), .A1 (nx8638)) ;
    nor03_2x ix8643 (.Y (nx8642), .A0 (gen_22_cmp_mReg_4), .A1 (nx9429), .A2 (
             nx11031)) ;
    nor03_2x ix8639 (.Y (nx8638), .A0 (nx8349), .A1 (nx11037), .A2 (nx11047)) ;
    nor02_2x ix8360 (.Y (nx8359), .A0 (nx8634), .A1 (nx8632)) ;
    nor03_2x ix8635 (.Y (nx8634), .A0 (nx8363), .A1 (nx9425), .A2 (nx11055)) ;
    dffr gen_22_cmp_mRegCmp_reg_Q_5 (.Q (gen_22_cmp_mReg_5), .QB (nx8363), .D (
         window_22__5), .CLK (start), .R (rst)) ;
    nor03_2x ix8633 (.Y (nx8632), .A0 (gen_22_cmp_mReg_5), .A1 (nx10131), .A2 (
             nx11063)) ;
    nand02 ix8669 (.Y (gen_22_cmp_BSCmp_op2_6), .A0 (nx8367), .A1 (nx8373)) ;
    nor02_2x ix8368 (.Y (nx8367), .A0 (nx8664), .A1 (nx8660)) ;
    nor03_2x ix8665 (.Y (nx8664), .A0 (gen_22_cmp_mReg_5), .A1 (nx9431), .A2 (
             nx11031)) ;
    nor03_2x ix8661 (.Y (nx8660), .A0 (nx8363), .A1 (nx11037), .A2 (nx11047)) ;
    nor02_2x ix8374 (.Y (nx8373), .A0 (nx8656), .A1 (nx8654)) ;
    nor03_2x ix8657 (.Y (nx8656), .A0 (nx8376), .A1 (nx9425), .A2 (nx11055)) ;
    dffr gen_22_cmp_mRegCmp_reg_Q_6 (.Q (gen_22_cmp_mReg_6), .QB (nx8376), .D (
         window_22__6), .CLK (start), .R (rst)) ;
    nor03_2x ix8655 (.Y (nx8654), .A0 (gen_22_cmp_mReg_6), .A1 (nx10131), .A2 (
             nx11063)) ;
    nand02 ix8691 (.Y (gen_22_cmp_BSCmp_op2_7), .A0 (nx8383), .A1 (nx8389)) ;
    nor02_2x ix8384 (.Y (nx8383), .A0 (nx8686), .A1 (nx8682)) ;
    nor03_2x ix8687 (.Y (nx8686), .A0 (gen_22_cmp_mReg_6), .A1 (nx9431), .A2 (
             nx11033)) ;
    nor03_2x ix8683 (.Y (nx8682), .A0 (nx8376), .A1 (nx11039), .A2 (nx11049)) ;
    nor02_2x ix8390 (.Y (nx8389), .A0 (nx8678), .A1 (nx8676)) ;
    nor03_2x ix8679 (.Y (nx8678), .A0 (nx8393), .A1 (nx9425), .A2 (nx11057)) ;
    dffr gen_22_cmp_mRegCmp_reg_Q_7 (.Q (gen_22_cmp_mReg_7), .QB (nx8393), .D (
         window_22__7), .CLK (start), .R (rst)) ;
    nor03_2x ix8677 (.Y (nx8676), .A0 (gen_22_cmp_mReg_7), .A1 (nx10131), .A2 (
             nx11065)) ;
    nand02 ix8713 (.Y (gen_22_cmp_BSCmp_op2_8), .A0 (nx8397), .A1 (nx8403)) ;
    nor02_2x ix8398 (.Y (nx8397), .A0 (nx8708), .A1 (nx8704)) ;
    nor03_2x ix8709 (.Y (nx8708), .A0 (gen_22_cmp_mReg_7), .A1 (nx9431), .A2 (
             nx11033)) ;
    nor03_2x ix8705 (.Y (nx8704), .A0 (nx8393), .A1 (nx11039), .A2 (nx11049)) ;
    nor02_2x ix8404 (.Y (nx8403), .A0 (nx8700), .A1 (nx8698)) ;
    nor03_2x ix8701 (.Y (nx8700), .A0 (nx8407), .A1 (nx9425), .A2 (nx11057)) ;
    dffr gen_22_cmp_mRegCmp_reg_Q_8 (.Q (gen_22_cmp_mReg_8), .QB (nx8407), .D (
         window_22__8), .CLK (start), .R (rst)) ;
    nor03_2x ix8699 (.Y (nx8698), .A0 (gen_22_cmp_mReg_8), .A1 (nx10133), .A2 (
             nx11065)) ;
    nand02 ix8735 (.Y (gen_22_cmp_BSCmp_op2_9), .A0 (nx8411), .A1 (nx8417)) ;
    nor02_2x ix8412 (.Y (nx8411), .A0 (nx8730), .A1 (nx8726)) ;
    nor03_2x ix8731 (.Y (nx8730), .A0 (gen_22_cmp_mReg_8), .A1 (nx9431), .A2 (
             nx11033)) ;
    nor03_2x ix8727 (.Y (nx8726), .A0 (nx8407), .A1 (nx11039), .A2 (nx11049)) ;
    nor02_2x ix8418 (.Y (nx8417), .A0 (nx8722), .A1 (nx8720)) ;
    nor03_2x ix8723 (.Y (nx8722), .A0 (nx8420), .A1 (nx9425), .A2 (nx11057)) ;
    dffr gen_22_cmp_mRegCmp_reg_Q_9 (.Q (gen_22_cmp_mReg_9), .QB (nx8420), .D (
         window_22__9), .CLK (start), .R (rst)) ;
    nor03_2x ix8721 (.Y (nx8720), .A0 (gen_22_cmp_mReg_9), .A1 (nx10133), .A2 (
             nx11065)) ;
    nand02 ix8757 (.Y (gen_22_cmp_BSCmp_op2_10), .A0 (nx8427), .A1 (nx8433)) ;
    nor02_2x ix8428 (.Y (nx8427), .A0 (nx8752), .A1 (nx8748)) ;
    nor03_2x ix8753 (.Y (nx8752), .A0 (gen_22_cmp_mReg_9), .A1 (nx9431), .A2 (
             nx11033)) ;
    nor03_2x ix8749 (.Y (nx8748), .A0 (nx8420), .A1 (nx11039), .A2 (nx11049)) ;
    nor02_2x ix8434 (.Y (nx8433), .A0 (nx8744), .A1 (nx8742)) ;
    nor03_2x ix8745 (.Y (nx8744), .A0 (nx8437), .A1 (nx9425), .A2 (nx11057)) ;
    dffr gen_22_cmp_mRegCmp_reg_Q_10 (.Q (gen_22_cmp_mReg_10), .QB (nx8437), .D (
         window_22__10), .CLK (start), .R (rst)) ;
    nor03_2x ix8743 (.Y (nx8742), .A0 (gen_22_cmp_mReg_10), .A1 (nx10133), .A2 (
             nx11065)) ;
    nand02 ix8779 (.Y (gen_22_cmp_BSCmp_op2_11), .A0 (nx8441), .A1 (nx8447)) ;
    nor02_2x ix8442 (.Y (nx8441), .A0 (nx8774), .A1 (nx8770)) ;
    nor03_2x ix8775 (.Y (nx8774), .A0 (gen_22_cmp_mReg_10), .A1 (nx9431), .A2 (
             nx11033)) ;
    nor03_2x ix8771 (.Y (nx8770), .A0 (nx8437), .A1 (nx11039), .A2 (nx11049)) ;
    nor02_2x ix8448 (.Y (nx8447), .A0 (nx8766), .A1 (nx8764)) ;
    nor03_2x ix8767 (.Y (nx8766), .A0 (nx8451), .A1 (nx9425), .A2 (nx11057)) ;
    dffr gen_22_cmp_mRegCmp_reg_Q_11 (.Q (gen_22_cmp_mReg_11), .QB (nx8451), .D (
         window_22__11), .CLK (start), .R (rst)) ;
    nor03_2x ix8765 (.Y (nx8764), .A0 (gen_22_cmp_mReg_11), .A1 (nx10133), .A2 (
             nx11065)) ;
    nand02 ix8801 (.Y (gen_22_cmp_BSCmp_op2_12), .A0 (nx8455), .A1 (nx8461)) ;
    nor02_2x ix8456 (.Y (nx8455), .A0 (nx8796), .A1 (nx8792)) ;
    nor03_2x ix8797 (.Y (nx8796), .A0 (gen_22_cmp_mReg_11), .A1 (nx9431), .A2 (
             nx11033)) ;
    nor03_2x ix8793 (.Y (nx8792), .A0 (nx8451), .A1 (nx11039), .A2 (nx11049)) ;
    nor02_2x ix8462 (.Y (nx8461), .A0 (nx8788), .A1 (nx8786)) ;
    nor03_2x ix8789 (.Y (nx8788), .A0 (nx8464), .A1 (nx9427), .A2 (nx11057)) ;
    dffr gen_22_cmp_mRegCmp_reg_Q_12 (.Q (gen_22_cmp_mReg_12), .QB (nx8464), .D (
         window_22__12), .CLK (start), .R (rst)) ;
    nor03_2x ix8787 (.Y (nx8786), .A0 (gen_22_cmp_mReg_12), .A1 (nx10133), .A2 (
             nx11065)) ;
    nand02 ix8823 (.Y (gen_22_cmp_BSCmp_op2_13), .A0 (nx8471), .A1 (nx8477)) ;
    nor02_2x ix8472 (.Y (nx8471), .A0 (nx8818), .A1 (nx8814)) ;
    nor03_2x ix8819 (.Y (nx8818), .A0 (gen_22_cmp_mReg_12), .A1 (nx9433), .A2 (
             nx11035)) ;
    nor03_2x ix8815 (.Y (nx8814), .A0 (nx8464), .A1 (nx11039), .A2 (nx11051)) ;
    nor02_2x ix8478 (.Y (nx8477), .A0 (nx8810), .A1 (nx8808)) ;
    nor03_2x ix8811 (.Y (nx8810), .A0 (nx8481), .A1 (nx9427), .A2 (nx11059)) ;
    dffr gen_22_cmp_mRegCmp_reg_Q_13 (.Q (gen_22_cmp_mReg_13), .QB (nx8481), .D (
         window_22__13), .CLK (start), .R (rst)) ;
    nor03_2x ix8809 (.Y (nx8808), .A0 (gen_22_cmp_mReg_13), .A1 (nx10133), .A2 (
             nx11067)) ;
    nand02 ix8845 (.Y (gen_22_cmp_BSCmp_op2_14), .A0 (nx8487), .A1 (nx8493)) ;
    nor02_2x ix8488 (.Y (nx8487), .A0 (nx8840), .A1 (nx8836)) ;
    nor03_2x ix8841 (.Y (nx8840), .A0 (gen_22_cmp_mReg_13), .A1 (nx9433), .A2 (
             nx11035)) ;
    nor03_2x ix8837 (.Y (nx8836), .A0 (nx8481), .A1 (nx11041), .A2 (nx11051)) ;
    nor02_2x ix8494 (.Y (nx8493), .A0 (nx8832), .A1 (nx8830)) ;
    nor03_2x ix8833 (.Y (nx8832), .A0 (nx8497), .A1 (nx9427), .A2 (nx11059)) ;
    dffr gen_22_cmp_mRegCmp_reg_Q_14 (.Q (gen_22_cmp_mReg_14), .QB (nx8497), .D (
         window_22__14), .CLK (start), .R (rst)) ;
    nor03_2x ix8831 (.Y (nx8830), .A0 (gen_22_cmp_mReg_14), .A1 (nx10133), .A2 (
             nx11067)) ;
    nand02 ix8867 (.Y (gen_22_cmp_BSCmp_op2_15), .A0 (nx8502), .A1 (nx8506)) ;
    nor02_2x ix8503 (.Y (nx8502), .A0 (nx8862), .A1 (nx8858)) ;
    nor03_2x ix8863 (.Y (nx8862), .A0 (gen_22_cmp_mReg_14), .A1 (nx9433), .A2 (
             nx11035)) ;
    nor03_2x ix8859 (.Y (nx8858), .A0 (nx8497), .A1 (nx11041), .A2 (nx11051)) ;
    nor02_2x ix8507 (.Y (nx8506), .A0 (nx8854), .A1 (nx8852)) ;
    nor03_2x ix8855 (.Y (nx8854), .A0 (nx8509), .A1 (nx9427), .A2 (nx11059)) ;
    dffr gen_22_cmp_mRegCmp_reg_Q_15 (.Q (gen_22_cmp_mReg_15), .QB (nx8509), .D (
         window_22__15), .CLK (start), .R (rst)) ;
    nor03_2x ix8853 (.Y (nx8852), .A0 (gen_22_cmp_mReg_15), .A1 (nx10135), .A2 (
             nx11067)) ;
    nand02 ix8877 (.Y (gen_22_cmp_BSCmp_op2_16), .A0 (nx8515), .A1 (nx8506)) ;
    nor02_2x ix8516 (.Y (nx8515), .A0 (nx8872), .A1 (nx8868)) ;
    nor03_2x ix8873 (.Y (nx8872), .A0 (gen_22_cmp_mReg_15), .A1 (nx9433), .A2 (
             nx11035)) ;
    nor03_2x ix8869 (.Y (nx8868), .A0 (nx8509), .A1 (nx11041), .A2 (nx11051)) ;
    nand02 ix8945 (.Y (gen_23_cmp_BSCmp_op2_1), .A0 (nx8523), .A1 (nx8543)) ;
    nor02_2x ix8524 (.Y (nx8523), .A0 (nx8940), .A1 (nx8936)) ;
    nor03_2x ix8941 (.Y (nx8940), .A0 (gen_23_cmp_mReg_0), .A1 (nx9417), .A2 (
             nx11071)) ;
    dffr gen_23_cmp_mRegCmp_reg_Q_0 (.Q (gen_23_cmp_mReg_0), .QB (nx8529), .D (
         window_23__0), .CLK (start), .R (rst)) ;
    inv01 ix8534 (.Y (nx8533), .A (gen_23_cmp_pMux_0)) ;
    nor03_2x ix8937 (.Y (nx8936), .A0 (nx8529), .A1 (nx11077), .A2 (nx11087)) ;
    inv02 ix8542 (.Y (nx8541), .A (gen_23_cmp_pMux_2)) ;
    nor02_2x ix8544 (.Y (nx8543), .A0 (nx8926), .A1 (nx8924)) ;
    nor03_2x ix8927 (.Y (nx8926), .A0 (nx8547), .A1 (nx9411), .A2 (nx11095)) ;
    dffr gen_23_cmp_mRegCmp_reg_Q_1 (.Q (gen_23_cmp_mReg_1), .QB (nx8547), .D (
         window_23__1), .CLK (start), .R (rst)) ;
    nor03_2x ix8925 (.Y (nx8924), .A0 (gen_23_cmp_mReg_1), .A1 (nx10137), .A2 (
             nx11103)) ;
    nor03_2x ix8885 (.Y (nx8884), .A0 (nx9417), .A1 (nx8541), .A2 (
             gen_23_cmp_pMux_0)) ;
    nand02 ix8967 (.Y (gen_23_cmp_BSCmp_op2_2), .A0 (nx8559), .A1 (nx8563)) ;
    nor02_2x ix8560 (.Y (nx8559), .A0 (nx8962), .A1 (nx8958)) ;
    nor03_2x ix8963 (.Y (nx8962), .A0 (gen_23_cmp_mReg_1), .A1 (nx9417), .A2 (
             nx11071)) ;
    nor03_2x ix8959 (.Y (nx8958), .A0 (nx8547), .A1 (nx11077), .A2 (nx11087)) ;
    nor02_2x ix8564 (.Y (nx8563), .A0 (nx8954), .A1 (nx8952)) ;
    nor03_2x ix8955 (.Y (nx8954), .A0 (nx8567), .A1 (nx9411), .A2 (nx11095)) ;
    dffr gen_23_cmp_mRegCmp_reg_Q_2 (.Q (gen_23_cmp_mReg_2), .QB (nx8567), .D (
         window_23__2), .CLK (start), .R (rst)) ;
    nor03_2x ix8953 (.Y (nx8952), .A0 (gen_23_cmp_mReg_2), .A1 (nx10137), .A2 (
             nx11103)) ;
    nand02 ix8989 (.Y (gen_23_cmp_BSCmp_op2_3), .A0 (nx8573), .A1 (nx8577)) ;
    nor02_2x ix8574 (.Y (nx8573), .A0 (nx8984), .A1 (nx8980)) ;
    nor03_2x ix8985 (.Y (nx8984), .A0 (gen_23_cmp_mReg_2), .A1 (nx9417), .A2 (
             nx11071)) ;
    nor03_2x ix8981 (.Y (nx8980), .A0 (nx8567), .A1 (nx11077), .A2 (nx11087)) ;
    nor02_2x ix8578 (.Y (nx8577), .A0 (nx8976), .A1 (nx8974)) ;
    nor03_2x ix8977 (.Y (nx8976), .A0 (nx8581), .A1 (nx9411), .A2 (nx11095)) ;
    dffr gen_23_cmp_mRegCmp_reg_Q_3 (.Q (gen_23_cmp_mReg_3), .QB (nx8581), .D (
         window_23__3), .CLK (start), .R (rst)) ;
    nor03_2x ix8975 (.Y (nx8974), .A0 (gen_23_cmp_mReg_3), .A1 (nx10137), .A2 (
             nx11103)) ;
    nand02 ix9011 (.Y (gen_23_cmp_BSCmp_op2_4), .A0 (nx8585), .A1 (nx8591)) ;
    nor02_2x ix8586 (.Y (nx8585), .A0 (nx9006), .A1 (nx9002)) ;
    nor03_2x ix9007 (.Y (nx9006), .A0 (gen_23_cmp_mReg_3), .A1 (nx9417), .A2 (
             nx11071)) ;
    nor03_2x ix9003 (.Y (nx9002), .A0 (nx8581), .A1 (nx11077), .A2 (nx11087)) ;
    nor02_2x ix8592 (.Y (nx8591), .A0 (nx8998), .A1 (nx8996)) ;
    nor03_2x ix8999 (.Y (nx8998), .A0 (nx8595), .A1 (nx9411), .A2 (nx11095)) ;
    dffr gen_23_cmp_mRegCmp_reg_Q_4 (.Q (gen_23_cmp_mReg_4), .QB (nx8595), .D (
         window_23__4), .CLK (start), .R (rst)) ;
    nor03_2x ix8997 (.Y (nx8996), .A0 (gen_23_cmp_mReg_4), .A1 (nx10137), .A2 (
             nx11103)) ;
    nand02 ix9033 (.Y (gen_23_cmp_BSCmp_op2_5), .A0 (nx8599), .A1 (nx8605)) ;
    nor02_2x ix8600 (.Y (nx8599), .A0 (nx9028), .A1 (nx9024)) ;
    nor03_2x ix9029 (.Y (nx9028), .A0 (gen_23_cmp_mReg_4), .A1 (nx9417), .A2 (
             nx11071)) ;
    nor03_2x ix9025 (.Y (nx9024), .A0 (nx8595), .A1 (nx11077), .A2 (nx11087)) ;
    nor02_2x ix8606 (.Y (nx8605), .A0 (nx9020), .A1 (nx9018)) ;
    nor03_2x ix9021 (.Y (nx9020), .A0 (nx8608), .A1 (nx9413), .A2 (nx11095)) ;
    dffr gen_23_cmp_mRegCmp_reg_Q_5 (.Q (gen_23_cmp_mReg_5), .QB (nx8608), .D (
         window_23__5), .CLK (start), .R (rst)) ;
    nor03_2x ix9019 (.Y (nx9018), .A0 (gen_23_cmp_mReg_5), .A1 (nx10137), .A2 (
             nx11103)) ;
    nand02 ix9055 (.Y (gen_23_cmp_BSCmp_op2_6), .A0 (nx8615), .A1 (nx8621)) ;
    nor02_2x ix8616 (.Y (nx8615), .A0 (nx9050), .A1 (nx9046)) ;
    nor03_2x ix9051 (.Y (nx9050), .A0 (gen_23_cmp_mReg_5), .A1 (nx9419), .A2 (
             nx11071)) ;
    nor03_2x ix9047 (.Y (nx9046), .A0 (nx8608), .A1 (nx11077), .A2 (nx11087)) ;
    nor02_2x ix8622 (.Y (nx8621), .A0 (nx9042), .A1 (nx9040)) ;
    nor03_2x ix9043 (.Y (nx9042), .A0 (nx8625), .A1 (nx9413), .A2 (nx11095)) ;
    dffr gen_23_cmp_mRegCmp_reg_Q_6 (.Q (gen_23_cmp_mReg_6), .QB (nx8625), .D (
         window_23__6), .CLK (start), .R (rst)) ;
    nor03_2x ix9041 (.Y (nx9040), .A0 (gen_23_cmp_mReg_6), .A1 (nx10137), .A2 (
             nx11103)) ;
    nand02 ix9077 (.Y (gen_23_cmp_BSCmp_op2_7), .A0 (nx8629), .A1 (nx8635)) ;
    nor02_2x ix8630 (.Y (nx8629), .A0 (nx9072), .A1 (nx9068)) ;
    nor03_2x ix9073 (.Y (nx9072), .A0 (gen_23_cmp_mReg_6), .A1 (nx9419), .A2 (
             nx11073)) ;
    nor03_2x ix9069 (.Y (nx9068), .A0 (nx8625), .A1 (nx11079), .A2 (nx11089)) ;
    nor02_2x ix8636 (.Y (nx8635), .A0 (nx9064), .A1 (nx9062)) ;
    nor03_2x ix9065 (.Y (nx9064), .A0 (nx8639), .A1 (nx9413), .A2 (nx11097)) ;
    dffr gen_23_cmp_mRegCmp_reg_Q_7 (.Q (gen_23_cmp_mReg_7), .QB (nx8639), .D (
         window_23__7), .CLK (start), .R (rst)) ;
    nor03_2x ix9063 (.Y (nx9062), .A0 (gen_23_cmp_mReg_7), .A1 (nx10137), .A2 (
             nx11105)) ;
    nand02 ix9099 (.Y (gen_23_cmp_BSCmp_op2_8), .A0 (nx8643), .A1 (nx8649)) ;
    nor02_2x ix8644 (.Y (nx8643), .A0 (nx9094), .A1 (nx9090)) ;
    nor03_2x ix9095 (.Y (nx9094), .A0 (gen_23_cmp_mReg_7), .A1 (nx9419), .A2 (
             nx11073)) ;
    nor03_2x ix9091 (.Y (nx9090), .A0 (nx8639), .A1 (nx11079), .A2 (nx11089)) ;
    nor02_2x ix8650 (.Y (nx8649), .A0 (nx9086), .A1 (nx9084)) ;
    nor03_2x ix9087 (.Y (nx9086), .A0 (nx8652), .A1 (nx9413), .A2 (nx11097)) ;
    dffr gen_23_cmp_mRegCmp_reg_Q_8 (.Q (gen_23_cmp_mReg_8), .QB (nx8652), .D (
         window_23__8), .CLK (start), .R (rst)) ;
    nor03_2x ix9085 (.Y (nx9084), .A0 (gen_23_cmp_mReg_8), .A1 (nx10139), .A2 (
             nx11105)) ;
    nand02 ix9121 (.Y (gen_23_cmp_BSCmp_op2_9), .A0 (nx8659), .A1 (nx8665)) ;
    nor02_2x ix8660 (.Y (nx8659), .A0 (nx9116), .A1 (nx9112)) ;
    nor03_2x ix9117 (.Y (nx9116), .A0 (gen_23_cmp_mReg_8), .A1 (nx9419), .A2 (
             nx11073)) ;
    nor03_2x ix9113 (.Y (nx9112), .A0 (nx8652), .A1 (nx11079), .A2 (nx11089)) ;
    nor02_2x ix8666 (.Y (nx8665), .A0 (nx9108), .A1 (nx9106)) ;
    nor03_2x ix9109 (.Y (nx9108), .A0 (nx8669), .A1 (nx9413), .A2 (nx11097)) ;
    dffr gen_23_cmp_mRegCmp_reg_Q_9 (.Q (gen_23_cmp_mReg_9), .QB (nx8669), .D (
         window_23__9), .CLK (start), .R (rst)) ;
    nor03_2x ix9107 (.Y (nx9106), .A0 (gen_23_cmp_mReg_9), .A1 (nx10139), .A2 (
             nx11105)) ;
    nand02 ix9143 (.Y (gen_23_cmp_BSCmp_op2_10), .A0 (nx8673), .A1 (nx8679)) ;
    nor02_2x ix8674 (.Y (nx8673), .A0 (nx9138), .A1 (nx9134)) ;
    nor03_2x ix9139 (.Y (nx9138), .A0 (gen_23_cmp_mReg_9), .A1 (nx9419), .A2 (
             nx11073)) ;
    nor03_2x ix9135 (.Y (nx9134), .A0 (nx8669), .A1 (nx11079), .A2 (nx11089)) ;
    nor02_2x ix8680 (.Y (nx8679), .A0 (nx9130), .A1 (nx9128)) ;
    nor03_2x ix9131 (.Y (nx9130), .A0 (nx8683), .A1 (nx9413), .A2 (nx11097)) ;
    dffr gen_23_cmp_mRegCmp_reg_Q_10 (.Q (gen_23_cmp_mReg_10), .QB (nx8683), .D (
         window_23__10), .CLK (start), .R (rst)) ;
    nor03_2x ix9129 (.Y (nx9128), .A0 (gen_23_cmp_mReg_10), .A1 (nx10139), .A2 (
             nx11105)) ;
    nand02 ix9165 (.Y (gen_23_cmp_BSCmp_op2_11), .A0 (nx8687), .A1 (nx8693)) ;
    nor02_2x ix8688 (.Y (nx8687), .A0 (nx9160), .A1 (nx9156)) ;
    nor03_2x ix9161 (.Y (nx9160), .A0 (gen_23_cmp_mReg_10), .A1 (nx9419), .A2 (
             nx11073)) ;
    nor03_2x ix9157 (.Y (nx9156), .A0 (nx8683), .A1 (nx11079), .A2 (nx11089)) ;
    nor02_2x ix8694 (.Y (nx8693), .A0 (nx9152), .A1 (nx9150)) ;
    nor03_2x ix9153 (.Y (nx9152), .A0 (nx8696), .A1 (nx9413), .A2 (nx11097)) ;
    dffr gen_23_cmp_mRegCmp_reg_Q_11 (.Q (gen_23_cmp_mReg_11), .QB (nx8696), .D (
         window_23__11), .CLK (start), .R (rst)) ;
    nor03_2x ix9151 (.Y (nx9150), .A0 (gen_23_cmp_mReg_11), .A1 (nx10139), .A2 (
             nx11105)) ;
    nand02 ix9187 (.Y (gen_23_cmp_BSCmp_op2_12), .A0 (nx8703), .A1 (nx8709)) ;
    nor02_2x ix8704 (.Y (nx8703), .A0 (nx9182), .A1 (nx9178)) ;
    nor03_2x ix9183 (.Y (nx9182), .A0 (gen_23_cmp_mReg_11), .A1 (nx9419), .A2 (
             nx11073)) ;
    nor03_2x ix9179 (.Y (nx9178), .A0 (nx8696), .A1 (nx11079), .A2 (nx11089)) ;
    nor02_2x ix8710 (.Y (nx8709), .A0 (nx9174), .A1 (nx9172)) ;
    nor03_2x ix9175 (.Y (nx9174), .A0 (nx8713), .A1 (nx9415), .A2 (nx11097)) ;
    dffr gen_23_cmp_mRegCmp_reg_Q_12 (.Q (gen_23_cmp_mReg_12), .QB (nx8713), .D (
         window_23__12), .CLK (start), .R (rst)) ;
    nor03_2x ix9173 (.Y (nx9172), .A0 (gen_23_cmp_mReg_12), .A1 (nx10139), .A2 (
             nx11105)) ;
    nand02 ix9209 (.Y (gen_23_cmp_BSCmp_op2_13), .A0 (nx8717), .A1 (nx8723)) ;
    nor02_2x ix8718 (.Y (nx8717), .A0 (nx9204), .A1 (nx9200)) ;
    nor03_2x ix9205 (.Y (nx9204), .A0 (gen_23_cmp_mReg_12), .A1 (nx9421), .A2 (
             nx11075)) ;
    nor03_2x ix9201 (.Y (nx9200), .A0 (nx8713), .A1 (nx11079), .A2 (nx11091)) ;
    nor02_2x ix8724 (.Y (nx8723), .A0 (nx9196), .A1 (nx9194)) ;
    nor03_2x ix9197 (.Y (nx9196), .A0 (nx8727), .A1 (nx9415), .A2 (nx11099)) ;
    dffr gen_23_cmp_mRegCmp_reg_Q_13 (.Q (gen_23_cmp_mReg_13), .QB (nx8727), .D (
         window_23__13), .CLK (start), .R (rst)) ;
    nor03_2x ix9195 (.Y (nx9194), .A0 (gen_23_cmp_mReg_13), .A1 (nx10139), .A2 (
             nx11107)) ;
    nand02 ix9231 (.Y (gen_23_cmp_BSCmp_op2_14), .A0 (nx8731), .A1 (nx8737)) ;
    nor02_2x ix8732 (.Y (nx8731), .A0 (nx9226), .A1 (nx9222)) ;
    nor03_2x ix9227 (.Y (nx9226), .A0 (gen_23_cmp_mReg_13), .A1 (nx9421), .A2 (
             nx11075)) ;
    nor03_2x ix9223 (.Y (nx9222), .A0 (nx8727), .A1 (nx11081), .A2 (nx11091)) ;
    nor02_2x ix8738 (.Y (nx8737), .A0 (nx9218), .A1 (nx9216)) ;
    nor03_2x ix9219 (.Y (nx9218), .A0 (nx8740), .A1 (nx9415), .A2 (nx11099)) ;
    dffr gen_23_cmp_mRegCmp_reg_Q_14 (.Q (gen_23_cmp_mReg_14), .QB (nx8740), .D (
         window_23__14), .CLK (start), .R (rst)) ;
    nor03_2x ix9217 (.Y (nx9216), .A0 (gen_23_cmp_mReg_14), .A1 (nx10139), .A2 (
             nx11107)) ;
    nand02 ix9253 (.Y (gen_23_cmp_BSCmp_op2_15), .A0 (nx8747), .A1 (nx8753)) ;
    nor02_2x ix8748 (.Y (nx8747), .A0 (nx9248), .A1 (nx9244)) ;
    nor03_2x ix9249 (.Y (nx9248), .A0 (gen_23_cmp_mReg_14), .A1 (nx9421), .A2 (
             nx11075)) ;
    nor03_2x ix9245 (.Y (nx9244), .A0 (nx8740), .A1 (nx11081), .A2 (nx11091)) ;
    nor02_2x ix8754 (.Y (nx8753), .A0 (nx9240), .A1 (nx9238)) ;
    nor03_2x ix9241 (.Y (nx9240), .A0 (nx8757), .A1 (nx9415), .A2 (nx11099)) ;
    dffr gen_23_cmp_mRegCmp_reg_Q_15 (.Q (gen_23_cmp_mReg_15), .QB (nx8757), .D (
         window_23__15), .CLK (start), .R (rst)) ;
    nor03_2x ix9239 (.Y (nx9238), .A0 (gen_23_cmp_mReg_15), .A1 (nx10141), .A2 (
             nx11107)) ;
    nand02 ix9263 (.Y (gen_23_cmp_BSCmp_op2_16), .A0 (nx8761), .A1 (nx8753)) ;
    nor02_2x ix8762 (.Y (nx8761), .A0 (nx9258), .A1 (nx9254)) ;
    nor03_2x ix9259 (.Y (nx9258), .A0 (gen_23_cmp_mReg_15), .A1 (nx9421), .A2 (
             nx11075)) ;
    nor03_2x ix9255 (.Y (nx9254), .A0 (nx8757), .A1 (nx11081), .A2 (nx11091)) ;
    nand02 ix9331 (.Y (gen_24_cmp_BSCmp_op2_1), .A0 (nx8769), .A1 (nx8789)) ;
    nor02_2x ix8770 (.Y (nx8769), .A0 (nx9326), .A1 (nx9322)) ;
    nor03_2x ix9327 (.Y (nx9326), .A0 (gen_24_cmp_mReg_0), .A1 (nx9405), .A2 (
             nx11111)) ;
    dffr gen_24_cmp_mRegCmp_reg_Q_0 (.Q (gen_24_cmp_mReg_0), .QB (nx8775), .D (
         window_24__0), .CLK (start), .R (rst)) ;
    inv01 ix8780 (.Y (nx8779), .A (gen_24_cmp_pMux_0)) ;
    nor03_2x ix9323 (.Y (nx9322), .A0 (nx8775), .A1 (nx11117), .A2 (nx11127)) ;
    inv02 ix8788 (.Y (nx8787), .A (gen_24_cmp_pMux_2)) ;
    nor02_2x ix8790 (.Y (nx8789), .A0 (nx9312), .A1 (nx9310)) ;
    nor03_2x ix9313 (.Y (nx9312), .A0 (nx8793), .A1 (nx9399), .A2 (nx11135)) ;
    dffr gen_24_cmp_mRegCmp_reg_Q_1 (.Q (gen_24_cmp_mReg_1), .QB (nx8793), .D (
         window_24__1), .CLK (start), .R (rst)) ;
    nor03_2x ix9311 (.Y (nx9310), .A0 (gen_24_cmp_mReg_1), .A1 (nx10143), .A2 (
             nx11143)) ;
    nor03_2x ix9271 (.Y (nx9270), .A0 (nx9405), .A1 (nx8787), .A2 (
             gen_24_cmp_pMux_0)) ;
    nand02 ix9353 (.Y (gen_24_cmp_BSCmp_op2_2), .A0 (nx8804), .A1 (nx8809)) ;
    nor02_2x ix8805 (.Y (nx8804), .A0 (nx9348), .A1 (nx9344)) ;
    nor03_2x ix9349 (.Y (nx9348), .A0 (gen_24_cmp_mReg_1), .A1 (nx9405), .A2 (
             nx11111)) ;
    nor03_2x ix9345 (.Y (nx9344), .A0 (nx8793), .A1 (nx11117), .A2 (nx11127)) ;
    nor02_2x ix8810 (.Y (nx8809), .A0 (nx9340), .A1 (nx9338)) ;
    nor03_2x ix9341 (.Y (nx9340), .A0 (nx8813), .A1 (nx9399), .A2 (nx11135)) ;
    dffr gen_24_cmp_mRegCmp_reg_Q_2 (.Q (gen_24_cmp_mReg_2), .QB (nx8813), .D (
         window_24__2), .CLK (start), .R (rst)) ;
    nor03_2x ix9339 (.Y (nx9338), .A0 (gen_24_cmp_mReg_2), .A1 (nx10143), .A2 (
             nx11143)) ;
    nand02 ix9375 (.Y (gen_24_cmp_BSCmp_op2_3), .A0 (nx8819), .A1 (nx8825)) ;
    nor02_2x ix8820 (.Y (nx8819), .A0 (nx9370), .A1 (nx9366)) ;
    nor03_2x ix9371 (.Y (nx9370), .A0 (gen_24_cmp_mReg_2), .A1 (nx9405), .A2 (
             nx11111)) ;
    nor03_2x ix9367 (.Y (nx9366), .A0 (nx8813), .A1 (nx11117), .A2 (nx11127)) ;
    nor02_2x ix8826 (.Y (nx8825), .A0 (nx9362), .A1 (nx9360)) ;
    nor03_2x ix9363 (.Y (nx9362), .A0 (nx8828), .A1 (nx9399), .A2 (nx11135)) ;
    dffr gen_24_cmp_mRegCmp_reg_Q_3 (.Q (gen_24_cmp_mReg_3), .QB (nx8828), .D (
         window_24__3), .CLK (start), .R (rst)) ;
    nor03_2x ix9361 (.Y (nx9360), .A0 (gen_24_cmp_mReg_3), .A1 (nx10143), .A2 (
             nx11143)) ;
    nand02 ix9397 (.Y (gen_24_cmp_BSCmp_op2_4), .A0 (nx8835), .A1 (nx8841)) ;
    nor02_2x ix8836 (.Y (nx8835), .A0 (nx9392), .A1 (nx9388)) ;
    nor03_2x ix9393 (.Y (nx9392), .A0 (gen_24_cmp_mReg_3), .A1 (nx9405), .A2 (
             nx11111)) ;
    nor03_2x ix9389 (.Y (nx9388), .A0 (nx8828), .A1 (nx11117), .A2 (nx11127)) ;
    nor02_2x ix8842 (.Y (nx8841), .A0 (nx9384), .A1 (nx9382)) ;
    nor03_2x ix9385 (.Y (nx9384), .A0 (nx8845), .A1 (nx9399), .A2 (nx11135)) ;
    dffr gen_24_cmp_mRegCmp_reg_Q_4 (.Q (gen_24_cmp_mReg_4), .QB (nx8845), .D (
         window_24__4), .CLK (start), .R (rst)) ;
    nor03_2x ix9383 (.Y (nx9382), .A0 (gen_24_cmp_mReg_4), .A1 (nx10143), .A2 (
             nx11143)) ;
    nand02 ix9419 (.Y (gen_24_cmp_BSCmp_op2_5), .A0 (nx8849), .A1 (nx8855)) ;
    nor02_2x ix8850 (.Y (nx8849), .A0 (nx9414), .A1 (nx9410)) ;
    nor03_2x ix9415 (.Y (nx9414), .A0 (gen_24_cmp_mReg_4), .A1 (nx9405), .A2 (
             nx11111)) ;
    nor03_2x ix9411 (.Y (nx9410), .A0 (nx8845), .A1 (nx11117), .A2 (nx11127)) ;
    nor02_2x ix8856 (.Y (nx8855), .A0 (nx9406), .A1 (nx9404)) ;
    nor03_2x ix9407 (.Y (nx9406), .A0 (nx8859), .A1 (nx9401), .A2 (nx11135)) ;
    dffr gen_24_cmp_mRegCmp_reg_Q_5 (.Q (gen_24_cmp_mReg_5), .QB (nx8859), .D (
         window_24__5), .CLK (start), .R (rst)) ;
    nor03_2x ix9405 (.Y (nx9404), .A0 (gen_24_cmp_mReg_5), .A1 (nx10143), .A2 (
             nx11143)) ;
    nand02 ix9441 (.Y (gen_24_cmp_BSCmp_op2_6), .A0 (nx8863), .A1 (nx8869)) ;
    nor02_2x ix8864 (.Y (nx8863), .A0 (nx9436), .A1 (nx9432)) ;
    nor03_2x ix9437 (.Y (nx9436), .A0 (gen_24_cmp_mReg_5), .A1 (nx9407), .A2 (
             nx11111)) ;
    nor03_2x ix9433 (.Y (nx9432), .A0 (nx8859), .A1 (nx11117), .A2 (nx11127)) ;
    nor02_2x ix8870 (.Y (nx8869), .A0 (nx9428), .A1 (nx9426)) ;
    nor03_2x ix9429 (.Y (nx9428), .A0 (nx8873), .A1 (nx9401), .A2 (nx11135)) ;
    dffr gen_24_cmp_mRegCmp_reg_Q_6 (.Q (gen_24_cmp_mReg_6), .QB (nx8873), .D (
         window_24__6), .CLK (start), .R (rst)) ;
    nor03_2x ix9427 (.Y (nx9426), .A0 (gen_24_cmp_mReg_6), .A1 (nx10143), .A2 (
             nx11143)) ;
    nand02 ix9463 (.Y (gen_24_cmp_BSCmp_op2_7), .A0 (nx8879), .A1 (nx8885)) ;
    nor02_2x ix8880 (.Y (nx8879), .A0 (nx9458), .A1 (nx9454)) ;
    nor03_2x ix9459 (.Y (nx9458), .A0 (gen_24_cmp_mReg_6), .A1 (nx9407), .A2 (
             nx11113)) ;
    nor03_2x ix9455 (.Y (nx9454), .A0 (nx8873), .A1 (nx11119), .A2 (nx11129)) ;
    nor02_2x ix8886 (.Y (nx8885), .A0 (nx9450), .A1 (nx9448)) ;
    nor03_2x ix9451 (.Y (nx9450), .A0 (nx8888), .A1 (nx9401), .A2 (nx11137)) ;
    dffr gen_24_cmp_mRegCmp_reg_Q_7 (.Q (gen_24_cmp_mReg_7), .QB (nx8888), .D (
         window_24__7), .CLK (start), .R (rst)) ;
    nor03_2x ix9449 (.Y (nx9448), .A0 (gen_24_cmp_mReg_7), .A1 (nx10143), .A2 (
             nx11145)) ;
    nand02 ix9485 (.Y (gen_24_cmp_BSCmp_op2_8), .A0 (nx8892), .A1 (nx8897)) ;
    nor02_2x ix8893 (.Y (nx8892), .A0 (nx9480), .A1 (nx9476)) ;
    nor03_2x ix9481 (.Y (nx9480), .A0 (gen_24_cmp_mReg_7), .A1 (nx9407), .A2 (
             nx11113)) ;
    nor03_2x ix9477 (.Y (nx9476), .A0 (nx8888), .A1 (nx11119), .A2 (nx11129)) ;
    nor02_2x ix8898 (.Y (nx8897), .A0 (nx9472), .A1 (nx9470)) ;
    nor03_2x ix9473 (.Y (nx9472), .A0 (nx8901), .A1 (nx9401), .A2 (nx11137)) ;
    dffr gen_24_cmp_mRegCmp_reg_Q_8 (.Q (gen_24_cmp_mReg_8), .QB (nx8901), .D (
         window_24__8), .CLK (start), .R (rst)) ;
    nor03_2x ix9471 (.Y (nx9470), .A0 (gen_24_cmp_mReg_8), .A1 (nx10145), .A2 (
             nx11145)) ;
    nand02 ix9507 (.Y (gen_24_cmp_BSCmp_op2_9), .A0 (nx8907), .A1 (nx8913)) ;
    nor02_2x ix8908 (.Y (nx8907), .A0 (nx9502), .A1 (nx9498)) ;
    nor03_2x ix9503 (.Y (nx9502), .A0 (gen_24_cmp_mReg_8), .A1 (nx9407), .A2 (
             nx11113)) ;
    nor03_2x ix9499 (.Y (nx9498), .A0 (nx8901), .A1 (nx11119), .A2 (nx11129)) ;
    nor02_2x ix8914 (.Y (nx8913), .A0 (nx9494), .A1 (nx9492)) ;
    nor03_2x ix9495 (.Y (nx9494), .A0 (nx8917), .A1 (nx9401), .A2 (nx11137)) ;
    dffr gen_24_cmp_mRegCmp_reg_Q_9 (.Q (gen_24_cmp_mReg_9), .QB (nx8917), .D (
         window_24__9), .CLK (start), .R (rst)) ;
    nor03_2x ix9493 (.Y (nx9492), .A0 (gen_24_cmp_mReg_9), .A1 (nx10145), .A2 (
             nx11145)) ;
    nand02 ix9529 (.Y (gen_24_cmp_BSCmp_op2_10), .A0 (nx8921), .A1 (nx8927)) ;
    nor02_2x ix8922 (.Y (nx8921), .A0 (nx9524), .A1 (nx9520)) ;
    nor03_2x ix9525 (.Y (nx9524), .A0 (gen_24_cmp_mReg_9), .A1 (nx9407), .A2 (
             nx11113)) ;
    nor03_2x ix9521 (.Y (nx9520), .A0 (nx8917), .A1 (nx11119), .A2 (nx11129)) ;
    nor02_2x ix8928 (.Y (nx8927), .A0 (nx9516), .A1 (nx9514)) ;
    nor03_2x ix9517 (.Y (nx9516), .A0 (nx8931), .A1 (nx9401), .A2 (nx11137)) ;
    dffr gen_24_cmp_mRegCmp_reg_Q_10 (.Q (gen_24_cmp_mReg_10), .QB (nx8931), .D (
         window_24__10), .CLK (start), .R (rst)) ;
    nor03_2x ix9515 (.Y (nx9514), .A0 (gen_24_cmp_mReg_10), .A1 (nx10145), .A2 (
             nx11145)) ;
    nand02 ix9551 (.Y (gen_24_cmp_BSCmp_op2_11), .A0 (nx8937), .A1 (nx8941)) ;
    nor02_2x ix8938 (.Y (nx8937), .A0 (nx9546), .A1 (nx9542)) ;
    nor03_2x ix9547 (.Y (nx9546), .A0 (gen_24_cmp_mReg_10), .A1 (nx9407), .A2 (
             nx11113)) ;
    nor03_2x ix9543 (.Y (nx9542), .A0 (nx8931), .A1 (nx11119), .A2 (nx11129)) ;
    nor02_2x ix8942 (.Y (nx8941), .A0 (nx9538), .A1 (nx9536)) ;
    nor03_2x ix9539 (.Y (nx9538), .A0 (nx8945), .A1 (nx9401), .A2 (nx11137)) ;
    dffr gen_24_cmp_mRegCmp_reg_Q_11 (.Q (gen_24_cmp_mReg_11), .QB (nx8945), .D (
         window_24__11), .CLK (start), .R (rst)) ;
    nor03_2x ix9537 (.Y (nx9536), .A0 (gen_24_cmp_mReg_11), .A1 (nx10145), .A2 (
             nx11145)) ;
    nand02 ix9573 (.Y (gen_24_cmp_BSCmp_op2_12), .A0 (nx8949), .A1 (nx8955)) ;
    nor02_2x ix8950 (.Y (nx8949), .A0 (nx9568), .A1 (nx9564)) ;
    nor03_2x ix9569 (.Y (nx9568), .A0 (gen_24_cmp_mReg_11), .A1 (nx9407), .A2 (
             nx11113)) ;
    nor03_2x ix9565 (.Y (nx9564), .A0 (nx8945), .A1 (nx11119), .A2 (nx11129)) ;
    nor02_2x ix8956 (.Y (nx8955), .A0 (nx9560), .A1 (nx9558)) ;
    nor03_2x ix9561 (.Y (nx9560), .A0 (nx8959), .A1 (nx9403), .A2 (nx11137)) ;
    dffr gen_24_cmp_mRegCmp_reg_Q_12 (.Q (gen_24_cmp_mReg_12), .QB (nx8959), .D (
         window_24__12), .CLK (start), .R (rst)) ;
    nor03_2x ix9559 (.Y (nx9558), .A0 (gen_24_cmp_mReg_12), .A1 (nx10145), .A2 (
             nx11145)) ;
    nand02 ix9595 (.Y (gen_24_cmp_BSCmp_op2_13), .A0 (nx8963), .A1 (nx8969)) ;
    nor02_2x ix8964 (.Y (nx8963), .A0 (nx9590), .A1 (nx9586)) ;
    nor03_2x ix9591 (.Y (nx9590), .A0 (gen_24_cmp_mReg_12), .A1 (nx9409), .A2 (
             nx11115)) ;
    nor03_2x ix9587 (.Y (nx9586), .A0 (nx8959), .A1 (nx11119), .A2 (nx11131)) ;
    nor02_2x ix8970 (.Y (nx8969), .A0 (nx9582), .A1 (nx9580)) ;
    nor03_2x ix9583 (.Y (nx9582), .A0 (nx8972), .A1 (nx9403), .A2 (nx11139)) ;
    dffr gen_24_cmp_mRegCmp_reg_Q_13 (.Q (gen_24_cmp_mReg_13), .QB (nx8972), .D (
         window_24__13), .CLK (start), .R (rst)) ;
    nor03_2x ix9581 (.Y (nx9580), .A0 (gen_24_cmp_mReg_13), .A1 (nx10145), .A2 (
             nx11147)) ;
    nand02 ix9617 (.Y (gen_24_cmp_BSCmp_op2_14), .A0 (nx8979), .A1 (nx8985)) ;
    nor02_2x ix8980 (.Y (nx8979), .A0 (nx9612), .A1 (nx9608)) ;
    nor03_2x ix9613 (.Y (nx9612), .A0 (gen_24_cmp_mReg_13), .A1 (nx9409), .A2 (
             nx11115)) ;
    nor03_2x ix9609 (.Y (nx9608), .A0 (nx8972), .A1 (nx11121), .A2 (nx11131)) ;
    nor02_2x ix8986 (.Y (nx8985), .A0 (nx9604), .A1 (nx9602)) ;
    nor03_2x ix9605 (.Y (nx9604), .A0 (nx8989), .A1 (nx9403), .A2 (nx11139)) ;
    dffr gen_24_cmp_mRegCmp_reg_Q_14 (.Q (gen_24_cmp_mReg_14), .QB (nx8989), .D (
         window_24__14), .CLK (start), .R (rst)) ;
    nor03_2x ix9603 (.Y (nx9602), .A0 (gen_24_cmp_mReg_14), .A1 (nx10145), .A2 (
             nx11147)) ;
    nand02 ix9639 (.Y (gen_24_cmp_BSCmp_op2_15), .A0 (nx8993), .A1 (nx8999)) ;
    nor02_2x ix8994 (.Y (nx8993), .A0 (nx9634), .A1 (nx9630)) ;
    nor03_2x ix9635 (.Y (nx9634), .A0 (gen_24_cmp_mReg_14), .A1 (nx9409), .A2 (
             nx11115)) ;
    nor03_2x ix9631 (.Y (nx9630), .A0 (nx8989), .A1 (nx11121), .A2 (nx11131)) ;
    nor02_2x ix9000 (.Y (nx8999), .A0 (nx9626), .A1 (nx9624)) ;
    nor03_2x ix9627 (.Y (nx9626), .A0 (nx9003), .A1 (nx9403), .A2 (nx11139)) ;
    dffr gen_24_cmp_mRegCmp_reg_Q_15 (.Q (gen_24_cmp_mReg_15), .QB (nx9003), .D (
         window_24__15), .CLK (start), .R (rst)) ;
    nor03_2x ix9625 (.Y (nx9624), .A0 (gen_24_cmp_mReg_15), .A1 (nx10147), .A2 (
             nx11147)) ;
    nand02 ix9649 (.Y (gen_24_cmp_BSCmp_op2_16), .A0 (nx9007), .A1 (nx8999)) ;
    nor02_2x ix9008 (.Y (nx9007), .A0 (nx9644), .A1 (nx9640)) ;
    nor03_2x ix9645 (.Y (nx9644), .A0 (gen_24_cmp_mReg_15), .A1 (nx9409), .A2 (
             nx11115)) ;
    nor03_2x ix9641 (.Y (nx9640), .A0 (nx9003), .A1 (nx11121), .A2 (nx11131)) ;
    nor02_2x ix19 (.Y (gen_0_cmp_BSCmp_carryIn), .A0 (nx2871), .A1 (nx9014)) ;
    nor02_2x ix9015 (.Y (nx9014), .A0 (nx10161), .A1 (nx2862)) ;
    nand02 ix39 (.Y (gen_0_cmp_BSCmp_op2_0), .A0 (nx9017), .A1 (nx9023)) ;
    nor02_2x ix9018 (.Y (nx9017), .A0 (nx34), .A1 (nx26)) ;
    nor03_2x ix35 (.Y (nx34), .A0 (nx2859), .A1 (nx9691), .A2 (nx10179)) ;
    nor03_2x ix27 (.Y (nx26), .A0 (gen_0_cmp_mReg_0), .A1 (nx10003), .A2 (
             nx10187)) ;
    nand03 ix9024 (.Y (nx9023), .A0 (nx10161), .A1 (nx9691), .A2 (nx2862)) ;
    nor02_2x ix405 (.Y (gen_1_cmp_BSCmp_carryIn), .A0 (nx3115), .A1 (nx9027)) ;
    nor02_2x ix9028 (.Y (nx9027), .A0 (nx10201), .A1 (nx3107)) ;
    nand02 ix425 (.Y (gen_1_cmp_BSCmp_op2_0), .A0 (nx9031), .A1 (nx9036)) ;
    nor02_2x ix9032 (.Y (nx9031), .A0 (nx420), .A1 (nx412)) ;
    nor03_2x ix421 (.Y (nx420), .A0 (nx3103), .A1 (nx9679), .A2 (nx10219)) ;
    nor03_2x ix413 (.Y (nx412), .A0 (gen_1_cmp_mReg_0), .A1 (nx10009), .A2 (
             nx10227)) ;
    nand03 ix9037 (.Y (nx9036), .A0 (nx10201), .A1 (nx9679), .A2 (nx3107)) ;
    nor02_2x ix791 (.Y (gen_2_cmp_BSCmp_carryIn), .A0 (nx3363), .A1 (nx9039)) ;
    nor02_2x ix9040 (.Y (nx9039), .A0 (nx10241), .A1 (nx3356)) ;
    nand02 ix811 (.Y (gen_2_cmp_BSCmp_op2_0), .A0 (nx9043), .A1 (nx9049)) ;
    nor02_2x ix9044 (.Y (nx9043), .A0 (nx806), .A1 (nx798)) ;
    nor03_2x ix807 (.Y (nx806), .A0 (nx3353), .A1 (nx9667), .A2 (nx10259)) ;
    nor03_2x ix799 (.Y (nx798), .A0 (gen_2_cmp_mReg_0), .A1 (nx10015), .A2 (
             nx10267)) ;
    nand03 ix9050 (.Y (nx9049), .A0 (nx10241), .A1 (nx9667), .A2 (nx3356)) ;
    nor02_2x ix1177 (.Y (gen_3_cmp_BSCmp_carryIn), .A0 (nx3611), .A1 (nx9053)) ;
    nor02_2x ix9054 (.Y (nx9053), .A0 (nx10281), .A1 (nx3603)) ;
    nand02 ix1197 (.Y (gen_3_cmp_BSCmp_op2_0), .A0 (nx9057), .A1 (nx9061)) ;
    nor02_2x ix9058 (.Y (nx9057), .A0 (nx1192), .A1 (nx1184)) ;
    nor03_2x ix1193 (.Y (nx1192), .A0 (nx3599), .A1 (nx9655), .A2 (nx10299)) ;
    nor03_2x ix1185 (.Y (nx1184), .A0 (gen_3_cmp_mReg_0), .A1 (nx10021), .A2 (
             nx10307)) ;
    nand03 ix9062 (.Y (nx9061), .A0 (nx10281), .A1 (nx9655), .A2 (nx3603)) ;
    nor02_2x ix1563 (.Y (gen_4_cmp_BSCmp_carryIn), .A0 (nx3857), .A1 (nx9065)) ;
    nor02_2x ix9066 (.Y (nx9065), .A0 (nx10321), .A1 (nx3849)) ;
    nand02 ix1583 (.Y (gen_4_cmp_BSCmp_op2_0), .A0 (nx9069), .A1 (nx9073)) ;
    nor02_2x ix9070 (.Y (nx9069), .A0 (nx1578), .A1 (nx1570)) ;
    nor03_2x ix1579 (.Y (nx1578), .A0 (nx3845), .A1 (nx9643), .A2 (nx10339)) ;
    nor03_2x ix1571 (.Y (nx1570), .A0 (gen_4_cmp_mReg_0), .A1 (nx10027), .A2 (
             nx10347)) ;
    nand03 ix9074 (.Y (nx9073), .A0 (nx10321), .A1 (nx9643), .A2 (nx3849)) ;
    nor02_2x ix1949 (.Y (gen_5_cmp_BSCmp_carryIn), .A0 (nx4101), .A1 (nx9077)) ;
    nor02_2x ix9078 (.Y (nx9077), .A0 (nx10361), .A1 (nx4093)) ;
    nand02 ix1969 (.Y (gen_5_cmp_BSCmp_op2_0), .A0 (nx9080), .A1 (nx9085)) ;
    nor02_2x ix9081 (.Y (nx9080), .A0 (nx1964), .A1 (nx1956)) ;
    nor03_2x ix1965 (.Y (nx1964), .A0 (nx4089), .A1 (nx9631), .A2 (nx10379)) ;
    nor03_2x ix1957 (.Y (nx1956), .A0 (gen_5_cmp_mReg_0), .A1 (nx10033), .A2 (
             nx10387)) ;
    nand03 ix9086 (.Y (nx9085), .A0 (nx10361), .A1 (nx9631), .A2 (nx4093)) ;
    nor02_2x ix2335 (.Y (gen_6_cmp_BSCmp_carryIn), .A0 (nx4349), .A1 (nx9089)) ;
    nor02_2x ix9090 (.Y (nx9089), .A0 (nx10401), .A1 (nx4340)) ;
    nand02 ix2355 (.Y (gen_6_cmp_BSCmp_op2_0), .A0 (nx9093), .A1 (nx9099)) ;
    nor02_2x ix9094 (.Y (nx9093), .A0 (nx2350), .A1 (nx2342)) ;
    nor03_2x ix2351 (.Y (nx2350), .A0 (nx4337), .A1 (nx9619), .A2 (nx10419)) ;
    nor03_2x ix2343 (.Y (nx2342), .A0 (gen_6_cmp_mReg_0), .A1 (nx10039), .A2 (
             nx10427)) ;
    nand03 ix9100 (.Y (nx9099), .A0 (nx10401), .A1 (nx9619), .A2 (nx4340)) ;
    nor02_2x ix2721 (.Y (gen_7_cmp_BSCmp_carryIn), .A0 (nx4595), .A1 (nx9102)) ;
    nor02_2x ix9103 (.Y (nx9102), .A0 (nx10441), .A1 (nx4587)) ;
    nand02 ix2741 (.Y (gen_7_cmp_BSCmp_op2_0), .A0 (nx9105), .A1 (nx9111)) ;
    nor02_2x ix9106 (.Y (nx9105), .A0 (nx2736), .A1 (nx2728)) ;
    nor03_2x ix2737 (.Y (nx2736), .A0 (nx4583), .A1 (nx9607), .A2 (nx10459)) ;
    nor03_2x ix2729 (.Y (nx2728), .A0 (gen_7_cmp_mReg_0), .A1 (nx10045), .A2 (
             nx10467)) ;
    nand03 ix9112 (.Y (nx9111), .A0 (nx10441), .A1 (nx9607), .A2 (nx4587)) ;
    nor02_2x ix3107 (.Y (gen_8_cmp_BSCmp_carryIn), .A0 (nx4841), .A1 (nx9115)) ;
    nor02_2x ix9116 (.Y (nx9115), .A0 (nx10481), .A1 (nx4834)) ;
    nand02 ix3127 (.Y (gen_8_cmp_BSCmp_op2_0), .A0 (nx9119), .A1 (nx9124)) ;
    nor02_2x ix9120 (.Y (nx9119), .A0 (nx3122), .A1 (nx3114)) ;
    nor03_2x ix3123 (.Y (nx3122), .A0 (nx4831), .A1 (nx9595), .A2 (nx10499)) ;
    nor03_2x ix3115 (.Y (nx3114), .A0 (gen_8_cmp_mReg_0), .A1 (nx10051), .A2 (
             nx10507)) ;
    nand03 ix9125 (.Y (nx9124), .A0 (nx10481), .A1 (nx9595), .A2 (nx4834)) ;
    nor02_2x ix3493 (.Y (gen_9_cmp_BSCmp_carryIn), .A0 (nx5085), .A1 (nx9127)) ;
    nor02_2x ix9128 (.Y (nx9127), .A0 (nx10521), .A1 (nx5077)) ;
    nand02 ix3513 (.Y (gen_9_cmp_BSCmp_op2_0), .A0 (nx9131), .A1 (nx9137)) ;
    nor02_2x ix9132 (.Y (nx9131), .A0 (nx3508), .A1 (nx3500)) ;
    nor03_2x ix3509 (.Y (nx3508), .A0 (nx5073), .A1 (nx9583), .A2 (nx10539)) ;
    nor03_2x ix3501 (.Y (nx3500), .A0 (gen_9_cmp_mReg_0), .A1 (nx10057), .A2 (
             nx10547)) ;
    nand03 ix9138 (.Y (nx9137), .A0 (nx10521), .A1 (nx9583), .A2 (nx5077)) ;
    nor02_2x ix3879 (.Y (gen_10_cmp_BSCmp_carryIn), .A0 (nx5335), .A1 (nx9141)
             ) ;
    nor02_2x ix9142 (.Y (nx9141), .A0 (nx10561), .A1 (nx5327)) ;
    nand02 ix3899 (.Y (gen_10_cmp_BSCmp_op2_0), .A0 (nx9145), .A1 (nx9149)) ;
    nor02_2x ix9146 (.Y (nx9145), .A0 (nx3894), .A1 (nx3886)) ;
    nor03_2x ix3895 (.Y (nx3894), .A0 (nx5323), .A1 (nx9571), .A2 (nx10579)) ;
    nor03_2x ix3887 (.Y (nx3886), .A0 (gen_10_cmp_mReg_0), .A1 (nx10063), .A2 (
             nx10587)) ;
    nand03 ix9150 (.Y (nx9149), .A0 (nx10561), .A1 (nx9571), .A2 (nx5327)) ;
    nor02_2x ix4265 (.Y (gen_11_cmp_BSCmp_carryIn), .A0 (nx5585), .A1 (nx9153)
             ) ;
    nor02_2x ix9154 (.Y (nx9153), .A0 (nx10601), .A1 (nx5577)) ;
    nand02 ix4285 (.Y (gen_11_cmp_BSCmp_op2_0), .A0 (nx9157), .A1 (nx9161)) ;
    nor02_2x ix9158 (.Y (nx9157), .A0 (nx4280), .A1 (nx4272)) ;
    nor03_2x ix4281 (.Y (nx4280), .A0 (nx5573), .A1 (nx9559), .A2 (nx10619)) ;
    nor03_2x ix4273 (.Y (nx4272), .A0 (gen_11_cmp_mReg_0), .A1 (nx10069), .A2 (
             nx10627)) ;
    nand03 ix9162 (.Y (nx9161), .A0 (nx10601), .A1 (nx9559), .A2 (nx5577)) ;
    nor02_2x ix4651 (.Y (gen_12_cmp_BSCmp_carryIn), .A0 (nx5829), .A1 (nx9165)
             ) ;
    nor02_2x ix9166 (.Y (nx9165), .A0 (nx10641), .A1 (nx5821)) ;
    nand02 ix4671 (.Y (gen_12_cmp_BSCmp_op2_0), .A0 (nx9168), .A1 (nx9173)) ;
    nor02_2x ix9169 (.Y (nx9168), .A0 (nx4666), .A1 (nx4658)) ;
    nor03_2x ix4667 (.Y (nx4666), .A0 (nx5817), .A1 (nx9547), .A2 (nx10659)) ;
    nor03_2x ix4659 (.Y (nx4658), .A0 (gen_12_cmp_mReg_0), .A1 (nx10075), .A2 (
             nx10667)) ;
    nand03 ix9174 (.Y (nx9173), .A0 (nx10641), .A1 (nx9547), .A2 (nx5821)) ;
    nor02_2x ix5037 (.Y (gen_13_cmp_BSCmp_carryIn), .A0 (nx6075), .A1 (nx9177)
             ) ;
    nor02_2x ix9178 (.Y (nx9177), .A0 (nx10681), .A1 (nx6067)) ;
    nand02 ix5057 (.Y (gen_13_cmp_BSCmp_op2_0), .A0 (nx9181), .A1 (nx9187)) ;
    nor02_2x ix9182 (.Y (nx9181), .A0 (nx5052), .A1 (nx5044)) ;
    nor03_2x ix5053 (.Y (nx5052), .A0 (nx6063), .A1 (nx9535), .A2 (nx10699)) ;
    nor03_2x ix5045 (.Y (nx5044), .A0 (gen_13_cmp_mReg_0), .A1 (nx10081), .A2 (
             nx10707)) ;
    nand03 ix9188 (.Y (nx9187), .A0 (nx10681), .A1 (nx9535), .A2 (nx6067)) ;
    nor02_2x ix5423 (.Y (gen_14_cmp_BSCmp_carryIn), .A0 (nx6323), .A1 (nx9190)
             ) ;
    nor02_2x ix9191 (.Y (nx9190), .A0 (nx10721), .A1 (nx6314)) ;
    nand02 ix5443 (.Y (gen_14_cmp_BSCmp_op2_0), .A0 (nx9193), .A1 (nx9199)) ;
    nor02_2x ix9194 (.Y (nx9193), .A0 (nx5438), .A1 (nx5430)) ;
    nor03_2x ix5439 (.Y (nx5438), .A0 (nx6311), .A1 (nx9523), .A2 (nx10739)) ;
    nor03_2x ix5431 (.Y (nx5430), .A0 (gen_14_cmp_mReg_0), .A1 (nx10087), .A2 (
             nx10747)) ;
    nand03 ix9200 (.Y (nx9199), .A0 (nx10721), .A1 (nx9523), .A2 (nx6314)) ;
    nor02_2x ix5809 (.Y (gen_15_cmp_BSCmp_carryIn), .A0 (nx6569), .A1 (nx9203)
             ) ;
    nor02_2x ix9204 (.Y (nx9203), .A0 (nx10761), .A1 (nx6561)) ;
    nand02 ix5829 (.Y (gen_15_cmp_BSCmp_op2_0), .A0 (nx9207), .A1 (nx9212)) ;
    nor02_2x ix9208 (.Y (nx9207), .A0 (nx5824), .A1 (nx5816)) ;
    nor03_2x ix5825 (.Y (nx5824), .A0 (nx6557), .A1 (nx9511), .A2 (nx10779)) ;
    nor03_2x ix5817 (.Y (nx5816), .A0 (gen_15_cmp_mReg_0), .A1 (nx10093), .A2 (
             nx10787)) ;
    nand03 ix9213 (.Y (nx9212), .A0 (nx10761), .A1 (nx9511), .A2 (nx6561)) ;
    nor02_2x ix6195 (.Y (gen_16_cmp_BSCmp_carryIn), .A0 (nx6815), .A1 (nx9215)
             ) ;
    nor02_2x ix9216 (.Y (nx9215), .A0 (nx10801), .A1 (nx6808)) ;
    nand02 ix6215 (.Y (gen_16_cmp_BSCmp_op2_0), .A0 (nx9219), .A1 (nx9225)) ;
    nor02_2x ix9220 (.Y (nx9219), .A0 (nx6210), .A1 (nx6202)) ;
    nor03_2x ix6211 (.Y (nx6210), .A0 (nx6805), .A1 (nx9499), .A2 (nx10819)) ;
    nor03_2x ix6203 (.Y (nx6202), .A0 (gen_16_cmp_mReg_0), .A1 (nx10099), .A2 (
             nx10827)) ;
    nand03 ix9226 (.Y (nx9225), .A0 (nx10801), .A1 (nx9499), .A2 (nx6808)) ;
    nor02_2x ix6581 (.Y (gen_17_cmp_BSCmp_carryIn), .A0 (nx7057), .A1 (nx9229)
             ) ;
    nor02_2x ix9230 (.Y (nx9229), .A0 (nx10841), .A1 (nx7049)) ;
    nand02 ix6601 (.Y (gen_17_cmp_BSCmp_op2_0), .A0 (nx9233), .A1 (nx9237)) ;
    nor02_2x ix9234 (.Y (nx9233), .A0 (nx6596), .A1 (nx6588)) ;
    nor03_2x ix6597 (.Y (nx6596), .A0 (nx7045), .A1 (nx9487), .A2 (nx10859)) ;
    nor03_2x ix6589 (.Y (nx6588), .A0 (gen_17_cmp_mReg_0), .A1 (nx10105), .A2 (
             nx10867)) ;
    nand03 ix9238 (.Y (nx9237), .A0 (nx10841), .A1 (nx9487), .A2 (nx7049)) ;
    nor02_2x ix6967 (.Y (gen_18_cmp_BSCmp_carryIn), .A0 (nx7305), .A1 (nx9241)
             ) ;
    nor02_2x ix9242 (.Y (nx9241), .A0 (nx10881), .A1 (nx7297)) ;
    nand02 ix6987 (.Y (gen_18_cmp_BSCmp_op2_0), .A0 (nx9245), .A1 (nx9249)) ;
    nor02_2x ix9246 (.Y (nx9245), .A0 (nx6982), .A1 (nx6974)) ;
    nor03_2x ix6983 (.Y (nx6982), .A0 (nx7293), .A1 (nx9475), .A2 (nx10899)) ;
    nor03_2x ix6975 (.Y (nx6974), .A0 (gen_18_cmp_mReg_0), .A1 (nx10111), .A2 (
             nx10907)) ;
    nand03 ix9250 (.Y (nx9249), .A0 (nx10881), .A1 (nx9475), .A2 (nx7297)) ;
    nor02_2x ix7353 (.Y (gen_19_cmp_BSCmp_carryIn), .A0 (nx7553), .A1 (nx9253)
             ) ;
    nor02_2x ix9254 (.Y (nx9253), .A0 (nx10921), .A1 (nx7545)) ;
    nand02 ix7373 (.Y (gen_19_cmp_BSCmp_op2_0), .A0 (nx9257), .A1 (nx9263)) ;
    nor02_2x ix9258 (.Y (nx9257), .A0 (nx7368), .A1 (nx7360)) ;
    nor03_2x ix7369 (.Y (nx7368), .A0 (nx7541), .A1 (nx9463), .A2 (nx10939)) ;
    nor03_2x ix7361 (.Y (nx7360), .A0 (gen_19_cmp_mReg_0), .A1 (nx10117), .A2 (
             nx10947)) ;
    nand03 ix9264 (.Y (nx9263), .A0 (nx10921), .A1 (nx9463), .A2 (nx7545)) ;
    nor02_2x ix7739 (.Y (gen_20_cmp_BSCmp_carryIn), .A0 (nx7801), .A1 (nx9267)
             ) ;
    nor02_2x ix9268 (.Y (nx9267), .A0 (nx10961), .A1 (nx7792)) ;
    nand02 ix7759 (.Y (gen_20_cmp_BSCmp_op2_0), .A0 (nx9271), .A1 (nx9275)) ;
    nor02_2x ix9272 (.Y (nx9271), .A0 (nx7754), .A1 (nx7746)) ;
    nor03_2x ix7755 (.Y (nx7754), .A0 (nx7789), .A1 (nx9451), .A2 (nx10979)) ;
    nor03_2x ix7747 (.Y (nx7746), .A0 (gen_20_cmp_mReg_0), .A1 (nx10123), .A2 (
             nx10987)) ;
    nand03 ix9276 (.Y (nx9275), .A0 (nx10961), .A1 (nx9451), .A2 (nx7792)) ;
    nor02_2x ix8125 (.Y (gen_21_cmp_BSCmp_carryIn), .A0 (nx8047), .A1 (nx9278)
             ) ;
    nor02_2x ix9279 (.Y (nx9278), .A0 (nx11001), .A1 (nx8039)) ;
    nand02 ix8145 (.Y (gen_21_cmp_BSCmp_op2_0), .A0 (nx9281), .A1 (nx9287)) ;
    nor02_2x ix9282 (.Y (nx9281), .A0 (nx8140), .A1 (nx8132)) ;
    nor03_2x ix8141 (.Y (nx8140), .A0 (nx8035), .A1 (nx9439), .A2 (nx11019)) ;
    nor03_2x ix8133 (.Y (nx8132), .A0 (gen_21_cmp_mReg_0), .A1 (nx10129), .A2 (
             nx11027)) ;
    nand03 ix9288 (.Y (nx9287), .A0 (nx11001), .A1 (nx9439), .A2 (nx8039)) ;
    nor02_2x ix8511 (.Y (gen_22_cmp_BSCmp_carryIn), .A0 (nx8291), .A1 (nx9291)
             ) ;
    nor02_2x ix9292 (.Y (nx9291), .A0 (nx11041), .A1 (nx8283)) ;
    nand02 ix8531 (.Y (gen_22_cmp_BSCmp_op2_0), .A0 (nx9295), .A1 (nx9301)) ;
    nor02_2x ix9296 (.Y (nx9295), .A0 (nx8526), .A1 (nx8518)) ;
    nor03_2x ix8527 (.Y (nx8526), .A0 (nx8279), .A1 (nx9427), .A2 (nx11059)) ;
    nor03_2x ix8519 (.Y (nx8518), .A0 (gen_22_cmp_mReg_0), .A1 (nx10135), .A2 (
             nx11067)) ;
    nand03 ix9302 (.Y (nx9301), .A0 (nx11041), .A1 (nx9427), .A2 (nx8283)) ;
    nor02_2x ix8897 (.Y (gen_23_cmp_BSCmp_carryIn), .A0 (nx8541), .A1 (nx9305)
             ) ;
    nor02_2x ix9306 (.Y (nx9305), .A0 (nx11081), .A1 (nx8533)) ;
    nand02 ix8917 (.Y (gen_23_cmp_BSCmp_op2_0), .A0 (nx9308), .A1 (nx9315)) ;
    nor02_2x ix9310 (.Y (nx9308), .A0 (nx8912), .A1 (nx8904)) ;
    nor03_2x ix8913 (.Y (nx8912), .A0 (nx8529), .A1 (nx9415), .A2 (nx11099)) ;
    nor03_2x ix8905 (.Y (nx8904), .A0 (gen_23_cmp_mReg_0), .A1 (nx10141), .A2 (
             nx11107)) ;
    nand03 ix9316 (.Y (nx9315), .A0 (nx11081), .A1 (nx9415), .A2 (nx8533)) ;
    nor02_2x ix9283 (.Y (gen_24_cmp_BSCmp_carryIn), .A0 (nx8787), .A1 (nx9319)
             ) ;
    nor02_2x ix9320 (.Y (nx9319), .A0 (nx11121), .A1 (nx8779)) ;
    nand02 ix9303 (.Y (gen_24_cmp_BSCmp_op2_0), .A0 (nx9323), .A1 (nx9327)) ;
    nor02_2x ix9324 (.Y (nx9323), .A0 (nx9298), .A1 (nx9290)) ;
    nor03_2x ix9299 (.Y (nx9298), .A0 (nx8775), .A1 (nx9403), .A2 (nx11139)) ;
    nor03_2x ix9291 (.Y (nx9290), .A0 (gen_24_cmp_mReg_0), .A1 (nx10147), .A2 (
             nx11147)) ;
    nand03 ix9328 (.Y (nx9327), .A0 (nx11121), .A1 (nx9403), .A2 (nx8779)) ;
    nor02_2x ix2840 (.Y (nx2839), .A0 (nx11197), .A1 (nx11171)) ;
    dffs_ni CounterCmp_reg_outp_0 (.Q (\$dummy [125]), .QB (nx9333), .D (nx2839)
            , .CLK (clk), .S (nx9670)) ;
    inv01 ix9671 (.Y (nx9670), .A (nx9336)) ;
    nor02_2x ix9338 (.Y (nx9336), .A0 (restartDetection), .A1 (rst)) ;
    dffr StartCaptuerCmp_reg_f (.Q (restartDetection), .QB (\$dummy [126]), .D (
         nx9650), .CLK (start), .R (nx9664)) ;
    inv01 ix9665 (.Y (nx9664), .A (nx9343)) ;
    nor02_2x ix9344 (.Y (nx9343), .A0 (StartCaptuerCmp_d), .A1 (rst)) ;
    dff StartCaptuerCmp_reg_d (.Q (StartCaptuerCmp_d), .QB (\$dummy [127]), .D (
        restartDetection), .CLK (nx9397)) ;
    dffr firtStartLachCmp_reg_Q_0 (.Q (\$dummy [128]), .QB (nx9353), .D (nx9650)
         , .CLK (start), .R (rst)) ;
    oai21 ix2834 (.Y (nx2833), .A0 (nx9357), .A1 (nx9353), .B0 (nx9365)) ;
    dffr CounterCmp_reg_outp_2 (.Q (\$dummy [129]), .QB (nx9357), .D (nx2823), .CLK (
         clk), .R (nx9670)) ;
    dffr CounterCmp_reg_outp_1 (.Q (\$dummy [130]), .QB (nx9361), .D (nx2813), .CLK (
         clk), .R (nx9670)) ;
    dffr CounterCmp_reg_outp_3 (.Q (done), .QB (nx9365), .D (nx2833), .CLK (clk)
         , .R (nx9670)) ;
    inv02 ix9374 (.Y (nx9375), .A (nx9373)) ;
    inv02 ix9376 (.Y (nx9377), .A (nx11201)) ;
    inv02 ix9378 (.Y (nx9379), .A (nx11201)) ;
    inv02 ix9380 (.Y (nx9381), .A (nx11201)) ;
    inv01 ix9388 (.Y (nx9389), .A (nx9333)) ;
    inv01 ix9390 (.Y (nx9391), .A (clk)) ;
    inv01 ix9392 (.Y (nx9393), .A (clk)) ;
    inv01 ix9394 (.Y (nx9395), .A (clk)) ;
    inv01 ix9396 (.Y (nx9397), .A (clk)) ;
    inv04 ix9398 (.Y (nx9399), .A (nx8787)) ;
    inv04 ix9400 (.Y (nx9401), .A (nx8787)) ;
    inv04 ix9402 (.Y (nx9403), .A (nx8787)) ;
    inv04 ix9404 (.Y (nx9405), .A (nx11121)) ;
    inv04 ix9406 (.Y (nx9407), .A (nx11121)) ;
    inv04 ix9408 (.Y (nx9409), .A (nx11123)) ;
    inv04 ix9410 (.Y (nx9411), .A (nx8541)) ;
    inv04 ix9412 (.Y (nx9413), .A (nx8541)) ;
    inv04 ix9414 (.Y (nx9415), .A (nx8541)) ;
    inv04 ix9416 (.Y (nx9417), .A (nx11081)) ;
    inv04 ix9418 (.Y (nx9419), .A (nx11081)) ;
    inv04 ix9420 (.Y (nx9421), .A (nx11083)) ;
    inv04 ix9422 (.Y (nx9423), .A (nx8291)) ;
    inv04 ix9424 (.Y (nx9425), .A (nx8291)) ;
    inv04 ix9426 (.Y (nx9427), .A (nx8291)) ;
    inv04 ix9428 (.Y (nx9429), .A (nx11041)) ;
    inv04 ix9430 (.Y (nx9431), .A (nx11041)) ;
    inv04 ix9432 (.Y (nx9433), .A (nx11043)) ;
    inv04 ix9434 (.Y (nx9435), .A (nx8047)) ;
    inv04 ix9436 (.Y (nx9437), .A (nx8047)) ;
    inv04 ix9438 (.Y (nx9439), .A (nx8047)) ;
    inv04 ix9440 (.Y (nx9441), .A (nx11001)) ;
    inv04 ix9442 (.Y (nx9443), .A (nx11001)) ;
    inv04 ix9444 (.Y (nx9445), .A (nx11003)) ;
    inv04 ix9446 (.Y (nx9447), .A (nx7801)) ;
    inv04 ix9448 (.Y (nx9449), .A (nx7801)) ;
    inv04 ix9450 (.Y (nx9451), .A (nx7801)) ;
    inv04 ix9452 (.Y (nx9453), .A (nx10961)) ;
    inv04 ix9454 (.Y (nx9455), .A (nx10961)) ;
    inv04 ix9456 (.Y (nx9457), .A (nx10963)) ;
    inv04 ix9458 (.Y (nx9459), .A (nx7553)) ;
    inv04 ix9460 (.Y (nx9461), .A (nx7553)) ;
    inv04 ix9462 (.Y (nx9463), .A (nx7553)) ;
    inv04 ix9464 (.Y (nx9465), .A (nx10921)) ;
    inv04 ix9466 (.Y (nx9467), .A (nx10921)) ;
    inv04 ix9468 (.Y (nx9469), .A (nx10923)) ;
    inv04 ix9470 (.Y (nx9471), .A (nx7305)) ;
    inv04 ix9472 (.Y (nx9473), .A (nx7305)) ;
    inv04 ix9474 (.Y (nx9475), .A (nx7305)) ;
    inv04 ix9476 (.Y (nx9477), .A (nx10881)) ;
    inv04 ix9478 (.Y (nx9479), .A (nx10881)) ;
    inv04 ix9480 (.Y (nx9481), .A (nx10883)) ;
    inv04 ix9482 (.Y (nx9483), .A (nx7057)) ;
    inv04 ix9484 (.Y (nx9485), .A (nx7057)) ;
    inv04 ix9486 (.Y (nx9487), .A (nx7057)) ;
    inv04 ix9488 (.Y (nx9489), .A (nx10841)) ;
    inv04 ix9490 (.Y (nx9491), .A (nx10841)) ;
    inv04 ix9492 (.Y (nx9493), .A (nx10843)) ;
    inv04 ix9494 (.Y (nx9495), .A (nx6815)) ;
    inv04 ix9496 (.Y (nx9497), .A (nx6815)) ;
    inv04 ix9498 (.Y (nx9499), .A (nx6815)) ;
    inv04 ix9500 (.Y (nx9501), .A (nx10801)) ;
    inv04 ix9502 (.Y (nx9503), .A (nx10801)) ;
    inv04 ix9504 (.Y (nx9505), .A (nx10803)) ;
    inv04 ix9506 (.Y (nx9507), .A (nx6569)) ;
    inv04 ix9508 (.Y (nx9509), .A (nx6569)) ;
    inv04 ix9510 (.Y (nx9511), .A (nx6569)) ;
    inv04 ix9512 (.Y (nx9513), .A (nx10761)) ;
    inv04 ix9514 (.Y (nx9515), .A (nx10761)) ;
    inv04 ix9516 (.Y (nx9517), .A (nx10763)) ;
    inv04 ix9518 (.Y (nx9519), .A (nx6323)) ;
    inv04 ix9520 (.Y (nx9521), .A (nx6323)) ;
    inv04 ix9522 (.Y (nx9523), .A (nx6323)) ;
    inv04 ix9524 (.Y (nx9525), .A (nx10721)) ;
    inv04 ix9526 (.Y (nx9527), .A (nx10721)) ;
    inv04 ix9528 (.Y (nx9529), .A (nx10723)) ;
    inv04 ix9530 (.Y (nx9531), .A (nx6075)) ;
    inv04 ix9532 (.Y (nx9533), .A (nx6075)) ;
    inv04 ix9534 (.Y (nx9535), .A (nx6075)) ;
    inv04 ix9536 (.Y (nx9537), .A (nx10681)) ;
    inv04 ix9538 (.Y (nx9539), .A (nx10681)) ;
    inv04 ix9540 (.Y (nx9541), .A (nx10683)) ;
    inv04 ix9542 (.Y (nx9543), .A (nx5829)) ;
    inv04 ix9544 (.Y (nx9545), .A (nx5829)) ;
    inv04 ix9546 (.Y (nx9547), .A (nx5829)) ;
    inv04 ix9548 (.Y (nx9549), .A (nx10641)) ;
    inv04 ix9550 (.Y (nx9551), .A (nx10641)) ;
    inv04 ix9552 (.Y (nx9553), .A (nx10643)) ;
    inv04 ix9554 (.Y (nx9555), .A (nx5585)) ;
    inv04 ix9556 (.Y (nx9557), .A (nx5585)) ;
    inv04 ix9558 (.Y (nx9559), .A (nx5585)) ;
    inv04 ix9560 (.Y (nx9561), .A (nx10601)) ;
    inv04 ix9562 (.Y (nx9563), .A (nx10601)) ;
    inv04 ix9564 (.Y (nx9565), .A (nx10603)) ;
    inv04 ix9566 (.Y (nx9567), .A (nx5335)) ;
    inv04 ix9568 (.Y (nx9569), .A (nx5335)) ;
    inv04 ix9570 (.Y (nx9571), .A (nx5335)) ;
    inv04 ix9572 (.Y (nx9573), .A (nx10561)) ;
    inv04 ix9574 (.Y (nx9575), .A (nx10561)) ;
    inv04 ix9576 (.Y (nx9577), .A (nx10563)) ;
    inv04 ix9578 (.Y (nx9579), .A (nx5085)) ;
    inv04 ix9580 (.Y (nx9581), .A (nx5085)) ;
    inv04 ix9582 (.Y (nx9583), .A (nx5085)) ;
    inv04 ix9584 (.Y (nx9585), .A (nx10521)) ;
    inv04 ix9586 (.Y (nx9587), .A (nx10521)) ;
    inv04 ix9588 (.Y (nx9589), .A (nx10523)) ;
    inv04 ix9590 (.Y (nx9591), .A (nx4841)) ;
    inv04 ix9592 (.Y (nx9593), .A (nx4841)) ;
    inv04 ix9594 (.Y (nx9595), .A (nx4841)) ;
    inv04 ix9596 (.Y (nx9597), .A (nx10481)) ;
    inv04 ix9598 (.Y (nx9599), .A (nx10481)) ;
    inv04 ix9600 (.Y (nx9601), .A (nx10483)) ;
    inv04 ix9602 (.Y (nx9603), .A (nx4595)) ;
    inv04 ix9604 (.Y (nx9605), .A (nx4595)) ;
    inv04 ix9606 (.Y (nx9607), .A (nx4595)) ;
    inv04 ix9608 (.Y (nx9609), .A (nx10441)) ;
    inv04 ix9610 (.Y (nx9611), .A (nx10441)) ;
    inv04 ix9612 (.Y (nx9613), .A (nx10443)) ;
    inv04 ix9614 (.Y (nx9615), .A (nx4349)) ;
    inv04 ix9616 (.Y (nx9617), .A (nx4349)) ;
    inv04 ix9618 (.Y (nx9619), .A (nx4349)) ;
    inv04 ix9620 (.Y (nx9621), .A (nx10401)) ;
    inv04 ix9622 (.Y (nx9623), .A (nx10401)) ;
    inv04 ix9624 (.Y (nx9625), .A (nx10403)) ;
    inv04 ix9626 (.Y (nx9627), .A (nx4101)) ;
    inv04 ix9628 (.Y (nx9629), .A (nx4101)) ;
    inv04 ix9630 (.Y (nx9631), .A (nx4101)) ;
    inv04 ix9632 (.Y (nx9633), .A (nx10361)) ;
    inv04 ix9634 (.Y (nx9635), .A (nx10361)) ;
    inv04 ix9636 (.Y (nx9637), .A (nx10363)) ;
    inv04 ix9638 (.Y (nx9639), .A (nx3857)) ;
    inv04 ix9640 (.Y (nx9641), .A (nx3857)) ;
    inv04 ix9642 (.Y (nx9643), .A (nx3857)) ;
    inv04 ix9644 (.Y (nx9645), .A (nx10321)) ;
    inv04 ix9646 (.Y (nx9647), .A (nx10321)) ;
    inv04 ix9648 (.Y (nx9649), .A (nx10323)) ;
    inv04 ix9650 (.Y (nx9651), .A (nx3611)) ;
    inv04 ix9652 (.Y (nx9653), .A (nx3611)) ;
    inv04 ix9654 (.Y (nx9655), .A (nx3611)) ;
    inv04 ix9656 (.Y (nx9657), .A (nx10281)) ;
    inv04 ix9658 (.Y (nx9659), .A (nx10281)) ;
    inv04 ix9660 (.Y (nx9661), .A (nx10283)) ;
    inv04 ix9662 (.Y (nx9663), .A (nx3363)) ;
    inv04 ix9664 (.Y (nx9665), .A (nx3363)) ;
    inv04 ix9666 (.Y (nx9667), .A (nx3363)) ;
    inv04 ix9668 (.Y (nx9669), .A (nx10241)) ;
    inv04 ix9670 (.Y (nx9671), .A (nx10241)) ;
    inv04 ix9672 (.Y (nx9673), .A (nx10243)) ;
    inv04 ix9674 (.Y (nx9675), .A (nx3115)) ;
    inv04 ix9676 (.Y (nx9677), .A (nx3115)) ;
    inv04 ix9678 (.Y (nx9679), .A (nx3115)) ;
    inv04 ix9680 (.Y (nx9681), .A (nx10201)) ;
    inv04 ix9682 (.Y (nx9683), .A (nx10201)) ;
    inv04 ix9684 (.Y (nx9685), .A (nx10203)) ;
    inv04 ix9686 (.Y (nx9687), .A (nx2871)) ;
    inv04 ix9688 (.Y (nx9689), .A (nx2871)) ;
    inv04 ix9690 (.Y (nx9691), .A (nx2871)) ;
    inv04 ix9692 (.Y (nx9693), .A (nx10161)) ;
    inv04 ix9694 (.Y (nx9695), .A (nx10161)) ;
    inv04 ix9696 (.Y (nx9697), .A (nx10163)) ;
    inv01 ix9698 (.Y (nx9699), .A (gen_24_cmp_BSCmp_op2_16)) ;
    inv02 ix9700 (.Y (nx9701), .A (nx9699)) ;
    inv02 ix9702 (.Y (nx9703), .A (nx9699)) ;
    inv02 ix9704 (.Y (nx9705), .A (nx9699)) ;
    inv02 ix9706 (.Y (nx9707), .A (nx9699)) ;
    inv02 ix9708 (.Y (nx9709), .A (nx9699)) ;
    inv01 ix9710 (.Y (nx9711), .A (gen_23_cmp_BSCmp_op2_16)) ;
    inv02 ix9712 (.Y (nx9713), .A (nx9711)) ;
    inv02 ix9714 (.Y (nx9715), .A (nx9711)) ;
    inv02 ix9716 (.Y (nx9717), .A (nx9711)) ;
    inv02 ix9718 (.Y (nx9719), .A (nx9711)) ;
    inv02 ix9720 (.Y (nx9721), .A (nx9711)) ;
    inv01 ix9722 (.Y (nx9723), .A (gen_22_cmp_BSCmp_op2_16)) ;
    inv02 ix9724 (.Y (nx9725), .A (nx9723)) ;
    inv02 ix9726 (.Y (nx9727), .A (nx9723)) ;
    inv02 ix9728 (.Y (nx9729), .A (nx9723)) ;
    inv02 ix9730 (.Y (nx9731), .A (nx9723)) ;
    inv02 ix9732 (.Y (nx9733), .A (nx9723)) ;
    inv01 ix9734 (.Y (nx9735), .A (gen_21_cmp_BSCmp_op2_16)) ;
    inv02 ix9736 (.Y (nx9737), .A (nx9735)) ;
    inv02 ix9738 (.Y (nx9739), .A (nx9735)) ;
    inv02 ix9740 (.Y (nx9741), .A (nx9735)) ;
    inv02 ix9742 (.Y (nx9743), .A (nx9735)) ;
    inv02 ix9744 (.Y (nx9745), .A (nx9735)) ;
    inv01 ix9746 (.Y (nx9747), .A (gen_20_cmp_BSCmp_op2_16)) ;
    inv02 ix9748 (.Y (nx9749), .A (nx9747)) ;
    inv02 ix9750 (.Y (nx9751), .A (nx9747)) ;
    inv02 ix9752 (.Y (nx9753), .A (nx9747)) ;
    inv02 ix9754 (.Y (nx9755), .A (nx9747)) ;
    inv02 ix9756 (.Y (nx9757), .A (nx9747)) ;
    inv01 ix9758 (.Y (nx9759), .A (gen_19_cmp_BSCmp_op2_16)) ;
    inv02 ix9760 (.Y (nx9761), .A (nx9759)) ;
    inv02 ix9762 (.Y (nx9763), .A (nx9759)) ;
    inv02 ix9764 (.Y (nx9765), .A (nx9759)) ;
    inv02 ix9766 (.Y (nx9767), .A (nx9759)) ;
    inv02 ix9768 (.Y (nx9769), .A (nx9759)) ;
    inv01 ix9770 (.Y (nx9771), .A (gen_18_cmp_BSCmp_op2_16)) ;
    inv02 ix9772 (.Y (nx9773), .A (nx9771)) ;
    inv02 ix9774 (.Y (nx9775), .A (nx9771)) ;
    inv02 ix9776 (.Y (nx9777), .A (nx9771)) ;
    inv02 ix9778 (.Y (nx9779), .A (nx9771)) ;
    inv02 ix9780 (.Y (nx9781), .A (nx9771)) ;
    inv01 ix9782 (.Y (nx9783), .A (gen_17_cmp_BSCmp_op2_16)) ;
    inv02 ix9784 (.Y (nx9785), .A (nx9783)) ;
    inv02 ix9786 (.Y (nx9787), .A (nx9783)) ;
    inv02 ix9788 (.Y (nx9789), .A (nx9783)) ;
    inv02 ix9790 (.Y (nx9791), .A (nx9783)) ;
    inv02 ix9792 (.Y (nx9793), .A (nx9783)) ;
    inv01 ix9794 (.Y (nx9795), .A (gen_16_cmp_BSCmp_op2_16)) ;
    inv02 ix9796 (.Y (nx9797), .A (nx9795)) ;
    inv02 ix9798 (.Y (nx9799), .A (nx9795)) ;
    inv02 ix9800 (.Y (nx9801), .A (nx9795)) ;
    inv02 ix9802 (.Y (nx9803), .A (nx9795)) ;
    inv02 ix9804 (.Y (nx9805), .A (nx9795)) ;
    inv01 ix9806 (.Y (nx9807), .A (gen_15_cmp_BSCmp_op2_16)) ;
    inv02 ix9808 (.Y (nx9809), .A (nx9807)) ;
    inv02 ix9810 (.Y (nx9811), .A (nx9807)) ;
    inv02 ix9812 (.Y (nx9813), .A (nx9807)) ;
    inv02 ix9814 (.Y (nx9815), .A (nx9807)) ;
    inv02 ix9816 (.Y (nx9817), .A (nx9807)) ;
    inv01 ix9818 (.Y (nx9819), .A (gen_14_cmp_BSCmp_op2_16)) ;
    inv02 ix9820 (.Y (nx9821), .A (nx9819)) ;
    inv02 ix9822 (.Y (nx9823), .A (nx9819)) ;
    inv02 ix9824 (.Y (nx9825), .A (nx9819)) ;
    inv02 ix9826 (.Y (nx9827), .A (nx9819)) ;
    inv02 ix9828 (.Y (nx9829), .A (nx9819)) ;
    inv01 ix9830 (.Y (nx9831), .A (gen_13_cmp_BSCmp_op2_16)) ;
    inv02 ix9832 (.Y (nx9833), .A (nx9831)) ;
    inv02 ix9834 (.Y (nx9835), .A (nx9831)) ;
    inv02 ix9836 (.Y (nx9837), .A (nx9831)) ;
    inv02 ix9838 (.Y (nx9839), .A (nx9831)) ;
    inv02 ix9840 (.Y (nx9841), .A (nx9831)) ;
    inv01 ix9842 (.Y (nx9843), .A (gen_12_cmp_BSCmp_op2_16)) ;
    inv02 ix9844 (.Y (nx9845), .A (nx9843)) ;
    inv02 ix9846 (.Y (nx9847), .A (nx9843)) ;
    inv02 ix9848 (.Y (nx9849), .A (nx9843)) ;
    inv02 ix9850 (.Y (nx9851), .A (nx9843)) ;
    inv02 ix9852 (.Y (nx9853), .A (nx9843)) ;
    inv01 ix9854 (.Y (nx9855), .A (gen_11_cmp_BSCmp_op2_16)) ;
    inv02 ix9856 (.Y (nx9857), .A (nx9855)) ;
    inv02 ix9858 (.Y (nx9859), .A (nx9855)) ;
    inv02 ix9860 (.Y (nx9861), .A (nx9855)) ;
    inv02 ix9862 (.Y (nx9863), .A (nx9855)) ;
    inv02 ix9864 (.Y (nx9865), .A (nx9855)) ;
    inv01 ix9866 (.Y (nx9867), .A (gen_10_cmp_BSCmp_op2_16)) ;
    inv02 ix9868 (.Y (nx9869), .A (nx9867)) ;
    inv02 ix9870 (.Y (nx9871), .A (nx9867)) ;
    inv02 ix9872 (.Y (nx9873), .A (nx9867)) ;
    inv02 ix9874 (.Y (nx9875), .A (nx9867)) ;
    inv02 ix9876 (.Y (nx9877), .A (nx9867)) ;
    inv01 ix9878 (.Y (nx9879), .A (gen_9_cmp_BSCmp_op2_16)) ;
    inv02 ix9880 (.Y (nx9881), .A (nx9879)) ;
    inv02 ix9882 (.Y (nx9883), .A (nx9879)) ;
    inv02 ix9884 (.Y (nx9885), .A (nx9879)) ;
    inv02 ix9886 (.Y (nx9887), .A (nx9879)) ;
    inv02 ix9888 (.Y (nx9889), .A (nx9879)) ;
    inv01 ix9890 (.Y (nx9891), .A (gen_8_cmp_BSCmp_op2_16)) ;
    inv02 ix9892 (.Y (nx9893), .A (nx9891)) ;
    inv02 ix9894 (.Y (nx9895), .A (nx9891)) ;
    inv02 ix9896 (.Y (nx9897), .A (nx9891)) ;
    inv02 ix9898 (.Y (nx9899), .A (nx9891)) ;
    inv02 ix9900 (.Y (nx9901), .A (nx9891)) ;
    inv01 ix9902 (.Y (nx9903), .A (gen_7_cmp_BSCmp_op2_16)) ;
    inv02 ix9904 (.Y (nx9905), .A (nx9903)) ;
    inv02 ix9906 (.Y (nx9907), .A (nx9903)) ;
    inv02 ix9908 (.Y (nx9909), .A (nx9903)) ;
    inv02 ix9910 (.Y (nx9911), .A (nx9903)) ;
    inv02 ix9912 (.Y (nx9913), .A (nx9903)) ;
    inv01 ix9914 (.Y (nx9915), .A (gen_6_cmp_BSCmp_op2_16)) ;
    inv02 ix9916 (.Y (nx9917), .A (nx9915)) ;
    inv02 ix9918 (.Y (nx9919), .A (nx9915)) ;
    inv02 ix9920 (.Y (nx9921), .A (nx9915)) ;
    inv02 ix9922 (.Y (nx9923), .A (nx9915)) ;
    inv02 ix9924 (.Y (nx9925), .A (nx9915)) ;
    inv01 ix9926 (.Y (nx9927), .A (gen_5_cmp_BSCmp_op2_16)) ;
    inv02 ix9928 (.Y (nx9929), .A (nx9927)) ;
    inv02 ix9930 (.Y (nx9931), .A (nx9927)) ;
    inv02 ix9932 (.Y (nx9933), .A (nx9927)) ;
    inv02 ix9934 (.Y (nx9935), .A (nx9927)) ;
    inv02 ix9936 (.Y (nx9937), .A (nx9927)) ;
    inv01 ix9938 (.Y (nx9939), .A (gen_4_cmp_BSCmp_op2_16)) ;
    inv02 ix9940 (.Y (nx9941), .A (nx9939)) ;
    inv02 ix9942 (.Y (nx9943), .A (nx9939)) ;
    inv02 ix9944 (.Y (nx9945), .A (nx9939)) ;
    inv02 ix9946 (.Y (nx9947), .A (nx9939)) ;
    inv02 ix9948 (.Y (nx9949), .A (nx9939)) ;
    inv01 ix9950 (.Y (nx9951), .A (gen_3_cmp_BSCmp_op2_16)) ;
    inv02 ix9952 (.Y (nx9953), .A (nx9951)) ;
    inv02 ix9954 (.Y (nx9955), .A (nx9951)) ;
    inv02 ix9956 (.Y (nx9957), .A (nx9951)) ;
    inv02 ix9958 (.Y (nx9959), .A (nx9951)) ;
    inv02 ix9960 (.Y (nx9961), .A (nx9951)) ;
    inv01 ix9962 (.Y (nx9963), .A (gen_2_cmp_BSCmp_op2_16)) ;
    inv02 ix9964 (.Y (nx9965), .A (nx9963)) ;
    inv02 ix9966 (.Y (nx9967), .A (nx9963)) ;
    inv02 ix9968 (.Y (nx9969), .A (nx9963)) ;
    inv02 ix9970 (.Y (nx9971), .A (nx9963)) ;
    inv02 ix9972 (.Y (nx9973), .A (nx9963)) ;
    inv01 ix9974 (.Y (nx9975), .A (gen_1_cmp_BSCmp_op2_16)) ;
    inv02 ix9976 (.Y (nx9977), .A (nx9975)) ;
    inv02 ix9978 (.Y (nx9979), .A (nx9975)) ;
    inv02 ix9980 (.Y (nx9981), .A (nx9975)) ;
    inv02 ix9982 (.Y (nx9983), .A (nx9975)) ;
    inv02 ix9984 (.Y (nx9985), .A (nx9975)) ;
    inv01 ix9986 (.Y (nx9987), .A (gen_0_cmp_BSCmp_op2_16)) ;
    inv02 ix9988 (.Y (nx9989), .A (nx9987)) ;
    inv02 ix9990 (.Y (nx9991), .A (nx9987)) ;
    inv02 ix9992 (.Y (nx9993), .A (nx9987)) ;
    inv02 ix9994 (.Y (nx9995), .A (nx9987)) ;
    inv02 ix9996 (.Y (nx9997), .A (nx9987)) ;
    buf02 ix9998 (.Y (nx9999), .A (nx6)) ;
    buf02 ix10000 (.Y (nx10001), .A (nx6)) ;
    buf02 ix10002 (.Y (nx10003), .A (nx6)) ;
    buf02 ix10004 (.Y (nx10005), .A (nx392)) ;
    buf02 ix10006 (.Y (nx10007), .A (nx392)) ;
    buf02 ix10008 (.Y (nx10009), .A (nx392)) ;
    buf02 ix10010 (.Y (nx10011), .A (nx778)) ;
    buf02 ix10012 (.Y (nx10013), .A (nx778)) ;
    buf02 ix10014 (.Y (nx10015), .A (nx778)) ;
    buf02 ix10016 (.Y (nx10017), .A (nx1164)) ;
    buf02 ix10018 (.Y (nx10019), .A (nx1164)) ;
    buf02 ix10020 (.Y (nx10021), .A (nx1164)) ;
    buf02 ix10022 (.Y (nx10023), .A (nx1550)) ;
    buf02 ix10024 (.Y (nx10025), .A (nx1550)) ;
    buf02 ix10026 (.Y (nx10027), .A (nx1550)) ;
    buf02 ix10028 (.Y (nx10029), .A (nx1936)) ;
    buf02 ix10030 (.Y (nx10031), .A (nx1936)) ;
    buf02 ix10032 (.Y (nx10033), .A (nx1936)) ;
    buf02 ix10034 (.Y (nx10035), .A (nx2322)) ;
    buf02 ix10036 (.Y (nx10037), .A (nx2322)) ;
    buf02 ix10038 (.Y (nx10039), .A (nx2322)) ;
    buf02 ix10040 (.Y (nx10041), .A (nx2708)) ;
    buf02 ix10042 (.Y (nx10043), .A (nx2708)) ;
    buf02 ix10044 (.Y (nx10045), .A (nx2708)) ;
    buf02 ix10046 (.Y (nx10047), .A (nx3094)) ;
    buf02 ix10048 (.Y (nx10049), .A (nx3094)) ;
    buf02 ix10050 (.Y (nx10051), .A (nx3094)) ;
    buf02 ix10052 (.Y (nx10053), .A (nx3480)) ;
    buf02 ix10054 (.Y (nx10055), .A (nx3480)) ;
    buf02 ix10056 (.Y (nx10057), .A (nx3480)) ;
    buf02 ix10058 (.Y (nx10059), .A (nx3866)) ;
    buf02 ix10060 (.Y (nx10061), .A (nx3866)) ;
    buf02 ix10062 (.Y (nx10063), .A (nx3866)) ;
    buf02 ix10064 (.Y (nx10065), .A (nx4252)) ;
    buf02 ix10066 (.Y (nx10067), .A (nx4252)) ;
    buf02 ix10068 (.Y (nx10069), .A (nx4252)) ;
    buf02 ix10070 (.Y (nx10071), .A (nx4638)) ;
    buf02 ix10072 (.Y (nx10073), .A (nx4638)) ;
    buf02 ix10074 (.Y (nx10075), .A (nx4638)) ;
    buf02 ix10076 (.Y (nx10077), .A (nx5024)) ;
    buf02 ix10078 (.Y (nx10079), .A (nx5024)) ;
    buf02 ix10080 (.Y (nx10081), .A (nx5024)) ;
    buf02 ix10082 (.Y (nx10083), .A (nx5410)) ;
    buf02 ix10084 (.Y (nx10085), .A (nx5410)) ;
    buf02 ix10086 (.Y (nx10087), .A (nx5410)) ;
    buf02 ix10088 (.Y (nx10089), .A (nx5796)) ;
    buf02 ix10090 (.Y (nx10091), .A (nx5796)) ;
    buf02 ix10092 (.Y (nx10093), .A (nx5796)) ;
    buf02 ix10094 (.Y (nx10095), .A (nx6182)) ;
    buf02 ix10096 (.Y (nx10097), .A (nx6182)) ;
    buf02 ix10098 (.Y (nx10099), .A (nx6182)) ;
    buf02 ix10100 (.Y (nx10101), .A (nx6568)) ;
    buf02 ix10102 (.Y (nx10103), .A (nx6568)) ;
    buf02 ix10104 (.Y (nx10105), .A (nx6568)) ;
    buf02 ix10106 (.Y (nx10107), .A (nx6954)) ;
    buf02 ix10108 (.Y (nx10109), .A (nx6954)) ;
    buf02 ix10110 (.Y (nx10111), .A (nx6954)) ;
    buf02 ix10112 (.Y (nx10113), .A (nx7340)) ;
    buf02 ix10114 (.Y (nx10115), .A (nx7340)) ;
    buf02 ix10116 (.Y (nx10117), .A (nx7340)) ;
    buf02 ix10118 (.Y (nx10119), .A (nx7726)) ;
    buf02 ix10120 (.Y (nx10121), .A (nx7726)) ;
    buf02 ix10122 (.Y (nx10123), .A (nx7726)) ;
    buf02 ix10124 (.Y (nx10125), .A (nx8112)) ;
    buf02 ix10126 (.Y (nx10127), .A (nx8112)) ;
    buf02 ix10128 (.Y (nx10129), .A (nx8112)) ;
    buf02 ix10130 (.Y (nx10131), .A (nx8498)) ;
    buf02 ix10132 (.Y (nx10133), .A (nx8498)) ;
    buf02 ix10134 (.Y (nx10135), .A (nx8498)) ;
    buf02 ix10136 (.Y (nx10137), .A (nx8884)) ;
    buf02 ix10138 (.Y (nx10139), .A (nx8884)) ;
    buf02 ix10140 (.Y (nx10141), .A (nx8884)) ;
    buf02 ix10142 (.Y (nx10143), .A (nx9270)) ;
    buf02 ix10144 (.Y (nx10145), .A (nx9270)) ;
    buf02 ix10146 (.Y (nx10147), .A (nx9270)) ;
    inv02 ix10150 (.Y (nx10151), .A (nx10149)) ;
    inv02 ix10152 (.Y (nx10153), .A (nx10149)) ;
    inv02 ix10154 (.Y (nx10155), .A (nx10149)) ;
    inv04 ix10156 (.Y (nx10157), .A (gen_0_cmp_pMux_1)) ;
    inv04 ix10158 (.Y (nx10159), .A (gen_0_cmp_pMux_1)) ;
    inv04 ix10160 (.Y (nx10161), .A (gen_0_cmp_pMux_1)) ;
    inv04 ix10162 (.Y (nx10163), .A (gen_0_cmp_pMux_1)) ;
    inv02 ix10166 (.Y (nx10167), .A (nx10165)) ;
    inv02 ix10168 (.Y (nx10169), .A (nx10165)) ;
    inv02 ix10170 (.Y (nx10171), .A (nx10165)) ;
    inv02 ix10174 (.Y (nx10175), .A (nx10173)) ;
    inv02 ix10176 (.Y (nx10177), .A (nx10173)) ;
    inv02 ix10178 (.Y (nx10179), .A (nx10173)) ;
    inv02 ix10182 (.Y (nx10183), .A (nx10181)) ;
    inv02 ix10184 (.Y (nx10185), .A (nx10181)) ;
    inv02 ix10186 (.Y (nx10187), .A (nx10181)) ;
    inv02 ix10190 (.Y (nx10191), .A (nx10189)) ;
    inv02 ix10192 (.Y (nx10193), .A (nx10189)) ;
    inv02 ix10194 (.Y (nx10195), .A (nx10189)) ;
    inv04 ix10196 (.Y (nx10197), .A (gen_1_cmp_pMux_1)) ;
    inv04 ix10198 (.Y (nx10199), .A (gen_1_cmp_pMux_1)) ;
    inv04 ix10200 (.Y (nx10201), .A (gen_1_cmp_pMux_1)) ;
    inv04 ix10202 (.Y (nx10203), .A (gen_1_cmp_pMux_1)) ;
    inv02 ix10206 (.Y (nx10207), .A (nx10205)) ;
    inv02 ix10208 (.Y (nx10209), .A (nx10205)) ;
    inv02 ix10210 (.Y (nx10211), .A (nx10205)) ;
    inv02 ix10214 (.Y (nx10215), .A (nx10213)) ;
    inv02 ix10216 (.Y (nx10217), .A (nx10213)) ;
    inv02 ix10218 (.Y (nx10219), .A (nx10213)) ;
    inv02 ix10222 (.Y (nx10223), .A (nx10221)) ;
    inv02 ix10224 (.Y (nx10225), .A (nx10221)) ;
    inv02 ix10226 (.Y (nx10227), .A (nx10221)) ;
    inv02 ix10230 (.Y (nx10231), .A (nx10229)) ;
    inv02 ix10232 (.Y (nx10233), .A (nx10229)) ;
    inv02 ix10234 (.Y (nx10235), .A (nx10229)) ;
    inv04 ix10236 (.Y (nx10237), .A (gen_2_cmp_pMux_1)) ;
    inv04 ix10238 (.Y (nx10239), .A (gen_2_cmp_pMux_1)) ;
    inv04 ix10240 (.Y (nx10241), .A (gen_2_cmp_pMux_1)) ;
    inv04 ix10242 (.Y (nx10243), .A (gen_2_cmp_pMux_1)) ;
    inv02 ix10246 (.Y (nx10247), .A (nx10245)) ;
    inv02 ix10248 (.Y (nx10249), .A (nx10245)) ;
    inv02 ix10250 (.Y (nx10251), .A (nx10245)) ;
    inv02 ix10254 (.Y (nx10255), .A (nx10253)) ;
    inv02 ix10256 (.Y (nx10257), .A (nx10253)) ;
    inv02 ix10258 (.Y (nx10259), .A (nx10253)) ;
    inv02 ix10262 (.Y (nx10263), .A (nx10261)) ;
    inv02 ix10264 (.Y (nx10265), .A (nx10261)) ;
    inv02 ix10266 (.Y (nx10267), .A (nx10261)) ;
    inv02 ix10270 (.Y (nx10271), .A (nx10269)) ;
    inv02 ix10272 (.Y (nx10273), .A (nx10269)) ;
    inv02 ix10274 (.Y (nx10275), .A (nx10269)) ;
    inv04 ix10276 (.Y (nx10277), .A (gen_3_cmp_pMux_1)) ;
    inv04 ix10278 (.Y (nx10279), .A (gen_3_cmp_pMux_1)) ;
    inv04 ix10280 (.Y (nx10281), .A (gen_3_cmp_pMux_1)) ;
    inv04 ix10282 (.Y (nx10283), .A (gen_3_cmp_pMux_1)) ;
    inv02 ix10286 (.Y (nx10287), .A (nx10285)) ;
    inv02 ix10288 (.Y (nx10289), .A (nx10285)) ;
    inv02 ix10290 (.Y (nx10291), .A (nx10285)) ;
    inv02 ix10294 (.Y (nx10295), .A (nx10293)) ;
    inv02 ix10296 (.Y (nx10297), .A (nx10293)) ;
    inv02 ix10298 (.Y (nx10299), .A (nx10293)) ;
    inv02 ix10302 (.Y (nx10303), .A (nx10301)) ;
    inv02 ix10304 (.Y (nx10305), .A (nx10301)) ;
    inv02 ix10306 (.Y (nx10307), .A (nx10301)) ;
    inv02 ix10310 (.Y (nx10311), .A (nx10309)) ;
    inv02 ix10312 (.Y (nx10313), .A (nx10309)) ;
    inv02 ix10314 (.Y (nx10315), .A (nx10309)) ;
    inv04 ix10316 (.Y (nx10317), .A (gen_4_cmp_pMux_1)) ;
    inv04 ix10318 (.Y (nx10319), .A (gen_4_cmp_pMux_1)) ;
    inv04 ix10320 (.Y (nx10321), .A (gen_4_cmp_pMux_1)) ;
    inv04 ix10322 (.Y (nx10323), .A (gen_4_cmp_pMux_1)) ;
    inv02 ix10326 (.Y (nx10327), .A (nx10325)) ;
    inv02 ix10328 (.Y (nx10329), .A (nx10325)) ;
    inv02 ix10330 (.Y (nx10331), .A (nx10325)) ;
    inv02 ix10334 (.Y (nx10335), .A (nx10333)) ;
    inv02 ix10336 (.Y (nx10337), .A (nx10333)) ;
    inv02 ix10338 (.Y (nx10339), .A (nx10333)) ;
    inv02 ix10342 (.Y (nx10343), .A (nx10341)) ;
    inv02 ix10344 (.Y (nx10345), .A (nx10341)) ;
    inv02 ix10346 (.Y (nx10347), .A (nx10341)) ;
    inv02 ix10350 (.Y (nx10351), .A (nx10349)) ;
    inv02 ix10352 (.Y (nx10353), .A (nx10349)) ;
    inv02 ix10354 (.Y (nx10355), .A (nx10349)) ;
    inv04 ix10356 (.Y (nx10357), .A (gen_5_cmp_pMux_1)) ;
    inv04 ix10358 (.Y (nx10359), .A (gen_5_cmp_pMux_1)) ;
    inv04 ix10360 (.Y (nx10361), .A (gen_5_cmp_pMux_1)) ;
    inv04 ix10362 (.Y (nx10363), .A (gen_5_cmp_pMux_1)) ;
    inv02 ix10366 (.Y (nx10367), .A (nx10365)) ;
    inv02 ix10368 (.Y (nx10369), .A (nx10365)) ;
    inv02 ix10370 (.Y (nx10371), .A (nx10365)) ;
    inv02 ix10374 (.Y (nx10375), .A (nx10373)) ;
    inv02 ix10376 (.Y (nx10377), .A (nx10373)) ;
    inv02 ix10378 (.Y (nx10379), .A (nx10373)) ;
    inv02 ix10382 (.Y (nx10383), .A (nx10381)) ;
    inv02 ix10384 (.Y (nx10385), .A (nx10381)) ;
    inv02 ix10386 (.Y (nx10387), .A (nx10381)) ;
    inv02 ix10390 (.Y (nx10391), .A (nx10389)) ;
    inv02 ix10392 (.Y (nx10393), .A (nx10389)) ;
    inv02 ix10394 (.Y (nx10395), .A (nx10389)) ;
    inv04 ix10396 (.Y (nx10397), .A (gen_6_cmp_pMux_1)) ;
    inv04 ix10398 (.Y (nx10399), .A (gen_6_cmp_pMux_1)) ;
    inv04 ix10400 (.Y (nx10401), .A (gen_6_cmp_pMux_1)) ;
    inv04 ix10402 (.Y (nx10403), .A (gen_6_cmp_pMux_1)) ;
    inv02 ix10406 (.Y (nx10407), .A (nx10405)) ;
    inv02 ix10408 (.Y (nx10409), .A (nx10405)) ;
    inv02 ix10410 (.Y (nx10411), .A (nx10405)) ;
    inv02 ix10414 (.Y (nx10415), .A (nx10413)) ;
    inv02 ix10416 (.Y (nx10417), .A (nx10413)) ;
    inv02 ix10418 (.Y (nx10419), .A (nx10413)) ;
    inv02 ix10422 (.Y (nx10423), .A (nx10421)) ;
    inv02 ix10424 (.Y (nx10425), .A (nx10421)) ;
    inv02 ix10426 (.Y (nx10427), .A (nx10421)) ;
    inv02 ix10430 (.Y (nx10431), .A (nx10429)) ;
    inv02 ix10432 (.Y (nx10433), .A (nx10429)) ;
    inv02 ix10434 (.Y (nx10435), .A (nx10429)) ;
    inv04 ix10436 (.Y (nx10437), .A (gen_7_cmp_pMux_1)) ;
    inv04 ix10438 (.Y (nx10439), .A (gen_7_cmp_pMux_1)) ;
    inv04 ix10440 (.Y (nx10441), .A (gen_7_cmp_pMux_1)) ;
    inv04 ix10442 (.Y (nx10443), .A (gen_7_cmp_pMux_1)) ;
    inv02 ix10446 (.Y (nx10447), .A (nx10445)) ;
    inv02 ix10448 (.Y (nx10449), .A (nx10445)) ;
    inv02 ix10450 (.Y (nx10451), .A (nx10445)) ;
    inv02 ix10454 (.Y (nx10455), .A (nx10453)) ;
    inv02 ix10456 (.Y (nx10457), .A (nx10453)) ;
    inv02 ix10458 (.Y (nx10459), .A (nx10453)) ;
    inv02 ix10462 (.Y (nx10463), .A (nx10461)) ;
    inv02 ix10464 (.Y (nx10465), .A (nx10461)) ;
    inv02 ix10466 (.Y (nx10467), .A (nx10461)) ;
    inv02 ix10470 (.Y (nx10471), .A (nx10469)) ;
    inv02 ix10472 (.Y (nx10473), .A (nx10469)) ;
    inv02 ix10474 (.Y (nx10475), .A (nx10469)) ;
    inv04 ix10476 (.Y (nx10477), .A (gen_8_cmp_pMux_1)) ;
    inv04 ix10478 (.Y (nx10479), .A (gen_8_cmp_pMux_1)) ;
    inv04 ix10480 (.Y (nx10481), .A (gen_8_cmp_pMux_1)) ;
    inv04 ix10482 (.Y (nx10483), .A (gen_8_cmp_pMux_1)) ;
    inv02 ix10486 (.Y (nx10487), .A (nx10485)) ;
    inv02 ix10488 (.Y (nx10489), .A (nx10485)) ;
    inv02 ix10490 (.Y (nx10491), .A (nx10485)) ;
    inv02 ix10494 (.Y (nx10495), .A (nx10493)) ;
    inv02 ix10496 (.Y (nx10497), .A (nx10493)) ;
    inv02 ix10498 (.Y (nx10499), .A (nx10493)) ;
    inv02 ix10502 (.Y (nx10503), .A (nx10501)) ;
    inv02 ix10504 (.Y (nx10505), .A (nx10501)) ;
    inv02 ix10506 (.Y (nx10507), .A (nx10501)) ;
    inv02 ix10510 (.Y (nx10511), .A (nx10509)) ;
    inv02 ix10512 (.Y (nx10513), .A (nx10509)) ;
    inv02 ix10514 (.Y (nx10515), .A (nx10509)) ;
    inv04 ix10516 (.Y (nx10517), .A (gen_9_cmp_pMux_1)) ;
    inv04 ix10518 (.Y (nx10519), .A (gen_9_cmp_pMux_1)) ;
    inv04 ix10520 (.Y (nx10521), .A (gen_9_cmp_pMux_1)) ;
    inv04 ix10522 (.Y (nx10523), .A (gen_9_cmp_pMux_1)) ;
    inv02 ix10526 (.Y (nx10527), .A (nx10525)) ;
    inv02 ix10528 (.Y (nx10529), .A (nx10525)) ;
    inv02 ix10530 (.Y (nx10531), .A (nx10525)) ;
    inv02 ix10534 (.Y (nx10535), .A (nx10533)) ;
    inv02 ix10536 (.Y (nx10537), .A (nx10533)) ;
    inv02 ix10538 (.Y (nx10539), .A (nx10533)) ;
    inv02 ix10542 (.Y (nx10543), .A (nx10541)) ;
    inv02 ix10544 (.Y (nx10545), .A (nx10541)) ;
    inv02 ix10546 (.Y (nx10547), .A (nx10541)) ;
    inv02 ix10550 (.Y (nx10551), .A (nx10549)) ;
    inv02 ix10552 (.Y (nx10553), .A (nx10549)) ;
    inv02 ix10554 (.Y (nx10555), .A (nx10549)) ;
    inv04 ix10556 (.Y (nx10557), .A (gen_10_cmp_pMux_1)) ;
    inv04 ix10558 (.Y (nx10559), .A (gen_10_cmp_pMux_1)) ;
    inv04 ix10560 (.Y (nx10561), .A (gen_10_cmp_pMux_1)) ;
    inv04 ix10562 (.Y (nx10563), .A (gen_10_cmp_pMux_1)) ;
    inv02 ix10566 (.Y (nx10567), .A (nx10565)) ;
    inv02 ix10568 (.Y (nx10569), .A (nx10565)) ;
    inv02 ix10570 (.Y (nx10571), .A (nx10565)) ;
    inv02 ix10574 (.Y (nx10575), .A (nx10573)) ;
    inv02 ix10576 (.Y (nx10577), .A (nx10573)) ;
    inv02 ix10578 (.Y (nx10579), .A (nx10573)) ;
    inv02 ix10582 (.Y (nx10583), .A (nx10581)) ;
    inv02 ix10584 (.Y (nx10585), .A (nx10581)) ;
    inv02 ix10586 (.Y (nx10587), .A (nx10581)) ;
    inv02 ix10590 (.Y (nx10591), .A (nx10589)) ;
    inv02 ix10592 (.Y (nx10593), .A (nx10589)) ;
    inv02 ix10594 (.Y (nx10595), .A (nx10589)) ;
    inv04 ix10596 (.Y (nx10597), .A (gen_11_cmp_pMux_1)) ;
    inv04 ix10598 (.Y (nx10599), .A (gen_11_cmp_pMux_1)) ;
    inv04 ix10600 (.Y (nx10601), .A (gen_11_cmp_pMux_1)) ;
    inv04 ix10602 (.Y (nx10603), .A (gen_11_cmp_pMux_1)) ;
    inv02 ix10606 (.Y (nx10607), .A (nx10605)) ;
    inv02 ix10608 (.Y (nx10609), .A (nx10605)) ;
    inv02 ix10610 (.Y (nx10611), .A (nx10605)) ;
    inv02 ix10614 (.Y (nx10615), .A (nx10613)) ;
    inv02 ix10616 (.Y (nx10617), .A (nx10613)) ;
    inv02 ix10618 (.Y (nx10619), .A (nx10613)) ;
    inv02 ix10622 (.Y (nx10623), .A (nx10621)) ;
    inv02 ix10624 (.Y (nx10625), .A (nx10621)) ;
    inv02 ix10626 (.Y (nx10627), .A (nx10621)) ;
    inv02 ix10630 (.Y (nx10631), .A (nx10629)) ;
    inv02 ix10632 (.Y (nx10633), .A (nx10629)) ;
    inv02 ix10634 (.Y (nx10635), .A (nx10629)) ;
    inv04 ix10636 (.Y (nx10637), .A (gen_12_cmp_pMux_1)) ;
    inv04 ix10638 (.Y (nx10639), .A (gen_12_cmp_pMux_1)) ;
    inv04 ix10640 (.Y (nx10641), .A (gen_12_cmp_pMux_1)) ;
    inv04 ix10642 (.Y (nx10643), .A (gen_12_cmp_pMux_1)) ;
    inv02 ix10646 (.Y (nx10647), .A (nx10645)) ;
    inv02 ix10648 (.Y (nx10649), .A (nx10645)) ;
    inv02 ix10650 (.Y (nx10651), .A (nx10645)) ;
    inv02 ix10654 (.Y (nx10655), .A (nx10653)) ;
    inv02 ix10656 (.Y (nx10657), .A (nx10653)) ;
    inv02 ix10658 (.Y (nx10659), .A (nx10653)) ;
    inv02 ix10662 (.Y (nx10663), .A (nx10661)) ;
    inv02 ix10664 (.Y (nx10665), .A (nx10661)) ;
    inv02 ix10666 (.Y (nx10667), .A (nx10661)) ;
    inv02 ix10670 (.Y (nx10671), .A (nx10669)) ;
    inv02 ix10672 (.Y (nx10673), .A (nx10669)) ;
    inv02 ix10674 (.Y (nx10675), .A (nx10669)) ;
    inv04 ix10676 (.Y (nx10677), .A (gen_13_cmp_pMux_1)) ;
    inv04 ix10678 (.Y (nx10679), .A (gen_13_cmp_pMux_1)) ;
    inv04 ix10680 (.Y (nx10681), .A (gen_13_cmp_pMux_1)) ;
    inv04 ix10682 (.Y (nx10683), .A (gen_13_cmp_pMux_1)) ;
    inv02 ix10686 (.Y (nx10687), .A (nx10685)) ;
    inv02 ix10688 (.Y (nx10689), .A (nx10685)) ;
    inv02 ix10690 (.Y (nx10691), .A (nx10685)) ;
    inv02 ix10694 (.Y (nx10695), .A (nx10693)) ;
    inv02 ix10696 (.Y (nx10697), .A (nx10693)) ;
    inv02 ix10698 (.Y (nx10699), .A (nx10693)) ;
    inv02 ix10702 (.Y (nx10703), .A (nx10701)) ;
    inv02 ix10704 (.Y (nx10705), .A (nx10701)) ;
    inv02 ix10706 (.Y (nx10707), .A (nx10701)) ;
    inv02 ix10710 (.Y (nx10711), .A (nx10709)) ;
    inv02 ix10712 (.Y (nx10713), .A (nx10709)) ;
    inv02 ix10714 (.Y (nx10715), .A (nx10709)) ;
    inv04 ix10716 (.Y (nx10717), .A (gen_14_cmp_pMux_1)) ;
    inv04 ix10718 (.Y (nx10719), .A (gen_14_cmp_pMux_1)) ;
    inv04 ix10720 (.Y (nx10721), .A (gen_14_cmp_pMux_1)) ;
    inv04 ix10722 (.Y (nx10723), .A (gen_14_cmp_pMux_1)) ;
    inv02 ix10726 (.Y (nx10727), .A (nx10725)) ;
    inv02 ix10728 (.Y (nx10729), .A (nx10725)) ;
    inv02 ix10730 (.Y (nx10731), .A (nx10725)) ;
    inv02 ix10734 (.Y (nx10735), .A (nx10733)) ;
    inv02 ix10736 (.Y (nx10737), .A (nx10733)) ;
    inv02 ix10738 (.Y (nx10739), .A (nx10733)) ;
    inv02 ix10742 (.Y (nx10743), .A (nx10741)) ;
    inv02 ix10744 (.Y (nx10745), .A (nx10741)) ;
    inv02 ix10746 (.Y (nx10747), .A (nx10741)) ;
    inv02 ix10750 (.Y (nx10751), .A (nx10749)) ;
    inv02 ix10752 (.Y (nx10753), .A (nx10749)) ;
    inv02 ix10754 (.Y (nx10755), .A (nx10749)) ;
    inv04 ix10756 (.Y (nx10757), .A (gen_15_cmp_pMux_1)) ;
    inv04 ix10758 (.Y (nx10759), .A (gen_15_cmp_pMux_1)) ;
    inv04 ix10760 (.Y (nx10761), .A (gen_15_cmp_pMux_1)) ;
    inv04 ix10762 (.Y (nx10763), .A (gen_15_cmp_pMux_1)) ;
    inv02 ix10766 (.Y (nx10767), .A (nx10765)) ;
    inv02 ix10768 (.Y (nx10769), .A (nx10765)) ;
    inv02 ix10770 (.Y (nx10771), .A (nx10765)) ;
    inv02 ix10774 (.Y (nx10775), .A (nx10773)) ;
    inv02 ix10776 (.Y (nx10777), .A (nx10773)) ;
    inv02 ix10778 (.Y (nx10779), .A (nx10773)) ;
    inv02 ix10782 (.Y (nx10783), .A (nx10781)) ;
    inv02 ix10784 (.Y (nx10785), .A (nx10781)) ;
    inv02 ix10786 (.Y (nx10787), .A (nx10781)) ;
    inv02 ix10790 (.Y (nx10791), .A (nx10789)) ;
    inv02 ix10792 (.Y (nx10793), .A (nx10789)) ;
    inv02 ix10794 (.Y (nx10795), .A (nx10789)) ;
    inv04 ix10796 (.Y (nx10797), .A (gen_16_cmp_pMux_1)) ;
    inv04 ix10798 (.Y (nx10799), .A (gen_16_cmp_pMux_1)) ;
    inv04 ix10800 (.Y (nx10801), .A (gen_16_cmp_pMux_1)) ;
    inv04 ix10802 (.Y (nx10803), .A (gen_16_cmp_pMux_1)) ;
    inv02 ix10806 (.Y (nx10807), .A (nx10805)) ;
    inv02 ix10808 (.Y (nx10809), .A (nx10805)) ;
    inv02 ix10810 (.Y (nx10811), .A (nx10805)) ;
    inv02 ix10814 (.Y (nx10815), .A (nx10813)) ;
    inv02 ix10816 (.Y (nx10817), .A (nx10813)) ;
    inv02 ix10818 (.Y (nx10819), .A (nx10813)) ;
    inv02 ix10822 (.Y (nx10823), .A (nx10821)) ;
    inv02 ix10824 (.Y (nx10825), .A (nx10821)) ;
    inv02 ix10826 (.Y (nx10827), .A (nx10821)) ;
    inv02 ix10830 (.Y (nx10831), .A (nx10829)) ;
    inv02 ix10832 (.Y (nx10833), .A (nx10829)) ;
    inv02 ix10834 (.Y (nx10835), .A (nx10829)) ;
    inv04 ix10836 (.Y (nx10837), .A (gen_17_cmp_pMux_1)) ;
    inv04 ix10838 (.Y (nx10839), .A (gen_17_cmp_pMux_1)) ;
    inv04 ix10840 (.Y (nx10841), .A (gen_17_cmp_pMux_1)) ;
    inv04 ix10842 (.Y (nx10843), .A (gen_17_cmp_pMux_1)) ;
    inv02 ix10846 (.Y (nx10847), .A (nx10845)) ;
    inv02 ix10848 (.Y (nx10849), .A (nx10845)) ;
    inv02 ix10850 (.Y (nx10851), .A (nx10845)) ;
    inv02 ix10854 (.Y (nx10855), .A (nx10853)) ;
    inv02 ix10856 (.Y (nx10857), .A (nx10853)) ;
    inv02 ix10858 (.Y (nx10859), .A (nx10853)) ;
    inv02 ix10862 (.Y (nx10863), .A (nx10861)) ;
    inv02 ix10864 (.Y (nx10865), .A (nx10861)) ;
    inv02 ix10866 (.Y (nx10867), .A (nx10861)) ;
    inv02 ix10870 (.Y (nx10871), .A (nx10869)) ;
    inv02 ix10872 (.Y (nx10873), .A (nx10869)) ;
    inv02 ix10874 (.Y (nx10875), .A (nx10869)) ;
    inv04 ix10876 (.Y (nx10877), .A (gen_18_cmp_pMux_1)) ;
    inv04 ix10878 (.Y (nx10879), .A (gen_18_cmp_pMux_1)) ;
    inv04 ix10880 (.Y (nx10881), .A (gen_18_cmp_pMux_1)) ;
    inv04 ix10882 (.Y (nx10883), .A (gen_18_cmp_pMux_1)) ;
    inv02 ix10886 (.Y (nx10887), .A (nx10885)) ;
    inv02 ix10888 (.Y (nx10889), .A (nx10885)) ;
    inv02 ix10890 (.Y (nx10891), .A (nx10885)) ;
    inv02 ix10894 (.Y (nx10895), .A (nx10893)) ;
    inv02 ix10896 (.Y (nx10897), .A (nx10893)) ;
    inv02 ix10898 (.Y (nx10899), .A (nx10893)) ;
    inv02 ix10902 (.Y (nx10903), .A (nx10901)) ;
    inv02 ix10904 (.Y (nx10905), .A (nx10901)) ;
    inv02 ix10906 (.Y (nx10907), .A (nx10901)) ;
    inv02 ix10910 (.Y (nx10911), .A (nx10909)) ;
    inv02 ix10912 (.Y (nx10913), .A (nx10909)) ;
    inv02 ix10914 (.Y (nx10915), .A (nx10909)) ;
    inv04 ix10916 (.Y (nx10917), .A (gen_19_cmp_pMux_1)) ;
    inv04 ix10918 (.Y (nx10919), .A (gen_19_cmp_pMux_1)) ;
    inv04 ix10920 (.Y (nx10921), .A (gen_19_cmp_pMux_1)) ;
    inv04 ix10922 (.Y (nx10923), .A (gen_19_cmp_pMux_1)) ;
    inv02 ix10926 (.Y (nx10927), .A (nx10925)) ;
    inv02 ix10928 (.Y (nx10929), .A (nx10925)) ;
    inv02 ix10930 (.Y (nx10931), .A (nx10925)) ;
    inv02 ix10934 (.Y (nx10935), .A (nx10933)) ;
    inv02 ix10936 (.Y (nx10937), .A (nx10933)) ;
    inv02 ix10938 (.Y (nx10939), .A (nx10933)) ;
    inv02 ix10942 (.Y (nx10943), .A (nx10941)) ;
    inv02 ix10944 (.Y (nx10945), .A (nx10941)) ;
    inv02 ix10946 (.Y (nx10947), .A (nx10941)) ;
    inv02 ix10950 (.Y (nx10951), .A (nx10949)) ;
    inv02 ix10952 (.Y (nx10953), .A (nx10949)) ;
    inv02 ix10954 (.Y (nx10955), .A (nx10949)) ;
    inv04 ix10956 (.Y (nx10957), .A (gen_20_cmp_pMux_1)) ;
    inv04 ix10958 (.Y (nx10959), .A (gen_20_cmp_pMux_1)) ;
    inv04 ix10960 (.Y (nx10961), .A (gen_20_cmp_pMux_1)) ;
    inv04 ix10962 (.Y (nx10963), .A (gen_20_cmp_pMux_1)) ;
    inv02 ix10966 (.Y (nx10967), .A (nx10965)) ;
    inv02 ix10968 (.Y (nx10969), .A (nx10965)) ;
    inv02 ix10970 (.Y (nx10971), .A (nx10965)) ;
    inv02 ix10974 (.Y (nx10975), .A (nx10973)) ;
    inv02 ix10976 (.Y (nx10977), .A (nx10973)) ;
    inv02 ix10978 (.Y (nx10979), .A (nx10973)) ;
    inv02 ix10982 (.Y (nx10983), .A (nx10981)) ;
    inv02 ix10984 (.Y (nx10985), .A (nx10981)) ;
    inv02 ix10986 (.Y (nx10987), .A (nx10981)) ;
    inv02 ix10990 (.Y (nx10991), .A (nx10989)) ;
    inv02 ix10992 (.Y (nx10993), .A (nx10989)) ;
    inv02 ix10994 (.Y (nx10995), .A (nx10989)) ;
    inv04 ix10996 (.Y (nx10997), .A (gen_21_cmp_pMux_1)) ;
    inv04 ix10998 (.Y (nx10999), .A (gen_21_cmp_pMux_1)) ;
    inv04 ix11000 (.Y (nx11001), .A (gen_21_cmp_pMux_1)) ;
    inv04 ix11002 (.Y (nx11003), .A (gen_21_cmp_pMux_1)) ;
    inv02 ix11006 (.Y (nx11007), .A (nx11005)) ;
    inv02 ix11008 (.Y (nx11009), .A (nx11005)) ;
    inv02 ix11010 (.Y (nx11011), .A (nx11005)) ;
    inv02 ix11014 (.Y (nx11015), .A (nx11013)) ;
    inv02 ix11016 (.Y (nx11017), .A (nx11013)) ;
    inv02 ix11018 (.Y (nx11019), .A (nx11013)) ;
    inv02 ix11022 (.Y (nx11023), .A (nx11021)) ;
    inv02 ix11024 (.Y (nx11025), .A (nx11021)) ;
    inv02 ix11026 (.Y (nx11027), .A (nx11021)) ;
    inv02 ix11030 (.Y (nx11031), .A (nx11029)) ;
    inv02 ix11032 (.Y (nx11033), .A (nx11029)) ;
    inv02 ix11034 (.Y (nx11035), .A (nx11029)) ;
    inv04 ix11036 (.Y (nx11037), .A (gen_22_cmp_pMux_1)) ;
    inv04 ix11038 (.Y (nx11039), .A (gen_22_cmp_pMux_1)) ;
    inv04 ix11040 (.Y (nx11041), .A (gen_22_cmp_pMux_1)) ;
    inv04 ix11042 (.Y (nx11043), .A (gen_22_cmp_pMux_1)) ;
    inv02 ix11046 (.Y (nx11047), .A (nx11045)) ;
    inv02 ix11048 (.Y (nx11049), .A (nx11045)) ;
    inv02 ix11050 (.Y (nx11051), .A (nx11045)) ;
    inv02 ix11054 (.Y (nx11055), .A (nx11053)) ;
    inv02 ix11056 (.Y (nx11057), .A (nx11053)) ;
    inv02 ix11058 (.Y (nx11059), .A (nx11053)) ;
    inv02 ix11062 (.Y (nx11063), .A (nx11061)) ;
    inv02 ix11064 (.Y (nx11065), .A (nx11061)) ;
    inv02 ix11066 (.Y (nx11067), .A (nx11061)) ;
    inv02 ix11070 (.Y (nx11071), .A (nx11069)) ;
    inv02 ix11072 (.Y (nx11073), .A (nx11069)) ;
    inv02 ix11074 (.Y (nx11075), .A (nx11069)) ;
    inv04 ix11076 (.Y (nx11077), .A (gen_23_cmp_pMux_1)) ;
    inv04 ix11078 (.Y (nx11079), .A (gen_23_cmp_pMux_1)) ;
    inv04 ix11080 (.Y (nx11081), .A (gen_23_cmp_pMux_1)) ;
    inv04 ix11082 (.Y (nx11083), .A (gen_23_cmp_pMux_1)) ;
    inv02 ix11086 (.Y (nx11087), .A (nx11085)) ;
    inv02 ix11088 (.Y (nx11089), .A (nx11085)) ;
    inv02 ix11090 (.Y (nx11091), .A (nx11085)) ;
    inv02 ix11094 (.Y (nx11095), .A (nx11093)) ;
    inv02 ix11096 (.Y (nx11097), .A (nx11093)) ;
    inv02 ix11098 (.Y (nx11099), .A (nx11093)) ;
    inv02 ix11102 (.Y (nx11103), .A (nx11101)) ;
    inv02 ix11104 (.Y (nx11105), .A (nx11101)) ;
    inv02 ix11106 (.Y (nx11107), .A (nx11101)) ;
    inv02 ix11110 (.Y (nx11111), .A (nx11109)) ;
    inv02 ix11112 (.Y (nx11113), .A (nx11109)) ;
    inv02 ix11114 (.Y (nx11115), .A (nx11109)) ;
    inv04 ix11116 (.Y (nx11117), .A (gen_24_cmp_pMux_1)) ;
    inv04 ix11118 (.Y (nx11119), .A (gen_24_cmp_pMux_1)) ;
    inv04 ix11120 (.Y (nx11121), .A (gen_24_cmp_pMux_1)) ;
    inv04 ix11122 (.Y (nx11123), .A (gen_24_cmp_pMux_1)) ;
    inv02 ix11126 (.Y (nx11127), .A (nx11125)) ;
    inv02 ix11128 (.Y (nx11129), .A (nx11125)) ;
    inv02 ix11130 (.Y (nx11131), .A (nx11125)) ;
    inv02 ix11134 (.Y (nx11135), .A (nx11133)) ;
    inv02 ix11136 (.Y (nx11137), .A (nx11133)) ;
    inv02 ix11138 (.Y (nx11139), .A (nx11133)) ;
    inv02 ix11142 (.Y (nx11143), .A (nx11141)) ;
    inv02 ix11144 (.Y (nx11145), .A (nx11141)) ;
    inv02 ix11146 (.Y (nx11147), .A (nx11141)) ;
    nor02_2x ix2861 (.Y (nx10149), .A0 (nx2871), .A1 (gen_0_cmp_pMux_0)) ;
    nor02_2x ix2870 (.Y (nx10165), .A0 (gen_0_cmp_pMux_2), .A1 (nx2862)) ;
    xnor2 ix2880 (.Y (nx10173), .A0 (gen_0_cmp_pMux_0), .A1 (nx10161)) ;
    aoi21 ix2884 (.Y (nx10181), .A0 (gen_0_cmp_pMux_1), .A1 (gen_0_cmp_pMux_0), 
          .B0 (nx2871)) ;
    nor02_2x ix3106 (.Y (nx10189), .A0 (nx3115), .A1 (gen_1_cmp_pMux_0)) ;
    nor02_2x ix3114 (.Y (nx10205), .A0 (gen_1_cmp_pMux_2), .A1 (nx3107)) ;
    xnor2 ix3124 (.Y (nx10213), .A0 (gen_1_cmp_pMux_0), .A1 (nx10201)) ;
    aoi21 ix3130 (.Y (nx10221), .A0 (gen_1_cmp_pMux_1), .A1 (gen_1_cmp_pMux_0), 
          .B0 (nx3115)) ;
    nor02_2x ix3355 (.Y (nx10229), .A0 (nx3363), .A1 (gen_2_cmp_pMux_0)) ;
    nor02_2x ix3362 (.Y (nx10245), .A0 (gen_2_cmp_pMux_2), .A1 (nx3356)) ;
    xnor2 ix3372 (.Y (nx10253), .A0 (gen_2_cmp_pMux_0), .A1 (nx10241)) ;
    aoi21 ix3378 (.Y (nx10261), .A0 (gen_2_cmp_pMux_1), .A1 (gen_2_cmp_pMux_0), 
          .B0 (nx3363)) ;
    nor02_2x ix3601 (.Y (nx10269), .A0 (nx3611), .A1 (gen_3_cmp_pMux_0)) ;
    nor02_2x ix3610 (.Y (nx10285), .A0 (gen_3_cmp_pMux_2), .A1 (nx3603)) ;
    xnor2 ix3620 (.Y (nx10293), .A0 (gen_3_cmp_pMux_0), .A1 (nx10281)) ;
    aoi21 ix3626 (.Y (nx10301), .A0 (gen_3_cmp_pMux_1), .A1 (gen_3_cmp_pMux_0), 
          .B0 (nx3611)) ;
    nor02_2x ix3848 (.Y (nx10309), .A0 (nx3857), .A1 (gen_4_cmp_pMux_0)) ;
    nor02_2x ix3856 (.Y (nx10325), .A0 (gen_4_cmp_pMux_2), .A1 (nx3849)) ;
    xnor2 ix3866 (.Y (nx10333), .A0 (gen_4_cmp_pMux_0), .A1 (nx10321)) ;
    aoi21 ix3871 (.Y (nx10341), .A0 (gen_4_cmp_pMux_1), .A1 (gen_4_cmp_pMux_0), 
          .B0 (nx3857)) ;
    nor02_2x ix4092 (.Y (nx10349), .A0 (nx4101), .A1 (gen_5_cmp_pMux_0)) ;
    nor02_2x ix4100 (.Y (nx10365), .A0 (gen_5_cmp_pMux_2), .A1 (nx4093)) ;
    xnor2 ix4110 (.Y (nx10373), .A0 (gen_5_cmp_pMux_0), .A1 (nx10361)) ;
    aoi21 ix4116 (.Y (nx10381), .A0 (gen_5_cmp_pMux_1), .A1 (gen_5_cmp_pMux_0), 
          .B0 (nx4101)) ;
    nor02_2x ix4339 (.Y (nx10389), .A0 (nx4349), .A1 (gen_6_cmp_pMux_0)) ;
    nor02_2x ix4348 (.Y (nx10405), .A0 (gen_6_cmp_pMux_2), .A1 (nx4340)) ;
    xnor2 ix4358 (.Y (nx10413), .A0 (gen_6_cmp_pMux_0), .A1 (nx10401)) ;
    aoi21 ix4362 (.Y (nx10421), .A0 (gen_6_cmp_pMux_1), .A1 (gen_6_cmp_pMux_0), 
          .B0 (nx4349)) ;
    nor02_2x ix4586 (.Y (nx10429), .A0 (nx4595), .A1 (gen_7_cmp_pMux_0)) ;
    nor02_2x ix4594 (.Y (nx10445), .A0 (gen_7_cmp_pMux_2), .A1 (nx4587)) ;
    xnor2 ix4604 (.Y (nx10453), .A0 (gen_7_cmp_pMux_0), .A1 (nx10441)) ;
    aoi21 ix4610 (.Y (nx10461), .A0 (gen_7_cmp_pMux_1), .A1 (gen_7_cmp_pMux_0), 
          .B0 (nx4595)) ;
    nor02_2x ix4833 (.Y (nx10469), .A0 (nx4841), .A1 (gen_8_cmp_pMux_0)) ;
    nor02_2x ix4840 (.Y (nx10485), .A0 (gen_8_cmp_pMux_2), .A1 (nx4834)) ;
    xnor2 ix4850 (.Y (nx10493), .A0 (gen_8_cmp_pMux_0), .A1 (nx10481)) ;
    aoi21 ix4856 (.Y (nx10501), .A0 (gen_8_cmp_pMux_1), .A1 (gen_8_cmp_pMux_0), 
          .B0 (nx4841)) ;
    nor02_2x ix5076 (.Y (nx10509), .A0 (nx5085), .A1 (gen_9_cmp_pMux_0)) ;
    nor02_2x ix5084 (.Y (nx10525), .A0 (gen_9_cmp_pMux_2), .A1 (nx5077)) ;
    xnor2 ix5094 (.Y (nx10533), .A0 (gen_9_cmp_pMux_0), .A1 (nx10521)) ;
    aoi21 ix5100 (.Y (nx10541), .A0 (gen_9_cmp_pMux_1), .A1 (gen_9_cmp_pMux_0), 
          .B0 (nx5085)) ;
    nor02_2x ix5326 (.Y (nx10549), .A0 (nx5335), .A1 (gen_10_cmp_pMux_0)) ;
    nor02_2x ix5334 (.Y (nx10565), .A0 (gen_10_cmp_pMux_2), .A1 (nx5327)) ;
    xnor2 ix5344 (.Y (nx10573), .A0 (gen_10_cmp_pMux_0), .A1 (nx10561)) ;
    aoi21 ix5350 (.Y (nx10581), .A0 (gen_10_cmp_pMux_1), .A1 (gen_10_cmp_pMux_0)
          , .B0 (nx5335)) ;
    nor02_2x ix5575 (.Y (nx10589), .A0 (nx5585), .A1 (gen_11_cmp_pMux_0)) ;
    nor02_2x ix5584 (.Y (nx10605), .A0 (gen_11_cmp_pMux_2), .A1 (nx5577)) ;
    xnor2 ix5594 (.Y (nx10613), .A0 (gen_11_cmp_pMux_0), .A1 (nx10601)) ;
    aoi21 ix5600 (.Y (nx10621), .A0 (gen_11_cmp_pMux_1), .A1 (gen_11_cmp_pMux_0)
          , .B0 (nx5585)) ;
    nor02_2x ix5820 (.Y (nx10629), .A0 (nx5829), .A1 (gen_12_cmp_pMux_0)) ;
    nor02_2x ix5828 (.Y (nx10645), .A0 (gen_12_cmp_pMux_2), .A1 (nx5821)) ;
    xnor2 ix5838 (.Y (nx10653), .A0 (gen_12_cmp_pMux_0), .A1 (nx10641)) ;
    aoi21 ix5844 (.Y (nx10661), .A0 (gen_12_cmp_pMux_1), .A1 (gen_12_cmp_pMux_0)
          , .B0 (nx5829)) ;
    nor02_2x ix6066 (.Y (nx10669), .A0 (nx6075), .A1 (gen_13_cmp_pMux_0)) ;
    nor02_2x ix6074 (.Y (nx10685), .A0 (gen_13_cmp_pMux_2), .A1 (nx6067)) ;
    xnor2 ix6084 (.Y (nx10693), .A0 (gen_13_cmp_pMux_0), .A1 (nx10681)) ;
    aoi21 ix6090 (.Y (nx10701), .A0 (gen_13_cmp_pMux_1), .A1 (gen_13_cmp_pMux_0)
          , .B0 (nx6075)) ;
    nor02_2x ix6313 (.Y (nx10709), .A0 (nx6323), .A1 (gen_14_cmp_pMux_0)) ;
    nor02_2x ix6322 (.Y (nx10725), .A0 (gen_14_cmp_pMux_2), .A1 (nx6314)) ;
    xnor2 ix6332 (.Y (nx10733), .A0 (gen_14_cmp_pMux_0), .A1 (nx10721)) ;
    aoi21 ix6336 (.Y (nx10741), .A0 (gen_14_cmp_pMux_1), .A1 (gen_14_cmp_pMux_0)
          , .B0 (nx6323)) ;
    nor02_2x ix6560 (.Y (nx10749), .A0 (nx6569), .A1 (gen_15_cmp_pMux_0)) ;
    nor02_2x ix6568 (.Y (nx10765), .A0 (gen_15_cmp_pMux_2), .A1 (nx6561)) ;
    xnor2 ix6577 (.Y (nx10773), .A0 (gen_15_cmp_pMux_0), .A1 (nx10761)) ;
    aoi21 ix6582 (.Y (nx10781), .A0 (gen_15_cmp_pMux_1), .A1 (gen_15_cmp_pMux_0)
          , .B0 (nx6569)) ;
    nor02_2x ix6807 (.Y (nx10789), .A0 (nx6815), .A1 (gen_16_cmp_pMux_0)) ;
    nor02_2x ix6814 (.Y (nx10805), .A0 (gen_16_cmp_pMux_2), .A1 (nx6808)) ;
    xnor2 ix6824 (.Y (nx10813), .A0 (gen_16_cmp_pMux_0), .A1 (nx10801)) ;
    aoi21 ix6830 (.Y (nx10821), .A0 (gen_16_cmp_pMux_1), .A1 (gen_16_cmp_pMux_0)
          , .B0 (nx6815)) ;
    nor02_2x ix7048 (.Y (nx10829), .A0 (nx7057), .A1 (gen_17_cmp_pMux_0)) ;
    nor02_2x ix7056 (.Y (nx10845), .A0 (gen_17_cmp_pMux_2), .A1 (nx7049)) ;
    xnor2 ix7066 (.Y (nx10853), .A0 (gen_17_cmp_pMux_0), .A1 (nx10841)) ;
    aoi21 ix7072 (.Y (nx10861), .A0 (gen_17_cmp_pMux_1), .A1 (gen_17_cmp_pMux_0)
          , .B0 (nx7057)) ;
    nor02_2x ix7295 (.Y (nx10869), .A0 (nx7305), .A1 (gen_18_cmp_pMux_0)) ;
    nor02_2x ix7304 (.Y (nx10885), .A0 (gen_18_cmp_pMux_2), .A1 (nx7297)) ;
    xnor2 ix7314 (.Y (nx10893), .A0 (gen_18_cmp_pMux_0), .A1 (nx10881)) ;
    aoi21 ix7320 (.Y (nx10901), .A0 (gen_18_cmp_pMux_1), .A1 (gen_18_cmp_pMux_0)
          , .B0 (nx7305)) ;
    nor02_2x ix7544 (.Y (nx10909), .A0 (nx7553), .A1 (gen_19_cmp_pMux_0)) ;
    nor02_2x ix7552 (.Y (nx10925), .A0 (gen_19_cmp_pMux_2), .A1 (nx7545)) ;
    xnor2 ix7562 (.Y (nx10933), .A0 (gen_19_cmp_pMux_0), .A1 (nx10921)) ;
    aoi21 ix7568 (.Y (nx10941), .A0 (gen_19_cmp_pMux_1), .A1 (gen_19_cmp_pMux_0)
          , .B0 (nx7553)) ;
    nor02_2x ix7791 (.Y (nx10949), .A0 (nx7801), .A1 (gen_20_cmp_pMux_0)) ;
    nor02_2x ix7800 (.Y (nx10965), .A0 (gen_20_cmp_pMux_2), .A1 (nx7792)) ;
    xnor2 ix7810 (.Y (nx10973), .A0 (gen_20_cmp_pMux_0), .A1 (nx10961)) ;
    aoi21 ix7814 (.Y (nx10981), .A0 (gen_20_cmp_pMux_1), .A1 (gen_20_cmp_pMux_0)
          , .B0 (nx7801)) ;
    nor02_2x ix8038 (.Y (nx10989), .A0 (nx8047), .A1 (gen_21_cmp_pMux_0)) ;
    nor02_2x ix8046 (.Y (nx11005), .A0 (gen_21_cmp_pMux_2), .A1 (nx8039)) ;
    xnor2 ix8056 (.Y (nx11013), .A0 (gen_21_cmp_pMux_0), .A1 (nx11001)) ;
    aoi21 ix8062 (.Y (nx11021), .A0 (gen_21_cmp_pMux_1), .A1 (gen_21_cmp_pMux_0)
          , .B0 (nx8047)) ;
    nor02_2x ix8282 (.Y (nx11029), .A0 (nx8291), .A1 (gen_22_cmp_pMux_0)) ;
    nor02_2x ix8290 (.Y (nx11045), .A0 (gen_22_cmp_pMux_2), .A1 (nx8283)) ;
    xnor2 ix8300 (.Y (nx11053), .A0 (gen_22_cmp_pMux_0), .A1 (nx11041)) ;
    aoi21 ix8306 (.Y (nx11061), .A0 (gen_22_cmp_pMux_1), .A1 (gen_22_cmp_pMux_0)
          , .B0 (nx8291)) ;
    nor02_2x ix8532 (.Y (nx11069), .A0 (nx8541), .A1 (gen_23_cmp_pMux_0)) ;
    nor02_2x ix8540 (.Y (nx11085), .A0 (gen_23_cmp_pMux_2), .A1 (nx8533)) ;
    xnor2 ix8550 (.Y (nx11093), .A0 (gen_23_cmp_pMux_0), .A1 (nx11081)) ;
    aoi21 ix8556 (.Y (nx11101), .A0 (gen_23_cmp_pMux_1), .A1 (gen_23_cmp_pMux_0)
          , .B0 (nx8541)) ;
    nor02_2x ix8778 (.Y (nx11109), .A0 (nx8787), .A1 (gen_24_cmp_pMux_0)) ;
    nor02_2x ix8786 (.Y (nx11125), .A0 (gen_24_cmp_pMux_2), .A1 (nx8779)) ;
    xnor2 ix8796 (.Y (nx11133), .A0 (gen_24_cmp_pMux_0), .A1 (nx11121)) ;
    aoi21 ix8802 (.Y (nx11141), .A0 (gen_24_cmp_pMux_1), .A1 (gen_24_cmp_pMux_0)
          , .B0 (nx8787)) ;
    nand02 ix9687 (.Y (nx9373), .A0 (nx11157), .A1 (nx9365)) ;
    inv01 ix11156 (.Y (nx11157), .A (nx9353)) ;
    mux21 ix2824 (.Y (nx2823), .A0 (nx9361), .A1 (nx9357), .S0 (nx11201)) ;
    mux21 ix2814 (.Y (nx2813), .A0 (nx11197), .A1 (nx9361), .S0 (nx11201)) ;
    inv02 ix11158 (.Y (nx11159), .A (nx11201)) ;
    inv02 ix11160 (.Y (nx11161), .A (nx11201)) ;
    inv02 ix11162 (.Y (nx11163), .A (nx11203)) ;
    inv02 ix11164 (.Y (nx11165), .A (nx11203)) ;
    inv02 ix11166 (.Y (nx11167), .A (nx11203)) ;
    inv02 ix11168 (.Y (nx11169), .A (nx11203)) ;
    inv02 ix11170 (.Y (nx11171), .A (nx11203)) ;
    inv02 ix11172 (.Y (nx11173), .A (nx11197)) ;
    inv02 ix11174 (.Y (nx11175), .A (nx11197)) ;
    inv02 ix11176 (.Y (nx11177), .A (nx11197)) ;
    inv02 ix11178 (.Y (nx11179), .A (nx11197)) ;
    inv02 ix11180 (.Y (nx11181), .A (nx11197)) ;
    inv02 ix11182 (.Y (nx11183), .A (nx11199)) ;
    inv02 ix11184 (.Y (nx11185), .A (nx11199)) ;
    inv02 ix11186 (.Y (nx11187), .A (nx11199)) ;
    inv02 ix11188 (.Y (nx11189), .A (nx11199)) ;
    inv01 ix11190 (.Y (nx11191), .A (nx11199)) ;
    inv02 ix11196 (.Y (nx11197), .A (nx9389)) ;
    inv02 ix11198 (.Y (nx11199), .A (nx9389)) ;
    inv02 ix11200 (.Y (nx11201), .A (nx9375)) ;
    inv02 ix11202 (.Y (nx11203), .A (nx9375)) ;
endmodule


module NBitAdder_24 ( a, b, carryIn, sum, carryOut ) ;

    input [23:0]a ;
    input [23:0]b ;
    input carryIn ;
    output [23:0]sum ;
    output carryOut ;

    wire nx6, nx8, nx16, nx18, nx22, nx24, nx30, nx32, nx38, nx40, nx46, nx48, 
         nx54, nx56, nx62, nx64, nx70, nx72, nx78, nx80, nx86, nx88, nx94, nx96, 
         nx102, nx104, nx110, nx112, nx118, nx120, nx126, nx128, nx134, nx136, 
         nx142, nx144, nx150, nx152, nx158, nx160, nx166, nx168, nx170, nx172, 
         nx103, nx109, nx111, nx113, nx115, nx119, nx123, nx127, nx133, nx135, 
         nx137, nx141, nx145, nx149, nx155, nx157, nx159, nx163, nx167, nx171, 
         nx177, nx179, nx181, nx185, nx189, nx193, nx199, nx201, nx203, nx207, 
         nx211, nx215, nx221, nx223, nx225, nx229, nx232, nx235, nx239, nx241, 
         nx243, nx246, nx249, nx252, nx256, nx258, nx260, nx263, nx266, nx269, 
         nx273, nx275, nx277, nx280, nx283, nx286, nx290, nx292, nx294, nx297, 
         nx300, nx303, nx307, nx309, nx311, nx314, nx317, nx320, nx323, nx326, 
         nx329, nx332, nx335, nx338, nx341, nx344, nx347, nx350, nx353, nx356, 
         nx358, nx360, nx362, nx364, nx366, nx368, nx370, nx372;



    fake_gnd ix44 (.Y (carryOut)) ;
    xnor2 ix229 (.Y (sum[0]), .A0 (carryIn), .A1 (nx103)) ;
    xnor2 ix104 (.Y (nx103), .A0 (a[0]), .A1 (b[0])) ;
    xnor2 ix227 (.Y (sum[1]), .A0 (nx6), .A1 (nx115)) ;
    oai22 ix7 (.Y (nx6), .A0 (nx109), .A1 (nx103), .B0 (nx111), .B1 (nx113)) ;
    inv01 ix110 (.Y (nx109), .A (carryIn)) ;
    inv01 ix112 (.Y (nx111), .A (b[0])) ;
    inv01 ix114 (.Y (nx113), .A (a[0])) ;
    xnor2 ix116 (.Y (nx115), .A0 (a[1]), .A1 (b[1])) ;
    xnor2 ix225 (.Y (sum[2]), .A0 (nx119), .A1 (nx16)) ;
    aoi22 ix120 (.Y (nx119), .A0 (b[1]), .A1 (a[1]), .B0 (nx6), .B1 (nx8)) ;
    xnor2 ix9 (.Y (nx8), .A0 (a[1]), .A1 (nx123)) ;
    inv01 ix124 (.Y (nx123), .A (b[1])) ;
    xnor2 ix17 (.Y (nx16), .A0 (a[2]), .A1 (nx127)) ;
    inv01 ix128 (.Y (nx127), .A (b[2])) ;
    xnor2 ix223 (.Y (sum[3]), .A0 (nx22), .A1 (nx137)) ;
    oai21 ix23 (.Y (nx22), .A0 (nx119), .A1 (nx133), .B0 (nx135)) ;
    xnor2 ix134 (.Y (nx133), .A0 (a[2]), .A1 (b[2])) ;
    nand02 ix136 (.Y (nx135), .A0 (b[2]), .A1 (a[2])) ;
    xnor2 ix138 (.Y (nx137), .A0 (a[3]), .A1 (b[3])) ;
    xnor2 ix221 (.Y (sum[4]), .A0 (nx141), .A1 (nx32)) ;
    aoi22 ix142 (.Y (nx141), .A0 (b[3]), .A1 (a[3]), .B0 (nx22), .B1 (nx24)) ;
    xnor2 ix25 (.Y (nx24), .A0 (a[3]), .A1 (nx145)) ;
    inv01 ix146 (.Y (nx145), .A (b[3])) ;
    xnor2 ix33 (.Y (nx32), .A0 (a[4]), .A1 (nx149)) ;
    inv01 ix150 (.Y (nx149), .A (b[4])) ;
    xnor2 ix219 (.Y (sum[5]), .A0 (nx38), .A1 (nx159)) ;
    oai21 ix39 (.Y (nx38), .A0 (nx141), .A1 (nx155), .B0 (nx157)) ;
    xnor2 ix156 (.Y (nx155), .A0 (a[4]), .A1 (b[4])) ;
    nand02 ix158 (.Y (nx157), .A0 (b[4]), .A1 (a[4])) ;
    xnor2 ix160 (.Y (nx159), .A0 (a[5]), .A1 (b[5])) ;
    xnor2 ix217 (.Y (sum[6]), .A0 (nx163), .A1 (nx48)) ;
    aoi22 ix164 (.Y (nx163), .A0 (b[5]), .A1 (a[5]), .B0 (nx38), .B1 (nx40)) ;
    xnor2 ix41 (.Y (nx40), .A0 (a[5]), .A1 (nx167)) ;
    inv01 ix168 (.Y (nx167), .A (b[5])) ;
    xnor2 ix49 (.Y (nx48), .A0 (a[6]), .A1 (nx171)) ;
    inv01 ix172 (.Y (nx171), .A (b[6])) ;
    xnor2 ix215 (.Y (sum[7]), .A0 (nx54), .A1 (nx181)) ;
    oai21 ix55 (.Y (nx54), .A0 (nx163), .A1 (nx177), .B0 (nx179)) ;
    xnor2 ix178 (.Y (nx177), .A0 (a[6]), .A1 (b[6])) ;
    nand02 ix180 (.Y (nx179), .A0 (b[6]), .A1 (a[6])) ;
    xnor2 ix182 (.Y (nx181), .A0 (a[7]), .A1 (b[7])) ;
    xnor2 ix213 (.Y (sum[8]), .A0 (nx185), .A1 (nx64)) ;
    aoi22 ix186 (.Y (nx185), .A0 (b[7]), .A1 (a[7]), .B0 (nx54), .B1 (nx56)) ;
    xnor2 ix57 (.Y (nx56), .A0 (a[7]), .A1 (nx189)) ;
    inv01 ix190 (.Y (nx189), .A (b[7])) ;
    xnor2 ix65 (.Y (nx64), .A0 (a[8]), .A1 (nx193)) ;
    inv01 ix194 (.Y (nx193), .A (b[8])) ;
    xnor2 ix211 (.Y (sum[9]), .A0 (nx70), .A1 (nx203)) ;
    oai21 ix71 (.Y (nx70), .A0 (nx185), .A1 (nx199), .B0 (nx201)) ;
    xnor2 ix200 (.Y (nx199), .A0 (a[8]), .A1 (b[8])) ;
    nand02 ix202 (.Y (nx201), .A0 (b[8]), .A1 (a[8])) ;
    xnor2 ix204 (.Y (nx203), .A0 (a[9]), .A1 (b[9])) ;
    xnor2 ix209 (.Y (sum[10]), .A0 (nx207), .A1 (nx80)) ;
    aoi22 ix208 (.Y (nx207), .A0 (b[9]), .A1 (a[9]), .B0 (nx70), .B1 (nx72)) ;
    xnor2 ix73 (.Y (nx72), .A0 (a[9]), .A1 (nx211)) ;
    inv01 ix212 (.Y (nx211), .A (b[9])) ;
    xnor2 ix81 (.Y (nx80), .A0 (a[10]), .A1 (nx215)) ;
    inv01 ix216 (.Y (nx215), .A (b[10])) ;
    xnor2 ix207 (.Y (sum[11]), .A0 (nx86), .A1 (nx225)) ;
    oai21 ix87 (.Y (nx86), .A0 (nx207), .A1 (nx221), .B0 (nx223)) ;
    xnor2 ix222 (.Y (nx221), .A0 (a[10]), .A1 (b[10])) ;
    nand02 ix224 (.Y (nx223), .A0 (b[10]), .A1 (a[10])) ;
    xnor2 ix226 (.Y (nx225), .A0 (a[11]), .A1 (b[11])) ;
    xnor2 ix205 (.Y (sum[12]), .A0 (nx229), .A1 (nx96)) ;
    aoi22 ix230 (.Y (nx229), .A0 (b[11]), .A1 (a[11]), .B0 (nx86), .B1 (nx88)) ;
    xnor2 ix89 (.Y (nx88), .A0 (a[11]), .A1 (nx232)) ;
    inv01 ix233 (.Y (nx232), .A (b[11])) ;
    xnor2 ix97 (.Y (nx96), .A0 (a[12]), .A1 (nx235)) ;
    inv01 ix236 (.Y (nx235), .A (b[12])) ;
    xnor2 ix203 (.Y (sum[13]), .A0 (nx102), .A1 (nx243)) ;
    oai21 ix103 (.Y (nx102), .A0 (nx229), .A1 (nx239), .B0 (nx241)) ;
    xnor2 ix240 (.Y (nx239), .A0 (a[12]), .A1 (b[12])) ;
    nand02 ix242 (.Y (nx241), .A0 (b[12]), .A1 (a[12])) ;
    xnor2 ix244 (.Y (nx243), .A0 (a[13]), .A1 (b[13])) ;
    xnor2 ix201 (.Y (sum[14]), .A0 (nx246), .A1 (nx112)) ;
    aoi22 ix247 (.Y (nx246), .A0 (b[13]), .A1 (a[13]), .B0 (nx102), .B1 (nx104)
          ) ;
    xnor2 ix105 (.Y (nx104), .A0 (a[13]), .A1 (nx249)) ;
    inv01 ix250 (.Y (nx249), .A (b[13])) ;
    xnor2 ix113 (.Y (nx112), .A0 (a[14]), .A1 (nx252)) ;
    inv01 ix253 (.Y (nx252), .A (b[14])) ;
    xnor2 ix199 (.Y (sum[15]), .A0 (nx118), .A1 (nx260)) ;
    oai21 ix119 (.Y (nx118), .A0 (nx246), .A1 (nx256), .B0 (nx258)) ;
    xnor2 ix257 (.Y (nx256), .A0 (a[14]), .A1 (b[14])) ;
    nand02 ix259 (.Y (nx258), .A0 (b[14]), .A1 (a[14])) ;
    xnor2 ix261 (.Y (nx260), .A0 (a[15]), .A1 (b[15])) ;
    xnor2 ix197 (.Y (sum[16]), .A0 (nx263), .A1 (nx128)) ;
    aoi22 ix264 (.Y (nx263), .A0 (b[15]), .A1 (a[15]), .B0 (nx118), .B1 (nx120)
          ) ;
    xnor2 ix121 (.Y (nx120), .A0 (a[15]), .A1 (nx266)) ;
    inv01 ix267 (.Y (nx266), .A (b[15])) ;
    xnor2 ix129 (.Y (nx128), .A0 (a[16]), .A1 (nx269)) ;
    inv01 ix270 (.Y (nx269), .A (b[16])) ;
    xnor2 ix195 (.Y (sum[17]), .A0 (nx134), .A1 (nx277)) ;
    oai21 ix135 (.Y (nx134), .A0 (nx263), .A1 (nx273), .B0 (nx275)) ;
    xnor2 ix274 (.Y (nx273), .A0 (a[16]), .A1 (b[16])) ;
    nand02 ix276 (.Y (nx275), .A0 (b[16]), .A1 (a[16])) ;
    xnor2 ix278 (.Y (nx277), .A0 (a[17]), .A1 (b[17])) ;
    xnor2 ix193 (.Y (sum[18]), .A0 (nx280), .A1 (nx144)) ;
    aoi22 ix281 (.Y (nx280), .A0 (b[17]), .A1 (a[17]), .B0 (nx134), .B1 (nx136)
          ) ;
    xnor2 ix137 (.Y (nx136), .A0 (a[17]), .A1 (nx283)) ;
    inv01 ix284 (.Y (nx283), .A (b[17])) ;
    xnor2 ix145 (.Y (nx144), .A0 (a[18]), .A1 (nx286)) ;
    inv01 ix287 (.Y (nx286), .A (b[18])) ;
    xnor2 ix191 (.Y (sum[19]), .A0 (nx150), .A1 (nx294)) ;
    oai21 ix151 (.Y (nx150), .A0 (nx280), .A1 (nx290), .B0 (nx292)) ;
    xnor2 ix291 (.Y (nx290), .A0 (a[18]), .A1 (b[18])) ;
    nand02 ix293 (.Y (nx292), .A0 (b[18]), .A1 (a[18])) ;
    xnor2 ix295 (.Y (nx294), .A0 (a[19]), .A1 (b[19])) ;
    xnor2 ix189 (.Y (sum[20]), .A0 (nx297), .A1 (nx160)) ;
    aoi22 ix298 (.Y (nx297), .A0 (b[19]), .A1 (a[19]), .B0 (nx150), .B1 (nx152)
          ) ;
    xnor2 ix153 (.Y (nx152), .A0 (a[19]), .A1 (nx300)) ;
    inv01 ix301 (.Y (nx300), .A (b[19])) ;
    xnor2 ix161 (.Y (nx160), .A0 (a[20]), .A1 (nx303)) ;
    inv01 ix304 (.Y (nx303), .A (b[20])) ;
    xnor2 ix187 (.Y (sum[21]), .A0 (nx166), .A1 (nx311)) ;
    oai21 ix167 (.Y (nx166), .A0 (nx297), .A1 (nx307), .B0 (nx309)) ;
    xnor2 ix308 (.Y (nx307), .A0 (a[20]), .A1 (b[20])) ;
    nand02 ix310 (.Y (nx309), .A0 (b[20]), .A1 (a[20])) ;
    xnor2 ix312 (.Y (nx311), .A0 (a[21]), .A1 (b[21])) ;
    xnor2 ix185 (.Y (sum[22]), .A0 (b[22]), .A1 (nx314)) ;
    aoi22 ix315 (.Y (nx314), .A0 (b[21]), .A1 (a[21]), .B0 (nx166), .B1 (nx168)
          ) ;
    xnor2 ix169 (.Y (nx168), .A0 (a[21]), .A1 (nx317)) ;
    inv01 ix318 (.Y (nx317), .A (b[21])) ;
    xnor2 ix179 (.Y (sum[23]), .A0 (b[23]), .A1 (nx320)) ;
    oai21 ix321 (.Y (nx320), .A0 (nx172), .A1 (nx170), .B0 (b[22])) ;
    nor02_2x ix173 (.Y (nx172), .A0 (nx317), .A1 (nx323)) ;
    inv01 ix324 (.Y (nx323), .A (a[21])) ;
    nor02ii ix171 (.Y (nx170), .A0 (nx326), .A1 (nx168)) ;
    aoi22 ix327 (.Y (nx326), .A0 (b[20]), .A1 (a[20]), .B0 (nx158), .B1 (nx160)
          ) ;
    oai21 ix159 (.Y (nx158), .A0 (nx329), .A1 (nx294), .B0 (nx372)) ;
    aoi22 ix330 (.Y (nx329), .A0 (b[18]), .A1 (a[18]), .B0 (nx142), .B1 (nx144)
          ) ;
    oai21 ix143 (.Y (nx142), .A0 (nx332), .A1 (nx277), .B0 (nx370)) ;
    aoi22 ix333 (.Y (nx332), .A0 (b[16]), .A1 (a[16]), .B0 (nx126), .B1 (nx128)
          ) ;
    oai21 ix127 (.Y (nx126), .A0 (nx335), .A1 (nx260), .B0 (nx368)) ;
    aoi22 ix336 (.Y (nx335), .A0 (b[14]), .A1 (a[14]), .B0 (nx110), .B1 (nx112)
          ) ;
    oai21 ix111 (.Y (nx110), .A0 (nx338), .A1 (nx243), .B0 (nx366)) ;
    aoi22 ix339 (.Y (nx338), .A0 (b[12]), .A1 (a[12]), .B0 (nx94), .B1 (nx96)) ;
    oai21 ix95 (.Y (nx94), .A0 (nx341), .A1 (nx225), .B0 (nx364)) ;
    aoi22 ix342 (.Y (nx341), .A0 (b[10]), .A1 (a[10]), .B0 (nx78), .B1 (nx80)) ;
    oai21 ix79 (.Y (nx78), .A0 (nx344), .A1 (nx203), .B0 (nx362)) ;
    aoi22 ix345 (.Y (nx344), .A0 (b[8]), .A1 (a[8]), .B0 (nx62), .B1 (nx64)) ;
    oai21 ix63 (.Y (nx62), .A0 (nx347), .A1 (nx181), .B0 (nx360)) ;
    aoi22 ix348 (.Y (nx347), .A0 (b[6]), .A1 (a[6]), .B0 (nx46), .B1 (nx48)) ;
    oai21 ix47 (.Y (nx46), .A0 (nx350), .A1 (nx159), .B0 (nx358)) ;
    aoi22 ix351 (.Y (nx350), .A0 (b[4]), .A1 (a[4]), .B0 (nx30), .B1 (nx32)) ;
    oai21 ix31 (.Y (nx30), .A0 (nx353), .A1 (nx137), .B0 (nx356)) ;
    aoi21 ix354 (.Y (nx353), .A0 (b[2]), .A1 (a[2]), .B0 (nx18)) ;
    nor02ii ix19 (.Y (nx18), .A0 (nx119), .A1 (nx16)) ;
    nand02 ix357 (.Y (nx356), .A0 (b[3]), .A1 (a[3])) ;
    nand02 ix359 (.Y (nx358), .A0 (b[5]), .A1 (a[5])) ;
    nand02 ix361 (.Y (nx360), .A0 (b[7]), .A1 (a[7])) ;
    nand02 ix363 (.Y (nx362), .A0 (b[9]), .A1 (a[9])) ;
    nand02 ix365 (.Y (nx364), .A0 (b[11]), .A1 (a[11])) ;
    nand02 ix367 (.Y (nx366), .A0 (b[13]), .A1 (a[13])) ;
    nand02 ix369 (.Y (nx368), .A0 (b[15]), .A1 (a[15])) ;
    nand02 ix371 (.Y (nx370), .A0 (b[17]), .A1 (a[17])) ;
    nand02 ix373 (.Y (nx372), .A0 (b[19]), .A1 (a[19])) ;
endmodule


module BinaryMux_33 ( a, b, sel, f ) ;

    input [32:0]a ;
    input [32:0]b ;
    input sel ;
    output [32:0]f ;

    wire nx93, nx97, nx99, nx105, nx107, nx111, nx113, nx117, nx119, nx123, 
         nx125, nx129, nx131, nx135, nx137, nx141, nx143, nx147, nx151, nx155, 
         nx158, nx161, nx164, nx167, nx170, nx173, nx176, nx179, nx182, nx185, 
         nx188, nx191, nx194, nx197, nx200, nx203, nx206, nx209, nx212, nx219, 
         nx221, nx223, nx225, nx227, nx229, nx231;



    assign f[31] = f[32] ;
    fake_gnd ix44 (.Y (f[32])) ;
    nor02_2x ix3 (.Y (f[0]), .A0 (nx93), .A1 (nx219)) ;
    inv01 ix94 (.Y (nx93), .A (a[0])) ;
    nand02_2x ix99 (.Y (f[1]), .A0 (nx97), .A1 (nx99)) ;
    nand02 ix98 (.Y (nx97), .A0 (b[1]), .A1 (nx219)) ;
    nand02 ix100 (.Y (nx99), .A0 (a[1]), .A1 (nx229)) ;
    nand02 ix107 (.Y (f[2]), .A0 (nx105), .A1 (nx107)) ;
    nand02 ix106 (.Y (nx105), .A0 (b[2]), .A1 (nx219)) ;
    nand02 ix108 (.Y (nx107), .A0 (a[2]), .A1 (nx229)) ;
    nand02 ix115 (.Y (f[3]), .A0 (nx111), .A1 (nx113)) ;
    nand02 ix112 (.Y (nx111), .A0 (b[3]), .A1 (nx219)) ;
    nand02 ix114 (.Y (nx113), .A0 (a[3]), .A1 (nx229)) ;
    nand02 ix123 (.Y (f[4]), .A0 (nx117), .A1 (nx119)) ;
    nand02 ix118 (.Y (nx117), .A0 (b[4]), .A1 (nx219)) ;
    nand02 ix120 (.Y (nx119), .A0 (a[4]), .A1 (nx229)) ;
    nand02 ix131 (.Y (f[5]), .A0 (nx123), .A1 (nx125)) ;
    nand02 ix124 (.Y (nx123), .A0 (b[5]), .A1 (nx219)) ;
    nand02 ix126 (.Y (nx125), .A0 (a[5]), .A1 (nx229)) ;
    nand02 ix139 (.Y (f[6]), .A0 (nx129), .A1 (nx131)) ;
    nand02 ix130 (.Y (nx129), .A0 (b[6]), .A1 (nx219)) ;
    nand02 ix132 (.Y (nx131), .A0 (a[6]), .A1 (nx229)) ;
    nand02 ix147 (.Y (f[7]), .A0 (nx135), .A1 (nx137)) ;
    nand02 ix136 (.Y (nx135), .A0 (b[7]), .A1 (nx221)) ;
    nand02 ix138 (.Y (nx137), .A0 (a[7]), .A1 (nx229)) ;
    nand02 ix155 (.Y (f[8]), .A0 (nx141), .A1 (nx143)) ;
    nand02 ix142 (.Y (nx141), .A0 (nx221), .A1 (b[8])) ;
    nand02 ix144 (.Y (nx143), .A0 (nx231), .A1 (a[8])) ;
    nor02_2x ix7 (.Y (f[9]), .A0 (nx147), .A1 (nx221)) ;
    inv01 ix148 (.Y (nx147), .A (a[9])) ;
    nor02_2x ix11 (.Y (f[10]), .A0 (nx151), .A1 (nx221)) ;
    inv01 ix152 (.Y (nx151), .A (a[10])) ;
    nor02_2x ix15 (.Y (f[11]), .A0 (nx155), .A1 (nx221)) ;
    inv01 ix156 (.Y (nx155), .A (a[11])) ;
    nor02_2x ix19 (.Y (f[12]), .A0 (nx158), .A1 (nx221)) ;
    inv01 ix159 (.Y (nx158), .A (a[12])) ;
    nor02_2x ix23 (.Y (f[13]), .A0 (nx161), .A1 (nx221)) ;
    inv01 ix162 (.Y (nx161), .A (a[13])) ;
    nor02_2x ix27 (.Y (f[14]), .A0 (nx164), .A1 (nx223)) ;
    inv01 ix165 (.Y (nx164), .A (a[14])) ;
    nor02_2x ix31 (.Y (f[15]), .A0 (nx167), .A1 (nx223)) ;
    inv01 ix168 (.Y (nx167), .A (a[15])) ;
    nor02_2x ix35 (.Y (f[16]), .A0 (nx170), .A1 (nx223)) ;
    inv01 ix171 (.Y (nx170), .A (a[16])) ;
    nor02_2x ix39 (.Y (f[17]), .A0 (nx173), .A1 (nx223)) ;
    inv01 ix174 (.Y (nx173), .A (a[17])) ;
    nor02_2x ix43 (.Y (f[18]), .A0 (nx176), .A1 (nx223)) ;
    inv01 ix177 (.Y (nx176), .A (a[18])) ;
    nor02_2x ix47 (.Y (f[19]), .A0 (nx179), .A1 (nx223)) ;
    inv01 ix180 (.Y (nx179), .A (a[19])) ;
    nor02_2x ix51 (.Y (f[20]), .A0 (nx182), .A1 (nx223)) ;
    inv01 ix183 (.Y (nx182), .A (a[20])) ;
    nor02_2x ix55 (.Y (f[21]), .A0 (nx185), .A1 (nx225)) ;
    inv01 ix186 (.Y (nx185), .A (a[21])) ;
    nor02_2x ix59 (.Y (f[22]), .A0 (nx188), .A1 (nx225)) ;
    inv01 ix189 (.Y (nx188), .A (a[22])) ;
    nor02_2x ix63 (.Y (f[23]), .A0 (nx191), .A1 (nx225)) ;
    inv01 ix192 (.Y (nx191), .A (a[23])) ;
    nor02_2x ix67 (.Y (f[24]), .A0 (nx194), .A1 (nx225)) ;
    inv01 ix195 (.Y (nx194), .A (a[24])) ;
    nor02_2x ix71 (.Y (f[25]), .A0 (nx197), .A1 (nx225)) ;
    inv01 ix198 (.Y (nx197), .A (a[25])) ;
    nor02_2x ix75 (.Y (f[26]), .A0 (nx200), .A1 (nx225)) ;
    inv01 ix201 (.Y (nx200), .A (a[26])) ;
    nor02_2x ix79 (.Y (f[27]), .A0 (nx203), .A1 (nx225)) ;
    inv01 ix204 (.Y (nx203), .A (a[27])) ;
    nor02_2x ix83 (.Y (f[28]), .A0 (nx206), .A1 (nx227)) ;
    inv01 ix207 (.Y (nx206), .A (a[28])) ;
    nor02_2x ix87 (.Y (f[29]), .A0 (nx209), .A1 (nx227)) ;
    inv01 ix210 (.Y (nx209), .A (a[29])) ;
    nor02_2x ix91 (.Y (f[30]), .A0 (nx212), .A1 (nx227)) ;
    inv01 ix213 (.Y (nx212), .A (a[30])) ;
    inv02 ix218 (.Y (nx219), .A (nx231)) ;
    inv02 ix220 (.Y (nx221), .A (nx231)) ;
    inv02 ix222 (.Y (nx223), .A (nx231)) ;
    inv02 ix224 (.Y (nx225), .A (nx231)) ;
    inv02 ix226 (.Y (nx227), .A (nx231)) ;
    inv02 ix228 (.Y (nx229), .A (sel)) ;
    inv02 ix230 (.Y (nx231), .A (sel)) ;
endmodule


module Reg_33 ( D, en, clk, rst, Q ) ;

    input [32:0]D ;
    input en ;
    input clk ;
    input rst ;
    output [32:0]Q ;

    wire nx115, nx125, nx135, nx145, nx155, nx165, nx175, nx185, nx195, nx205, 
         nx215, nx225, nx235, nx245, nx255, nx265, nx275, nx285, nx295, nx305, 
         nx315, nx325, nx335, nx345, nx355, nx365, nx375, nx385, nx395, nx405, 
         nx415, nx427, nx431, nx436, nx438, nx443, nx445, nx450, nx452, nx457, 
         nx459, nx464, nx466, nx471, nx473, nx478, nx480, nx485, nx487, nx492, 
         nx494, nx499, nx501, nx506, nx508, nx513, nx515, nx520, nx522, nx527, 
         nx529, nx534, nx536, nx541, nx543, nx548, nx550, nx555, nx557, nx562, 
         nx564, nx569, nx571, nx576, nx578, nx583, nx585, nx590, nx592, nx597, 
         nx599, nx604, nx606, nx611, nx613, nx618, nx620, nx625, nx627, nx632, 
         nx634, nx639, nx641, nx649, nx651, nx653, nx655, nx657, nx663, nx665, 
         nx667, nx669, nx671, nx673, nx675, nx677, nx679, nx681, nx683, nx685;
    wire [30:0] \$dummy ;




    assign Q[31] = Q[32] ;
    fake_gnd ix43 (.Y (Q[32])) ;
    dffr reg_Q_0 (.Q (Q[0]), .QB (\$dummy [0]), .D (nx115), .CLK (nx675), .R (
         rst)) ;
    nand02 ix116 (.Y (nx115), .A0 (nx427), .A1 (nx431)) ;
    nand02 ix428 (.Y (nx427), .A0 (Q[0]), .A1 (nx685)) ;
    nand02 ix432 (.Y (nx431), .A0 (D[0]), .A1 (nx663)) ;
    dffr reg_Q_1 (.Q (Q[1]), .QB (\$dummy [1]), .D (nx125), .CLK (nx675), .R (
         rst)) ;
    nand02 ix126 (.Y (nx125), .A0 (nx436), .A1 (nx438)) ;
    nand02 ix437 (.Y (nx436), .A0 (Q[1]), .A1 (nx685)) ;
    nand02 ix439 (.Y (nx438), .A0 (D[1]), .A1 (nx663)) ;
    dffr reg_Q_2 (.Q (Q[2]), .QB (\$dummy [2]), .D (nx135), .CLK (nx675), .R (
         rst)) ;
    nand02 ix136 (.Y (nx135), .A0 (nx443), .A1 (nx445)) ;
    nand02 ix444 (.Y (nx443), .A0 (Q[2]), .A1 (nx685)) ;
    nand02 ix446 (.Y (nx445), .A0 (D[2]), .A1 (nx663)) ;
    dffr reg_Q_3 (.Q (Q[3]), .QB (\$dummy [3]), .D (nx145), .CLK (nx675), .R (
         rst)) ;
    nand02 ix146 (.Y (nx145), .A0 (nx450), .A1 (nx452)) ;
    nand02 ix451 (.Y (nx450), .A0 (Q[3]), .A1 (nx685)) ;
    nand02 ix453 (.Y (nx452), .A0 (D[3]), .A1 (nx663)) ;
    dffr reg_Q_4 (.Q (Q[4]), .QB (\$dummy [4]), .D (nx155), .CLK (nx675), .R (
         rst)) ;
    nand02 ix156 (.Y (nx155), .A0 (nx457), .A1 (nx459)) ;
    nand02 ix458 (.Y (nx457), .A0 (Q[4]), .A1 (nx685)) ;
    nand02 ix460 (.Y (nx459), .A0 (D[4]), .A1 (nx663)) ;
    dffr reg_Q_5 (.Q (Q[5]), .QB (\$dummy [5]), .D (nx165), .CLK (nx675), .R (
         rst)) ;
    nand02 ix166 (.Y (nx165), .A0 (nx464), .A1 (nx466)) ;
    nand02 ix465 (.Y (nx464), .A0 (Q[5]), .A1 (nx685)) ;
    nand02 ix467 (.Y (nx466), .A0 (D[5]), .A1 (nx663)) ;
    dffr reg_Q_6 (.Q (Q[6]), .QB (\$dummy [6]), .D (nx175), .CLK (nx675), .R (
         rst)) ;
    nand02 ix176 (.Y (nx175), .A0 (nx471), .A1 (nx473)) ;
    nand02 ix472 (.Y (nx471), .A0 (Q[6]), .A1 (nx685)) ;
    nand02 ix474 (.Y (nx473), .A0 (D[6]), .A1 (nx663)) ;
    dffr reg_Q_7 (.Q (Q[7]), .QB (\$dummy [7]), .D (nx185), .CLK (nx677), .R (
         rst)) ;
    nand02 ix186 (.Y (nx185), .A0 (nx478), .A1 (nx480)) ;
    nand02 ix479 (.Y (nx478), .A0 (Q[7]), .A1 (nx651)) ;
    nand02 ix481 (.Y (nx480), .A0 (D[7]), .A1 (nx665)) ;
    dffr reg_Q_8 (.Q (Q[8]), .QB (\$dummy [8]), .D (nx195), .CLK (nx677), .R (
         rst)) ;
    nand02 ix196 (.Y (nx195), .A0 (nx485), .A1 (nx487)) ;
    nand02 ix486 (.Y (nx485), .A0 (Q[8]), .A1 (nx651)) ;
    nand02 ix488 (.Y (nx487), .A0 (D[8]), .A1 (nx665)) ;
    dffr reg_Q_9 (.Q (Q[9]), .QB (\$dummy [9]), .D (nx205), .CLK (nx677), .R (
         rst)) ;
    nand02 ix206 (.Y (nx205), .A0 (nx492), .A1 (nx494)) ;
    nand02 ix493 (.Y (nx492), .A0 (Q[9]), .A1 (nx651)) ;
    nand02 ix495 (.Y (nx494), .A0 (D[9]), .A1 (nx665)) ;
    dffr reg_Q_10 (.Q (Q[10]), .QB (\$dummy [10]), .D (nx215), .CLK (nx677), .R (
         rst)) ;
    nand02 ix216 (.Y (nx215), .A0 (nx499), .A1 (nx501)) ;
    nand02 ix500 (.Y (nx499), .A0 (Q[10]), .A1 (nx651)) ;
    nand02 ix502 (.Y (nx501), .A0 (D[10]), .A1 (nx665)) ;
    dffr reg_Q_11 (.Q (Q[11]), .QB (\$dummy [11]), .D (nx225), .CLK (nx677), .R (
         rst)) ;
    nand02 ix226 (.Y (nx225), .A0 (nx506), .A1 (nx508)) ;
    nand02 ix507 (.Y (nx506), .A0 (Q[11]), .A1 (nx651)) ;
    nand02 ix509 (.Y (nx508), .A0 (D[11]), .A1 (nx665)) ;
    dffr reg_Q_12 (.Q (Q[12]), .QB (\$dummy [12]), .D (nx235), .CLK (nx677), .R (
         rst)) ;
    nand02 ix236 (.Y (nx235), .A0 (nx513), .A1 (nx515)) ;
    nand02 ix514 (.Y (nx513), .A0 (Q[12]), .A1 (nx651)) ;
    nand02 ix516 (.Y (nx515), .A0 (D[12]), .A1 (nx665)) ;
    dffr reg_Q_13 (.Q (Q[13]), .QB (\$dummy [13]), .D (nx245), .CLK (nx677), .R (
         rst)) ;
    nand02 ix246 (.Y (nx245), .A0 (nx520), .A1 (nx522)) ;
    nand02 ix521 (.Y (nx520), .A0 (Q[13]), .A1 (nx651)) ;
    nand02 ix523 (.Y (nx522), .A0 (D[13]), .A1 (nx665)) ;
    dffr reg_Q_14 (.Q (Q[14]), .QB (\$dummy [14]), .D (nx255), .CLK (nx679), .R (
         rst)) ;
    nand02 ix256 (.Y (nx255), .A0 (nx527), .A1 (nx529)) ;
    nand02 ix528 (.Y (nx527), .A0 (Q[14]), .A1 (nx653)) ;
    nand02 ix530 (.Y (nx529), .A0 (D[14]), .A1 (nx667)) ;
    dffr reg_Q_15 (.Q (Q[15]), .QB (\$dummy [15]), .D (nx265), .CLK (nx679), .R (
         rst)) ;
    nand02 ix266 (.Y (nx265), .A0 (nx534), .A1 (nx536)) ;
    nand02 ix535 (.Y (nx534), .A0 (Q[15]), .A1 (nx653)) ;
    nand02 ix537 (.Y (nx536), .A0 (D[15]), .A1 (nx667)) ;
    dffr reg_Q_16 (.Q (Q[16]), .QB (\$dummy [16]), .D (nx275), .CLK (nx679), .R (
         rst)) ;
    nand02 ix276 (.Y (nx275), .A0 (nx541), .A1 (nx543)) ;
    nand02 ix542 (.Y (nx541), .A0 (Q[16]), .A1 (nx653)) ;
    nand02 ix544 (.Y (nx543), .A0 (D[16]), .A1 (nx667)) ;
    dffr reg_Q_17 (.Q (Q[17]), .QB (\$dummy [17]), .D (nx285), .CLK (nx679), .R (
         rst)) ;
    nand02 ix286 (.Y (nx285), .A0 (nx548), .A1 (nx550)) ;
    nand02 ix549 (.Y (nx548), .A0 (Q[17]), .A1 (nx653)) ;
    nand02 ix551 (.Y (nx550), .A0 (D[17]), .A1 (nx667)) ;
    dffr reg_Q_18 (.Q (Q[18]), .QB (\$dummy [18]), .D (nx295), .CLK (nx679), .R (
         rst)) ;
    nand02 ix296 (.Y (nx295), .A0 (nx555), .A1 (nx557)) ;
    nand02 ix556 (.Y (nx555), .A0 (Q[18]), .A1 (nx653)) ;
    nand02 ix558 (.Y (nx557), .A0 (D[18]), .A1 (nx667)) ;
    dffr reg_Q_19 (.Q (Q[19]), .QB (\$dummy [19]), .D (nx305), .CLK (nx679), .R (
         rst)) ;
    nand02 ix306 (.Y (nx305), .A0 (nx562), .A1 (nx564)) ;
    nand02 ix563 (.Y (nx562), .A0 (Q[19]), .A1 (nx653)) ;
    nand02 ix565 (.Y (nx564), .A0 (D[19]), .A1 (nx667)) ;
    dffr reg_Q_20 (.Q (Q[20]), .QB (\$dummy [20]), .D (nx315), .CLK (nx679), .R (
         rst)) ;
    nand02 ix316 (.Y (nx315), .A0 (nx569), .A1 (nx571)) ;
    nand02 ix570 (.Y (nx569), .A0 (Q[20]), .A1 (nx653)) ;
    nand02 ix572 (.Y (nx571), .A0 (D[20]), .A1 (nx667)) ;
    dffr reg_Q_21 (.Q (Q[21]), .QB (\$dummy [21]), .D (nx325), .CLK (nx681), .R (
         rst)) ;
    nand02 ix326 (.Y (nx325), .A0 (nx576), .A1 (nx578)) ;
    nand02 ix577 (.Y (nx576), .A0 (Q[21]), .A1 (nx655)) ;
    nand02 ix579 (.Y (nx578), .A0 (D[21]), .A1 (nx669)) ;
    dffr reg_Q_22 (.Q (Q[22]), .QB (\$dummy [22]), .D (nx335), .CLK (nx681), .R (
         rst)) ;
    nand02 ix336 (.Y (nx335), .A0 (nx583), .A1 (nx585)) ;
    nand02 ix584 (.Y (nx583), .A0 (Q[22]), .A1 (nx655)) ;
    nand02 ix586 (.Y (nx585), .A0 (D[22]), .A1 (nx669)) ;
    dffr reg_Q_23 (.Q (Q[23]), .QB (\$dummy [23]), .D (nx345), .CLK (nx681), .R (
         rst)) ;
    nand02 ix346 (.Y (nx345), .A0 (nx590), .A1 (nx592)) ;
    nand02 ix591 (.Y (nx590), .A0 (Q[23]), .A1 (nx655)) ;
    nand02 ix593 (.Y (nx592), .A0 (D[23]), .A1 (nx669)) ;
    dffr reg_Q_24 (.Q (Q[24]), .QB (\$dummy [24]), .D (nx355), .CLK (nx681), .R (
         rst)) ;
    nand02 ix356 (.Y (nx355), .A0 (nx597), .A1 (nx599)) ;
    nand02 ix598 (.Y (nx597), .A0 (Q[24]), .A1 (nx655)) ;
    nand02 ix600 (.Y (nx599), .A0 (D[24]), .A1 (nx669)) ;
    dffr reg_Q_25 (.Q (Q[25]), .QB (\$dummy [25]), .D (nx365), .CLK (nx681), .R (
         rst)) ;
    nand02 ix366 (.Y (nx365), .A0 (nx604), .A1 (nx606)) ;
    nand02 ix605 (.Y (nx604), .A0 (Q[25]), .A1 (nx655)) ;
    nand02 ix607 (.Y (nx606), .A0 (D[25]), .A1 (nx669)) ;
    dffr reg_Q_26 (.Q (Q[26]), .QB (\$dummy [26]), .D (nx375), .CLK (nx681), .R (
         rst)) ;
    nand02 ix376 (.Y (nx375), .A0 (nx611), .A1 (nx613)) ;
    nand02 ix612 (.Y (nx611), .A0 (Q[26]), .A1 (nx655)) ;
    nand02 ix614 (.Y (nx613), .A0 (D[26]), .A1 (nx669)) ;
    dffr reg_Q_27 (.Q (Q[27]), .QB (\$dummy [27]), .D (nx385), .CLK (nx681), .R (
         rst)) ;
    nand02 ix386 (.Y (nx385), .A0 (nx618), .A1 (nx620)) ;
    nand02 ix619 (.Y (nx618), .A0 (Q[27]), .A1 (nx655)) ;
    nand02 ix621 (.Y (nx620), .A0 (D[27]), .A1 (nx669)) ;
    dffr reg_Q_28 (.Q (Q[28]), .QB (\$dummy [28]), .D (nx395), .CLK (nx683), .R (
         rst)) ;
    nand02 ix396 (.Y (nx395), .A0 (nx625), .A1 (nx627)) ;
    nand02 ix626 (.Y (nx625), .A0 (Q[28]), .A1 (nx657)) ;
    nand02 ix628 (.Y (nx627), .A0 (D[28]), .A1 (nx671)) ;
    dffr reg_Q_29 (.Q (Q[29]), .QB (\$dummy [29]), .D (nx405), .CLK (nx683), .R (
         rst)) ;
    nand02 ix406 (.Y (nx405), .A0 (nx632), .A1 (nx634)) ;
    nand02 ix633 (.Y (nx632), .A0 (Q[29]), .A1 (nx657)) ;
    nand02 ix635 (.Y (nx634), .A0 (D[29]), .A1 (nx671)) ;
    dffr reg_Q_30 (.Q (Q[30]), .QB (\$dummy [30]), .D (nx415), .CLK (nx683), .R (
         rst)) ;
    nand02 ix416 (.Y (nx415), .A0 (nx639), .A1 (nx641)) ;
    nand02 ix640 (.Y (nx639), .A0 (Q[30]), .A1 (nx657)) ;
    nand02 ix642 (.Y (nx641), .A0 (D[30]), .A1 (nx671)) ;
    inv02 ix648 (.Y (nx649), .A (en)) ;
    inv02 ix650 (.Y (nx651), .A (nx671)) ;
    inv02 ix652 (.Y (nx653), .A (nx671)) ;
    inv02 ix654 (.Y (nx655), .A (nx671)) ;
    inv02 ix656 (.Y (nx657), .A (nx671)) ;
    inv02 ix662 (.Y (nx663), .A (nx649)) ;
    inv02 ix664 (.Y (nx665), .A (nx649)) ;
    inv02 ix666 (.Y (nx667), .A (nx649)) ;
    inv02 ix668 (.Y (nx669), .A (nx649)) ;
    inv02 ix670 (.Y (nx671), .A (nx649)) ;
    inv01 ix672 (.Y (nx673), .A (clk)) ;
    inv02 ix674 (.Y (nx675), .A (nx673)) ;
    inv02 ix676 (.Y (nx677), .A (nx673)) ;
    inv02 ix678 (.Y (nx679), .A (nx673)) ;
    inv02 ix680 (.Y (nx681), .A (nx673)) ;
    inv02 ix682 (.Y (nx683), .A (nx673)) ;
    inv02 ix684 (.Y (nx685), .A (en)) ;
endmodule

